magic
tech sky130B
magscale 1 2
timestamp 1662734359
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 484394 700680 484400 700732
rect 484452 700720 484458 700732
rect 543458 700720 543464 700732
rect 484452 700692 543464 700720
rect 484452 700680 484458 700692
rect 543458 700680 543464 700692
rect 543516 700680 543522 700732
rect 283834 700612 283840 700664
rect 283892 700652 283898 700664
rect 381538 700652 381544 700664
rect 283892 700624 381544 700652
rect 283892 700612 283898 700624
rect 381538 700612 381544 700624
rect 381596 700612 381602 700664
rect 400122 700612 400128 700664
rect 400180 700652 400186 700664
rect 527174 700652 527180 700664
rect 400180 700624 527180 700652
rect 400180 700612 400186 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 218974 700544 218980 700596
rect 219032 700584 219038 700596
rect 347222 700584 347228 700596
rect 219032 700556 347228 700584
rect 219032 700544 219038 700556
rect 347222 700544 347228 700556
rect 347280 700544 347286 700596
rect 413646 700544 413652 700596
rect 413704 700584 413710 700596
rect 551278 700584 551284 700596
rect 413704 700556 551284 700584
rect 413704 700544 413710 700556
rect 551278 700544 551284 700556
rect 551336 700544 551342 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 347130 700516 347136 700528
rect 105504 700488 347136 700516
rect 105504 700476 105510 700488
rect 347130 700476 347136 700488
rect 347188 700476 347194 700528
rect 404998 700476 405004 700528
rect 405056 700516 405062 700528
rect 559650 700516 559656 700528
rect 405056 700488 559656 700516
rect 405056 700476 405062 700488
rect 559650 700476 559656 700488
rect 559708 700476 559714 700528
rect 202782 700408 202788 700460
rect 202840 700448 202846 700460
rect 498194 700448 498200 700460
rect 202840 700420 498200 700448
rect 202840 700408 202846 700420
rect 498194 700408 498200 700420
rect 498252 700408 498258 700460
rect 267642 700340 267648 700392
rect 267700 700380 267706 700392
rect 564710 700380 564716 700392
rect 267700 700352 564716 700380
rect 267700 700340 267706 700352
rect 564710 700340 564716 700352
rect 564768 700340 564774 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 567194 700312 567200 700324
rect 24360 700284 567200 700312
rect 24360 700272 24366 700284
rect 567194 700272 567200 700284
rect 567252 700272 567258 700324
rect 137830 698912 137836 698964
rect 137888 698952 137894 698964
rect 374822 698952 374828 698964
rect 137888 698924 374828 698952
rect 137888 698912 137894 698924
rect 374822 698912 374828 698924
rect 374880 698912 374886 698964
rect 429838 698912 429844 698964
rect 429896 698952 429902 698964
rect 550910 698952 550916 698964
rect 429896 698924 550916 698952
rect 429896 698912 429902 698924
rect 550910 698912 550916 698924
rect 550968 698912 550974 698964
rect 153194 694764 153200 694816
rect 153252 694804 153258 694816
rect 552934 694804 552940 694816
rect 153252 694776 552940 694804
rect 153252 694764 153258 694776
rect 552934 694764 552940 694776
rect 552992 694764 552998 694816
rect 71774 690616 71780 690668
rect 71832 690656 71838 690668
rect 399938 690656 399944 690668
rect 71832 690628 399944 690656
rect 71832 690616 71838 690628
rect 399938 690616 399944 690628
rect 399996 690616 400002 690668
rect 462314 690616 462320 690668
rect 462372 690656 462378 690668
rect 550266 690656 550272 690668
rect 462372 690628 550272 690656
rect 462372 690616 462378 690628
rect 550266 690616 550272 690628
rect 550324 690616 550330 690668
rect 331214 689324 331220 689376
rect 331272 689364 331278 689376
rect 400858 689364 400864 689376
rect 331272 689336 400864 689364
rect 331272 689324 331278 689336
rect 400858 689324 400864 689336
rect 400916 689324 400922 689376
rect 364334 689256 364340 689308
rect 364392 689296 364398 689308
rect 550358 689296 550364 689308
rect 364392 689268 550364 689296
rect 364392 689256 364398 689268
rect 550358 689256 550364 689268
rect 550416 689256 550422 689308
rect 299474 687964 299480 688016
rect 299532 688004 299538 688016
rect 551094 688004 551100 688016
rect 299532 687976 551100 688004
rect 299532 687964 299538 687976
rect 551094 687964 551100 687976
rect 551152 687964 551158 688016
rect 234614 687896 234620 687948
rect 234672 687936 234678 687948
rect 538214 687936 538220 687948
rect 234672 687908 538220 687936
rect 234672 687896 234678 687908
rect 538214 687896 538220 687908
rect 538272 687896 538278 687948
rect 405090 687488 405096 687540
rect 405148 687528 405154 687540
rect 554130 687528 554136 687540
rect 405148 687500 554136 687528
rect 405148 687488 405154 687500
rect 554130 687488 554136 687500
rect 554188 687488 554194 687540
rect 403986 687420 403992 687472
rect 404044 687460 404050 687472
rect 553946 687460 553952 687472
rect 404044 687432 553952 687460
rect 404044 687420 404050 687432
rect 553946 687420 553952 687432
rect 554004 687420 554010 687472
rect 396902 687352 396908 687404
rect 396960 687392 396966 687404
rect 554222 687392 554228 687404
rect 396960 687364 554228 687392
rect 396960 687352 396966 687364
rect 554222 687352 554228 687364
rect 554280 687352 554286 687404
rect 407022 687284 407028 687336
rect 407080 687324 407086 687336
rect 569954 687324 569960 687336
rect 407080 687296 569960 687324
rect 407080 687284 407086 687296
rect 569954 687284 569960 687296
rect 570012 687284 570018 687336
rect 413462 687216 413468 687268
rect 413520 687256 413526 687268
rect 582374 687256 582380 687268
rect 413520 687228 582380 687256
rect 413520 687216 413526 687228
rect 582374 687216 582380 687228
rect 582432 687216 582438 687268
rect 347774 686536 347780 686588
rect 347832 686576 347838 686588
rect 568758 686576 568764 686588
rect 347832 686548 568764 686576
rect 347832 686536 347838 686548
rect 568758 686536 568764 686548
rect 568816 686536 568822 686588
rect 6914 686468 6920 686520
rect 6972 686508 6978 686520
rect 549990 686508 549996 686520
rect 6972 686480 549996 686508
rect 6972 686468 6978 686480
rect 549990 686468 549996 686480
rect 550048 686468 550054 686520
rect 384942 686128 384948 686180
rect 385000 686168 385006 686180
rect 446398 686168 446404 686180
rect 385000 686140 446404 686168
rect 385000 686128 385006 686140
rect 446398 686128 446404 686140
rect 446456 686128 446462 686180
rect 407666 686060 407672 686112
rect 407724 686100 407730 686112
rect 553762 686100 553768 686112
rect 407724 686072 553768 686100
rect 407724 686060 407730 686072
rect 553762 686060 553768 686072
rect 553820 686060 553826 686112
rect 402790 685992 402796 686044
rect 402848 686032 402854 686044
rect 554038 686032 554044 686044
rect 402848 686004 554044 686032
rect 402848 685992 402854 686004
rect 554038 685992 554044 686004
rect 554096 685992 554102 686044
rect 363598 685924 363604 685976
rect 363656 685964 363662 685976
rect 528830 685964 528836 685976
rect 363656 685936 528836 685964
rect 363656 685924 363662 685936
rect 528830 685924 528836 685936
rect 528888 685924 528894 685976
rect 405182 685856 405188 685908
rect 405240 685896 405246 685908
rect 580902 685896 580908 685908
rect 405240 685868 580908 685896
rect 405240 685856 405246 685868
rect 580902 685856 580908 685868
rect 580960 685856 580966 685908
rect 402330 685516 402336 685568
rect 402388 685556 402394 685568
rect 468386 685556 468392 685568
rect 402388 685528 468392 685556
rect 402388 685516 402394 685528
rect 468386 685516 468392 685528
rect 468444 685516 468450 685568
rect 407574 685448 407580 685500
rect 407632 685488 407638 685500
rect 456794 685488 456800 685500
rect 407632 685460 456800 685488
rect 407632 685448 407638 685460
rect 456794 685448 456800 685460
rect 456852 685448 456858 685500
rect 173158 685380 173164 685432
rect 173216 685420 173222 685432
rect 514754 685420 514760 685432
rect 173216 685392 514760 685420
rect 173216 685380 173222 685392
rect 514754 685380 514760 685392
rect 514812 685380 514818 685432
rect 409690 685312 409696 685364
rect 409748 685352 409754 685364
rect 450262 685352 450268 685364
rect 409748 685324 450268 685352
rect 409748 685312 409754 685324
rect 450262 685312 450268 685324
rect 450320 685312 450326 685364
rect 409046 685244 409052 685296
rect 409104 685284 409110 685296
rect 454218 685284 454224 685296
rect 409104 685256 454224 685284
rect 409104 685244 409110 685256
rect 454218 685244 454224 685256
rect 454276 685244 454282 685296
rect 407758 685176 407764 685228
rect 407816 685216 407822 685228
rect 470870 685216 470876 685228
rect 407816 685188 470876 685216
rect 407816 685176 407822 685188
rect 470870 685176 470876 685188
rect 470928 685176 470934 685228
rect 407850 685108 407856 685160
rect 407908 685148 407914 685160
rect 509234 685148 509240 685160
rect 407908 685120 509240 685148
rect 407908 685108 407914 685120
rect 509234 685108 509240 685120
rect 509292 685108 509298 685160
rect 468294 685040 468300 685092
rect 468352 685080 468358 685092
rect 571334 685080 571340 685092
rect 468352 685052 571340 685080
rect 468352 685040 468358 685052
rect 571334 685040 571340 685052
rect 571392 685040 571398 685092
rect 362218 684972 362224 685024
rect 362276 685012 362282 685024
rect 473538 685012 473544 685024
rect 362276 684984 473544 685012
rect 362276 684972 362282 684984
rect 473538 684972 473544 684984
rect 473596 684972 473602 685024
rect 487614 684972 487620 685024
rect 487672 685012 487678 685024
rect 582466 685012 582472 685024
rect 487672 684984 582472 685012
rect 487672 684972 487678 684984
rect 582466 684972 582472 684984
rect 582524 684972 582530 685024
rect 359458 684904 359464 684956
rect 359516 684944 359522 684956
rect 470594 684944 470600 684956
rect 359516 684916 470600 684944
rect 359516 684904 359522 684916
rect 470594 684904 470600 684916
rect 470652 684904 470658 684956
rect 476482 684904 476488 684956
rect 476540 684944 476546 684956
rect 581086 684944 581092 684956
rect 476540 684916 581092 684944
rect 476540 684904 476546 684916
rect 581086 684904 581092 684916
rect 581144 684904 581150 684956
rect 409138 684836 409144 684888
rect 409196 684876 409202 684888
rect 523034 684876 523040 684888
rect 409196 684848 523040 684876
rect 409196 684836 409202 684848
rect 523034 684836 523040 684848
rect 523092 684836 523098 684888
rect 453850 684768 453856 684820
rect 453908 684808 453914 684820
rect 576854 684808 576860 684820
rect 453908 684780 576860 684808
rect 453908 684768 453914 684780
rect 576854 684768 576860 684780
rect 576912 684768 576918 684820
rect 409322 684700 409328 684752
rect 409380 684740 409386 684752
rect 535454 684740 535460 684752
rect 409380 684712 535460 684740
rect 409380 684700 409386 684712
rect 535454 684700 535460 684712
rect 535512 684700 535518 684752
rect 406654 684632 406660 684684
rect 406712 684672 406718 684684
rect 552474 684672 552480 684684
rect 406712 684644 552480 684672
rect 406712 684632 406718 684644
rect 552474 684632 552480 684644
rect 552532 684632 552538 684684
rect 388714 684564 388720 684616
rect 388772 684604 388778 684616
rect 539134 684604 539140 684616
rect 388772 684576 539140 684604
rect 388772 684564 388778 684576
rect 539134 684564 539140 684576
rect 539192 684564 539198 684616
rect 405274 684496 405280 684548
rect 405332 684536 405338 684548
rect 437566 684536 437572 684548
rect 405332 684508 437572 684536
rect 405332 684496 405338 684508
rect 437566 684496 437572 684508
rect 437624 684496 437630 684548
rect 489546 684496 489552 684548
rect 489604 684536 489610 684548
rect 580994 684536 581000 684548
rect 489604 684508 581000 684536
rect 489604 684496 489610 684508
rect 580994 684496 581000 684508
rect 581052 684496 581058 684548
rect 21358 684020 21364 684072
rect 21416 684060 21422 684072
rect 502518 684060 502524 684072
rect 21416 684032 502524 684060
rect 21416 684020 21422 684032
rect 502518 684020 502524 684032
rect 502576 684020 502582 684072
rect 409230 683952 409236 684004
rect 409288 683992 409294 684004
rect 497274 683992 497280 684004
rect 409288 683964 497280 683992
rect 409288 683952 409294 683964
rect 497274 683952 497280 683964
rect 497332 683952 497338 684004
rect 400030 683884 400036 683936
rect 400088 683924 400094 683936
rect 521838 683924 521844 683936
rect 400088 683896 521844 683924
rect 400088 683884 400094 683896
rect 521838 683884 521844 683896
rect 521896 683884 521902 683936
rect 407942 683816 407948 683868
rect 408000 683856 408006 683868
rect 436094 683856 436100 683868
rect 408000 683828 436100 683856
rect 408000 683816 408006 683828
rect 436094 683816 436100 683828
rect 436152 683816 436158 683868
rect 438670 683816 438676 683868
rect 438728 683856 438734 683868
rect 567930 683856 567936 683868
rect 438728 683828 567936 683856
rect 438728 683816 438734 683828
rect 567930 683816 567936 683828
rect 567988 683816 567994 683868
rect 429010 683748 429016 683800
rect 429068 683788 429074 683800
rect 563698 683788 563704 683800
rect 429068 683760 563704 683788
rect 429068 683748 429074 683760
rect 563698 683748 563704 683760
rect 563756 683748 563762 683800
rect 392578 683680 392584 683732
rect 392636 683720 392642 683732
rect 429654 683720 429660 683732
rect 392636 683692 429660 683720
rect 392636 683680 392642 683692
rect 429654 683680 429660 683692
rect 429712 683680 429718 683732
rect 435450 683680 435456 683732
rect 435508 683720 435514 683732
rect 572806 683720 572812 683732
rect 435508 683692 572812 683720
rect 435508 683680 435514 683692
rect 572806 683680 572812 683692
rect 572864 683680 572870 683732
rect 408126 683612 408132 683664
rect 408184 683652 408190 683664
rect 550634 683652 550640 683664
rect 408184 683624 550640 683652
rect 408184 683612 408190 683624
rect 550634 683612 550640 683624
rect 550692 683612 550698 683664
rect 398098 683544 398104 683596
rect 398156 683584 398162 683596
rect 545574 683584 545580 683596
rect 398156 683556 545580 683584
rect 398156 683544 398162 683556
rect 545574 683544 545580 683556
rect 545632 683544 545638 683596
rect 404262 683476 404268 683528
rect 404320 683516 404326 683528
rect 555234 683516 555240 683528
rect 404320 683488 555240 683516
rect 404320 683476 404326 683488
rect 555234 683476 555240 683488
rect 555292 683476 555298 683528
rect 416682 683408 416688 683460
rect 416740 683448 416746 683460
rect 573634 683448 573640 683460
rect 416740 683420 573640 683448
rect 416740 683408 416746 683420
rect 573634 683408 573640 683420
rect 573692 683408 573698 683460
rect 408310 683340 408316 683392
rect 408368 683380 408374 683392
rect 581178 683380 581184 683392
rect 408368 683352 581184 683380
rect 408368 683340 408374 683352
rect 581178 683340 581184 683352
rect 581236 683340 581242 683392
rect 406838 683272 406844 683324
rect 406896 683312 406902 683324
rect 580350 683312 580356 683324
rect 406896 683284 580356 683312
rect 406896 683272 406902 683284
rect 580350 683272 580356 683284
rect 580408 683272 580414 683324
rect 31018 683204 31024 683256
rect 31076 683244 31082 683256
rect 509510 683244 509516 683256
rect 31076 683216 509516 683244
rect 31076 683204 31082 683216
rect 509510 683204 509516 683216
rect 509568 683204 509574 683256
rect 409414 683136 409420 683188
rect 409472 683176 409478 683188
rect 424594 683176 424600 683188
rect 409472 683148 424600 683176
rect 409472 683136 409478 683148
rect 424594 683136 424600 683148
rect 424652 683136 424658 683188
rect 510522 683136 510528 683188
rect 510580 683176 510586 683188
rect 579154 683176 579160 683188
rect 510580 683148 579160 683176
rect 510580 683136 510586 683148
rect 579154 683136 579160 683148
rect 579212 683136 579218 683188
rect 3418 682660 3424 682712
rect 3476 682700 3482 682712
rect 550450 682700 550456 682712
rect 3476 682672 550456 682700
rect 3476 682660 3482 682672
rect 550450 682660 550456 682672
rect 550508 682660 550514 682712
rect 529658 682592 529664 682644
rect 529716 682632 529722 682644
rect 551462 682632 551468 682644
rect 529716 682604 551468 682632
rect 529716 682592 529722 682604
rect 551462 682592 551468 682604
rect 551520 682592 551526 682644
rect 26142 682524 26148 682576
rect 26200 682564 26206 682576
rect 532694 682564 532700 682576
rect 26200 682536 532700 682564
rect 26200 682524 26206 682536
rect 532694 682524 532700 682536
rect 532752 682524 532758 682576
rect 495158 682456 495164 682508
rect 495216 682496 495222 682508
rect 551554 682496 551560 682508
rect 495216 682468 551560 682496
rect 495216 682456 495222 682468
rect 551554 682456 551560 682468
rect 551612 682456 551618 682508
rect 402238 682388 402244 682440
rect 402296 682428 402302 682440
rect 440418 682428 440424 682440
rect 402296 682400 440424 682428
rect 402296 682388 402302 682400
rect 440418 682388 440424 682400
rect 440476 682388 440482 682440
rect 477494 682388 477500 682440
rect 477552 682428 477558 682440
rect 567286 682428 567292 682440
rect 477552 682400 567292 682428
rect 477552 682388 477558 682400
rect 567286 682388 567292 682400
rect 567344 682388 567350 682440
rect 382918 682320 382924 682372
rect 382976 682360 382982 682372
rect 422386 682360 422392 682372
rect 382976 682332 422392 682360
rect 382976 682320 382982 682332
rect 422386 682320 422392 682332
rect 422444 682320 422450 682372
rect 502242 682320 502248 682372
rect 502300 682360 502306 682372
rect 561030 682360 561036 682372
rect 502300 682332 561036 682360
rect 502300 682320 502306 682332
rect 561030 682320 561036 682332
rect 561088 682320 561094 682372
rect 389818 682252 389824 682304
rect 389876 682292 389882 682304
rect 480346 682292 480352 682304
rect 389876 682264 480352 682292
rect 389876 682252 389882 682264
rect 480346 682252 480352 682264
rect 480404 682252 480410 682304
rect 484854 682252 484860 682304
rect 484912 682292 484918 682304
rect 575474 682292 575480 682304
rect 484912 682264 575480 682292
rect 484912 682252 484918 682264
rect 575474 682252 575480 682264
rect 575532 682252 575538 682304
rect 397362 682184 397368 682236
rect 397420 682224 397426 682236
rect 442258 682224 442264 682236
rect 397420 682196 442264 682224
rect 397420 682184 397426 682196
rect 442258 682184 442264 682196
rect 442316 682184 442322 682236
rect 458174 682184 458180 682236
rect 458232 682224 458238 682236
rect 554866 682224 554872 682236
rect 458232 682196 554872 682224
rect 458232 682184 458238 682196
rect 554866 682184 554872 682196
rect 554924 682184 554930 682236
rect 373902 682116 373908 682168
rect 373960 682156 373966 682168
rect 416590 682156 416596 682168
rect 373960 682128 416596 682156
rect 373960 682116 373966 682128
rect 416590 682116 416596 682128
rect 416648 682116 416654 682168
rect 432874 682116 432880 682168
rect 432932 682156 432938 682168
rect 570598 682156 570604 682168
rect 432932 682128 570604 682156
rect 432932 682116 432938 682128
rect 570598 682116 570604 682128
rect 570656 682116 570662 682168
rect 408034 682048 408040 682100
rect 408092 682088 408098 682100
rect 547782 682088 547788 682100
rect 408092 682060 547788 682088
rect 408092 682048 408098 682060
rect 547782 682048 547788 682060
rect 547840 682048 547846 682100
rect 549898 682048 549904 682100
rect 549956 682088 549962 682100
rect 574094 682088 574100 682100
rect 549956 682060 574100 682088
rect 549956 682048 549962 682060
rect 574094 682048 574100 682060
rect 574152 682048 574158 682100
rect 384390 681980 384396 682032
rect 384448 682020 384454 682032
rect 530118 682020 530124 682032
rect 384448 681992 530124 682020
rect 384448 681980 384454 681992
rect 530118 681980 530124 681992
rect 530176 681980 530182 682032
rect 537846 681980 537852 682032
rect 537904 682020 537910 682032
rect 565906 682020 565912 682032
rect 537904 681992 565912 682020
rect 537904 681980 537910 681992
rect 565906 681980 565912 681992
rect 565964 681980 565970 682032
rect 380158 681912 380164 681964
rect 380216 681952 380222 681964
rect 545114 681952 545120 681964
rect 380216 681924 545120 681952
rect 380216 681912 380222 681924
rect 545114 681912 545120 681924
rect 545172 681912 545178 681964
rect 548794 681912 548800 681964
rect 548852 681952 548858 681964
rect 576946 681952 576952 681964
rect 548852 681924 576952 681952
rect 548852 681912 548858 681924
rect 576946 681912 576952 681924
rect 577004 681912 577010 681964
rect 409506 681844 409512 681896
rect 409564 681884 409570 681896
rect 580442 681884 580448 681896
rect 409564 681856 580448 681884
rect 409564 681844 409570 681856
rect 580442 681844 580448 681856
rect 580500 681844 580506 681896
rect 17770 681776 17776 681828
rect 17828 681816 17834 681828
rect 411622 681816 411628 681828
rect 17828 681788 411628 681816
rect 17828 681776 17834 681788
rect 411622 681776 411628 681788
rect 411680 681776 411686 681828
rect 512730 681776 512736 681828
rect 512788 681816 512794 681828
rect 577222 681816 577228 681828
rect 512788 681788 577228 681816
rect 512788 681776 512794 681788
rect 577222 681776 577228 681788
rect 577280 681776 577286 681828
rect 389082 681708 389088 681760
rect 389140 681748 389146 681760
rect 412910 681748 412916 681760
rect 389140 681720 412916 681748
rect 389140 681708 389146 681720
rect 412910 681708 412916 681720
rect 412968 681708 412974 681760
rect 440050 681708 440056 681760
rect 440108 681748 440114 681760
rect 458174 681748 458180 681760
rect 440108 681720 458180 681748
rect 440108 681708 440114 681720
rect 458174 681708 458180 681720
rect 458232 681708 458238 681760
rect 541710 681708 541716 681760
rect 541768 681748 541774 681760
rect 577498 681748 577504 681760
rect 541768 681720 577504 681748
rect 541768 681708 541774 681720
rect 577498 681708 577504 681720
rect 577556 681708 577562 681760
rect 8938 681300 8944 681352
rect 8996 681340 9002 681352
rect 552106 681340 552112 681352
rect 8996 681312 552112 681340
rect 8996 681300 9002 681312
rect 552106 681300 552112 681312
rect 552164 681300 552170 681352
rect 406562 681232 406568 681284
rect 406620 681272 406626 681284
rect 457346 681272 457352 681284
rect 406620 681244 457352 681272
rect 406620 681232 406626 681244
rect 457346 681232 457352 681244
rect 457404 681232 457410 681284
rect 501782 681232 501788 681284
rect 501840 681272 501846 681284
rect 574738 681272 574744 681284
rect 501840 681244 574744 681272
rect 501840 681232 501846 681244
rect 574738 681232 574744 681244
rect 574796 681232 574802 681284
rect 377398 681164 377404 681216
rect 377456 681204 377462 681216
rect 419994 681204 420000 681216
rect 377456 681176 420000 681204
rect 377456 681164 377462 681176
rect 419994 681164 420000 681176
rect 420052 681164 420058 681216
rect 427814 681164 427820 681216
rect 427872 681204 427878 681216
rect 504358 681204 504364 681216
rect 427872 681176 504364 681204
rect 427872 681164 427878 681176
rect 504358 681164 504364 681176
rect 504416 681164 504422 681216
rect 517238 681164 517244 681216
rect 517296 681204 517302 681216
rect 572898 681204 572904 681216
rect 517296 681176 572904 681204
rect 517296 681164 517302 681176
rect 572898 681164 572904 681176
rect 572956 681164 572962 681216
rect 403710 681096 403716 681148
rect 403768 681136 403774 681148
rect 463786 681136 463792 681148
rect 403768 681108 463792 681136
rect 403768 681096 403774 681108
rect 463786 681096 463792 681108
rect 463844 681096 463850 681148
rect 499206 681096 499212 681148
rect 499264 681136 499270 681148
rect 580258 681136 580264 681148
rect 499264 681108 580264 681136
rect 499264 681096 499270 681108
rect 580258 681096 580264 681108
rect 580316 681096 580322 681148
rect 408218 681028 408224 681080
rect 408276 681068 408282 681080
rect 408276 681040 431954 681068
rect 408276 681028 408282 681040
rect 400950 680960 400956 681012
rect 401008 681000 401014 681012
rect 427906 681000 427912 681012
rect 401008 680972 427912 681000
rect 401008 680960 401014 680972
rect 427906 680960 427912 680972
rect 427964 680960 427970 681012
rect 431926 681000 431954 681040
rect 439314 681028 439320 681080
rect 439372 681068 439378 681080
rect 439372 681040 440188 681068
rect 439372 681028 439378 681040
rect 440050 681000 440056 681012
rect 431926 680972 440056 681000
rect 440050 680960 440056 680972
rect 440108 680960 440114 681012
rect 440160 681000 440188 681040
rect 440326 681028 440332 681080
rect 440384 681068 440390 681080
rect 524414 681068 524420 681080
rect 440384 681040 524420 681068
rect 440384 681028 440390 681040
rect 524414 681028 524420 681040
rect 524472 681028 524478 681080
rect 547782 681028 547788 681080
rect 547840 681068 547846 681080
rect 555326 681068 555332 681080
rect 547840 681040 555332 681068
rect 547840 681028 547846 681040
rect 555326 681028 555332 681040
rect 555384 681028 555390 681080
rect 551002 681000 551008 681012
rect 440160 680972 551008 681000
rect 551002 680960 551008 680972
rect 551060 680960 551066 681012
rect 347038 680892 347044 680944
rect 347096 680932 347102 680944
rect 432046 680932 432052 680944
rect 347096 680904 432052 680932
rect 347096 680892 347102 680904
rect 432046 680892 432052 680904
rect 432104 680892 432110 680944
rect 434622 680892 434628 680944
rect 434680 680932 434686 680944
rect 550726 680932 550732 680944
rect 434680 680904 550732 680932
rect 434680 680892 434686 680904
rect 550726 680892 550732 680904
rect 550784 680892 550790 680944
rect 409598 680824 409604 680876
rect 409656 680864 409662 680876
rect 552382 680864 552388 680876
rect 409656 680836 552388 680864
rect 409656 680824 409662 680836
rect 552382 680824 552388 680836
rect 552440 680824 552446 680876
rect 408954 680756 408960 680808
rect 409012 680796 409018 680808
rect 552198 680796 552204 680808
rect 409012 680768 552204 680796
rect 409012 680756 409018 680768
rect 552198 680756 552204 680768
rect 552256 680756 552262 680808
rect 409874 680688 409880 680740
rect 409932 680728 409938 680740
rect 553486 680728 553492 680740
rect 409932 680700 553492 680728
rect 409932 680688 409938 680700
rect 553486 680688 553492 680700
rect 553544 680688 553550 680740
rect 403802 680620 403808 680672
rect 403860 680660 403866 680672
rect 553394 680660 553400 680672
rect 403860 680632 553400 680660
rect 403860 680620 403866 680632
rect 553394 680620 553400 680632
rect 553452 680620 553458 680672
rect 405458 680552 405464 680604
rect 405516 680592 405522 680604
rect 580626 680592 580632 680604
rect 405516 680564 580632 680592
rect 405516 680552 405522 680564
rect 580626 680552 580632 680564
rect 580684 680552 580690 680604
rect 402514 680484 402520 680536
rect 402572 680524 402578 680536
rect 580718 680524 580724 680536
rect 402572 680496 580724 680524
rect 402572 680484 402578 680496
rect 580718 680484 580724 680496
rect 580776 680484 580782 680536
rect 173250 680416 173256 680468
rect 173308 680456 173314 680468
rect 461210 680456 461216 680468
rect 173308 680428 461216 680456
rect 173308 680416 173314 680428
rect 461210 680416 461216 680428
rect 461268 680416 461274 680468
rect 496630 680416 496636 680468
rect 496688 680456 496694 680468
rect 577130 680456 577136 680468
rect 496688 680428 577136 680456
rect 496688 680416 496694 680428
rect 577130 680416 577136 680428
rect 577188 680416 577194 680468
rect 427078 680348 427084 680400
rect 427136 680388 427142 680400
rect 440142 680388 440148 680400
rect 427136 680360 440148 680388
rect 427136 680348 427142 680360
rect 440142 680348 440148 680360
rect 440200 680348 440206 680400
rect 402422 679600 402428 679652
rect 402480 679640 402486 679652
rect 427078 679640 427084 679652
rect 402480 679612 427084 679640
rect 402480 679600 402486 679612
rect 427078 679600 427084 679612
rect 427136 679600 427142 679652
rect 440142 679600 440148 679652
rect 440200 679640 440206 679652
rect 580534 679640 580540 679652
rect 440200 679612 580540 679640
rect 440200 679600 440206 679612
rect 580534 679600 580540 679612
rect 580592 679600 580598 679652
rect 399478 679532 399484 679584
rect 399536 679572 399542 679584
rect 553670 679572 553676 679584
rect 399536 679544 553676 679572
rect 399536 679532 399542 679544
rect 553670 679532 553676 679544
rect 553728 679532 553734 679584
rect 409782 679464 409788 679516
rect 409840 679504 409846 679516
rect 449802 679504 449808 679516
rect 409840 679476 449808 679504
rect 409840 679464 409846 679476
rect 449802 679464 449808 679476
rect 449860 679464 449866 679516
rect 511442 679464 511448 679516
rect 511500 679504 511506 679516
rect 577038 679504 577044 679516
rect 511500 679476 577044 679504
rect 511500 679464 511506 679476
rect 577038 679464 577044 679476
rect 577096 679464 577102 679516
rect 408402 679396 408408 679448
rect 408460 679436 408466 679448
rect 553118 679436 553124 679448
rect 408460 679408 553124 679436
rect 408460 679396 408466 679408
rect 553118 679396 553124 679408
rect 553176 679396 553182 679448
rect 406470 679328 406476 679380
rect 406528 679368 406534 679380
rect 551922 679368 551928 679380
rect 406528 679340 551928 679368
rect 406528 679328 406534 679340
rect 551922 679328 551928 679340
rect 551980 679328 551986 679380
rect 405550 679260 405556 679312
rect 405608 679300 405614 679312
rect 551186 679300 551192 679312
rect 405608 679272 551192 679300
rect 405608 679260 405614 679272
rect 551186 679260 551192 679272
rect 551244 679260 551250 679312
rect 404906 679192 404912 679244
rect 404964 679232 404970 679244
rect 552566 679232 552572 679244
rect 404964 679204 552572 679232
rect 404964 679192 404970 679204
rect 552566 679192 552572 679204
rect 552624 679192 552630 679244
rect 402606 679124 402612 679176
rect 402664 679164 402670 679176
rect 553854 679164 553860 679176
rect 402664 679136 553860 679164
rect 402664 679124 402670 679136
rect 553854 679124 553860 679136
rect 553912 679124 553918 679176
rect 552014 679056 552020 679108
rect 552072 679096 552078 679108
rect 582834 679096 582840 679108
rect 552072 679068 582840 679096
rect 552072 679056 552078 679068
rect 582834 679056 582840 679068
rect 582892 679056 582898 679108
rect 395430 678988 395436 679040
rect 395488 679028 395494 679040
rect 580810 679028 580816 679040
rect 395488 679000 580816 679028
rect 395488 678988 395494 679000
rect 580810 678988 580816 679000
rect 580868 678988 580874 679040
rect 408034 678512 408040 678564
rect 408092 678552 408098 678564
rect 408310 678552 408316 678564
rect 408092 678524 408316 678552
rect 408092 678512 408098 678524
rect 408310 678512 408316 678524
rect 408368 678512 408374 678564
rect 407850 678376 407856 678428
rect 407908 678416 407914 678428
rect 408034 678416 408040 678428
rect 407908 678388 408040 678416
rect 407908 678376 407914 678388
rect 408034 678376 408040 678388
rect 408092 678376 408098 678428
rect 399846 678240 399852 678292
rect 399904 678280 399910 678292
rect 409874 678280 409880 678292
rect 399904 678252 409880 678280
rect 399904 678240 399910 678252
rect 409874 678240 409880 678252
rect 409932 678240 409938 678292
rect 407574 678172 407580 678224
rect 407632 678212 407638 678224
rect 407758 678212 407764 678224
rect 407632 678184 407764 678212
rect 407632 678172 407638 678184
rect 407758 678172 407764 678184
rect 407816 678172 407822 678224
rect 552014 678104 552020 678156
rect 552072 678144 552078 678156
rect 552290 678144 552296 678156
rect 552072 678116 552296 678144
rect 552072 678104 552078 678116
rect 552290 678104 552296 678116
rect 552348 678104 552354 678156
rect 7558 677560 7564 677612
rect 7616 677600 7622 677612
rect 407114 677600 407120 677612
rect 7616 677572 407120 677600
rect 7616 677560 7622 677572
rect 407114 677560 407120 677572
rect 407172 677560 407178 677612
rect 552014 677560 552020 677612
rect 552072 677600 552078 677612
rect 579614 677600 579620 677612
rect 552072 677572 579620 677600
rect 552072 677560 552078 677572
rect 579614 677560 579620 677572
rect 579672 677560 579678 677612
rect 40034 676812 40040 676864
rect 40092 676852 40098 676864
rect 396994 676852 397000 676864
rect 40092 676824 397000 676852
rect 40092 676812 40098 676824
rect 396994 676812 397000 676824
rect 397052 676812 397058 676864
rect 551554 676540 551560 676592
rect 551612 676580 551618 676592
rect 552750 676580 552756 676592
rect 551612 676552 552756 676580
rect 551612 676540 551618 676552
rect 552750 676540 552756 676552
rect 552808 676540 552814 676592
rect 166902 676132 166908 676184
rect 166960 676172 166966 676184
rect 169754 676172 169760 676184
rect 166960 676144 169760 676172
rect 166960 676132 166966 676144
rect 169754 676132 169760 676144
rect 169812 676172 169818 676184
rect 340874 676172 340880 676184
rect 169812 676144 340880 676172
rect 169812 676132 169818 676144
rect 340874 676132 340880 676144
rect 340932 676132 340938 676184
rect 340874 674976 340880 675028
rect 340932 675016 340938 675028
rect 351178 675016 351184 675028
rect 340932 674988 351184 675016
rect 340932 674976 340938 674988
rect 351178 674976 351184 674988
rect 351236 674976 351242 675028
rect 328546 674908 328552 674960
rect 328604 674948 328610 674960
rect 347774 674948 347780 674960
rect 328604 674920 347780 674948
rect 328604 674908 328610 674920
rect 347774 674908 347780 674920
rect 347832 674908 347838 674960
rect 154482 674840 154488 674892
rect 154540 674880 154546 674892
rect 172698 674880 172704 674892
rect 154540 674852 172704 674880
rect 154540 674840 154546 674852
rect 172698 674840 172704 674852
rect 172756 674840 172762 674892
rect 329742 674840 329748 674892
rect 329800 674880 329806 674892
rect 361574 674880 361580 674892
rect 329800 674852 361580 674880
rect 329800 674840 329806 674852
rect 361574 674840 361580 674852
rect 361632 674840 361638 674892
rect 552014 674840 552020 674892
rect 552072 674880 552078 674892
rect 575658 674880 575664 674892
rect 552072 674852 575664 674880
rect 552072 674840 552078 674852
rect 575658 674840 575664 674852
rect 575716 674840 575722 674892
rect 552198 674160 552204 674212
rect 552256 674160 552262 674212
rect 550174 674092 550180 674144
rect 550232 674132 550238 674144
rect 550450 674132 550456 674144
rect 550232 674104 550456 674132
rect 550232 674092 550238 674104
rect 550450 674092 550456 674104
rect 550508 674092 550514 674144
rect 550818 674092 550824 674144
rect 550876 674132 550882 674144
rect 551370 674132 551376 674144
rect 550876 674104 551376 674132
rect 550876 674092 550882 674104
rect 551370 674092 551376 674104
rect 551428 674092 551434 674144
rect 552216 674008 552244 674160
rect 552198 673956 552204 674008
rect 552256 673956 552262 674008
rect 552014 672052 552020 672104
rect 552072 672092 552078 672104
rect 571610 672092 571616 672104
rect 552072 672064 571616 672092
rect 552072 672052 552078 672064
rect 571610 672052 571616 672064
rect 571668 672052 571674 672104
rect 347222 670624 347228 670676
rect 347280 670664 347286 670676
rect 407114 670664 407120 670676
rect 347280 670636 407120 670664
rect 347280 670624 347286 670636
rect 407114 670624 407120 670636
rect 407172 670624 407178 670676
rect 383010 667904 383016 667956
rect 383068 667944 383074 667956
rect 407114 667944 407120 667956
rect 383068 667916 407120 667944
rect 383068 667904 383074 667916
rect 407114 667904 407120 667916
rect 407172 667904 407178 667956
rect 553302 666544 553308 666596
rect 553360 666584 553366 666596
rect 566734 666584 566740 666596
rect 553360 666556 566740 666584
rect 553360 666544 553366 666556
rect 566734 666544 566740 666556
rect 566792 666544 566798 666596
rect 385678 665184 385684 665236
rect 385736 665224 385742 665236
rect 407114 665224 407120 665236
rect 385736 665196 407120 665224
rect 385736 665184 385742 665196
rect 407114 665184 407120 665196
rect 407172 665184 407178 665236
rect 397454 663688 397460 663740
rect 397512 663728 397518 663740
rect 407206 663728 407212 663740
rect 397512 663700 407212 663728
rect 397512 663688 397518 663700
rect 407206 663688 407212 663700
rect 407264 663688 407270 663740
rect 393958 661172 393964 661224
rect 394016 661212 394022 661224
rect 407298 661212 407304 661224
rect 394016 661184 407304 661212
rect 394016 661172 394022 661184
rect 407298 661172 407304 661184
rect 407356 661172 407362 661224
rect 387242 661104 387248 661156
rect 387300 661144 387306 661156
rect 407206 661144 407212 661156
rect 387300 661116 407212 661144
rect 387300 661104 387306 661116
rect 407206 661104 407212 661116
rect 407264 661104 407270 661156
rect 348786 661036 348792 661088
rect 348844 661076 348850 661088
rect 407390 661076 407396 661088
rect 348844 661048 407396 661076
rect 348844 661036 348850 661048
rect 407390 661036 407396 661048
rect 407448 661036 407454 661088
rect 404722 658248 404728 658300
rect 404780 658288 404786 658300
rect 407298 658288 407304 658300
rect 404780 658260 407304 658288
rect 404780 658248 404786 658260
rect 407298 658248 407304 658260
rect 407356 658248 407362 658300
rect 3326 658180 3332 658232
rect 3384 658220 3390 658232
rect 8938 658220 8944 658232
rect 3384 658192 8944 658220
rect 3384 658180 3390 658192
rect 8938 658180 8944 658192
rect 8996 658180 9002 658232
rect 553302 656888 553308 656940
rect 553360 656928 553366 656940
rect 558914 656928 558920 656940
rect 553360 656900 558920 656928
rect 553360 656888 553366 656900
rect 558914 656888 558920 656900
rect 558972 656888 558978 656940
rect 347130 655460 347136 655512
rect 347188 655500 347194 655512
rect 407206 655500 407212 655512
rect 347188 655472 407212 655500
rect 347188 655460 347194 655472
rect 407206 655460 407212 655472
rect 407264 655460 407270 655512
rect 404078 654168 404084 654220
rect 404136 654208 404142 654220
rect 407206 654208 407212 654220
rect 404136 654180 407212 654208
rect 404136 654168 404142 654180
rect 407206 654168 407212 654180
rect 407264 654168 407270 654220
rect 552106 653216 552112 653268
rect 552164 653256 552170 653268
rect 554958 653256 554964 653268
rect 552164 653228 554964 653256
rect 552164 653216 552170 653228
rect 554958 653216 554964 653228
rect 555016 653216 555022 653268
rect 376018 652740 376024 652792
rect 376076 652780 376082 652792
rect 407206 652780 407212 652792
rect 376076 652752 407212 652780
rect 376076 652740 376082 652752
rect 407206 652740 407212 652752
rect 407264 652740 407270 652792
rect 351178 650632 351184 650684
rect 351236 650672 351242 650684
rect 402698 650672 402704 650684
rect 351236 650644 402704 650672
rect 351236 650632 351242 650644
rect 402698 650632 402704 650644
rect 402756 650672 402762 650684
rect 407206 650672 407212 650684
rect 402756 650644 407212 650672
rect 402756 650632 402762 650644
rect 407206 650632 407212 650644
rect 407264 650632 407270 650684
rect 367830 648592 367836 648644
rect 367888 648632 367894 648644
rect 407206 648632 407212 648644
rect 367888 648604 407212 648632
rect 367888 648592 367894 648604
rect 407206 648592 407212 648604
rect 407264 648592 407270 648644
rect 553302 648592 553308 648644
rect 553360 648632 553366 648644
rect 564526 648632 564532 648644
rect 553360 648604 564532 648632
rect 553360 648592 553366 648604
rect 564526 648592 564532 648604
rect 564584 648592 564590 648644
rect 552566 645872 552572 645924
rect 552624 645912 552630 645924
rect 556430 645912 556436 645924
rect 552624 645884 556436 645912
rect 552624 645872 552630 645884
rect 556430 645872 556436 645884
rect 556488 645872 556494 645924
rect 553210 644648 553216 644700
rect 553268 644688 553274 644700
rect 556798 644688 556804 644700
rect 553268 644660 556804 644688
rect 553268 644648 553274 644660
rect 556798 644648 556804 644660
rect 556856 644648 556862 644700
rect 402882 644444 402888 644496
rect 402940 644484 402946 644496
rect 407206 644484 407212 644496
rect 402940 644456 407212 644484
rect 402940 644444 402946 644456
rect 407206 644444 407212 644456
rect 407264 644444 407270 644496
rect 552106 644444 552112 644496
rect 552164 644484 552170 644496
rect 565262 644484 565268 644496
rect 552164 644456 565268 644484
rect 552164 644444 552170 644456
rect 565262 644444 565268 644456
rect 565320 644444 565326 644496
rect 570690 643084 570696 643136
rect 570748 643124 570754 643136
rect 579982 643124 579988 643136
rect 570748 643096 579988 643124
rect 570748 643084 570754 643096
rect 579982 643084 579988 643096
rect 580040 643084 580046 643136
rect 552014 642540 552020 642592
rect 552072 642580 552078 642592
rect 554222 642580 554228 642592
rect 552072 642552 554228 642580
rect 552072 642540 552078 642552
rect 554222 642540 554228 642552
rect 554280 642540 554286 642592
rect 347130 641724 347136 641776
rect 347188 641764 347194 641776
rect 407206 641764 407212 641776
rect 347188 641736 407212 641764
rect 347188 641724 347194 641736
rect 407206 641724 407212 641736
rect 407264 641724 407270 641776
rect 358078 640296 358084 640348
rect 358136 640336 358142 640348
rect 407206 640336 407212 640348
rect 358136 640308 407212 640336
rect 358136 640296 358142 640308
rect 407206 640296 407212 640308
rect 407264 640296 407270 640348
rect 553302 640296 553308 640348
rect 553360 640336 553366 640348
rect 574278 640336 574284 640348
rect 553360 640308 574284 640336
rect 553360 640296 553366 640308
rect 574278 640296 574284 640308
rect 574336 640296 574342 640348
rect 552106 637848 552112 637900
rect 552164 637888 552170 637900
rect 557810 637888 557816 637900
rect 552164 637860 557816 637888
rect 552164 637848 552170 637860
rect 557810 637848 557816 637860
rect 557868 637848 557874 637900
rect 404170 637644 404176 637696
rect 404228 637684 404234 637696
rect 407298 637684 407304 637696
rect 404228 637656 407304 637684
rect 404228 637644 404234 637656
rect 407298 637644 407304 637656
rect 407356 637644 407362 637696
rect 393222 637576 393228 637628
rect 393280 637616 393286 637628
rect 407206 637616 407212 637628
rect 393280 637588 407212 637616
rect 393280 637576 393286 637588
rect 407206 637576 407212 637588
rect 407264 637576 407270 637628
rect 552014 637576 552020 637628
rect 552072 637616 552078 637628
rect 562594 637616 562600 637628
rect 552072 637588 562600 637616
rect 552072 637576 552078 637588
rect 562594 637576 562600 637588
rect 562652 637576 562658 637628
rect 383562 636216 383568 636268
rect 383620 636256 383626 636268
rect 407206 636256 407212 636268
rect 383620 636228 407212 636256
rect 383620 636216 383626 636228
rect 407206 636216 407212 636228
rect 407264 636216 407270 636268
rect 408310 635536 408316 635588
rect 408368 635536 408374 635588
rect 408328 635384 408356 635536
rect 408310 635332 408316 635384
rect 408368 635332 408374 635384
rect 367738 633428 367744 633480
rect 367796 633468 367802 633480
rect 407206 633468 407212 633480
rect 367796 633440 407212 633468
rect 367796 633428 367802 633440
rect 407206 633428 407212 633440
rect 407264 633428 407270 633480
rect 360838 632068 360844 632120
rect 360896 632108 360902 632120
rect 407206 632108 407212 632120
rect 360896 632080 407212 632108
rect 360896 632068 360902 632080
rect 407206 632068 407212 632080
rect 407264 632068 407270 632120
rect 556798 632000 556804 632052
rect 556856 632040 556862 632052
rect 580166 632040 580172 632052
rect 556856 632012 580172 632040
rect 556856 632000 556862 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 552014 631184 552020 631236
rect 552072 631224 552078 631236
rect 554222 631224 554228 631236
rect 552072 631196 554228 631224
rect 552072 631184 552078 631196
rect 554222 631184 554228 631196
rect 554280 631184 554286 631236
rect 408218 628600 408224 628652
rect 408276 628640 408282 628652
rect 408402 628640 408408 628652
rect 408276 628612 408408 628640
rect 408276 628600 408282 628612
rect 408402 628600 408408 628612
rect 408460 628600 408466 628652
rect 395338 627920 395344 627972
rect 395396 627960 395402 627972
rect 407206 627960 407212 627972
rect 395396 627932 407212 627960
rect 395396 627920 395402 627932
rect 407206 627920 407212 627932
rect 407264 627920 407270 627972
rect 552014 625336 552020 625388
rect 552072 625376 552078 625388
rect 557074 625376 557080 625388
rect 552072 625348 557080 625376
rect 552072 625336 552078 625348
rect 557074 625336 557080 625348
rect 557132 625336 557138 625388
rect 552014 623772 552020 623824
rect 552072 623812 552078 623824
rect 582650 623812 582656 623824
rect 552072 623784 582656 623812
rect 552072 623772 552078 623784
rect 582650 623772 582656 623784
rect 582708 623772 582714 623824
rect 552566 619624 552572 619676
rect 552624 619664 552630 619676
rect 576118 619664 576124 619676
rect 552624 619636 576124 619664
rect 552624 619624 552630 619636
rect 576118 619624 576124 619636
rect 576176 619624 576182 619676
rect 396718 618332 396724 618384
rect 396776 618372 396782 618384
rect 407298 618372 407304 618384
rect 396776 618344 407304 618372
rect 396776 618332 396782 618344
rect 407298 618332 407304 618344
rect 407356 618332 407362 618384
rect 387426 618264 387432 618316
rect 387484 618304 387490 618316
rect 407206 618304 407212 618316
rect 387484 618276 407212 618304
rect 387484 618264 387490 618276
rect 407206 618264 407212 618276
rect 407264 618264 407270 618316
rect 553302 616836 553308 616888
rect 553360 616876 553366 616888
rect 576302 616876 576308 616888
rect 553360 616848 576308 616876
rect 553360 616836 553366 616848
rect 576302 616836 576308 616848
rect 576360 616836 576366 616888
rect 371878 615476 371884 615528
rect 371936 615516 371942 615528
rect 407298 615516 407304 615528
rect 371936 615488 407304 615516
rect 371936 615476 371942 615488
rect 407298 615476 407304 615488
rect 407356 615476 407362 615528
rect 553302 612824 553308 612876
rect 553360 612864 553366 612876
rect 558546 612864 558552 612876
rect 553360 612836 558552 612864
rect 553360 612824 553366 612836
rect 558546 612824 558552 612836
rect 558604 612824 558610 612876
rect 399754 612756 399760 612808
rect 399812 612796 399818 612808
rect 407206 612796 407212 612808
rect 399812 612768 407212 612796
rect 399812 612756 399818 612768
rect 407206 612756 407212 612768
rect 407264 612756 407270 612808
rect 553210 612756 553216 612808
rect 553268 612796 553274 612808
rect 578878 612796 578884 612808
rect 553268 612768 578884 612796
rect 553268 612756 553274 612768
rect 578878 612756 578884 612768
rect 578936 612756 578942 612808
rect 553302 611328 553308 611380
rect 553360 611368 553366 611380
rect 569402 611368 569408 611380
rect 553360 611340 569408 611368
rect 553360 611328 553366 611340
rect 569402 611328 569408 611340
rect 569460 611328 569466 611380
rect 553302 609968 553308 610020
rect 553360 610008 553366 610020
rect 571978 610008 571984 610020
rect 553360 609980 571984 610008
rect 553360 609968 553366 609980
rect 571978 609968 571984 609980
rect 572036 609968 572042 610020
rect 350442 608608 350448 608660
rect 350500 608648 350506 608660
rect 368474 608648 368480 608660
rect 350500 608620 368480 608648
rect 350500 608608 350506 608620
rect 368474 608608 368480 608620
rect 368532 608608 368538 608660
rect 381630 608608 381636 608660
rect 381688 608648 381694 608660
rect 407206 608648 407212 608660
rect 381688 608620 407212 608648
rect 381688 608608 381694 608620
rect 407206 608608 407212 608620
rect 407264 608608 407270 608660
rect 552474 608608 552480 608660
rect 552532 608648 552538 608660
rect 555694 608648 555700 608660
rect 552532 608620 555700 608648
rect 552532 608608 552538 608620
rect 555694 608608 555700 608620
rect 555752 608608 555758 608660
rect 552198 607248 552204 607300
rect 552256 607288 552262 607300
rect 555050 607288 555056 607300
rect 552256 607260 555056 607288
rect 552256 607248 552262 607260
rect 555050 607248 555056 607260
rect 555108 607248 555114 607300
rect 176562 607180 176568 607232
rect 176620 607220 176626 607232
rect 209038 607220 209044 607232
rect 176620 607192 209044 607220
rect 176620 607180 176626 607192
rect 209038 607180 209044 607192
rect 209096 607180 209102 607232
rect 176562 605820 176568 605872
rect 176620 605860 176626 605872
rect 203518 605860 203524 605872
rect 176620 605832 203524 605860
rect 176620 605820 176626 605832
rect 203518 605820 203524 605832
rect 203576 605820 203582 605872
rect 350442 605820 350448 605872
rect 350500 605860 350506 605872
rect 371234 605860 371240 605872
rect 350500 605832 371240 605860
rect 350500 605820 350506 605832
rect 371234 605820 371240 605832
rect 371292 605820 371298 605872
rect 350442 604460 350448 604512
rect 350500 604500 350506 604512
rect 364334 604500 364340 604512
rect 350500 604472 364340 604500
rect 350500 604460 350506 604472
rect 364334 604460 364340 604472
rect 364392 604460 364398 604512
rect 552014 603916 552020 603968
rect 552072 603956 552078 603968
rect 554866 603956 554872 603968
rect 552072 603928 554872 603956
rect 552072 603916 552078 603928
rect 554866 603916 554872 603928
rect 554924 603916 554930 603968
rect 553302 603100 553308 603152
rect 553360 603140 553366 603152
rect 582558 603140 582564 603152
rect 553360 603112 582564 603140
rect 553360 603100 553366 603112
rect 582558 603100 582564 603112
rect 582616 603100 582622 603152
rect 404262 603032 404268 603084
rect 404320 603072 404326 603084
rect 407298 603072 407304 603084
rect 404320 603044 407304 603072
rect 404320 603032 404326 603044
rect 407298 603032 407304 603044
rect 407356 603032 407362 603084
rect 366358 601672 366364 601724
rect 366416 601712 366422 601724
rect 407298 601712 407304 601724
rect 366416 601684 407304 601712
rect 366416 601672 366422 601684
rect 407298 601672 407304 601684
rect 407356 601672 407362 601724
rect 174538 598952 174544 599004
rect 174596 598992 174602 599004
rect 207014 598992 207020 599004
rect 174596 598964 207020 598992
rect 174596 598952 174602 598964
rect 207014 598952 207020 598964
rect 207072 598952 207078 599004
rect 374638 598952 374644 599004
rect 374696 598992 374702 599004
rect 407298 598992 407304 599004
rect 374696 598964 407304 598992
rect 374696 598952 374702 598964
rect 407298 598952 407304 598964
rect 407356 598952 407362 599004
rect 553302 598952 553308 599004
rect 553360 598992 553366 599004
rect 560478 598992 560484 599004
rect 553360 598964 560484 598992
rect 553360 598952 553366 598964
rect 560478 598952 560484 598964
rect 560536 598952 560542 599004
rect 394602 596164 394608 596216
rect 394660 596204 394666 596216
rect 407298 596204 407304 596216
rect 394660 596176 407304 596204
rect 394660 596164 394666 596176
rect 407298 596164 407304 596176
rect 407356 596164 407362 596216
rect 398742 594804 398748 594856
rect 398800 594844 398806 594856
rect 407298 594844 407304 594856
rect 398800 594816 407304 594844
rect 398800 594804 398806 594816
rect 407298 594804 407304 594816
rect 407356 594804 407362 594856
rect 34146 593512 34152 593564
rect 34204 593552 34210 593564
rect 34330 593552 34336 593564
rect 34204 593524 34336 593552
rect 34204 593512 34210 593524
rect 34330 593512 34336 593524
rect 34388 593512 34394 593564
rect 404262 592016 404268 592068
rect 404320 592056 404326 592068
rect 407298 592056 407304 592068
rect 404320 592028 407304 592056
rect 404320 592016 404326 592028
rect 407298 592016 407304 592028
rect 407356 592016 407362 592068
rect 404814 590860 404820 590912
rect 404872 590900 404878 590912
rect 405182 590900 405188 590912
rect 404872 590872 405188 590900
rect 404872 590860 404878 590872
rect 405182 590860 405188 590872
rect 405240 590860 405246 590912
rect 405182 590724 405188 590776
rect 405240 590764 405246 590776
rect 407390 590764 407396 590776
rect 405240 590736 407396 590764
rect 405240 590724 405246 590736
rect 407390 590724 407396 590736
rect 407448 590724 407454 590776
rect 401502 590656 401508 590708
rect 401560 590696 401566 590708
rect 407298 590696 407304 590708
rect 401560 590668 407304 590696
rect 401560 590656 401566 590668
rect 407298 590656 407304 590668
rect 407356 590656 407362 590708
rect 34146 589976 34152 590028
rect 34204 590016 34210 590028
rect 209130 590016 209136 590028
rect 34204 589988 209136 590016
rect 34204 589976 34210 589988
rect 209130 589976 209136 589988
rect 209188 589976 209194 590028
rect 34054 589908 34060 589960
rect 34112 589948 34118 589960
rect 36446 589948 36452 589960
rect 34112 589920 36452 589948
rect 34112 589908 34118 589920
rect 36446 589908 36452 589920
rect 36504 589908 36510 589960
rect 33962 589840 33968 589892
rect 34020 589880 34026 589892
rect 36538 589880 36544 589892
rect 34020 589852 36544 589880
rect 34020 589840 34026 589852
rect 36538 589840 36544 589852
rect 36596 589840 36602 589892
rect 47578 589228 47584 589280
rect 47636 589268 47642 589280
rect 207750 589268 207756 589280
rect 47636 589240 207756 589268
rect 47636 589228 47642 589240
rect 207750 589228 207756 589240
rect 207808 589228 207814 589280
rect 239306 589228 239312 589280
rect 239364 589268 239370 589280
rect 402330 589268 402336 589280
rect 239364 589240 402336 589268
rect 239364 589228 239370 589240
rect 402330 589228 402336 589240
rect 402388 589228 402394 589280
rect 39850 589160 39856 589212
rect 39908 589200 39914 589212
rect 207658 589200 207664 589212
rect 39908 589172 207664 589200
rect 39908 589160 39914 589172
rect 207658 589160 207664 589172
rect 207716 589160 207722 589212
rect 225138 589160 225144 589212
rect 225196 589200 225202 589212
rect 404906 589200 404912 589212
rect 225196 589172 404912 589200
rect 225196 589160 225202 589172
rect 404906 589160 404912 589172
rect 404964 589160 404970 589212
rect 140774 589092 140780 589144
rect 140832 589132 140838 589144
rect 349338 589132 349344 589144
rect 140832 589104 349344 589132
rect 140832 589092 140838 589104
rect 349338 589092 349344 589104
rect 349396 589092 349402 589144
rect 35618 589024 35624 589076
rect 35676 589064 35682 589076
rect 78858 589064 78864 589076
rect 35676 589036 78864 589064
rect 35676 589024 35682 589036
rect 78858 589024 78864 589036
rect 78916 589024 78922 589076
rect 86034 589024 86040 589076
rect 86092 589064 86098 589076
rect 402606 589064 402612 589076
rect 86092 589036 402612 589064
rect 86092 589024 86098 589036
rect 402606 589024 402612 589036
rect 402664 589024 402670 589076
rect 39390 588956 39396 589008
rect 39448 588996 39454 589008
rect 402422 588996 402428 589008
rect 39448 588968 402428 588996
rect 39448 588956 39454 588968
rect 402422 588956 402428 588968
rect 402480 588956 402486 589008
rect 552106 588956 552112 589008
rect 552164 588996 552170 589008
rect 554130 588996 554136 589008
rect 552164 588968 554136 588996
rect 552164 588956 552170 588968
rect 554130 588956 554136 588968
rect 554188 588956 554194 589008
rect 42058 588888 42064 588940
rect 42116 588928 42122 588940
rect 405274 588928 405280 588940
rect 42116 588900 405280 588928
rect 42116 588888 42122 588900
rect 405274 588888 405280 588900
rect 405332 588888 405338 588940
rect 40770 588820 40776 588872
rect 40828 588860 40834 588872
rect 405090 588860 405096 588872
rect 40828 588832 405096 588860
rect 40828 588820 40834 588832
rect 405090 588820 405096 588832
rect 405148 588820 405154 588872
rect 40862 588752 40868 588804
rect 40920 588792 40926 588804
rect 405550 588792 405556 588804
rect 40920 588764 405556 588792
rect 40920 588752 40926 588764
rect 405550 588752 405556 588764
rect 405608 588752 405614 588804
rect 35342 588684 35348 588736
rect 35400 588724 35406 588736
rect 405182 588724 405188 588736
rect 35400 588696 405188 588724
rect 35400 588684 35406 588696
rect 405182 588684 405188 588696
rect 405240 588684 405246 588736
rect 32766 588616 32772 588668
rect 32824 588656 32830 588668
rect 406746 588656 406752 588668
rect 32824 588628 406752 588656
rect 32824 588616 32830 588628
rect 406746 588616 406752 588628
rect 406804 588616 406810 588668
rect 3510 588548 3516 588600
rect 3568 588588 3574 588600
rect 399662 588588 399668 588600
rect 3568 588560 399668 588588
rect 3568 588548 3574 588560
rect 399662 588548 399668 588560
rect 399720 588548 399726 588600
rect 43714 588480 43720 588532
rect 43772 588520 43778 588532
rect 172698 588520 172704 588532
rect 43772 588492 172704 588520
rect 43772 588480 43778 588492
rect 172698 588480 172704 588492
rect 172756 588480 172762 588532
rect 292758 588480 292764 588532
rect 292816 588520 292822 588532
rect 399478 588520 399484 588532
rect 292816 588492 399484 588520
rect 292816 588480 292822 588492
rect 399478 588480 399484 588492
rect 399536 588480 399542 588532
rect 317414 588412 317420 588464
rect 317472 588452 317478 588464
rect 347774 588452 347780 588464
rect 317472 588424 347780 588452
rect 317472 588412 317478 588424
rect 347774 588412 347780 588424
rect 347832 588412 347838 588464
rect 393130 587868 393136 587920
rect 393188 587908 393194 587920
rect 407298 587908 407304 587920
rect 393188 587880 407304 587908
rect 393188 587868 393194 587880
rect 407298 587868 407304 587880
rect 407356 587868 407362 587920
rect 44726 587528 44732 587580
rect 44784 587568 44790 587580
rect 264422 587568 264428 587580
rect 44784 587540 264428 587568
rect 44784 587528 44790 587540
rect 264422 587528 264428 587540
rect 264480 587528 264486 587580
rect 42518 587460 42524 587512
rect 42576 587500 42582 587512
rect 407298 587500 407304 587512
rect 42576 587472 407304 587500
rect 42576 587460 42582 587472
rect 407298 587460 407304 587472
rect 407356 587460 407362 587512
rect 57882 587392 57888 587444
rect 57940 587432 57946 587444
rect 82078 587432 82084 587444
rect 57940 587404 82084 587432
rect 57940 587392 57946 587404
rect 82078 587392 82084 587404
rect 82136 587392 82142 587444
rect 49050 587324 49056 587376
rect 49108 587364 49114 587376
rect 78674 587364 78680 587376
rect 49108 587336 78680 587364
rect 49108 587324 49114 587336
rect 78674 587324 78680 587336
rect 78732 587324 78738 587376
rect 316034 587324 316040 587376
rect 316092 587364 316098 587376
rect 350534 587364 350540 587376
rect 316092 587336 350540 587364
rect 316092 587324 316098 587336
rect 350534 587324 350540 587336
rect 350592 587324 350598 587376
rect 33042 587256 33048 587308
rect 33100 587296 33106 587308
rect 71774 587296 71780 587308
rect 33100 587268 71780 587296
rect 33100 587256 33106 587268
rect 71774 587256 71780 587268
rect 71832 587256 71838 587308
rect 308490 587256 308496 587308
rect 308548 587296 308554 587308
rect 354766 587296 354772 587308
rect 308548 587268 354772 587296
rect 308548 587256 308554 587268
rect 354766 587256 354772 587268
rect 354824 587256 354830 587308
rect 37182 587188 37188 587240
rect 37240 587228 37246 587240
rect 81894 587228 81900 587240
rect 37240 587200 81900 587228
rect 37240 587188 37246 587200
rect 81894 587188 81900 587200
rect 81952 587188 81958 587240
rect 291010 587188 291016 587240
rect 291068 587228 291074 587240
rect 352006 587228 352012 587240
rect 291068 587200 352012 587228
rect 291068 587188 291074 587200
rect 352006 587188 352012 587200
rect 352064 587188 352070 587240
rect 45370 587120 45376 587172
rect 45428 587160 45434 587172
rect 95234 587160 95240 587172
rect 45428 587132 95240 587160
rect 45428 587120 45434 587132
rect 95234 587120 95240 587132
rect 95292 587120 95298 587172
rect 286318 587120 286324 587172
rect 286376 587160 286382 587172
rect 348418 587160 348424 587172
rect 286376 587132 348424 587160
rect 286376 587120 286382 587132
rect 348418 587120 348424 587132
rect 348476 587120 348482 587172
rect 34238 587052 34244 587104
rect 34296 587092 34302 587104
rect 101950 587092 101956 587104
rect 34296 587064 101956 587092
rect 34296 587052 34302 587064
rect 101950 587052 101956 587064
rect 102008 587052 102014 587104
rect 281074 587052 281080 587104
rect 281132 587092 281138 587104
rect 350626 587092 350632 587104
rect 281132 587064 350632 587092
rect 281132 587052 281138 587064
rect 350626 587052 350632 587064
rect 350684 587052 350690 587104
rect 22830 586984 22836 587036
rect 22888 587024 22894 587036
rect 106918 587024 106924 587036
rect 22888 586996 106924 587024
rect 22888 586984 22894 586996
rect 106918 586984 106924 586996
rect 106976 586984 106982 587036
rect 261018 586984 261024 587036
rect 261076 587024 261082 587036
rect 356514 587024 356520 587036
rect 261076 586996 356520 587024
rect 261076 586984 261082 586996
rect 356514 586984 356520 586996
rect 356572 586984 356578 587036
rect 45002 586916 45008 586968
rect 45060 586956 45066 586968
rect 131758 586956 131764 586968
rect 45060 586928 131764 586956
rect 45060 586916 45066 586928
rect 131758 586916 131764 586928
rect 131816 586916 131822 586968
rect 248138 586916 248144 586968
rect 248196 586956 248202 586968
rect 348694 586956 348700 586968
rect 248196 586928 348700 586956
rect 248196 586916 248202 586928
rect 348694 586916 348700 586928
rect 348752 586916 348758 586968
rect 41322 586848 41328 586900
rect 41380 586888 41386 586900
rect 139394 586888 139400 586900
rect 41380 586860 139400 586888
rect 41380 586848 41386 586860
rect 139394 586848 139400 586860
rect 139452 586848 139458 586900
rect 141970 586848 141976 586900
rect 142028 586888 142034 586900
rect 163958 586888 163964 586900
rect 142028 586860 163964 586888
rect 142028 586848 142034 586860
rect 163958 586848 163964 586860
rect 164016 586848 164022 586900
rect 256602 586848 256608 586900
rect 256660 586888 256666 586900
rect 359274 586888 359280 586900
rect 256660 586860 359280 586888
rect 256660 586848 256666 586860
rect 359274 586848 359280 586860
rect 359332 586848 359338 586900
rect 22922 586780 22928 586832
rect 22980 586820 22986 586832
rect 124398 586820 124404 586832
rect 22980 586792 124404 586820
rect 22980 586780 22986 586792
rect 124398 586780 124404 586792
rect 124456 586780 124462 586832
rect 124858 586780 124864 586832
rect 124916 586820 124922 586832
rect 133966 586820 133972 586832
rect 124916 586792 133972 586820
rect 124916 586780 124922 586792
rect 133966 586780 133972 586792
rect 134024 586780 134030 586832
rect 153838 586780 153844 586832
rect 153896 586820 153902 586832
rect 227806 586820 227812 586832
rect 153896 586792 227812 586820
rect 153896 586780 153902 586792
rect 227806 586780 227812 586792
rect 227864 586780 227870 586832
rect 240778 586780 240784 586832
rect 240836 586820 240842 586832
rect 348510 586820 348516 586832
rect 240836 586792 348516 586820
rect 240836 586780 240842 586792
rect 348510 586780 348516 586792
rect 348568 586780 348574 586832
rect 77202 586712 77208 586764
rect 77260 586752 77266 586764
rect 180058 586752 180064 586764
rect 77260 586724 180064 586752
rect 77260 586712 77266 586724
rect 180058 586712 180064 586724
rect 180116 586712 180122 586764
rect 209774 586712 209780 586764
rect 209832 586752 209838 586764
rect 238754 586752 238760 586764
rect 209832 586724 238760 586752
rect 209832 586712 209838 586724
rect 238754 586712 238760 586724
rect 238812 586712 238818 586764
rect 242434 586712 242440 586764
rect 242492 586752 242498 586764
rect 357710 586752 357716 586764
rect 242492 586724 357716 586752
rect 242492 586712 242498 586724
rect 357710 586712 357716 586724
rect 357768 586712 357774 586764
rect 245562 586644 245568 586696
rect 245620 586684 245626 586696
rect 361850 586684 361856 586696
rect 245620 586656 361856 586684
rect 245620 586644 245626 586656
rect 361850 586644 361856 586656
rect 361908 586644 361914 586696
rect 48958 586576 48964 586628
rect 49016 586616 49022 586628
rect 245838 586616 245844 586628
rect 49016 586588 245844 586616
rect 49016 586576 49022 586588
rect 245838 586576 245844 586588
rect 245896 586576 245902 586628
rect 260650 586576 260656 586628
rect 260708 586616 260714 586628
rect 361758 586616 361764 586628
rect 260708 586588 361764 586616
rect 260708 586576 260714 586588
rect 361758 586576 361764 586588
rect 361816 586576 361822 586628
rect 31570 586508 31576 586560
rect 31628 586548 31634 586560
rect 81158 586548 81164 586560
rect 31628 586520 81164 586548
rect 31628 586508 31634 586520
rect 81158 586508 81164 586520
rect 81216 586508 81222 586560
rect 333882 586508 333888 586560
rect 333940 586548 333946 586560
rect 348602 586548 348608 586560
rect 333940 586520 348608 586548
rect 333940 586508 333946 586520
rect 348602 586508 348608 586520
rect 348660 586508 348666 586560
rect 553302 586508 553308 586560
rect 553360 586548 553366 586560
rect 578970 586548 578976 586560
rect 553360 586520 578976 586548
rect 553360 586508 553366 586520
rect 578970 586508 578976 586520
rect 579028 586508 579034 586560
rect 273530 586032 273536 586084
rect 273588 586072 273594 586084
rect 306926 586072 306932 586084
rect 273588 586044 306932 586072
rect 273588 586032 273594 586044
rect 306926 586032 306932 586044
rect 306984 586032 306990 586084
rect 47210 585964 47216 586016
rect 47268 586004 47274 586016
rect 240502 586004 240508 586016
rect 47268 585976 240508 586004
rect 47268 585964 47274 585976
rect 240502 585964 240508 585976
rect 240560 585964 240566 586016
rect 265066 585964 265072 586016
rect 265124 586004 265130 586016
rect 298094 586004 298100 586016
rect 265124 585976 298100 586004
rect 265124 585964 265130 585976
rect 298094 585964 298100 585976
rect 298152 585964 298158 586016
rect 320450 585964 320456 586016
rect 320508 586004 320514 586016
rect 348786 586004 348792 586016
rect 320508 585976 348792 586004
rect 320508 585964 320514 585976
rect 348786 585964 348792 585976
rect 348844 585964 348850 586016
rect 81802 585896 81808 585948
rect 81860 585936 81866 585948
rect 349706 585936 349712 585948
rect 81860 585908 349712 585936
rect 81860 585896 81866 585908
rect 349706 585896 349712 585908
rect 349764 585896 349770 585948
rect 66346 585828 66352 585880
rect 66404 585868 66410 585880
rect 356422 585868 356428 585880
rect 66404 585840 356428 585868
rect 66404 585828 66410 585840
rect 356422 585828 356428 585840
rect 356480 585828 356486 585880
rect 100846 585760 100852 585812
rect 100904 585800 100910 585812
rect 405366 585800 405372 585812
rect 100904 585772 405372 585800
rect 100904 585760 100910 585772
rect 405366 585760 405372 585772
rect 405424 585760 405430 585812
rect 200666 585148 200672 585200
rect 200724 585188 200730 585200
rect 376110 585188 376116 585200
rect 200724 585160 376116 585188
rect 200724 585148 200730 585160
rect 376110 585148 376116 585160
rect 376168 585148 376174 585200
rect 552566 585148 552572 585200
rect 552624 585188 552630 585200
rect 571426 585188 571432 585200
rect 552624 585160 571432 585188
rect 552624 585148 552630 585160
rect 571426 585148 571432 585160
rect 571484 585148 571490 585200
rect 215478 584604 215484 584656
rect 215536 584644 215542 584656
rect 282914 584644 282920 584656
rect 215536 584616 282920 584644
rect 215536 584604 215542 584616
rect 282914 584604 282920 584616
rect 282972 584604 282978 584656
rect 307754 584604 307760 584656
rect 307812 584644 307818 584656
rect 349154 584644 349160 584656
rect 307812 584616 349160 584644
rect 307812 584604 307818 584616
rect 349154 584604 349160 584616
rect 349212 584604 349218 584656
rect 115198 584536 115204 584588
rect 115256 584576 115262 584588
rect 211614 584576 211620 584588
rect 115256 584548 211620 584576
rect 115256 584536 115262 584548
rect 211614 584536 211620 584548
rect 211672 584536 211678 584588
rect 269758 584536 269764 584588
rect 269816 584576 269822 584588
rect 346854 584576 346860 584588
rect 269816 584548 346860 584576
rect 269816 584536 269822 584548
rect 346854 584536 346860 584548
rect 346912 584536 346918 584588
rect 79778 584468 79784 584520
rect 79836 584508 79842 584520
rect 350718 584508 350724 584520
rect 79836 584480 350724 584508
rect 79836 584468 79842 584480
rect 350718 584468 350724 584480
rect 350776 584468 350782 584520
rect 40954 584400 40960 584452
rect 41012 584440 41018 584452
rect 349246 584440 349252 584452
rect 41012 584412 349252 584440
rect 41012 584400 41018 584412
rect 349246 584400 349252 584412
rect 349304 584400 349310 584452
rect 377490 583720 377496 583772
rect 377548 583760 377554 583772
rect 407298 583760 407304 583772
rect 377548 583732 407304 583760
rect 377548 583720 377554 583732
rect 407298 583720 407304 583732
rect 407356 583720 407362 583772
rect 552934 583720 552940 583772
rect 552992 583760 552998 583772
rect 560386 583760 560392 583772
rect 552992 583732 560392 583760
rect 552992 583720 552998 583732
rect 560386 583720 560392 583732
rect 560444 583720 560450 583772
rect 43898 583040 43904 583092
rect 43956 583080 43962 583092
rect 87138 583080 87144 583092
rect 43956 583052 87144 583080
rect 43956 583040 43962 583052
rect 87138 583040 87144 583052
rect 87196 583040 87202 583092
rect 159082 583040 159088 583092
rect 159140 583080 159146 583092
rect 270218 583080 270224 583092
rect 159140 583052 270224 583080
rect 159140 583040 159146 583052
rect 270218 583040 270224 583052
rect 270276 583040 270282 583092
rect 84378 582972 84384 583024
rect 84436 583012 84442 583024
rect 349614 583012 349620 583024
rect 84436 582984 349620 583012
rect 84436 582972 84442 582984
rect 349614 582972 349620 582984
rect 349672 582972 349678 583024
rect 243538 581884 243544 581936
rect 243596 581924 243602 581936
rect 349246 581924 349252 581936
rect 243596 581896 349252 581924
rect 243596 581884 243602 581896
rect 349246 581884 349252 581896
rect 349304 581884 349310 581936
rect 147214 581816 147220 581868
rect 147272 581856 147278 581868
rect 274634 581856 274640 581868
rect 147272 581828 274640 581856
rect 147272 581816 147278 581828
rect 274634 581816 274640 581828
rect 274692 581816 274698 581868
rect 87322 581748 87328 581800
rect 87380 581788 87386 581800
rect 248414 581788 248420 581800
rect 87380 581760 248420 581788
rect 87380 581748 87386 581760
rect 248414 581748 248420 581760
rect 248472 581748 248478 581800
rect 46750 581680 46756 581732
rect 46808 581720 46814 581732
rect 253934 581720 253940 581732
rect 46808 581692 253940 581720
rect 46808 581680 46814 581692
rect 253934 581680 253940 581692
rect 253992 581680 253998 581732
rect 109034 581612 109040 581664
rect 109092 581652 109098 581664
rect 330110 581652 330116 581664
rect 109092 581624 330116 581652
rect 109092 581612 109098 581624
rect 330110 581612 330116 581624
rect 330168 581612 330174 581664
rect 209130 580456 209136 580508
rect 209188 580496 209194 580508
rect 250438 580496 250444 580508
rect 209188 580468 250444 580496
rect 209188 580456 209194 580468
rect 250438 580456 250444 580468
rect 250496 580456 250502 580508
rect 160094 580388 160100 580440
rect 160152 580428 160158 580440
rect 258166 580428 258172 580440
rect 160152 580400 258172 580428
rect 160152 580388 160158 580400
rect 258166 580388 258172 580400
rect 258224 580388 258230 580440
rect 297910 580388 297916 580440
rect 297968 580428 297974 580440
rect 367830 580428 367836 580440
rect 297968 580400 367836 580428
rect 297968 580388 297974 580400
rect 367830 580388 367836 580400
rect 367888 580388 367894 580440
rect 46198 580320 46204 580372
rect 46256 580360 46262 580372
rect 209774 580360 209780 580372
rect 46256 580332 209780 580360
rect 46256 580320 46262 580332
rect 209774 580320 209780 580332
rect 209832 580320 209838 580372
rect 245746 580320 245752 580372
rect 245804 580360 245810 580372
rect 347130 580360 347136 580372
rect 245804 580332 347136 580360
rect 245804 580320 245810 580332
rect 347130 580320 347136 580332
rect 347188 580320 347194 580372
rect 99466 580252 99472 580304
rect 99524 580292 99530 580304
rect 355134 580292 355140 580304
rect 99524 580264 355140 580292
rect 99524 580252 99530 580264
rect 355134 580252 355140 580264
rect 355192 580252 355198 580304
rect 383378 579640 383384 579692
rect 383436 579680 383442 579692
rect 407298 579680 407304 579692
rect 383436 579652 407304 579680
rect 383436 579640 383442 579652
rect 407298 579640 407304 579652
rect 407356 579640 407362 579692
rect 171686 579096 171692 579148
rect 171744 579136 171750 579148
rect 238846 579136 238852 579148
rect 171744 579108 238852 579136
rect 171744 579096 171750 579108
rect 238846 579096 238852 579108
rect 238904 579096 238910 579148
rect 208026 579028 208032 579080
rect 208084 579068 208090 579080
rect 347958 579068 347964 579080
rect 208084 579040 347964 579068
rect 208084 579028 208090 579040
rect 347958 579028 347964 579040
rect 348016 579028 348022 579080
rect 46474 578960 46480 579012
rect 46532 579000 46538 579012
rect 302234 579000 302240 579012
rect 46532 578972 302240 579000
rect 46532 578960 46538 578972
rect 302234 578960 302240 578972
rect 302292 578960 302298 579012
rect 35434 578892 35440 578944
rect 35492 578932 35498 578944
rect 306282 578932 306288 578944
rect 35492 578904 306288 578932
rect 35492 578892 35498 578904
rect 306282 578892 306288 578904
rect 306340 578892 306346 578944
rect 111794 577600 111800 577652
rect 111852 577640 111858 577652
rect 219986 577640 219992 577652
rect 111852 577612 219992 577640
rect 111852 577600 111858 577612
rect 219986 577600 219992 577612
rect 220044 577600 220050 577652
rect 231670 577600 231676 577652
rect 231728 577640 231734 577652
rect 355042 577640 355048 577652
rect 231728 577612 355048 577640
rect 231728 577600 231734 577612
rect 355042 577600 355048 577612
rect 355100 577600 355106 577652
rect 107654 577532 107660 577584
rect 107712 577572 107718 577584
rect 234614 577572 234620 577584
rect 107712 577544 234620 577572
rect 107712 577532 107718 577544
rect 234614 577532 234620 577544
rect 234672 577532 234678 577584
rect 246942 577532 246948 577584
rect 247000 577572 247006 577584
rect 281810 577572 281816 577584
rect 247000 577544 281816 577572
rect 247000 577532 247006 577544
rect 281810 577532 281816 577544
rect 281868 577532 281874 577584
rect 41230 577464 41236 577516
rect 41288 577504 41294 577516
rect 53834 577504 53840 577516
rect 41288 577476 53840 577504
rect 41288 577464 41294 577476
rect 53834 577464 53840 577476
rect 53892 577464 53898 577516
rect 74442 577464 74448 577516
rect 74500 577504 74506 577516
rect 351086 577504 351092 577516
rect 74500 577476 351092 577504
rect 74500 577464 74506 577476
rect 351086 577464 351092 577476
rect 351144 577464 351150 577516
rect 553302 577192 553308 577244
rect 553360 577232 553366 577244
rect 557626 577232 557632 577244
rect 553360 577204 557632 577232
rect 553360 577192 553366 577204
rect 557626 577192 557632 577204
rect 557684 577192 557690 577244
rect 388438 576852 388444 576904
rect 388496 576892 388502 576904
rect 407298 576892 407304 576904
rect 388496 576864 407304 576892
rect 388496 576852 388502 576864
rect 407298 576852 407304 576864
rect 407356 576852 407362 576904
rect 150526 576240 150532 576292
rect 150584 576280 150590 576292
rect 172606 576280 172612 576292
rect 150584 576252 172612 576280
rect 150584 576240 150590 576252
rect 172606 576240 172612 576252
rect 172664 576240 172670 576292
rect 244182 576240 244188 576292
rect 244240 576280 244246 576292
rect 350810 576280 350816 576292
rect 244240 576252 350816 576280
rect 244240 576240 244246 576252
rect 350810 576240 350816 576252
rect 350868 576240 350874 576292
rect 49142 576172 49148 576224
rect 49200 576212 49206 576224
rect 224954 576212 224960 576224
rect 49200 576184 224960 576212
rect 49200 576172 49206 576184
rect 224954 576172 224960 576184
rect 225012 576172 225018 576224
rect 238662 576172 238668 576224
rect 238720 576212 238726 576224
rect 348234 576212 348240 576224
rect 238720 576184 348240 576212
rect 238720 576172 238726 576184
rect 348234 576172 348240 576184
rect 348292 576172 348298 576224
rect 43806 576104 43812 576156
rect 43864 576144 43870 576156
rect 63586 576144 63592 576156
rect 43864 576116 63592 576144
rect 43864 576104 43870 576116
rect 63586 576104 63592 576116
rect 63644 576104 63650 576156
rect 89622 576104 89628 576156
rect 89680 576144 89686 576156
rect 350350 576144 350356 576156
rect 89680 576116 350356 576144
rect 89680 576104 89686 576116
rect 350350 576104 350356 576116
rect 350408 576104 350414 576156
rect 550174 575968 550180 576020
rect 550232 576008 550238 576020
rect 550450 576008 550456 576020
rect 550232 575980 550456 576008
rect 550232 575968 550238 575980
rect 550450 575968 550456 575980
rect 550508 575968 550514 576020
rect 403894 575492 403900 575544
rect 403952 575532 403958 575544
rect 407298 575532 407304 575544
rect 403952 575504 407304 575532
rect 403952 575492 403958 575504
rect 407298 575492 407304 575504
rect 407356 575492 407362 575544
rect 553302 575492 553308 575544
rect 553360 575532 553366 575544
rect 560662 575532 560668 575544
rect 553360 575504 560668 575532
rect 553360 575492 553366 575504
rect 560662 575492 560668 575504
rect 560720 575492 560726 575544
rect 117314 574948 117320 575000
rect 117372 574988 117378 575000
rect 237374 574988 237380 575000
rect 117372 574960 237380 574988
rect 117372 574948 117378 574960
rect 237374 574948 237380 574960
rect 237432 574948 237438 575000
rect 45278 574880 45284 574932
rect 45336 574920 45342 574932
rect 136634 574920 136640 574932
rect 45336 574892 136640 574920
rect 45336 574880 45342 574892
rect 136634 574880 136640 574892
rect 136692 574880 136698 574932
rect 209038 574880 209044 574932
rect 209096 574920 209102 574932
rect 349890 574920 349896 574932
rect 209096 574892 349896 574920
rect 209096 574880 209102 574892
rect 349890 574880 349896 574892
rect 349948 574880 349954 574932
rect 62022 574812 62028 574864
rect 62080 574852 62086 574864
rect 350902 574852 350908 574864
rect 62080 574824 350908 574852
rect 62080 574812 62086 574824
rect 350902 574812 350908 574824
rect 350960 574812 350966 574864
rect 3602 574744 3608 574796
rect 3660 574784 3666 574796
rect 365070 574784 365076 574796
rect 3660 574756 365076 574784
rect 3660 574744 3666 574756
rect 365070 574744 365076 574756
rect 365128 574744 365134 574796
rect 403986 573996 403992 574048
rect 404044 574036 404050 574048
rect 407298 574036 407304 574048
rect 404044 574008 407304 574036
rect 404044 573996 404050 574008
rect 407298 573996 407304 574008
rect 407356 573996 407362 574048
rect 552106 573996 552112 574048
rect 552164 574036 552170 574048
rect 554038 574036 554044 574048
rect 552164 574008 554044 574036
rect 552164 573996 552170 574008
rect 554038 573996 554044 574008
rect 554096 573996 554102 574048
rect 163406 573656 163412 573708
rect 163464 573696 163470 573708
rect 235994 573696 236000 573708
rect 163464 573668 236000 573696
rect 163464 573656 163470 573668
rect 235994 573656 236000 573668
rect 236052 573656 236058 573708
rect 85482 573588 85488 573640
rect 85540 573628 85546 573640
rect 147950 573628 147956 573640
rect 85540 573600 147956 573628
rect 85540 573588 85546 573600
rect 147950 573588 147956 573600
rect 148008 573588 148014 573640
rect 160002 573588 160008 573640
rect 160060 573628 160066 573640
rect 349338 573628 349344 573640
rect 160060 573600 349344 573628
rect 160060 573588 160066 573600
rect 349338 573588 349344 573600
rect 349396 573588 349402 573640
rect 46658 573520 46664 573572
rect 46716 573560 46722 573572
rect 264974 573560 264980 573572
rect 46716 573532 264980 573560
rect 46716 573520 46722 573532
rect 264974 573520 264980 573532
rect 265032 573520 265038 573572
rect 97902 573452 97908 573504
rect 97960 573492 97966 573504
rect 331490 573492 331496 573504
rect 97960 573464 331496 573492
rect 97960 573452 97966 573464
rect 331490 573452 331496 573464
rect 331548 573452 331554 573504
rect 35526 573384 35532 573436
rect 35584 573424 35590 573436
rect 349154 573424 349160 573436
rect 35584 573396 349160 573424
rect 35584 573384 35590 573396
rect 349154 573384 349160 573396
rect 349212 573384 349218 573436
rect 52638 573316 52644 573368
rect 52696 573356 52702 573368
rect 404998 573356 405004 573368
rect 52696 573328 405004 573356
rect 52696 573316 52702 573328
rect 404998 573316 405004 573328
rect 405056 573316 405062 573368
rect 403986 572704 403992 572756
rect 404044 572744 404050 572756
rect 407298 572744 407304 572756
rect 404044 572716 407304 572744
rect 404044 572704 404050 572716
rect 407298 572704 407304 572716
rect 407356 572704 407362 572756
rect 551370 572704 551376 572756
rect 551428 572744 551434 572756
rect 552014 572744 552020 572756
rect 551428 572716 552020 572744
rect 551428 572704 551434 572716
rect 552014 572704 552020 572716
rect 552072 572704 552078 572756
rect 209682 572160 209688 572212
rect 209740 572200 209746 572212
rect 278682 572200 278688 572212
rect 209740 572172 278688 572200
rect 209740 572160 209746 572172
rect 278682 572160 278688 572172
rect 278740 572160 278746 572212
rect 45094 572092 45100 572144
rect 45152 572132 45158 572144
rect 91094 572132 91100 572144
rect 45152 572104 91100 572132
rect 45152 572092 45158 572104
rect 91094 572092 91100 572104
rect 91152 572092 91158 572144
rect 155218 572092 155224 572144
rect 155276 572132 155282 572144
rect 255314 572132 255320 572144
rect 155276 572104 255320 572132
rect 155276 572092 155282 572104
rect 255314 572092 255320 572104
rect 255372 572092 255378 572144
rect 86862 572024 86868 572076
rect 86920 572064 86926 572076
rect 237374 572064 237380 572076
rect 86920 572036 237380 572064
rect 86920 572024 86926 572036
rect 237374 572024 237380 572036
rect 237432 572024 237438 572076
rect 268930 572024 268936 572076
rect 268988 572064 268994 572076
rect 354950 572064 354956 572076
rect 268988 572036 354956 572064
rect 268988 572024 268994 572036
rect 354950 572024 354956 572036
rect 355008 572024 355014 572076
rect 45738 571956 45744 572008
rect 45796 571996 45802 572008
rect 300854 571996 300860 572008
rect 45796 571968 300860 571996
rect 45796 571956 45802 571968
rect 300854 571956 300860 571968
rect 300912 571956 300918 572008
rect 366450 571344 366456 571396
rect 366508 571384 366514 571396
rect 407298 571384 407304 571396
rect 366508 571356 407304 571384
rect 366508 571344 366514 571356
rect 407298 571344 407304 571356
rect 407356 571344 407362 571396
rect 207934 570868 207940 570920
rect 207992 570908 207998 570920
rect 350994 570908 351000 570920
rect 207992 570880 351000 570908
rect 207992 570868 207998 570880
rect 350994 570868 351000 570880
rect 351052 570868 351058 570920
rect 208118 570800 208124 570852
rect 208176 570840 208182 570852
rect 356146 570840 356152 570852
rect 208176 570812 356152 570840
rect 208176 570800 208182 570812
rect 356146 570800 356152 570812
rect 356204 570800 356210 570852
rect 208302 570732 208308 570784
rect 208360 570772 208366 570784
rect 363138 570772 363144 570784
rect 208360 570744 363144 570772
rect 208360 570732 208366 570744
rect 363138 570732 363144 570744
rect 363196 570732 363202 570784
rect 47762 570664 47768 570716
rect 47820 570704 47826 570716
rect 258074 570704 258080 570716
rect 47820 570676 258080 570704
rect 47820 570664 47826 570676
rect 258074 570664 258080 570676
rect 258132 570664 258138 570716
rect 263502 570664 263508 570716
rect 263560 570704 263566 570716
rect 353294 570704 353300 570716
rect 263560 570676 353300 570704
rect 263560 570664 263566 570676
rect 353294 570664 353300 570676
rect 353352 570664 353358 570716
rect 67542 570596 67548 570648
rect 67600 570636 67606 570648
rect 353846 570636 353852 570648
rect 67600 570608 353852 570636
rect 67600 570596 67606 570608
rect 353846 570596 353852 570608
rect 353904 570596 353910 570648
rect 266262 569508 266268 569560
rect 266320 569548 266326 569560
rect 347774 569548 347780 569560
rect 266320 569520 347780 569548
rect 266320 569508 266326 569520
rect 347774 569508 347780 569520
rect 347832 569508 347838 569560
rect 252462 569440 252468 569492
rect 252520 569480 252526 569492
rect 353754 569480 353760 569492
rect 252520 569452 353760 569480
rect 252520 569440 252526 569452
rect 353754 569440 353760 569452
rect 353812 569440 353818 569492
rect 234522 569372 234528 569424
rect 234580 569412 234586 569424
rect 352374 569412 352380 569424
rect 234580 569384 352380 569412
rect 234580 569372 234586 569384
rect 352374 569372 352380 569384
rect 352432 569372 352438 569424
rect 231762 569304 231768 569356
rect 231820 569344 231826 569356
rect 354858 569344 354864 569356
rect 231820 569316 354864 569344
rect 231820 569304 231826 569316
rect 354858 569304 354864 569316
rect 354916 569304 354922 569356
rect 122742 569236 122748 569288
rect 122800 569276 122806 569288
rect 352466 569276 352472 569288
rect 122800 569248 352472 569276
rect 122800 569236 122806 569248
rect 352466 569236 352472 569248
rect 352524 569236 352530 569288
rect 117222 569168 117228 569220
rect 117280 569208 117286 569220
rect 353386 569208 353392 569220
rect 117280 569180 353392 569208
rect 117280 569168 117286 569180
rect 353386 569168 353392 569180
rect 353444 569168 353450 569220
rect 272886 568896 272892 568948
rect 272944 568936 272950 568948
rect 370498 568936 370504 568948
rect 272944 568908 370504 568936
rect 272944 568896 272950 568908
rect 370498 568896 370504 568908
rect 370556 568896 370562 568948
rect 234890 568828 234896 568880
rect 234948 568868 234954 568880
rect 357618 568868 357624 568880
rect 234948 568840 357624 568868
rect 234948 568828 234954 568840
rect 357618 568828 357624 568840
rect 357676 568828 357682 568880
rect 244550 568760 244556 568812
rect 244608 568800 244614 568812
rect 373994 568800 374000 568812
rect 244608 568772 374000 568800
rect 244608 568760 244614 568772
rect 373994 568760 374000 568772
rect 374052 568760 374058 568812
rect 222010 568692 222016 568744
rect 222068 568732 222074 568744
rect 361666 568732 361672 568744
rect 222068 568704 361672 568732
rect 222068 568692 222074 568704
rect 361666 568692 361672 568704
rect 361724 568692 361730 568744
rect 217502 568624 217508 568676
rect 217560 568664 217566 568676
rect 357434 568664 357440 568676
rect 217560 568636 357440 568664
rect 217560 568624 217566 568636
rect 357434 568624 357440 568636
rect 357492 568624 357498 568676
rect 35066 568556 35072 568608
rect 35124 568596 35130 568608
rect 407298 568596 407304 568608
rect 35124 568568 407304 568596
rect 35124 568556 35130 568568
rect 407298 568556 407304 568568
rect 407356 568556 407362 568608
rect 552566 568556 552572 568608
rect 552624 568596 552630 568608
rect 574186 568596 574192 568608
rect 552624 568568 574192 568596
rect 552624 568556 552630 568568
rect 574186 568556 574192 568568
rect 574244 568556 574250 568608
rect 296622 568148 296628 568200
rect 296680 568188 296686 568200
rect 348142 568188 348148 568200
rect 296680 568160 348148 568188
rect 296680 568148 296686 568160
rect 348142 568148 348148 568160
rect 348200 568148 348206 568200
rect 269022 568080 269028 568132
rect 269080 568120 269086 568132
rect 351178 568120 351184 568132
rect 269080 568092 351184 568120
rect 269080 568080 269086 568092
rect 351178 568080 351184 568092
rect 351236 568080 351242 568132
rect 249702 568012 249708 568064
rect 249760 568052 249766 568064
rect 351914 568052 351920 568064
rect 249760 568024 351920 568052
rect 249760 568012 249766 568024
rect 351914 568012 351920 568024
rect 351972 568012 351978 568064
rect 267642 567944 267648 567996
rect 267700 567984 267706 567996
rect 369946 567984 369952 567996
rect 267700 567956 369952 567984
rect 267700 567944 267706 567956
rect 369946 567944 369952 567956
rect 370004 567944 370010 567996
rect 233142 567876 233148 567928
rect 233200 567916 233206 567928
rect 352190 567916 352196 567928
rect 233200 567888 352196 567916
rect 233200 567876 233206 567888
rect 352190 567876 352196 567888
rect 352248 567876 352254 567928
rect 43530 567808 43536 567860
rect 43588 567848 43594 567860
rect 128354 567848 128360 567860
rect 43588 567820 128360 567848
rect 43588 567808 43594 567820
rect 128354 567808 128360 567820
rect 128412 567808 128418 567860
rect 208210 567808 208216 567860
rect 208268 567848 208274 567860
rect 360378 567848 360384 567860
rect 208268 567820 360384 567848
rect 208268 567808 208274 567820
rect 360378 567808 360384 567820
rect 360436 567808 360442 567860
rect 254854 567536 254860 567588
rect 254912 567576 254918 567588
rect 365162 567576 365168 567588
rect 254912 567548 365168 567576
rect 254912 567536 254918 567548
rect 365162 567536 365168 567548
rect 365220 567536 365226 567588
rect 243262 567468 243268 567520
rect 243320 567508 243326 567520
rect 385954 567508 385960 567520
rect 243320 567480 385960 567508
rect 243320 567468 243326 567480
rect 385954 567468 385960 567480
rect 386012 567468 386018 567520
rect 140222 567400 140228 567452
rect 140280 567440 140286 567452
rect 359550 567440 359556 567452
rect 140280 567412 359556 567440
rect 140280 567400 140286 567412
rect 359550 567400 359556 567412
rect 359608 567400 359614 567452
rect 131206 567332 131212 567384
rect 131264 567372 131270 567384
rect 353938 567372 353944 567384
rect 131264 567344 353944 567372
rect 131264 567332 131270 567344
rect 353938 567332 353944 567344
rect 353996 567332 354002 567384
rect 375098 567332 375104 567384
rect 375156 567372 375162 567384
rect 407298 567372 407304 567384
rect 375156 567344 407304 567372
rect 375156 567332 375162 567344
rect 407298 567332 407304 567344
rect 407356 567332 407362 567384
rect 143442 567264 143448 567316
rect 143500 567304 143506 567316
rect 384482 567304 384488 567316
rect 143500 567276 384488 567304
rect 143500 567264 143506 567276
rect 384482 567264 384488 567276
rect 384540 567264 384546 567316
rect 553302 567264 553308 567316
rect 553360 567304 553366 567316
rect 560570 567304 560576 567316
rect 553360 567276 560576 567304
rect 553360 567264 553366 567276
rect 560570 567264 560576 567276
rect 560628 567264 560634 567316
rect 116394 567196 116400 567248
rect 116452 567236 116458 567248
rect 401042 567236 401048 567248
rect 116452 567208 401048 567236
rect 116452 567196 116458 567208
rect 401042 567196 401048 567208
rect 401100 567196 401106 567248
rect 552474 567196 552480 567248
rect 552532 567236 552538 567248
rect 563330 567236 563336 567248
rect 552532 567208 563336 567236
rect 552532 567196 552538 567208
rect 563330 567196 563336 567208
rect 563388 567196 563394 567248
rect 293862 566720 293868 566772
rect 293920 566760 293926 566772
rect 350258 566760 350264 566772
rect 293920 566732 350264 566760
rect 293920 566720 293926 566732
rect 350258 566720 350264 566732
rect 350316 566720 350322 566772
rect 45922 566652 45928 566704
rect 45980 566692 45986 566704
rect 174538 566692 174544 566704
rect 45980 566664 174544 566692
rect 45980 566652 45986 566664
rect 174538 566652 174544 566664
rect 174596 566652 174602 566704
rect 262030 566652 262036 566704
rect 262088 566692 262094 566704
rect 348050 566692 348056 566704
rect 262088 566664 348056 566692
rect 262088 566652 262094 566664
rect 348050 566652 348056 566664
rect 348108 566652 348114 566704
rect 82078 566584 82084 566636
rect 82136 566624 82142 566636
rect 226886 566624 226892 566636
rect 82136 566596 226892 566624
rect 82136 566584 82142 566596
rect 226886 566584 226892 566596
rect 226944 566584 226950 566636
rect 257982 566584 257988 566636
rect 258040 566624 258046 566636
rect 349522 566624 349528 566636
rect 258040 566596 349528 566624
rect 258040 566584 258046 566596
rect 349522 566584 349528 566596
rect 349580 566584 349586 566636
rect 47026 566516 47032 566568
rect 47084 566556 47090 566568
rect 118694 566556 118700 566568
rect 47084 566528 118700 566556
rect 47084 566516 47090 566528
rect 118694 566516 118700 566528
rect 118752 566516 118758 566568
rect 128262 566516 128268 566568
rect 128320 566556 128326 566568
rect 359182 566556 359188 566568
rect 128320 566528 359188 566556
rect 128320 566516 128326 566528
rect 359182 566516 359188 566528
rect 359240 566516 359246 566568
rect 104802 566448 104808 566500
rect 104860 566488 104866 566500
rect 349430 566488 349436 566500
rect 104860 566460 349436 566488
rect 104860 566448 104866 566460
rect 349430 566448 349436 566460
rect 349488 566448 349494 566500
rect 317782 566380 317788 566432
rect 317840 566420 317846 566432
rect 367186 566420 367192 566432
rect 317840 566392 367192 566420
rect 317840 566380 317846 566392
rect 367186 566380 367192 566392
rect 367244 566380 367250 566432
rect 314930 566312 314936 566364
rect 314988 566352 314994 566364
rect 373258 566352 373264 566364
rect 314988 566324 373264 566352
rect 314988 566312 314994 566324
rect 373258 566312 373264 566324
rect 373316 566312 373322 566364
rect 275002 566244 275008 566296
rect 275060 566284 275066 566296
rect 392670 566284 392676 566296
rect 275060 566256 392676 566284
rect 275060 566244 275066 566256
rect 392670 566244 392676 566256
rect 392728 566244 392734 566296
rect 240962 566176 240968 566228
rect 241020 566216 241026 566228
rect 358814 566216 358820 566228
rect 241020 566188 358820 566216
rect 241020 566176 241026 566188
rect 358814 566176 358820 566188
rect 358872 566176 358878 566228
rect 198458 566108 198464 566160
rect 198516 566148 198522 566160
rect 357158 566148 357164 566160
rect 198516 566120 357164 566148
rect 198516 566108 198522 566120
rect 357158 566108 357164 566120
rect 357216 566108 357222 566160
rect 20622 566040 20628 566092
rect 20680 566080 20686 566092
rect 121546 566080 121552 566092
rect 20680 566052 121552 566080
rect 20680 566040 20686 566052
rect 121546 566040 121552 566052
rect 121604 566040 121610 566092
rect 217042 566040 217048 566092
rect 217100 566080 217106 566092
rect 381722 566080 381728 566092
rect 217100 566052 381728 566080
rect 217100 566040 217106 566052
rect 381722 566040 381728 566052
rect 381780 566040 381786 566092
rect 36814 565972 36820 566024
rect 36872 566012 36878 566024
rect 376478 566012 376484 566024
rect 36872 565984 376484 566012
rect 36872 565972 36878 565984
rect 376478 565972 376484 565984
rect 376536 565972 376542 566024
rect 32582 565904 32588 565956
rect 32640 565944 32646 565956
rect 405090 565944 405096 565956
rect 32640 565916 405096 565944
rect 32640 565904 32646 565916
rect 405090 565904 405096 565916
rect 405148 565904 405154 565956
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 17218 565876 17224 565888
rect 3292 565848 17224 565876
rect 3292 565836 3298 565848
rect 17218 565836 17224 565848
rect 17276 565836 17282 565888
rect 31294 565836 31300 565888
rect 31352 565876 31358 565888
rect 404998 565876 405004 565888
rect 31352 565848 405004 565876
rect 31352 565836 31358 565848
rect 404998 565836 405004 565848
rect 405056 565836 405062 565888
rect 25958 565564 25964 565616
rect 26016 565604 26022 565616
rect 311158 565604 311164 565616
rect 26016 565576 311164 565604
rect 26016 565564 26022 565576
rect 311158 565564 311164 565576
rect 311216 565564 311222 565616
rect 130746 565496 130752 565548
rect 130804 565536 130810 565548
rect 353570 565536 353576 565548
rect 130804 565508 353576 565536
rect 130804 565496 130810 565508
rect 353570 565496 353576 565508
rect 353628 565496 353634 565548
rect 203518 565428 203524 565480
rect 203576 565468 203582 565480
rect 243446 565468 243452 565480
rect 203576 565440 243452 565468
rect 203576 565428 203582 565440
rect 243446 565428 243452 565440
rect 243504 565428 243510 565480
rect 32950 565360 32956 565412
rect 33008 565400 33014 565412
rect 93854 565400 93860 565412
rect 33008 565372 93860 565400
rect 33008 565360 33014 565372
rect 93854 565360 93860 565372
rect 93912 565360 93918 565412
rect 135898 565360 135904 565412
rect 135956 565400 135962 565412
rect 252554 565400 252560 565412
rect 135956 565372 252560 565400
rect 135956 565360 135962 565372
rect 252554 565360 252560 565372
rect 252612 565360 252618 565412
rect 45186 565292 45192 565344
rect 45244 565332 45250 565344
rect 175366 565332 175372 565344
rect 45244 565304 175372 565332
rect 45244 565292 45250 565304
rect 175366 565292 175372 565304
rect 175424 565292 175430 565344
rect 180058 565292 180064 565344
rect 180116 565332 180122 565344
rect 225414 565332 225420 565344
rect 180116 565304 225420 565332
rect 180116 565292 180122 565304
rect 225414 565292 225420 565304
rect 225472 565292 225478 565344
rect 230382 565292 230388 565344
rect 230440 565332 230446 565344
rect 310514 565332 310520 565344
rect 230440 565304 310520 565332
rect 230440 565292 230446 565304
rect 310514 565292 310520 565304
rect 310572 565292 310578 565344
rect 44634 565224 44640 565276
rect 44692 565264 44698 565276
rect 78766 565264 78772 565276
rect 44692 565236 78772 565264
rect 44692 565224 44698 565236
rect 78766 565224 78772 565236
rect 78824 565224 78830 565276
rect 91002 565224 91008 565276
rect 91060 565264 91066 565276
rect 253934 565264 253940 565276
rect 91060 565236 253940 565264
rect 91060 565224 91066 565236
rect 253934 565224 253940 565236
rect 253992 565224 253998 565276
rect 333790 565224 333796 565276
rect 333848 565264 333854 565276
rect 347866 565264 347872 565276
rect 333848 565236 347872 565264
rect 333848 565224 333854 565236
rect 347866 565224 347872 565236
rect 347924 565224 347930 565276
rect 64782 565156 64788 565208
rect 64840 565196 64846 565208
rect 249794 565196 249800 565208
rect 64840 565168 249800 565196
rect 64840 565156 64846 565168
rect 249794 565156 249800 565168
rect 249852 565156 249858 565208
rect 324682 565156 324688 565208
rect 324740 565196 324746 565208
rect 354674 565196 354680 565208
rect 324740 565168 354680 565196
rect 324740 565156 324746 565168
rect 354674 565156 354680 565168
rect 354732 565156 354738 565208
rect 77110 565088 77116 565140
rect 77168 565128 77174 565140
rect 295702 565128 295708 565140
rect 77168 565100 295708 565128
rect 77168 565088 77174 565100
rect 295702 565088 295708 565100
rect 295760 565088 295766 565140
rect 315942 565088 315948 565140
rect 316000 565128 316006 565140
rect 374730 565128 374736 565140
rect 316000 565100 374736 565128
rect 316000 565088 316006 565100
rect 374730 565088 374736 565100
rect 374788 565088 374794 565140
rect 265986 565020 265992 565072
rect 266044 565060 266050 565072
rect 358906 565060 358912 565072
rect 266044 565032 358912 565060
rect 266044 565020 266050 565032
rect 358906 565020 358912 565032
rect 358964 565020 358970 565072
rect 23382 564952 23388 565004
rect 23440 564992 23446 565004
rect 82814 564992 82820 565004
rect 23440 564964 82820 564992
rect 23440 564952 23446 564964
rect 82814 564952 82820 564964
rect 82872 564952 82878 565004
rect 263410 564952 263416 565004
rect 263468 564992 263474 565004
rect 360194 564992 360200 565004
rect 263468 564964 360200 564992
rect 263468 564952 263474 564964
rect 360194 564952 360200 564964
rect 360252 564952 360258 565004
rect 42426 564884 42432 564936
rect 42484 564924 42490 564936
rect 104342 564924 104348 564936
rect 42484 564896 104348 564924
rect 42484 564884 42490 564896
rect 104342 564884 104348 564896
rect 104400 564884 104406 564936
rect 238662 564884 238668 564936
rect 238720 564924 238726 564936
rect 360286 564924 360292 564936
rect 238720 564896 360292 564924
rect 238720 564884 238726 564896
rect 360286 564884 360292 564896
rect 360344 564884 360350 564936
rect 36906 564816 36912 564868
rect 36964 564856 36970 564868
rect 111886 564856 111892 564868
rect 36964 564828 111892 564856
rect 36964 564816 36970 564828
rect 111886 564816 111892 564828
rect 111944 564816 111950 564868
rect 251818 564816 251824 564868
rect 251876 564856 251882 564868
rect 379146 564856 379152 564868
rect 251876 564828 379152 564856
rect 251876 564816 251882 564828
rect 379146 564816 379152 564828
rect 379204 564816 379210 564868
rect 39298 564748 39304 564800
rect 39356 564788 39362 564800
rect 168558 564788 168564 564800
rect 39356 564760 168564 564788
rect 39356 564748 39362 564760
rect 168558 564748 168564 564760
rect 168616 564748 168622 564800
rect 269850 564748 269856 564800
rect 269908 564788 269914 564800
rect 399570 564788 399576 564800
rect 269908 564760 399576 564788
rect 269908 564748 269914 564760
rect 399570 564748 399576 564760
rect 399628 564748 399634 564800
rect 38102 564680 38108 564732
rect 38160 564720 38166 564732
rect 191374 564720 191380 564732
rect 38160 564692 191380 564720
rect 38160 564680 38166 564692
rect 191374 564680 191380 564692
rect 191432 564680 191438 564732
rect 232498 564680 232504 564732
rect 232556 564720 232562 564732
rect 368658 564720 368664 564732
rect 232556 564692 368664 564720
rect 232556 564680 232562 564692
rect 368658 564680 368664 564692
rect 368716 564680 368722 564732
rect 33962 564612 33968 564664
rect 34020 564652 34026 564664
rect 244734 564652 244740 564664
rect 34020 564624 244740 564652
rect 34020 564612 34026 564624
rect 244734 564612 244740 564624
rect 244792 564612 244798 564664
rect 248322 564612 248328 564664
rect 248380 564652 248386 564664
rect 396810 564652 396816 564664
rect 248380 564624 396816 564652
rect 248380 564612 248386 564624
rect 396810 564612 396816 564624
rect 396868 564612 396874 564664
rect 40586 564544 40592 564596
rect 40644 564584 40650 564596
rect 124950 564584 124956 564596
rect 40644 564556 124956 564584
rect 40644 564544 40650 564556
rect 124950 564544 124956 564556
rect 125008 564544 125014 564596
rect 340138 564544 340144 564596
rect 340196 564584 340202 564596
rect 383102 564584 383108 564596
rect 340196 564556 383108 564584
rect 340196 564544 340202 564556
rect 383102 564544 383108 564556
rect 383160 564544 383166 564596
rect 298922 564476 298928 564528
rect 298980 564516 298986 564528
rect 402422 564516 402428 564528
rect 298980 564488 402428 564516
rect 298980 564476 298986 564488
rect 402422 564476 402428 564488
rect 402480 564476 402486 564528
rect 41046 564408 41052 564460
rect 41104 564448 41110 564460
rect 382182 564448 382188 564460
rect 41104 564420 382188 564448
rect 41104 564408 41110 564420
rect 382182 564408 382188 564420
rect 382240 564408 382246 564460
rect 405550 564408 405556 564460
rect 405608 564448 405614 564460
rect 407390 564448 407396 564460
rect 405608 564420 407396 564448
rect 405608 564408 405614 564420
rect 407390 564408 407396 564420
rect 407448 564408 407454 564460
rect 31386 564068 31392 564120
rect 31444 564108 31450 564120
rect 339126 564108 339132 564120
rect 31444 564080 339132 564108
rect 31444 564068 31450 564080
rect 339126 564068 339132 564080
rect 339184 564068 339190 564120
rect 23198 564000 23204 564052
rect 23256 564040 23262 564052
rect 255774 564040 255780 564052
rect 23256 564012 255780 564040
rect 23256 564000 23262 564012
rect 255774 564000 255780 564012
rect 255832 564000 255838 564052
rect 24302 563932 24308 563984
rect 24360 563972 24366 563984
rect 56594 563972 56600 563984
rect 24360 563944 56600 563972
rect 24360 563932 24366 563944
rect 56594 563932 56600 563944
rect 56652 563932 56658 563984
rect 327810 563932 327816 563984
rect 327868 563972 327874 563984
rect 352834 563972 352840 563984
rect 327868 563944 352840 563972
rect 327868 563932 327874 563944
rect 352834 563932 352840 563944
rect 352892 563932 352898 563984
rect 41874 563864 41880 563916
rect 41932 563904 41938 563916
rect 74626 563904 74632 563916
rect 41932 563876 74632 563904
rect 41932 563864 41938 563876
rect 74626 563864 74632 563876
rect 74684 563864 74690 563916
rect 204162 563864 204168 563916
rect 204220 563904 204226 563916
rect 247034 563904 247040 563916
rect 204220 563876 247040 563904
rect 204220 563864 204226 563876
rect 247034 563864 247040 563876
rect 247092 563864 247098 563916
rect 264882 563864 264888 563916
rect 264940 563904 264946 563916
rect 343726 563904 343732 563916
rect 264940 563876 343732 563904
rect 264940 563864 264946 563876
rect 343726 563864 343732 563876
rect 343784 563864 343790 563916
rect 44818 563796 44824 563848
rect 44876 563836 44882 563848
rect 88334 563836 88340 563848
rect 44876 563808 88340 563836
rect 44876 563796 44882 563808
rect 88334 563796 88340 563808
rect 88392 563796 88398 563848
rect 153930 563796 153936 563848
rect 153988 563836 153994 563848
rect 175458 563836 175464 563848
rect 153988 563808 175464 563836
rect 153988 563796 153994 563808
rect 175458 563796 175464 563808
rect 175516 563796 175522 563848
rect 179690 563796 179696 563848
rect 179748 563836 179754 563848
rect 262214 563836 262220 563848
rect 179748 563808 262220 563836
rect 179748 563796 179754 563808
rect 262214 563796 262220 563808
rect 262272 563796 262278 563848
rect 299382 563796 299388 563848
rect 299440 563836 299446 563848
rect 389910 563836 389916 563848
rect 299440 563808 389916 563836
rect 299440 563796 299446 563808
rect 389910 563796 389916 563808
rect 389968 563796 389974 563848
rect 40678 563728 40684 563780
rect 40736 563768 40742 563780
rect 87046 563768 87052 563780
rect 40736 563740 87052 563768
rect 40736 563728 40742 563740
rect 87046 563728 87052 563740
rect 87104 563728 87110 563780
rect 95142 563728 95148 563780
rect 95200 563768 95206 563780
rect 222194 563768 222200 563780
rect 95200 563740 222200 563768
rect 95200 563728 95206 563740
rect 222194 563728 222200 563740
rect 222252 563728 222258 563780
rect 224770 563728 224776 563780
rect 224828 563768 224834 563780
rect 355318 563768 355324 563780
rect 224828 563740 355324 563768
rect 224828 563728 224834 563740
rect 355318 563728 355324 563740
rect 355376 563728 355382 563780
rect 46382 563660 46388 563712
rect 46440 563700 46446 563712
rect 175274 563700 175280 563712
rect 46440 563672 175280 563700
rect 46440 563660 46446 563672
rect 175274 563660 175280 563672
rect 175332 563660 175338 563712
rect 208026 563660 208032 563712
rect 208084 563700 208090 563712
rect 353662 563700 353668 563712
rect 208084 563672 353668 563700
rect 208084 563660 208090 563672
rect 353662 563660 353668 563672
rect 353720 563660 353726 563712
rect 224218 563592 224224 563644
rect 224276 563632 224282 563644
rect 398282 563632 398288 563644
rect 224276 563604 398288 563632
rect 224276 563592 224282 563604
rect 398282 563592 398288 563604
rect 398340 563592 398346 563644
rect 43438 563524 43444 563576
rect 43496 563564 43502 563576
rect 162302 563564 162308 563576
rect 43496 563536 162308 563564
rect 43496 563524 43502 563536
rect 162302 563524 162308 563536
rect 162360 563524 162366 563576
rect 180702 563524 180708 563576
rect 180760 563564 180766 563576
rect 378778 563564 378784 563576
rect 180760 563536 378784 563564
rect 180760 563524 180766 563536
rect 378778 563524 378784 563536
rect 378836 563524 378842 563576
rect 179138 563456 179144 563508
rect 179196 563496 179202 563508
rect 385770 563496 385776 563508
rect 179196 563468 385776 563496
rect 179196 563456 179202 563468
rect 385770 563456 385776 563468
rect 385828 563456 385834 563508
rect 39206 563388 39212 563440
rect 39264 563428 39270 563440
rect 181070 563428 181076 563440
rect 39264 563400 181076 563428
rect 39264 563388 39270 563400
rect 181070 563388 181076 563400
rect 181128 563388 181134 563440
rect 249702 563388 249708 563440
rect 249760 563428 249766 563440
rect 389174 563428 389180 563440
rect 249760 563400 389180 563428
rect 249760 563388 249766 563400
rect 389174 563388 389180 563400
rect 389232 563388 389238 563440
rect 22002 563320 22008 563372
rect 22060 563360 22066 563372
rect 301406 563360 301412 563372
rect 22060 563332 301412 563360
rect 22060 563320 22066 563332
rect 301406 563320 301412 563332
rect 301464 563320 301470 563372
rect 307662 563320 307668 563372
rect 307720 563360 307726 563372
rect 402330 563360 402336 563372
rect 307720 563332 402336 563360
rect 307720 563320 307726 563332
rect 402330 563320 402336 563332
rect 402388 563320 402394 563372
rect 24762 563252 24768 563304
rect 24820 563292 24826 563304
rect 325970 563292 325976 563304
rect 24820 563264 325976 563292
rect 24820 563252 24826 563264
rect 325970 563252 325976 563264
rect 326028 563252 326034 563304
rect 338758 563252 338764 563304
rect 338816 563292 338822 563304
rect 365714 563292 365720 563304
rect 338816 563264 365720 563292
rect 338816 563252 338822 563264
rect 365714 563252 365720 563264
rect 365772 563252 365778 563304
rect 336642 563184 336648 563236
rect 336700 563224 336706 563236
rect 364426 563224 364432 563236
rect 336700 563196 364432 563224
rect 336700 563184 336706 563196
rect 364426 563184 364432 563196
rect 364484 563184 364490 563236
rect 38470 563116 38476 563168
rect 38528 563156 38534 563168
rect 401134 563156 401140 563168
rect 38528 563128 401140 563156
rect 38528 563116 38534 563128
rect 401134 563116 401140 563128
rect 401192 563116 401198 563168
rect 31110 563048 31116 563100
rect 31168 563088 31174 563100
rect 395522 563088 395528 563100
rect 31168 563060 395528 563088
rect 31168 563048 31174 563060
rect 395522 563048 395528 563060
rect 395580 563048 395586 563100
rect 48222 562980 48228 563032
rect 48280 563020 48286 563032
rect 49142 563020 49148 563032
rect 48280 562992 49148 563020
rect 48280 562980 48286 562992
rect 49142 562980 49148 562992
rect 49200 562980 49206 563032
rect 23014 562708 23020 562760
rect 23072 562748 23078 562760
rect 113450 562748 113456 562760
rect 23072 562720 113456 562748
rect 23072 562708 23078 562720
rect 113450 562708 113456 562720
rect 113508 562708 113514 562760
rect 203610 562708 203616 562760
rect 203668 562748 203674 562760
rect 340782 562748 340788 562760
rect 203668 562720 340788 562748
rect 203668 562708 203674 562720
rect 340782 562708 340788 562720
rect 340840 562708 340846 562760
rect 43346 562640 43352 562692
rect 43404 562680 43410 562692
rect 405182 562680 405188 562692
rect 43404 562652 405188 562680
rect 43404 562640 43410 562652
rect 405182 562640 405188 562652
rect 405240 562640 405246 562692
rect 23106 562572 23112 562624
rect 23164 562612 23170 562624
rect 65702 562612 65708 562624
rect 23164 562584 65708 562612
rect 23164 562572 23170 562584
rect 65702 562572 65708 562584
rect 65760 562572 65766 562624
rect 73062 562572 73068 562624
rect 73120 562612 73126 562624
rect 91278 562612 91284 562624
rect 73120 562584 91284 562612
rect 73120 562572 73126 562584
rect 91278 562572 91284 562584
rect 91336 562572 91342 562624
rect 338022 562572 338028 562624
rect 338080 562612 338086 562624
rect 347038 562612 347044 562624
rect 338080 562584 347044 562612
rect 338080 562572 338086 562584
rect 347038 562572 347044 562584
rect 347096 562572 347102 562624
rect 75822 562504 75828 562556
rect 75880 562544 75886 562556
rect 124858 562544 124864 562556
rect 75880 562516 124864 562544
rect 75880 562504 75886 562516
rect 124858 562504 124864 562516
rect 124916 562504 124922 562556
rect 214466 562504 214472 562556
rect 214524 562544 214530 562556
rect 249702 562544 249708 562556
rect 214524 562516 249708 562544
rect 214524 562504 214530 562516
rect 249702 562504 249708 562516
rect 249760 562504 249766 562556
rect 304074 562504 304080 562556
rect 304132 562544 304138 562556
rect 369118 562544 369124 562556
rect 304132 562516 369124 562544
rect 304132 562504 304138 562516
rect 369118 562504 369124 562516
rect 369176 562504 369182 562556
rect 39758 562436 39764 562488
rect 39816 562476 39822 562488
rect 81618 562476 81624 562488
rect 39816 562448 81624 562476
rect 39816 562436 39822 562448
rect 81618 562436 81624 562448
rect 81676 562436 81682 562488
rect 82814 562436 82820 562488
rect 82872 562476 82878 562488
rect 148134 562476 148140 562488
rect 82872 562448 148140 562476
rect 82872 562436 82878 562448
rect 148134 562436 148140 562448
rect 148192 562436 148198 562488
rect 208762 562436 208768 562488
rect 208820 562476 208826 562488
rect 338758 562476 338764 562488
rect 208820 562448 338764 562476
rect 208820 562436 208826 562448
rect 338758 562436 338764 562448
rect 338816 562436 338822 562488
rect 36998 562368 37004 562420
rect 37056 562408 37062 562420
rect 83734 562408 83740 562420
rect 37056 562380 83740 562408
rect 37056 562368 37062 562380
rect 83734 562368 83740 562380
rect 83792 562368 83798 562420
rect 90818 562368 90824 562420
rect 90876 562408 90882 562420
rect 173158 562408 173164 562420
rect 90876 562380 173164 562408
rect 90876 562368 90882 562380
rect 173158 562368 173164 562380
rect 173216 562368 173222 562420
rect 186866 562368 186872 562420
rect 186924 562408 186930 562420
rect 335354 562408 335360 562420
rect 186924 562380 335360 562408
rect 186924 562368 186930 562380
rect 335354 562368 335360 562380
rect 335412 562368 335418 562420
rect 339126 562368 339132 562420
rect 339184 562408 339190 562420
rect 381998 562408 382004 562420
rect 339184 562380 382004 562408
rect 339184 562368 339190 562380
rect 381998 562368 382004 562380
rect 382056 562368 382062 562420
rect 552014 562368 552020 562420
rect 552072 562408 552078 562420
rect 556614 562408 556620 562420
rect 552072 562380 556620 562408
rect 552072 562368 552078 562380
rect 556614 562368 556620 562380
rect 556672 562368 556678 562420
rect 47394 562300 47400 562352
rect 47452 562340 47458 562352
rect 74534 562340 74540 562352
rect 47452 562312 74540 562340
rect 47452 562300 47458 562312
rect 74534 562300 74540 562312
rect 74592 562300 74598 562352
rect 76650 562300 76656 562352
rect 76708 562340 76714 562352
rect 173250 562340 173256 562352
rect 76708 562312 173256 562340
rect 76708 562300 76714 562312
rect 173250 562300 173256 562312
rect 173308 562300 173314 562352
rect 226794 562300 226800 562352
rect 226852 562340 226858 562352
rect 406562 562340 406568 562352
rect 226852 562312 406568 562340
rect 226852 562300 226858 562312
rect 406562 562300 406568 562312
rect 406620 562300 406626 562352
rect 35526 562232 35532 562284
rect 35584 562272 35590 562284
rect 94774 562272 94780 562284
rect 35584 562244 94780 562272
rect 35584 562232 35590 562244
rect 94774 562232 94780 562244
rect 94832 562232 94838 562284
rect 278314 562232 278320 562284
rect 278372 562272 278378 562284
rect 346486 562272 346492 562284
rect 278372 562244 346492 562272
rect 278372 562232 278378 562244
rect 346486 562232 346492 562244
rect 346544 562232 346550 562284
rect 40494 562164 40500 562216
rect 40552 562204 40558 562216
rect 99374 562204 99380 562216
rect 40552 562176 99380 562204
rect 40552 562164 40558 562176
rect 99374 562164 99380 562176
rect 99432 562164 99438 562216
rect 236362 562164 236368 562216
rect 236420 562204 236426 562216
rect 336366 562204 336372 562216
rect 236420 562176 336372 562204
rect 236420 562164 236426 562176
rect 336366 562164 336372 562176
rect 336424 562164 336430 562216
rect 347682 562164 347688 562216
rect 347740 562204 347746 562216
rect 378870 562204 378876 562216
rect 347740 562176 378876 562204
rect 347740 562164 347746 562176
rect 378870 562164 378876 562176
rect 378928 562164 378934 562216
rect 38378 562096 38384 562148
rect 38436 562136 38442 562148
rect 105078 562136 105084 562148
rect 38436 562108 105084 562136
rect 38436 562096 38442 562108
rect 105078 562096 105084 562108
rect 105136 562096 105142 562148
rect 260282 562096 260288 562148
rect 260340 562136 260346 562148
rect 367922 562136 367928 562148
rect 260340 562108 367928 562136
rect 260340 562096 260346 562108
rect 367922 562096 367928 562108
rect 367980 562096 367986 562148
rect 27430 562028 27436 562080
rect 27488 562068 27494 562080
rect 51534 562068 51540 562080
rect 27488 562040 51540 562068
rect 27488 562028 27494 562040
rect 51534 562028 51540 562040
rect 51592 562028 51598 562080
rect 51626 562028 51632 562080
rect 51684 562068 51690 562080
rect 138014 562068 138020 562080
rect 51684 562040 138020 562068
rect 51684 562028 51690 562040
rect 138014 562028 138020 562040
rect 138072 562028 138078 562080
rect 250438 562028 250444 562080
rect 250496 562068 250502 562080
rect 372062 562068 372068 562080
rect 250496 562040 372068 562068
rect 250496 562028 250502 562040
rect 372062 562028 372068 562040
rect 372120 562028 372126 562080
rect 32858 561960 32864 562012
rect 32916 562000 32922 562012
rect 138566 562000 138572 562012
rect 32916 561972 138572 562000
rect 32916 561960 32922 561972
rect 138566 561960 138572 561972
rect 138624 561960 138630 562012
rect 336274 561960 336280 562012
rect 336332 562000 336338 562012
rect 381814 562000 381820 562012
rect 336332 561972 381820 562000
rect 336332 561960 336338 561972
rect 381814 561960 381820 561972
rect 381872 561960 381878 562012
rect 42334 561892 42340 561944
rect 42392 561932 42398 561944
rect 193858 561932 193864 561944
rect 42392 561904 193864 561932
rect 42392 561892 42398 561904
rect 193858 561892 193864 561904
rect 193916 561892 193922 561944
rect 201402 561892 201408 561944
rect 201460 561932 201466 561944
rect 366542 561932 366548 561944
rect 201460 561904 366548 561932
rect 201460 561892 201466 561904
rect 366542 561892 366548 561904
rect 366600 561892 366606 561944
rect 51074 561824 51080 561876
rect 51132 561864 51138 561876
rect 181622 561864 181628 561876
rect 51132 561836 181628 561864
rect 51132 561824 51138 561836
rect 181622 561824 181628 561836
rect 181680 561824 181686 561876
rect 184842 561824 184848 561876
rect 184900 561864 184906 561876
rect 368566 561864 368572 561876
rect 184900 561836 368572 561864
rect 184900 561824 184906 561836
rect 368566 561824 368572 561836
rect 368624 561824 368630 561876
rect 110138 561756 110144 561808
rect 110196 561796 110202 561808
rect 391474 561796 391480 561808
rect 110196 561768 391480 561796
rect 110196 561756 110202 561768
rect 391474 561756 391480 561768
rect 391532 561756 391538 561808
rect 19150 561688 19156 561740
rect 19208 561728 19214 561740
rect 50246 561728 50252 561740
rect 19208 561700 50252 561728
rect 19208 561688 19214 561700
rect 50246 561688 50252 561700
rect 50304 561688 50310 561740
rect 337562 561688 337568 561740
rect 337620 561728 337626 561740
rect 346394 561728 346400 561740
rect 337620 561700 346400 561728
rect 337620 561688 337626 561700
rect 346394 561688 346400 561700
rect 346452 561688 346458 561740
rect 32674 561620 32680 561672
rect 32732 561660 32738 561672
rect 407298 561660 407304 561672
rect 32732 561632 407304 561660
rect 32732 561620 32738 561632
rect 407298 561620 407304 561632
rect 407356 561620 407362 561672
rect 47118 561552 47124 561604
rect 47176 561592 47182 561604
rect 67634 561592 67640 561604
rect 47176 561564 67640 561592
rect 47176 561552 47182 561564
rect 67634 561552 67640 561564
rect 67692 561552 67698 561604
rect 25682 561484 25688 561536
rect 25740 561524 25746 561536
rect 52454 561524 52460 561536
rect 25740 561496 52460 561524
rect 25740 561484 25746 561496
rect 52454 561484 52460 561496
rect 52512 561484 52518 561536
rect 35434 561416 35440 561468
rect 35492 561456 35498 561468
rect 63678 561456 63684 561468
rect 35492 561428 63684 561456
rect 35492 561416 35498 561428
rect 63678 561416 63684 561428
rect 63736 561416 63742 561468
rect 47302 561348 47308 561400
rect 47360 561388 47366 561400
rect 77294 561388 77300 561400
rect 47360 561360 77300 561388
rect 47360 561348 47366 561360
rect 77294 561348 77300 561360
rect 77352 561348 77358 561400
rect 38194 561280 38200 561332
rect 38252 561320 38258 561332
rect 69014 561320 69020 561332
rect 38252 561292 69020 561320
rect 38252 561280 38258 561292
rect 69014 561280 69020 561292
rect 69072 561280 69078 561332
rect 27154 561212 27160 561264
rect 27212 561252 27218 561264
rect 59354 561252 59360 561264
rect 27212 561224 59360 561252
rect 27212 561212 27218 561224
rect 59354 561212 59360 561224
rect 59412 561212 59418 561264
rect 37090 561144 37096 561196
rect 37148 561184 37154 561196
rect 70394 561184 70400 561196
rect 37148 561156 70400 561184
rect 37148 561144 37154 561156
rect 70394 561144 70400 561156
rect 70452 561144 70458 561196
rect 30006 561076 30012 561128
rect 30064 561116 30070 561128
rect 63494 561116 63500 561128
rect 30064 561088 63500 561116
rect 30064 561076 30070 561088
rect 63494 561076 63500 561088
rect 63552 561076 63558 561128
rect 313090 561076 313096 561128
rect 313148 561116 313154 561128
rect 352558 561116 352564 561128
rect 313148 561088 352564 561116
rect 313148 561076 313154 561088
rect 352558 561076 352564 561088
rect 352616 561076 352622 561128
rect 38286 561008 38292 561060
rect 38344 561048 38350 561060
rect 82998 561048 83004 561060
rect 38344 561020 83004 561048
rect 38344 561008 38350 561020
rect 82998 561008 83004 561020
rect 83056 561008 83062 561060
rect 305914 561008 305920 561060
rect 305972 561048 305978 561060
rect 364978 561048 364984 561060
rect 305972 561020 364984 561048
rect 305972 561008 305978 561020
rect 364978 561008 364984 561020
rect 365036 561008 365042 561060
rect 39482 560940 39488 560992
rect 39540 560980 39546 560992
rect 86954 560980 86960 560992
rect 39540 560952 86960 560980
rect 39540 560940 39546 560952
rect 86954 560940 86960 560952
rect 87012 560940 87018 560992
rect 291194 560940 291200 560992
rect 291252 560980 291258 560992
rect 352282 560980 352288 560992
rect 291252 560952 352288 560980
rect 291252 560940 291258 560952
rect 352282 560940 352288 560952
rect 352340 560940 352346 560992
rect 47486 560872 47492 560924
rect 47544 560912 47550 560924
rect 62114 560912 62120 560924
rect 47544 560884 62120 560912
rect 47544 560872 47550 560884
rect 62114 560872 62120 560884
rect 62172 560872 62178 560924
rect 287882 560872 287888 560924
rect 287940 560912 287946 560924
rect 382274 560912 382280 560924
rect 287940 560884 382280 560912
rect 287940 560872 287946 560884
rect 382274 560872 382280 560884
rect 382332 560872 382338 560924
rect 255682 560804 255688 560856
rect 255740 560844 255746 560856
rect 358998 560844 359004 560856
rect 255740 560816 359004 560844
rect 255740 560804 255746 560816
rect 358998 560804 359004 560816
rect 359056 560804 359062 560856
rect 233786 560736 233792 560788
rect 233844 560776 233850 560788
rect 351270 560776 351276 560788
rect 233844 560748 351276 560776
rect 233844 560736 233850 560748
rect 351270 560736 351276 560748
rect 351328 560736 351334 560788
rect 235810 560668 235816 560720
rect 235868 560708 235874 560720
rect 399478 560708 399484 560720
rect 235868 560680 399484 560708
rect 235868 560668 235874 560680
rect 399478 560668 399484 560680
rect 399536 560668 399542 560720
rect 146202 560600 146208 560652
rect 146260 560640 146266 560652
rect 352650 560640 352656 560652
rect 146260 560612 352656 560640
rect 146260 560600 146266 560612
rect 352650 560600 352656 560612
rect 352708 560600 352714 560652
rect 183002 560532 183008 560584
rect 183060 560572 183066 560584
rect 403618 560572 403624 560584
rect 183060 560544 403624 560572
rect 183060 560532 183066 560544
rect 403618 560532 403624 560544
rect 403676 560532 403682 560584
rect 62482 560464 62488 560516
rect 62540 560504 62546 560516
rect 392762 560504 392768 560516
rect 62540 560476 392768 560504
rect 62540 560464 62546 560476
rect 392762 560464 392768 560476
rect 392820 560464 392826 560516
rect 43622 560396 43628 560448
rect 43680 560436 43686 560448
rect 405274 560436 405280 560448
rect 43680 560408 405280 560436
rect 43680 560396 43686 560408
rect 405274 560396 405280 560408
rect 405332 560396 405338 560448
rect 44082 560328 44088 560380
rect 44140 560368 44146 560380
rect 407758 560368 407764 560380
rect 44140 560340 407764 560368
rect 44140 560328 44146 560340
rect 407758 560328 407764 560340
rect 407816 560328 407822 560380
rect 552934 560328 552940 560380
rect 552992 560368 552998 560380
rect 569218 560368 569224 560380
rect 552992 560340 569224 560368
rect 552992 560328 552998 560340
rect 569218 560328 569224 560340
rect 569276 560328 569282 560380
rect 325602 560260 325608 560312
rect 325660 560300 325666 560312
rect 357526 560300 357532 560312
rect 325660 560272 357532 560300
rect 325660 560260 325666 560272
rect 357526 560260 357532 560272
rect 357584 560260 357590 560312
rect 553302 560260 553308 560312
rect 553360 560300 553366 560312
rect 582742 560300 582748 560312
rect 553360 560272 582748 560300
rect 553360 560260 553366 560272
rect 582742 560260 582748 560272
rect 582800 560260 582806 560312
rect 46842 560192 46848 560244
rect 46900 560232 46906 560244
rect 49050 560232 49056 560244
rect 46900 560204 49056 560232
rect 46900 560192 46906 560204
rect 49050 560192 49056 560204
rect 49108 560192 49114 560244
rect 49602 560192 49608 560244
rect 49660 560232 49666 560244
rect 59170 560232 59176 560244
rect 49660 560204 59176 560232
rect 49660 560192 49666 560204
rect 59170 560192 59176 560204
rect 59228 560192 59234 560244
rect 46566 560124 46572 560176
rect 46624 560164 46630 560176
rect 48866 560164 48872 560176
rect 46624 560136 48872 560164
rect 46624 560124 46630 560136
rect 48866 560124 48872 560136
rect 48924 560124 48930 560176
rect 294782 560096 294788 560108
rect 289786 560068 294788 560096
rect 142126 560000 151814 560028
rect 142126 559620 142154 560000
rect 148870 559960 148876 559972
rect 133846 559592 142154 559620
rect 142264 559932 148876 559960
rect 36630 559512 36636 559564
rect 36688 559552 36694 559564
rect 133846 559552 133874 559592
rect 36688 559524 133874 559552
rect 36688 559512 36694 559524
rect 39666 558900 39672 558952
rect 39724 558940 39730 558952
rect 142264 558940 142292 559932
rect 148870 559920 148876 559932
rect 148928 559920 148934 559972
rect 151786 559620 151814 560000
rect 277026 559920 277032 559972
rect 277084 559920 277090 559972
rect 153166 559728 154574 559756
rect 153166 559620 153194 559728
rect 151786 559592 153194 559620
rect 154546 559552 154574 559728
rect 277044 559552 277072 559920
rect 289786 559620 289814 560068
rect 294782 560056 294788 560068
rect 294840 560056 294846 560108
rect 281506 559592 289814 559620
rect 294662 560000 299474 560028
rect 281506 559552 281534 559592
rect 154546 559524 269114 559552
rect 277044 559524 281534 559552
rect 269086 559348 269114 559524
rect 269086 559320 276014 559348
rect 275986 559212 276014 559320
rect 294662 559280 294690 560000
rect 294782 559920 294788 559972
rect 294840 559920 294846 559972
rect 285784 559252 294690 559280
rect 275986 559184 285674 559212
rect 285646 559144 285674 559184
rect 285784 559144 285812 559252
rect 294800 559212 294828 559920
rect 299446 559892 299474 560000
rect 335326 560000 340644 560028
rect 334986 559920 334992 559972
rect 335044 559960 335050 559972
rect 335326 559960 335354 560000
rect 335044 559932 335354 559960
rect 335044 559920 335050 559932
rect 339402 559920 339408 559972
rect 339460 559920 339466 559972
rect 299446 559864 300854 559892
rect 300826 559484 300854 559864
rect 303586 559592 304994 559620
rect 300826 559456 302234 559484
rect 302206 559416 302234 559456
rect 303586 559416 303614 559592
rect 304966 559552 304994 559592
rect 339420 559552 339448 559920
rect 304966 559524 306374 559552
rect 306346 559484 306374 559524
rect 307726 559524 309134 559552
rect 307726 559484 307754 559524
rect 306346 559456 307754 559484
rect 309106 559484 309134 559524
rect 310486 559524 339448 559552
rect 310486 559484 310514 559524
rect 309106 559456 310514 559484
rect 340616 559416 340644 560000
rect 346486 559988 346492 560040
rect 346544 560028 346550 560040
rect 348326 560028 348332 560040
rect 346544 560000 348332 560028
rect 346544 559988 346550 560000
rect 348326 559988 348332 560000
rect 348384 559988 348390 560040
rect 340690 559920 340696 559972
rect 340748 559920 340754 559972
rect 340782 559920 340788 559972
rect 340840 559920 340846 559972
rect 346394 559920 346400 559972
rect 346452 559960 346458 559972
rect 346452 559932 347728 559960
rect 346452 559920 346458 559932
rect 340708 559484 340736 559920
rect 340800 559688 340828 559920
rect 347700 559904 347728 559932
rect 347682 559852 347688 559904
rect 347740 559852 347746 559904
rect 360562 559688 360568 559700
rect 340800 559660 360568 559688
rect 360562 559648 360568 559660
rect 360620 559648 360626 559700
rect 347682 559580 347688 559632
rect 347740 559620 347746 559632
rect 407942 559620 407948 559632
rect 347740 559592 407948 559620
rect 347740 559580 347746 559592
rect 407942 559580 407948 559592
rect 408000 559580 408006 559632
rect 348326 559512 348332 559564
rect 348384 559552 348390 559564
rect 407574 559552 407580 559564
rect 348384 559524 407580 559552
rect 348384 559512 348390 559524
rect 407574 559512 407580 559524
rect 407632 559512 407638 559564
rect 347682 559484 347688 559496
rect 340708 559456 347688 559484
rect 347682 559444 347688 559456
rect 347740 559444 347746 559496
rect 302206 559388 303614 559416
rect 307726 559388 309134 559416
rect 340616 559388 347774 559416
rect 307726 559348 307754 559388
rect 302206 559320 303614 559348
rect 302206 559280 302234 559320
rect 300826 559252 302234 559280
rect 300826 559212 300854 559252
rect 294800 559184 300854 559212
rect 303586 559212 303614 559320
rect 306346 559320 307754 559348
rect 309106 559348 309134 559388
rect 309106 559320 310514 559348
rect 306346 559280 306374 559320
rect 304966 559252 306374 559280
rect 304966 559212 304994 559252
rect 303586 559184 304994 559212
rect 285646 559116 285812 559144
rect 39724 558912 142292 558940
rect 310486 558940 310514 559320
rect 347746 559076 347774 559388
rect 365806 559076 365812 559088
rect 347746 559048 365812 559076
rect 365806 559036 365812 559048
rect 365864 559036 365870 559088
rect 347682 558968 347688 559020
rect 347740 559008 347746 559020
rect 391290 559008 391296 559020
rect 347740 558980 391296 559008
rect 347740 558968 347746 558980
rect 391290 558968 391296 558980
rect 391348 558968 391354 559020
rect 352098 558940 352104 558952
rect 310486 558912 352104 558940
rect 39724 558900 39730 558912
rect 352098 558900 352104 558912
rect 352156 558900 352162 558952
rect 349430 558152 349436 558204
rect 349488 558192 349494 558204
rect 349798 558192 349804 558204
rect 349488 558164 349804 558192
rect 349488 558152 349494 558164
rect 349798 558152 349804 558164
rect 349856 558152 349862 558204
rect 552934 557608 552940 557660
rect 552992 557648 552998 557660
rect 561858 557648 561864 557660
rect 552992 557620 561864 557648
rect 552992 557608 552998 557620
rect 561858 557608 561864 557620
rect 561916 557608 561922 557660
rect 553302 557540 553308 557592
rect 553360 557580 553366 557592
rect 568666 557580 568672 557592
rect 553360 557552 568672 557580
rect 553360 557540 553366 557552
rect 568666 557540 568672 557552
rect 568724 557540 568730 557592
rect 552014 556520 552020 556572
rect 552072 556560 552078 556572
rect 554866 556560 554872 556572
rect 552072 556532 554872 556560
rect 552072 556520 552078 556532
rect 554866 556520 554872 556532
rect 554924 556520 554930 556572
rect 44542 556180 44548 556232
rect 44600 556220 44606 556232
rect 46290 556220 46296 556232
rect 44600 556192 46296 556220
rect 44600 556180 44606 556192
rect 46290 556180 46296 556192
rect 46348 556180 46354 556232
rect 349430 554684 349436 554736
rect 349488 554724 349494 554736
rect 351914 554724 351920 554736
rect 349488 554696 351920 554724
rect 349488 554684 349494 554696
rect 351914 554684 351920 554696
rect 351972 554684 351978 554736
rect 552014 553800 552020 553852
rect 552072 553840 552078 553852
rect 553946 553840 553952 553852
rect 552072 553812 553952 553840
rect 552072 553800 552078 553812
rect 553946 553800 553952 553812
rect 554004 553800 554010 553852
rect 398558 552032 398564 552084
rect 398616 552072 398622 552084
rect 407298 552072 407304 552084
rect 398616 552044 407304 552072
rect 398616 552032 398622 552044
rect 407298 552032 407304 552044
rect 407356 552032 407362 552084
rect 552382 552032 552388 552084
rect 552440 552072 552446 552084
rect 579706 552072 579712 552084
rect 552440 552044 579712 552072
rect 552440 552032 552446 552044
rect 579706 552032 579712 552044
rect 579764 552032 579770 552084
rect 405274 551964 405280 552016
rect 405332 552004 405338 552016
rect 407390 552004 407396 552016
rect 405332 551976 407396 552004
rect 405332 551964 405338 551976
rect 407390 551964 407396 551976
rect 407448 551964 407454 552016
rect 42702 551080 42708 551132
rect 42760 551120 42766 551132
rect 46290 551120 46296 551132
rect 42760 551092 46296 551120
rect 42760 551080 42766 551092
rect 46290 551080 46296 551092
rect 46348 551080 46354 551132
rect 41138 550808 41144 550860
rect 41196 550848 41202 550860
rect 46290 550848 46296 550860
rect 41196 550820 46296 550848
rect 41196 550808 41202 550820
rect 46290 550808 46296 550820
rect 46348 550808 46354 550860
rect 553302 550808 553308 550860
rect 553360 550848 553366 550860
rect 559466 550848 559472 550860
rect 553360 550820 559472 550848
rect 553360 550808 553366 550820
rect 559466 550808 559472 550820
rect 559524 550808 559530 550860
rect 350442 550604 350448 550656
rect 350500 550644 350506 550656
rect 388530 550644 388536 550656
rect 350500 550616 388536 550644
rect 350500 550604 350506 550616
rect 388530 550604 388536 550616
rect 388588 550604 388594 550656
rect 398650 550604 398656 550656
rect 398708 550644 398714 550656
rect 407298 550644 407304 550656
rect 398708 550616 407304 550644
rect 398708 550604 398714 550616
rect 407298 550604 407304 550616
rect 407356 550604 407362 550656
rect 42610 549244 42616 549296
rect 42668 549284 42674 549296
rect 46290 549284 46296 549296
rect 42668 549256 46296 549284
rect 42668 549244 42674 549256
rect 46290 549244 46296 549256
rect 46348 549244 46354 549296
rect 358262 549244 358268 549296
rect 358320 549284 358326 549296
rect 407298 549284 407304 549296
rect 358320 549256 407304 549284
rect 358320 549244 358326 549256
rect 407298 549244 407304 549256
rect 407356 549244 407362 549296
rect 553302 549244 553308 549296
rect 553360 549284 553366 549296
rect 575566 549284 575572 549296
rect 553360 549256 575572 549284
rect 553360 549244 553366 549256
rect 575566 549244 575572 549256
rect 575624 549244 575630 549296
rect 46106 549108 46112 549160
rect 46164 549148 46170 549160
rect 46290 549148 46296 549160
rect 46164 549120 46296 549148
rect 46164 549108 46170 549120
rect 46290 549108 46296 549120
rect 46348 549108 46354 549160
rect 350166 546524 350172 546576
rect 350224 546564 350230 546576
rect 366634 546564 366640 546576
rect 350224 546536 366640 546564
rect 350224 546524 350230 546536
rect 366634 546524 366640 546536
rect 366692 546524 366698 546576
rect 377582 546524 377588 546576
rect 377640 546564 377646 546576
rect 407298 546564 407304 546576
rect 377640 546536 407304 546564
rect 377640 546524 377646 546536
rect 407298 546524 407304 546536
rect 407356 546524 407362 546576
rect 30190 546456 30196 546508
rect 30248 546496 30254 546508
rect 46106 546496 46112 546508
rect 30248 546468 46112 546496
rect 30248 546456 30254 546468
rect 46106 546456 46112 546468
rect 46164 546456 46170 546508
rect 350442 546456 350448 546508
rect 350500 546496 350506 546508
rect 388622 546496 388628 546508
rect 350500 546468 388628 546496
rect 350500 546456 350506 546468
rect 388622 546456 388628 546468
rect 388680 546456 388686 546508
rect 553302 546456 553308 546508
rect 553360 546496 553366 546508
rect 560754 546496 560760 546508
rect 553360 546468 560760 546496
rect 553360 546456 553366 546468
rect 560754 546456 560760 546468
rect 560812 546456 560818 546508
rect 551462 545300 551468 545352
rect 551520 545340 551526 545352
rect 552014 545340 552020 545352
rect 551520 545312 552020 545340
rect 551520 545300 551526 545312
rect 552014 545300 552020 545312
rect 552072 545300 552078 545352
rect 34054 545096 34060 545148
rect 34112 545136 34118 545148
rect 46014 545136 46020 545148
rect 34112 545108 46020 545136
rect 34112 545096 34118 545108
rect 46014 545096 46020 545108
rect 46072 545096 46078 545148
rect 405366 543804 405372 543856
rect 405424 543844 405430 543856
rect 407390 543844 407396 543856
rect 405424 543816 407396 543844
rect 405424 543804 405430 543816
rect 407390 543804 407396 543816
rect 407448 543804 407454 543856
rect 43162 543736 43168 543788
rect 43220 543776 43226 543788
rect 46106 543776 46112 543788
rect 43220 543748 46112 543776
rect 43220 543736 43226 543748
rect 46106 543736 46112 543748
rect 46164 543736 46170 543788
rect 377674 543736 377680 543788
rect 377732 543776 377738 543788
rect 407298 543776 407304 543788
rect 377732 543748 407304 543776
rect 377732 543736 377738 543748
rect 407298 543736 407304 543748
rect 407356 543736 407362 543788
rect 553302 543736 553308 543788
rect 553360 543776 553366 543788
rect 561950 543776 561956 543788
rect 553360 543748 561956 543776
rect 553360 543736 553366 543748
rect 561950 543736 561956 543748
rect 562008 543736 562014 543788
rect 350442 542376 350448 542428
rect 350500 542416 350506 542428
rect 363782 542416 363788 542428
rect 350500 542388 363788 542416
rect 350500 542376 350506 542388
rect 363782 542376 363788 542388
rect 363840 542376 363846 542428
rect 353938 542308 353944 542360
rect 353996 542348 354002 542360
rect 407298 542348 407304 542360
rect 353996 542320 407304 542348
rect 353996 542308 354002 542320
rect 407298 542308 407304 542320
rect 407356 542308 407362 542360
rect 21910 540948 21916 541000
rect 21968 540988 21974 541000
rect 46106 540988 46112 541000
rect 21968 540960 46112 540988
rect 21968 540948 21974 540960
rect 46106 540948 46112 540960
rect 46164 540948 46170 541000
rect 552566 539588 552572 539640
rect 552624 539628 552630 539640
rect 567378 539628 567384 539640
rect 552624 539600 567384 539628
rect 552624 539588 552630 539600
rect 567378 539588 567384 539600
rect 567436 539588 567442 539640
rect 350442 538228 350448 538280
rect 350500 538268 350506 538280
rect 367830 538268 367836 538280
rect 350500 538240 367836 538268
rect 350500 538228 350506 538240
rect 367830 538228 367836 538240
rect 367888 538228 367894 538280
rect 552566 538228 552572 538280
rect 552624 538268 552630 538280
rect 559558 538268 559564 538280
rect 552624 538240 559564 538268
rect 552624 538228 552630 538240
rect 559558 538228 559564 538240
rect 559616 538228 559622 538280
rect 44082 538160 44088 538212
rect 44140 538200 44146 538212
rect 46106 538200 46112 538212
rect 44140 538172 46112 538200
rect 44140 538160 44146 538172
rect 46106 538160 46112 538172
rect 46164 538160 46170 538212
rect 350442 536800 350448 536852
rect 350500 536840 350506 536852
rect 372614 536840 372620 536852
rect 350500 536812 372620 536840
rect 350500 536800 350506 536812
rect 372614 536800 372620 536812
rect 372672 536800 372678 536852
rect 553302 535848 553308 535900
rect 553360 535888 553366 535900
rect 559374 535888 559380 535900
rect 553360 535860 559380 535888
rect 553360 535848 553366 535860
rect 559374 535848 559380 535860
rect 559432 535848 559438 535900
rect 552382 534148 552388 534200
rect 552440 534188 552446 534200
rect 570138 534188 570144 534200
rect 552440 534160 570144 534188
rect 552440 534148 552446 534160
rect 570138 534148 570144 534160
rect 570196 534148 570202 534200
rect 350442 534080 350448 534132
rect 350500 534120 350506 534132
rect 380250 534120 380256 534132
rect 350500 534092 380256 534120
rect 350500 534080 350506 534092
rect 380250 534080 380256 534092
rect 380308 534080 380314 534132
rect 394142 534080 394148 534132
rect 394200 534120 394206 534132
rect 407298 534120 407304 534132
rect 394200 534092 407304 534120
rect 394200 534080 394206 534092
rect 407298 534080 407304 534092
rect 407356 534080 407362 534132
rect 553302 534080 553308 534132
rect 553360 534120 553366 534132
rect 581546 534120 581552 534132
rect 553360 534092 581552 534120
rect 553360 534080 553366 534092
rect 581546 534080 581552 534092
rect 581604 534080 581610 534132
rect 550174 533332 550180 533384
rect 550232 533372 550238 533384
rect 550450 533372 550456 533384
rect 550232 533344 550456 533372
rect 550232 533332 550238 533344
rect 550450 533332 550456 533344
rect 550508 533332 550514 533384
rect 350166 532788 350172 532840
rect 350224 532828 350230 532840
rect 359090 532828 359096 532840
rect 350224 532800 359096 532828
rect 350224 532788 350230 532800
rect 359090 532788 359096 532800
rect 359148 532788 359154 532840
rect 350442 532720 350448 532772
rect 350500 532760 350506 532772
rect 381906 532760 381912 532772
rect 350500 532732 381912 532760
rect 350500 532720 350506 532732
rect 381906 532720 381912 532732
rect 381964 532720 381970 532772
rect 552014 532516 552020 532568
rect 552072 532556 552078 532568
rect 553762 532556 553768 532568
rect 552072 532528 553768 532556
rect 552072 532516 552078 532528
rect 553762 532516 553768 532528
rect 553820 532516 553826 532568
rect 43070 531768 43076 531820
rect 43128 531808 43134 531820
rect 46014 531808 46020 531820
rect 43128 531780 46020 531808
rect 43128 531768 43134 531780
rect 46014 531768 46020 531780
rect 46072 531768 46078 531820
rect 349430 531292 349436 531344
rect 349488 531332 349494 531344
rect 351362 531332 351368 531344
rect 349488 531304 351368 531332
rect 349488 531292 349494 531304
rect 351362 531292 351368 531304
rect 351420 531292 351426 531344
rect 552014 530884 552020 530936
rect 552072 530924 552078 530936
rect 553854 530924 553860 530936
rect 552072 530896 553860 530924
rect 552072 530884 552078 530896
rect 553854 530884 553860 530896
rect 553912 530884 553918 530936
rect 39022 529932 39028 529984
rect 39080 529972 39086 529984
rect 46106 529972 46112 529984
rect 39080 529944 46112 529972
rect 39080 529932 39086 529944
rect 46106 529932 46112 529944
rect 46164 529932 46170 529984
rect 350442 529932 350448 529984
rect 350500 529972 350506 529984
rect 380434 529972 380440 529984
rect 350500 529944 380440 529972
rect 350500 529932 350506 529944
rect 380434 529932 380440 529944
rect 380492 529932 380498 529984
rect 552658 529932 552664 529984
rect 552716 529972 552722 529984
rect 563422 529972 563428 529984
rect 552716 529944 563428 529972
rect 552716 529932 552722 529944
rect 563422 529932 563428 529944
rect 563480 529932 563486 529984
rect 42242 528572 42248 528624
rect 42300 528612 42306 528624
rect 45830 528612 45836 528624
rect 42300 528584 45836 528612
rect 42300 528572 42306 528584
rect 45830 528572 45836 528584
rect 45888 528572 45894 528624
rect 370590 528572 370596 528624
rect 370648 528612 370654 528624
rect 407298 528612 407304 528624
rect 370648 528584 407304 528612
rect 370648 528572 370654 528584
rect 407298 528572 407304 528584
rect 407356 528572 407362 528624
rect 350442 527144 350448 527196
rect 350500 527184 350506 527196
rect 376294 527184 376300 527196
rect 350500 527156 376300 527184
rect 350500 527144 350506 527156
rect 376294 527144 376300 527156
rect 376352 527144 376358 527196
rect 553302 527144 553308 527196
rect 553360 527184 553366 527196
rect 564802 527184 564808 527196
rect 553360 527156 564808 527184
rect 553360 527144 553366 527156
rect 564802 527144 564808 527156
rect 564860 527144 564866 527196
rect 552014 526056 552020 526108
rect 552072 526096 552078 526108
rect 553762 526096 553768 526108
rect 552072 526068 553768 526096
rect 552072 526056 552078 526068
rect 553762 526056 553768 526068
rect 553820 526056 553826 526108
rect 350442 525920 350448 525972
rect 350500 525960 350506 525972
rect 356698 525960 356704 525972
rect 350500 525932 356704 525960
rect 350500 525920 350506 525932
rect 356698 525920 356704 525932
rect 356756 525920 356762 525972
rect 44726 525716 44732 525768
rect 44784 525756 44790 525768
rect 46106 525756 46112 525768
rect 44784 525728 46112 525756
rect 44784 525716 44790 525728
rect 46106 525716 46112 525728
rect 46164 525716 46170 525768
rect 552014 525716 552020 525768
rect 552072 525756 552078 525768
rect 553670 525756 553676 525768
rect 552072 525728 553676 525756
rect 552072 525716 552078 525728
rect 553670 525716 553676 525728
rect 553728 525716 553734 525768
rect 571978 525716 571984 525768
rect 572036 525756 572042 525768
rect 579798 525756 579804 525768
rect 572036 525728 579804 525756
rect 572036 525716 572042 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 40770 525648 40776 525700
rect 40828 525688 40834 525700
rect 45646 525688 45652 525700
rect 40828 525660 45652 525688
rect 40828 525648 40834 525660
rect 45646 525648 45652 525660
rect 45704 525648 45710 525700
rect 402606 525036 402612 525088
rect 402664 525076 402670 525088
rect 407298 525076 407304 525088
rect 402664 525048 407304 525076
rect 402664 525036 402670 525048
rect 407298 525036 407304 525048
rect 407356 525036 407362 525088
rect 390370 524424 390376 524476
rect 390428 524464 390434 524476
rect 407390 524464 407396 524476
rect 390428 524436 407396 524464
rect 390428 524424 390434 524436
rect 407390 524424 407396 524436
rect 407448 524424 407454 524476
rect 387334 523064 387340 523116
rect 387392 523104 387398 523116
rect 407298 523104 407304 523116
rect 387392 523076 407304 523104
rect 387392 523064 387398 523076
rect 407298 523064 407304 523076
rect 407356 523064 407362 523116
rect 350442 522996 350448 523048
rect 350500 523036 350506 523048
rect 378962 523036 378968 523048
rect 350500 523008 378968 523036
rect 350500 522996 350506 523008
rect 378962 522996 378968 523008
rect 379020 522996 379026 523048
rect 399938 522928 399944 522980
rect 399996 522968 400002 522980
rect 407298 522968 407304 522980
rect 399996 522940 407304 522968
rect 399996 522928 400002 522940
rect 407298 522928 407304 522940
rect 407356 522928 407362 522980
rect 401226 521704 401232 521756
rect 401284 521744 401290 521756
rect 407390 521744 407396 521756
rect 401284 521716 407396 521744
rect 401284 521704 401290 521716
rect 407390 521704 407396 521716
rect 407448 521704 407454 521756
rect 350074 521160 350080 521212
rect 350132 521200 350138 521212
rect 352098 521200 352104 521212
rect 350132 521172 352104 521200
rect 350132 521160 350138 521172
rect 352098 521160 352104 521172
rect 352156 521160 352162 521212
rect 23290 520276 23296 520328
rect 23348 520316 23354 520328
rect 46198 520316 46204 520328
rect 23348 520288 46204 520316
rect 23348 520276 23354 520288
rect 46198 520276 46204 520288
rect 46256 520276 46262 520328
rect 373534 520276 373540 520328
rect 373592 520316 373598 520328
rect 407298 520316 407304 520328
rect 373592 520288 407304 520316
rect 373592 520276 373598 520288
rect 407298 520276 407304 520288
rect 407356 520276 407362 520328
rect 552014 520276 552020 520328
rect 552072 520316 552078 520328
rect 571518 520316 571524 520328
rect 552072 520288 571524 520316
rect 552072 520276 552078 520288
rect 571518 520276 571524 520288
rect 571576 520276 571582 520328
rect 552014 519256 552020 519308
rect 552072 519296 552078 519308
rect 553670 519296 553676 519308
rect 552072 519268 553676 519296
rect 552072 519256 552078 519268
rect 553670 519256 553676 519268
rect 553728 519256 553734 519308
rect 552014 518916 552020 518968
rect 552072 518956 552078 518968
rect 564618 518956 564624 518968
rect 552072 518928 564624 518956
rect 552072 518916 552078 518928
rect 564618 518916 564624 518928
rect 564676 518916 564682 518968
rect 398466 517556 398472 517608
rect 398524 517596 398530 517608
rect 407298 517596 407304 517608
rect 398524 517568 407304 517596
rect 398524 517556 398530 517568
rect 407298 517556 407304 517568
rect 407356 517556 407362 517608
rect 350442 517488 350448 517540
rect 350500 517528 350506 517540
rect 383194 517528 383200 517540
rect 350500 517500 383200 517528
rect 350500 517488 350506 517500
rect 383194 517488 383200 517500
rect 383252 517488 383258 517540
rect 388990 517488 388996 517540
rect 389048 517528 389054 517540
rect 407390 517528 407396 517540
rect 389048 517500 407396 517528
rect 389048 517488 389054 517500
rect 407390 517488 407396 517500
rect 407448 517488 407454 517540
rect 350442 516264 350448 516316
rect 350500 516304 350506 516316
rect 367094 516304 367100 516316
rect 350500 516276 367100 516304
rect 350500 516264 350506 516276
rect 367094 516264 367100 516276
rect 367152 516264 367158 516316
rect 350074 516196 350080 516248
rect 350132 516236 350138 516248
rect 384666 516236 384672 516248
rect 350132 516208 384672 516236
rect 350132 516196 350138 516208
rect 384666 516196 384672 516208
rect 384724 516196 384730 516248
rect 394510 516196 394516 516248
rect 394568 516236 394574 516248
rect 407298 516236 407304 516248
rect 394568 516208 407304 516236
rect 394568 516196 394574 516208
rect 407298 516196 407304 516208
rect 407356 516196 407362 516248
rect 40402 516128 40408 516180
rect 40460 516168 40466 516180
rect 46014 516168 46020 516180
rect 40460 516140 46020 516168
rect 40460 516128 40466 516140
rect 46014 516128 46020 516140
rect 46072 516128 46078 516180
rect 358170 516128 358176 516180
rect 358228 516168 358234 516180
rect 407390 516168 407396 516180
rect 358228 516140 407396 516168
rect 358228 516128 358234 516140
rect 407390 516128 407396 516140
rect 407448 516128 407454 516180
rect 552014 516128 552020 516180
rect 552072 516168 552078 516180
rect 570874 516168 570880 516180
rect 552072 516140 570880 516168
rect 552072 516128 552078 516140
rect 570874 516128 570880 516140
rect 570932 516128 570938 516180
rect 405182 516060 405188 516112
rect 405240 516100 405246 516112
rect 407666 516100 407672 516112
rect 405240 516072 407672 516100
rect 405240 516060 405246 516072
rect 407666 516060 407672 516072
rect 407724 516060 407730 516112
rect 552014 514768 552020 514820
rect 552072 514808 552078 514820
rect 567562 514808 567568 514820
rect 552072 514780 567568 514808
rect 552072 514768 552078 514780
rect 567562 514768 567568 514780
rect 567620 514768 567626 514820
rect 350074 513408 350080 513460
rect 350132 513448 350138 513460
rect 354122 513448 354128 513460
rect 350132 513420 354128 513448
rect 350132 513408 350138 513420
rect 354122 513408 354128 513420
rect 354180 513408 354186 513460
rect 42150 513340 42156 513392
rect 42208 513380 42214 513392
rect 45922 513380 45928 513392
rect 42208 513352 45928 513380
rect 42208 513340 42214 513352
rect 45922 513340 45928 513352
rect 45980 513340 45986 513392
rect 350442 513340 350448 513392
rect 350500 513380 350506 513392
rect 368014 513380 368020 513392
rect 350500 513352 368020 513380
rect 350500 513340 350506 513352
rect 368014 513340 368020 513352
rect 368072 513340 368078 513392
rect 374822 513272 374828 513324
rect 374880 513312 374886 513324
rect 407298 513312 407304 513324
rect 374880 513284 407304 513312
rect 374880 513272 374886 513284
rect 407298 513272 407304 513284
rect 407356 513272 407362 513324
rect 373442 511980 373448 512032
rect 373500 512020 373506 512032
rect 407298 512020 407304 512032
rect 373500 511992 407304 512020
rect 373500 511980 373506 511992
rect 407298 511980 407304 511992
rect 407356 511980 407362 512032
rect 350442 511912 350448 511964
rect 350500 511952 350506 511964
rect 353294 511952 353300 511964
rect 350500 511924 353300 511952
rect 350500 511912 350506 511924
rect 353294 511912 353300 511924
rect 353352 511912 353358 511964
rect 43990 510552 43996 510604
rect 44048 510592 44054 510604
rect 46106 510592 46112 510604
rect 44048 510564 46112 510592
rect 44048 510552 44054 510564
rect 46106 510552 46112 510564
rect 46164 510552 46170 510604
rect 553302 509872 553308 509924
rect 553360 509912 553366 509924
rect 559098 509912 559104 509924
rect 553360 509884 559104 509912
rect 553360 509872 553366 509884
rect 559098 509872 559104 509884
rect 559156 509872 559162 509924
rect 40494 509260 40500 509312
rect 40552 509300 40558 509312
rect 46014 509300 46020 509312
rect 40552 509272 46020 509300
rect 40552 509260 40558 509272
rect 46014 509260 46020 509272
rect 46072 509260 46078 509312
rect 385862 509260 385868 509312
rect 385920 509300 385926 509312
rect 407298 509300 407304 509312
rect 385920 509272 407304 509300
rect 385920 509260 385926 509272
rect 407298 509260 407304 509272
rect 407356 509260 407362 509312
rect 350442 509192 350448 509244
rect 350500 509232 350506 509244
rect 399846 509232 399852 509244
rect 350500 509204 399852 509232
rect 350500 509192 350506 509204
rect 399846 509192 399852 509204
rect 399904 509192 399910 509244
rect 359550 509124 359556 509176
rect 359608 509164 359614 509176
rect 407298 509164 407304 509176
rect 359608 509136 407304 509164
rect 359608 509124 359614 509136
rect 407298 509124 407304 509136
rect 407356 509124 407362 509176
rect 349982 506540 349988 506592
rect 350040 506580 350046 506592
rect 352098 506580 352104 506592
rect 350040 506552 352104 506580
rect 350040 506540 350046 506552
rect 352098 506540 352104 506552
rect 352156 506540 352162 506592
rect 27522 506472 27528 506524
rect 27580 506512 27586 506524
rect 46106 506512 46112 506524
rect 27580 506484 46112 506512
rect 27580 506472 27586 506484
rect 46106 506472 46112 506484
rect 46164 506472 46170 506524
rect 349890 506472 349896 506524
rect 349948 506512 349954 506524
rect 351270 506512 351276 506524
rect 349948 506484 351276 506512
rect 349948 506472 349954 506484
rect 351270 506472 351276 506484
rect 351328 506472 351334 506524
rect 359550 506472 359556 506524
rect 359608 506512 359614 506524
rect 407298 506512 407304 506524
rect 359608 506484 407304 506512
rect 359608 506472 359614 506484
rect 407298 506472 407304 506484
rect 407356 506472 407362 506524
rect 350442 506404 350448 506456
rect 350500 506444 350506 506456
rect 403802 506444 403808 506456
rect 350500 506416 403808 506444
rect 350500 506404 350506 506416
rect 403802 506404 403808 506416
rect 403860 506404 403866 506456
rect 553118 506404 553124 506456
rect 553176 506444 553182 506456
rect 570690 506444 570696 506456
rect 553176 506416 570696 506444
rect 553176 506404 553182 506416
rect 570690 506404 570696 506416
rect 570748 506404 570754 506456
rect 21818 505112 21824 505164
rect 21876 505152 21882 505164
rect 46106 505152 46112 505164
rect 21876 505124 46112 505152
rect 21876 505112 21882 505124
rect 46106 505112 46112 505124
rect 46164 505112 46170 505164
rect 350074 505112 350080 505164
rect 350132 505152 350138 505164
rect 380618 505152 380624 505164
rect 350132 505124 380624 505152
rect 350132 505112 350138 505124
rect 380618 505112 380624 505124
rect 380676 505112 380682 505164
rect 553302 505112 553308 505164
rect 553360 505152 553366 505164
rect 572990 505152 572996 505164
rect 553360 505124 572996 505152
rect 553360 505112 553366 505124
rect 572990 505112 572996 505124
rect 573048 505112 573054 505164
rect 350442 503684 350448 503736
rect 350500 503724 350506 503736
rect 360470 503724 360476 503736
rect 350500 503696 360476 503724
rect 350500 503684 350506 503696
rect 360470 503684 360476 503696
rect 360528 503684 360534 503736
rect 553302 503684 553308 503736
rect 553360 503724 553366 503736
rect 566274 503724 566280 503736
rect 553360 503696 566280 503724
rect 553360 503684 553366 503696
rect 566274 503684 566280 503696
rect 566332 503684 566338 503736
rect 553302 502392 553308 502444
rect 553360 502432 553366 502444
rect 559006 502432 559012 502444
rect 553360 502404 559012 502432
rect 553360 502392 553366 502404
rect 559006 502392 559012 502404
rect 559064 502392 559070 502444
rect 39390 501848 39396 501900
rect 39448 501888 39454 501900
rect 46106 501888 46112 501900
rect 39448 501860 46112 501888
rect 39448 501848 39454 501860
rect 46106 501848 46112 501860
rect 46164 501848 46170 501900
rect 553118 501032 553124 501084
rect 553176 501072 553182 501084
rect 566182 501072 566188 501084
rect 553176 501044 566188 501072
rect 553176 501032 553182 501044
rect 566182 501032 566188 501044
rect 566240 501032 566246 501084
rect 397270 500964 397276 501016
rect 397328 501004 397334 501016
rect 407298 501004 407304 501016
rect 397328 500976 407304 501004
rect 397328 500964 397334 500976
rect 407298 500964 407304 500976
rect 407356 500964 407362 501016
rect 553302 500964 553308 501016
rect 553360 501004 553366 501016
rect 572070 501004 572076 501016
rect 553360 500976 572076 501004
rect 553360 500964 553366 500976
rect 572070 500964 572076 500976
rect 572128 500964 572134 501016
rect 39850 500896 39856 500948
rect 39908 500936 39914 500948
rect 45646 500936 45652 500948
rect 39908 500908 45652 500936
rect 39908 500896 39914 500908
rect 45646 500896 45652 500908
rect 45704 500896 45710 500948
rect 402146 500896 402152 500948
rect 402204 500936 402210 500948
rect 407390 500936 407396 500948
rect 402204 500908 407396 500936
rect 402204 500896 402210 500908
rect 407390 500896 407396 500908
rect 407448 500896 407454 500948
rect 553302 499808 553308 499860
rect 553360 499848 553366 499860
rect 557718 499848 557724 499860
rect 553360 499820 557724 499848
rect 553360 499808 553366 499820
rect 557718 499808 557724 499820
rect 557776 499808 557782 499860
rect 350442 499536 350448 499588
rect 350500 499576 350506 499588
rect 380526 499576 380532 499588
rect 350500 499548 380532 499576
rect 350500 499536 350506 499548
rect 380526 499536 380532 499548
rect 380584 499536 380590 499588
rect 348694 498516 348700 498568
rect 348752 498556 348758 498568
rect 349154 498556 349160 498568
rect 348752 498528 349160 498556
rect 348752 498516 348758 498528
rect 349154 498516 349160 498528
rect 349212 498516 349218 498568
rect 45922 498244 45928 498296
rect 45980 498284 45986 498296
rect 46474 498284 46480 498296
rect 45980 498256 46480 498284
rect 45980 498244 45986 498256
rect 46474 498244 46480 498256
rect 46532 498244 46538 498296
rect 350442 498176 350448 498228
rect 350500 498216 350506 498228
rect 355226 498216 355232 498228
rect 350500 498188 355232 498216
rect 350500 498176 350506 498188
rect 355226 498176 355232 498188
rect 355284 498176 355290 498228
rect 553302 498176 553308 498228
rect 553360 498216 553366 498228
rect 577314 498216 577320 498228
rect 553360 498188 577320 498216
rect 553360 498176 553366 498188
rect 577314 498176 577320 498188
rect 577372 498176 577378 498228
rect 42058 498108 42064 498160
rect 42116 498148 42122 498160
rect 46474 498148 46480 498160
rect 42116 498120 46480 498148
rect 42116 498108 42122 498120
rect 46474 498108 46480 498120
rect 46532 498108 46538 498160
rect 41046 496748 41052 496800
rect 41104 496788 41110 496800
rect 46474 496788 46480 496800
rect 41104 496760 46480 496788
rect 41104 496748 41110 496760
rect 46474 496748 46480 496760
rect 46532 496748 46538 496800
rect 552198 496544 552204 496596
rect 552256 496584 552262 496596
rect 555326 496584 555332 496596
rect 552256 496556 555332 496584
rect 552256 496544 552262 496556
rect 555326 496544 555332 496556
rect 555384 496544 555390 496596
rect 21726 495456 21732 495508
rect 21784 495496 21790 495508
rect 46106 495496 46112 495508
rect 21784 495468 46112 495496
rect 21784 495456 21790 495468
rect 46106 495456 46112 495468
rect 46164 495456 46170 495508
rect 350442 495456 350448 495508
rect 350500 495496 350506 495508
rect 387518 495496 387524 495508
rect 350500 495468 387524 495496
rect 350500 495456 350506 495468
rect 387518 495456 387524 495468
rect 387576 495456 387582 495508
rect 391842 495456 391848 495508
rect 391900 495496 391906 495508
rect 407298 495496 407304 495508
rect 391900 495468 407304 495496
rect 391900 495456 391906 495468
rect 407298 495456 407304 495468
rect 407356 495456 407362 495508
rect 553302 495456 553308 495508
rect 553360 495496 553366 495508
rect 563606 495496 563612 495508
rect 553360 495468 563612 495496
rect 553360 495456 553366 495468
rect 563606 495456 563612 495468
rect 563664 495456 563670 495508
rect 42518 495388 42524 495440
rect 42576 495428 42582 495440
rect 46474 495428 46480 495440
rect 42576 495400 46480 495428
rect 42576 495388 42582 495400
rect 46474 495388 46480 495400
rect 46532 495388 46538 495440
rect 350442 494504 350448 494556
rect 350500 494544 350506 494556
rect 355410 494544 355416 494556
rect 350500 494516 355416 494544
rect 350500 494504 350506 494516
rect 355410 494504 355416 494516
rect 355468 494504 355474 494556
rect 348602 493960 348608 494012
rect 348660 494000 348666 494012
rect 349430 494000 349436 494012
rect 348660 493972 349436 494000
rect 348660 493960 348666 493972
rect 349430 493960 349436 493972
rect 349488 493960 349494 494012
rect 24210 492668 24216 492720
rect 24268 492708 24274 492720
rect 46474 492708 46480 492720
rect 24268 492680 46480 492708
rect 24268 492668 24274 492680
rect 46474 492668 46480 492680
rect 46532 492668 46538 492720
rect 360930 492668 360936 492720
rect 360988 492708 360994 492720
rect 407298 492708 407304 492720
rect 360988 492680 407304 492708
rect 360988 492668 360994 492680
rect 407298 492668 407304 492680
rect 407356 492668 407362 492720
rect 552566 492668 552572 492720
rect 552624 492708 552630 492720
rect 581454 492708 581460 492720
rect 552624 492680 581460 492708
rect 552624 492668 552630 492680
rect 581454 492668 581460 492680
rect 581512 492668 581518 492720
rect 348970 491648 348976 491700
rect 349028 491688 349034 491700
rect 349890 491688 349896 491700
rect 349028 491660 349896 491688
rect 349028 491648 349034 491660
rect 349890 491648 349896 491660
rect 349948 491648 349954 491700
rect 350350 491376 350356 491428
rect 350408 491416 350414 491428
rect 353478 491416 353484 491428
rect 350408 491388 353484 491416
rect 350408 491376 350414 491388
rect 353478 491376 353484 491388
rect 353536 491376 353542 491428
rect 350442 491308 350448 491360
rect 350500 491348 350506 491360
rect 372430 491348 372436 491360
rect 350500 491320 372436 491348
rect 350500 491308 350506 491320
rect 372430 491308 372436 491320
rect 372488 491308 372494 491360
rect 350350 491240 350356 491292
rect 350408 491280 350414 491292
rect 352282 491280 352288 491292
rect 350408 491252 352288 491280
rect 350408 491240 350414 491252
rect 352282 491240 352288 491252
rect 352340 491240 352346 491292
rect 350442 489948 350448 490000
rect 350500 489988 350506 490000
rect 374822 489988 374828 490000
rect 350500 489960 374828 489988
rect 350500 489948 350506 489960
rect 374822 489948 374828 489960
rect 374880 489948 374886 490000
rect 28626 489880 28632 489932
rect 28684 489920 28690 489932
rect 46474 489920 46480 489932
rect 28684 489892 46480 489920
rect 28684 489880 28690 489892
rect 46474 489880 46480 489892
rect 46532 489880 46538 489932
rect 362310 489880 362316 489932
rect 362368 489920 362374 489932
rect 407298 489920 407304 489932
rect 362368 489892 407304 489920
rect 362368 489880 362374 489892
rect 407298 489880 407304 489892
rect 407356 489880 407362 489932
rect 348510 488860 348516 488912
rect 348568 488900 348574 488912
rect 349614 488900 349620 488912
rect 348568 488872 349620 488900
rect 348568 488860 348574 488872
rect 349614 488860 349620 488872
rect 349672 488860 349678 488912
rect 553302 488792 553308 488844
rect 553360 488832 553366 488844
rect 559190 488832 559196 488844
rect 553360 488804 559196 488832
rect 553360 488792 553366 488804
rect 559190 488792 559196 488804
rect 559248 488792 559254 488844
rect 391750 488520 391756 488572
rect 391808 488560 391814 488572
rect 407298 488560 407304 488572
rect 391808 488532 407304 488560
rect 391808 488520 391814 488532
rect 407298 488520 407304 488532
rect 407356 488520 407362 488572
rect 350442 488452 350448 488504
rect 350500 488492 350506 488504
rect 387426 488492 387432 488504
rect 350500 488464 387432 488492
rect 350500 488452 350506 488464
rect 387426 488452 387432 488464
rect 387484 488452 387490 488504
rect 39206 487772 39212 487824
rect 39264 487812 39270 487824
rect 45646 487812 45652 487824
rect 39264 487784 45652 487812
rect 39264 487772 39270 487784
rect 45646 487772 45652 487784
rect 45704 487772 45710 487824
rect 395982 487160 395988 487212
rect 396040 487200 396046 487212
rect 407298 487200 407304 487212
rect 396040 487172 407304 487200
rect 396040 487160 396046 487172
rect 407298 487160 407304 487172
rect 407356 487160 407362 487212
rect 553302 487160 553308 487212
rect 553360 487200 553366 487212
rect 573082 487200 573088 487212
rect 553360 487172 573088 487200
rect 553360 487160 553366 487172
rect 573082 487160 573088 487172
rect 573140 487160 573146 487212
rect 46474 486072 46480 486124
rect 46532 486112 46538 486124
rect 46750 486112 46756 486124
rect 46532 486084 46756 486112
rect 46532 486072 46538 486084
rect 46750 486072 46756 486084
rect 46808 486072 46814 486124
rect 19242 485800 19248 485852
rect 19300 485840 19306 485852
rect 46750 485840 46756 485852
rect 19300 485812 46756 485840
rect 19300 485800 19306 485812
rect 46750 485800 46756 485812
rect 46808 485800 46814 485852
rect 386322 485800 386328 485852
rect 386380 485840 386386 485852
rect 407298 485840 407304 485852
rect 386380 485812 407304 485840
rect 386380 485800 386386 485812
rect 407298 485800 407304 485812
rect 407356 485800 407362 485852
rect 405458 485732 405464 485784
rect 405516 485772 405522 485784
rect 407482 485772 407488 485784
rect 405516 485744 407488 485772
rect 405516 485732 405522 485744
rect 407482 485732 407488 485744
rect 407540 485732 407546 485784
rect 552842 484576 552848 484628
rect 552900 484616 552906 484628
rect 556246 484616 556252 484628
rect 552900 484588 556252 484616
rect 552900 484576 552906 484588
rect 556246 484576 556252 484588
rect 556304 484576 556310 484628
rect 42058 484440 42064 484492
rect 42116 484480 42122 484492
rect 46750 484480 46756 484492
rect 42116 484452 46756 484480
rect 42116 484440 42122 484452
rect 46750 484440 46756 484452
rect 46808 484440 46814 484492
rect 19058 484372 19064 484424
rect 19116 484412 19122 484424
rect 45830 484412 45836 484424
rect 19116 484384 45836 484412
rect 19116 484372 19122 484384
rect 45830 484372 45836 484384
rect 45888 484372 45894 484424
rect 349982 484372 349988 484424
rect 350040 484412 350046 484424
rect 352282 484412 352288 484424
rect 350040 484384 352288 484412
rect 350040 484372 350046 484384
rect 352282 484372 352288 484384
rect 352340 484372 352346 484424
rect 370682 484372 370688 484424
rect 370740 484412 370746 484424
rect 407298 484412 407304 484424
rect 370740 484384 407304 484412
rect 370740 484372 370746 484384
rect 407298 484372 407304 484384
rect 407356 484372 407362 484424
rect 551278 484304 551284 484356
rect 551336 484344 551342 484356
rect 552014 484344 552020 484356
rect 551336 484316 552020 484344
rect 551336 484304 551342 484316
rect 552014 484304 552020 484316
rect 552072 484304 552078 484356
rect 379054 483080 379060 483132
rect 379112 483120 379118 483132
rect 407298 483120 407304 483132
rect 379112 483092 407304 483120
rect 379112 483080 379118 483092
rect 407298 483080 407304 483092
rect 407356 483080 407362 483132
rect 350442 483012 350448 483064
rect 350500 483052 350506 483064
rect 386046 483052 386052 483064
rect 350500 483024 386052 483052
rect 350500 483012 350506 483024
rect 386046 483012 386052 483024
rect 386104 483012 386110 483064
rect 406010 483012 406016 483064
rect 406068 483052 406074 483064
rect 407850 483052 407856 483064
rect 406068 483024 407856 483052
rect 406068 483012 406074 483024
rect 407850 483012 407856 483024
rect 407908 483012 407914 483064
rect 552566 483012 552572 483064
rect 552624 483052 552630 483064
rect 575750 483052 575756 483064
rect 552624 483024 575756 483052
rect 552624 483012 552630 483024
rect 575750 483012 575756 483024
rect 575808 483012 575814 483064
rect 350442 481652 350448 481704
rect 350500 481692 350506 481704
rect 367278 481692 367284 481704
rect 350500 481664 367284 481692
rect 350500 481652 350506 481664
rect 367278 481652 367284 481664
rect 367336 481652 367342 481704
rect 384850 481652 384856 481704
rect 384908 481692 384914 481704
rect 407298 481692 407304 481704
rect 384908 481664 407304 481692
rect 384908 481652 384914 481664
rect 407298 481652 407304 481664
rect 407356 481652 407362 481704
rect 45002 481312 45008 481364
rect 45060 481352 45066 481364
rect 46474 481352 46480 481364
rect 45060 481324 46480 481352
rect 45060 481312 45066 481324
rect 46474 481312 46480 481324
rect 46532 481312 46538 481364
rect 40954 480632 40960 480684
rect 41012 480672 41018 480684
rect 46290 480672 46296 480684
rect 41012 480644 46296 480672
rect 41012 480632 41018 480644
rect 46290 480632 46296 480644
rect 46348 480632 46354 480684
rect 350074 480292 350080 480344
rect 350132 480332 350138 480344
rect 362954 480332 362960 480344
rect 350132 480304 362960 480332
rect 350132 480292 350138 480304
rect 362954 480292 362960 480304
rect 363012 480292 363018 480344
rect 38562 480224 38568 480276
rect 38620 480264 38626 480276
rect 46750 480264 46756 480276
rect 38620 480236 46756 480264
rect 38620 480224 38626 480236
rect 46750 480224 46756 480236
rect 46808 480224 46814 480276
rect 350442 480224 350448 480276
rect 350500 480264 350506 480276
rect 368750 480264 368756 480276
rect 350500 480236 368756 480264
rect 350500 480224 350506 480236
rect 368750 480224 368756 480236
rect 368808 480224 368814 480276
rect 553302 478864 553308 478916
rect 553360 478904 553366 478916
rect 577406 478904 577412 478916
rect 553360 478876 577412 478904
rect 553360 478864 553366 478876
rect 577406 478864 577412 478876
rect 577464 478864 577470 478916
rect 401410 477504 401416 477556
rect 401468 477544 401474 477556
rect 407298 477544 407304 477556
rect 401468 477516 407304 477544
rect 401468 477504 401474 477516
rect 407298 477504 407304 477516
rect 407356 477504 407362 477556
rect 552566 477504 552572 477556
rect 552624 477544 552630 477556
rect 563974 477544 563980 477556
rect 552624 477516 563980 477544
rect 552624 477504 552630 477516
rect 563974 477504 563980 477516
rect 564032 477504 564038 477556
rect 350074 476144 350080 476196
rect 350132 476184 350138 476196
rect 364518 476184 364524 476196
rect 350132 476156 364524 476184
rect 350132 476144 350138 476156
rect 364518 476144 364524 476156
rect 364576 476144 364582 476196
rect 350442 476076 350448 476128
rect 350500 476116 350506 476128
rect 377766 476116 377772 476128
rect 350500 476088 377772 476116
rect 350500 476076 350506 476088
rect 377766 476076 377772 476088
rect 377824 476076 377830 476128
rect 363874 474784 363880 474836
rect 363932 474824 363938 474836
rect 407298 474824 407304 474836
rect 363932 474796 407304 474824
rect 363932 474784 363938 474796
rect 407298 474784 407304 474796
rect 407356 474784 407362 474836
rect 553302 474784 553308 474836
rect 553360 474824 553366 474836
rect 563146 474824 563152 474836
rect 553360 474796 563152 474824
rect 553360 474784 553366 474796
rect 563146 474784 563152 474796
rect 563204 474784 563210 474836
rect 552934 474716 552940 474768
rect 552992 474756 552998 474768
rect 582926 474756 582932 474768
rect 552992 474728 582932 474756
rect 552992 474716 552998 474728
rect 582926 474716 582932 474728
rect 582984 474716 582990 474768
rect 43346 474648 43352 474700
rect 43404 474688 43410 474700
rect 46750 474688 46756 474700
rect 43404 474660 46756 474688
rect 43404 474648 43410 474660
rect 46750 474648 46756 474660
rect 46808 474648 46814 474700
rect 390462 473424 390468 473476
rect 390520 473464 390526 473476
rect 407298 473464 407304 473476
rect 390520 473436 407304 473464
rect 390520 473424 390526 473436
rect 407298 473424 407304 473436
rect 407356 473424 407362 473476
rect 350442 473356 350448 473408
rect 350500 473396 350506 473408
rect 356238 473396 356244 473408
rect 350500 473368 356244 473396
rect 350500 473356 350506 473368
rect 356238 473356 356244 473368
rect 356296 473356 356302 473408
rect 372246 473356 372252 473408
rect 372304 473396 372310 473408
rect 407390 473396 407396 473408
rect 372304 473368 407396 473396
rect 372304 473356 372310 473368
rect 407390 473356 407396 473368
rect 407448 473356 407454 473408
rect 384758 471996 384764 472048
rect 384816 472036 384822 472048
rect 407298 472036 407304 472048
rect 384816 472008 407304 472036
rect 384816 471996 384822 472008
rect 407298 471996 407304 472008
rect 407356 471996 407362 472048
rect 553302 470568 553308 470620
rect 553360 470608 553366 470620
rect 567838 470608 567844 470620
rect 553360 470580 567844 470608
rect 553360 470568 553366 470580
rect 567838 470568 567844 470580
rect 567896 470568 567902 470620
rect 570782 470568 570788 470620
rect 570840 470608 570846 470620
rect 580166 470608 580172 470620
rect 570840 470580 580172 470608
rect 570840 470568 570846 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 37642 469208 37648 469260
rect 37700 469248 37706 469260
rect 46750 469248 46756 469260
rect 37700 469220 46756 469248
rect 37700 469208 37706 469220
rect 46750 469208 46756 469220
rect 46808 469208 46814 469260
rect 365254 469208 365260 469260
rect 365312 469248 365318 469260
rect 407298 469248 407304 469260
rect 365312 469220 407304 469248
rect 365312 469208 365318 469220
rect 407298 469208 407304 469220
rect 407356 469208 407362 469260
rect 553302 469208 553308 469260
rect 553360 469248 553366 469260
rect 578326 469248 578332 469260
rect 553360 469220 578332 469248
rect 553360 469208 553366 469220
rect 578326 469208 578332 469220
rect 578384 469208 578390 469260
rect 39390 467916 39396 467968
rect 39448 467956 39454 467968
rect 46750 467956 46756 467968
rect 39448 467928 46756 467956
rect 39448 467916 39454 467928
rect 46750 467916 46756 467928
rect 46808 467916 46814 467968
rect 21634 467848 21640 467900
rect 21692 467888 21698 467900
rect 46658 467888 46664 467900
rect 21692 467860 46664 467888
rect 21692 467848 21698 467860
rect 46658 467848 46664 467860
rect 46716 467848 46722 467900
rect 386230 467848 386236 467900
rect 386288 467888 386294 467900
rect 407298 467888 407304 467900
rect 386288 467860 407304 467888
rect 386288 467848 386294 467860
rect 407298 467848 407304 467860
rect 407356 467848 407362 467900
rect 350442 466420 350448 466472
rect 350500 466460 350506 466472
rect 391198 466460 391204 466472
rect 350500 466432 391204 466460
rect 350500 466420 350506 466432
rect 391198 466420 391204 466432
rect 391256 466420 391262 466472
rect 553302 466420 553308 466472
rect 553360 466460 553366 466472
rect 567654 466460 567660 466472
rect 553360 466432 567660 466460
rect 553360 466420 553366 466432
rect 567654 466420 567660 466432
rect 567712 466420 567718 466472
rect 350074 466352 350080 466404
rect 350132 466392 350138 466404
rect 396902 466392 396908 466404
rect 350132 466364 396908 466392
rect 350132 466352 350138 466364
rect 396902 466352 396908 466364
rect 396960 466352 396966 466404
rect 350442 465060 350448 465112
rect 350500 465100 350506 465112
rect 371326 465100 371332 465112
rect 350500 465072 371332 465100
rect 350500 465060 350506 465072
rect 371326 465060 371332 465072
rect 371384 465060 371390 465112
rect 401318 465060 401324 465112
rect 401376 465100 401382 465112
rect 407298 465100 407304 465112
rect 401376 465072 407304 465100
rect 401376 465060 401382 465072
rect 407298 465060 407304 465072
rect 407356 465060 407362 465112
rect 552014 465060 552020 465112
rect 552072 465100 552078 465112
rect 574462 465100 574468 465112
rect 552072 465072 574468 465100
rect 552072 465060 552078 465072
rect 574462 465060 574468 465072
rect 574520 465060 574526 465112
rect 40954 464108 40960 464160
rect 41012 464148 41018 464160
rect 46750 464148 46756 464160
rect 41012 464120 46756 464148
rect 41012 464108 41018 464120
rect 46750 464108 46756 464120
rect 46808 464108 46814 464160
rect 552014 463904 552020 463956
rect 552072 463944 552078 463956
rect 556338 463944 556344 463956
rect 552072 463916 556344 463944
rect 552072 463904 552078 463916
rect 556338 463904 556344 463916
rect 556396 463904 556402 463956
rect 21542 463700 21548 463752
rect 21600 463740 21606 463752
rect 46750 463740 46756 463752
rect 21600 463712 46756 463740
rect 21600 463700 21606 463712
rect 46750 463700 46756 463712
rect 46808 463700 46814 463752
rect 383286 463700 383292 463752
rect 383344 463740 383350 463752
rect 407298 463740 407304 463752
rect 383344 463712 407304 463740
rect 383344 463700 383350 463712
rect 407298 463700 407304 463712
rect 407356 463700 407362 463752
rect 36814 463632 36820 463684
rect 36872 463672 36878 463684
rect 46658 463672 46664 463684
rect 36872 463644 46664 463672
rect 36872 463632 36878 463644
rect 46658 463632 46664 463644
rect 46716 463632 46722 463684
rect 350074 462408 350080 462460
rect 350132 462448 350138 462460
rect 369210 462448 369216 462460
rect 350132 462420 369216 462448
rect 350132 462408 350138 462420
rect 369210 462408 369216 462420
rect 369268 462408 369274 462460
rect 403802 462408 403808 462460
rect 403860 462448 403866 462460
rect 407390 462448 407396 462460
rect 403860 462420 407396 462448
rect 403860 462408 403866 462420
rect 407390 462408 407396 462420
rect 407448 462408 407454 462460
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 19978 462380 19984 462392
rect 3568 462352 19984 462380
rect 3568 462340 3574 462352
rect 19978 462340 19984 462352
rect 20036 462340 20042 462392
rect 350442 462340 350448 462392
rect 350500 462380 350506 462392
rect 386138 462380 386144 462392
rect 350500 462352 386144 462380
rect 350500 462340 350506 462352
rect 386138 462340 386144 462352
rect 386196 462340 386202 462392
rect 396902 462340 396908 462392
rect 396960 462380 396966 462392
rect 407298 462380 407304 462392
rect 396960 462352 407304 462380
rect 396960 462340 396966 462352
rect 407298 462340 407304 462352
rect 407356 462340 407362 462392
rect 552014 462340 552020 462392
rect 552072 462380 552078 462392
rect 574646 462380 574652 462392
rect 552072 462352 574652 462380
rect 552072 462340 552078 462352
rect 574646 462340 574652 462352
rect 574704 462340 574710 462392
rect 350442 460980 350448 461032
rect 350500 461020 350506 461032
rect 363046 461020 363052 461032
rect 350500 460992 363052 461020
rect 350500 460980 350506 460992
rect 363046 460980 363052 460992
rect 363104 460980 363110 461032
rect 24578 460912 24584 460964
rect 24636 460952 24642 460964
rect 46750 460952 46756 460964
rect 24636 460924 46756 460952
rect 24636 460912 24642 460924
rect 46750 460912 46756 460924
rect 46808 460912 46814 460964
rect 350074 460912 350080 460964
rect 350132 460952 350138 460964
rect 371418 460952 371424 460964
rect 350132 460924 371424 460952
rect 350132 460912 350138 460924
rect 371418 460912 371424 460924
rect 371476 460912 371482 460964
rect 38470 460844 38476 460896
rect 38528 460884 38534 460896
rect 46658 460884 46664 460896
rect 38528 460856 46664 460884
rect 38528 460844 38534 460856
rect 46658 460844 46664 460856
rect 46716 460844 46722 460896
rect 552198 459620 552204 459672
rect 552256 459660 552262 459672
rect 573266 459660 573272 459672
rect 552256 459632 573272 459660
rect 552256 459620 552262 459632
rect 573266 459620 573272 459632
rect 573324 459620 573330 459672
rect 350442 459552 350448 459604
rect 350500 459592 350506 459604
rect 373810 459592 373816 459604
rect 350500 459564 373816 459592
rect 350500 459552 350506 459564
rect 373810 459552 373816 459564
rect 373868 459552 373874 459604
rect 552014 459552 552020 459604
rect 552072 459592 552078 459604
rect 581270 459592 581276 459604
rect 552072 459564 581276 459592
rect 552072 459552 552078 459564
rect 581270 459552 581276 459564
rect 581328 459552 581334 459604
rect 552014 459008 552020 459060
rect 552072 459048 552078 459060
rect 553946 459048 553952 459060
rect 552072 459020 553952 459048
rect 552072 459008 552078 459020
rect 553946 459008 553952 459020
rect 554004 459008 554010 459060
rect 551278 458328 551284 458380
rect 551336 458368 551342 458380
rect 553026 458368 553032 458380
rect 551336 458340 553032 458368
rect 551336 458328 551342 458340
rect 553026 458328 553032 458340
rect 553084 458328 553090 458380
rect 402698 458192 402704 458244
rect 402756 458232 402762 458244
rect 407298 458232 407304 458244
rect 402756 458204 407304 458232
rect 402756 458192 402762 458204
rect 407298 458192 407304 458204
rect 407356 458192 407362 458244
rect 350442 457240 350448 457292
rect 350500 457280 350506 457292
rect 356330 457280 356336 457292
rect 350500 457252 356336 457280
rect 350500 457240 350506 457252
rect 356330 457240 356336 457252
rect 356388 457240 356394 457292
rect 372338 456764 372344 456816
rect 372396 456804 372402 456816
rect 407298 456804 407304 456816
rect 372396 456776 407304 456804
rect 372396 456764 372402 456776
rect 407298 456764 407304 456776
rect 407356 456764 407362 456816
rect 552014 456764 552020 456816
rect 552072 456804 552078 456816
rect 576210 456804 576216 456816
rect 552072 456776 576216 456804
rect 552072 456764 552078 456776
rect 576210 456764 576216 456776
rect 576268 456764 576274 456816
rect 43622 456696 43628 456748
rect 43680 456736 43686 456748
rect 46658 456736 46664 456748
rect 43680 456708 46664 456736
rect 43680 456696 43686 456708
rect 46658 456696 46664 456708
rect 46716 456696 46722 456748
rect 387518 456696 387524 456748
rect 387576 456736 387582 456748
rect 407390 456736 407396 456748
rect 387576 456708 407396 456736
rect 387576 456696 387582 456708
rect 407390 456696 407396 456708
rect 407448 456696 407454 456748
rect 40862 456628 40868 456680
rect 40920 456668 40926 456680
rect 46750 456668 46756 456680
rect 40920 456640 46756 456668
rect 40920 456628 40926 456640
rect 46750 456628 46756 456640
rect 46808 456628 46814 456680
rect 552014 456288 552020 456340
rect 552072 456328 552078 456340
rect 553854 456328 553860 456340
rect 552072 456300 553860 456328
rect 552072 456288 552078 456300
rect 553854 456288 553860 456300
rect 553912 456288 553918 456340
rect 349062 456084 349068 456136
rect 349120 456124 349126 456136
rect 352006 456124 352012 456136
rect 349120 456096 352012 456124
rect 349120 456084 349126 456096
rect 352006 456084 352012 456096
rect 352064 456084 352070 456136
rect 379146 455336 379152 455388
rect 379204 455376 379210 455388
rect 407390 455376 407396 455388
rect 379204 455348 407396 455376
rect 379204 455336 379210 455348
rect 407390 455336 407396 455348
rect 407448 455336 407454 455388
rect 350442 454112 350448 454164
rect 350500 454152 350506 454164
rect 380802 454152 380808 454164
rect 350500 454124 380808 454152
rect 350500 454112 350506 454124
rect 380802 454112 380808 454124
rect 380860 454112 380866 454164
rect 375282 454044 375288 454096
rect 375340 454084 375346 454096
rect 407298 454084 407304 454096
rect 375340 454056 407304 454084
rect 375340 454044 375346 454056
rect 407298 454044 407304 454056
rect 407356 454044 407362 454096
rect 552474 454044 552480 454096
rect 552532 454084 552538 454096
rect 565998 454084 566004 454096
rect 552532 454056 566004 454084
rect 552532 454044 552538 454056
rect 565998 454044 566004 454056
rect 566056 454044 566062 454096
rect 405458 452616 405464 452668
rect 405516 452656 405522 452668
rect 407666 452656 407672 452668
rect 405516 452628 407672 452656
rect 405516 452616 405522 452628
rect 407666 452616 407672 452628
rect 407724 452616 407730 452668
rect 552566 452616 552572 452668
rect 552624 452656 552630 452668
rect 559282 452656 559288 452668
rect 552624 452628 559288 452656
rect 552624 452616 552630 452628
rect 559282 452616 559288 452628
rect 559340 452616 559346 452668
rect 377858 451324 377864 451376
rect 377916 451364 377922 451376
rect 407298 451364 407304 451376
rect 377916 451336 407304 451364
rect 377916 451324 377922 451336
rect 407298 451324 407304 451336
rect 407356 451324 407362 451376
rect 350442 451256 350448 451308
rect 350500 451296 350506 451308
rect 380342 451296 380348 451308
rect 350500 451268 380348 451296
rect 350500 451256 350506 451268
rect 380342 451256 380348 451268
rect 380400 451256 380406 451308
rect 32582 451188 32588 451240
rect 32640 451228 32646 451240
rect 46750 451228 46756 451240
rect 32640 451200 46756 451228
rect 32640 451188 32646 451200
rect 46750 451188 46756 451200
rect 46808 451188 46814 451240
rect 350442 451120 350448 451172
rect 350500 451160 350506 451172
rect 353754 451160 353760 451172
rect 350500 451132 353760 451160
rect 350500 451120 350506 451132
rect 353754 451120 353760 451132
rect 353812 451120 353818 451172
rect 350442 449896 350448 449948
rect 350500 449936 350506 449948
rect 374546 449936 374552 449948
rect 350500 449908 374552 449936
rect 350500 449896 350506 449908
rect 374546 449896 374552 449908
rect 374604 449896 374610 449948
rect 553302 448604 553308 448656
rect 553360 448644 553366 448656
rect 561766 448644 561772 448656
rect 553360 448616 561772 448644
rect 553360 448604 553366 448616
rect 561766 448604 561772 448616
rect 561824 448604 561830 448656
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 20070 448576 20076 448588
rect 3200 448548 20076 448576
rect 3200 448536 3206 448548
rect 20070 448536 20076 448548
rect 20128 448536 20134 448588
rect 385586 448536 385592 448588
rect 385644 448576 385650 448588
rect 407298 448576 407304 448588
rect 385644 448548 407304 448576
rect 385644 448536 385650 448548
rect 407298 448536 407304 448548
rect 407356 448536 407362 448588
rect 553026 448536 553032 448588
rect 553084 448576 553090 448588
rect 570230 448576 570236 448588
rect 553084 448548 570236 448576
rect 553084 448536 553090 448548
rect 570230 448536 570236 448548
rect 570288 448536 570294 448588
rect 350442 447108 350448 447160
rect 350500 447148 350506 447160
rect 365898 447148 365904 447160
rect 350500 447120 365904 447148
rect 350500 447108 350506 447120
rect 365898 447108 365904 447120
rect 365956 447108 365962 447160
rect 379422 447108 379428 447160
rect 379480 447148 379486 447160
rect 407298 447148 407304 447160
rect 379480 447120 407304 447148
rect 379480 447108 379486 447120
rect 407298 447108 407304 447120
rect 407356 447108 407362 447160
rect 395522 447040 395528 447092
rect 395580 447080 395586 447092
rect 407390 447080 407396 447092
rect 395580 447052 407396 447080
rect 395580 447040 395586 447052
rect 407390 447040 407396 447052
rect 407448 447040 407454 447092
rect 350442 445816 350448 445868
rect 350500 445856 350506 445868
rect 366726 445856 366732 445868
rect 350500 445828 366732 445856
rect 350500 445816 350506 445828
rect 366726 445816 366732 445828
rect 366784 445816 366790 445868
rect 44726 445748 44732 445800
rect 44784 445788 44790 445800
rect 46474 445788 46480 445800
rect 44784 445760 46480 445788
rect 44784 445748 44790 445760
rect 46474 445748 46480 445760
rect 46532 445748 46538 445800
rect 350074 445748 350080 445800
rect 350132 445788 350138 445800
rect 375374 445788 375380 445800
rect 350132 445760 375380 445788
rect 350132 445748 350138 445760
rect 375374 445748 375380 445760
rect 375432 445748 375438 445800
rect 350442 445680 350448 445732
rect 350500 445720 350506 445732
rect 400950 445720 400956 445732
rect 350500 445692 400956 445720
rect 350500 445680 350506 445692
rect 400950 445680 400956 445692
rect 401008 445680 401014 445732
rect 396994 445612 397000 445664
rect 397052 445652 397058 445664
rect 407298 445652 407304 445664
rect 397052 445624 407304 445652
rect 397052 445612 397058 445624
rect 407298 445612 407304 445624
rect 407356 445612 407362 445664
rect 27062 444388 27068 444440
rect 27120 444428 27126 444440
rect 45922 444428 45928 444440
rect 27120 444400 45928 444428
rect 27120 444388 27126 444400
rect 45922 444388 45928 444400
rect 45980 444388 45986 444440
rect 552566 444388 552572 444440
rect 552624 444428 552630 444440
rect 583018 444428 583024 444440
rect 552624 444400 583024 444428
rect 552624 444388 552630 444400
rect 583018 444388 583024 444400
rect 583076 444388 583082 444440
rect 24486 442960 24492 443012
rect 24544 443000 24550 443012
rect 46750 443000 46756 443012
rect 24544 442972 46756 443000
rect 24544 442960 24550 442972
rect 46750 442960 46756 442972
rect 46808 442960 46814 443012
rect 553302 442960 553308 443012
rect 553360 443000 553366 443012
rect 573358 443000 573364 443012
rect 553360 442972 573364 443000
rect 553360 442960 553366 442972
rect 573358 442960 573364 442972
rect 573416 442960 573422 443012
rect 350442 441600 350448 441652
rect 350500 441640 350506 441652
rect 368842 441640 368848 441652
rect 350500 441612 368848 441640
rect 350500 441600 350506 441612
rect 368842 441600 368848 441612
rect 368900 441600 368906 441652
rect 370774 441600 370780 441652
rect 370832 441640 370838 441652
rect 407298 441640 407304 441652
rect 370832 441612 407304 441640
rect 370832 441600 370838 441612
rect 407298 441600 407304 441612
rect 407356 441600 407362 441652
rect 401134 441532 401140 441584
rect 401192 441572 401198 441584
rect 407390 441572 407396 441584
rect 401192 441544 407396 441572
rect 401192 441532 401198 441544
rect 407390 441532 407396 441544
rect 407448 441532 407454 441584
rect 350442 440240 350448 440292
rect 350500 440280 350506 440292
rect 382090 440280 382096 440292
rect 350500 440252 382096 440280
rect 350500 440240 350506 440252
rect 382090 440240 382096 440252
rect 382148 440240 382154 440292
rect 42518 438880 42524 438932
rect 42576 438920 42582 438932
rect 45922 438920 45928 438932
rect 42576 438892 45928 438920
rect 42576 438880 42582 438892
rect 45922 438880 45928 438892
rect 45980 438880 45986 438932
rect 374914 438880 374920 438932
rect 374972 438920 374978 438932
rect 407206 438920 407212 438932
rect 374972 438892 407212 438920
rect 374972 438880 374978 438892
rect 407206 438880 407212 438892
rect 407264 438880 407270 438932
rect 404998 438812 405004 438864
rect 405056 438852 405062 438864
rect 407482 438852 407488 438864
rect 405056 438824 407488 438852
rect 405056 438812 405062 438824
rect 407482 438812 407488 438824
rect 407540 438812 407546 438864
rect 553302 438064 553308 438116
rect 553360 438104 553366 438116
rect 557994 438104 558000 438116
rect 553360 438076 558000 438104
rect 553360 438064 553366 438076
rect 557994 438064 558000 438076
rect 558052 438064 558058 438116
rect 350074 437452 350080 437504
rect 350132 437492 350138 437504
rect 387610 437492 387616 437504
rect 350132 437464 387616 437492
rect 350132 437452 350138 437464
rect 387610 437452 387616 437464
rect 387668 437452 387674 437504
rect 393038 437452 393044 437504
rect 393096 437492 393102 437504
rect 407206 437492 407212 437504
rect 393096 437464 407212 437492
rect 393096 437452 393102 437464
rect 407206 437452 407212 437464
rect 407264 437452 407270 437504
rect 553302 437452 553308 437504
rect 553360 437492 553366 437504
rect 562226 437492 562232 437504
rect 553360 437464 562232 437492
rect 553360 437452 553366 437464
rect 562226 437452 562232 437464
rect 562284 437452 562290 437504
rect 350442 437384 350448 437436
rect 350500 437424 350506 437436
rect 403710 437424 403716 437436
rect 350500 437396 403716 437424
rect 350500 437384 350506 437396
rect 403710 437384 403716 437396
rect 403768 437384 403774 437436
rect 43622 436092 43628 436144
rect 43680 436132 43686 436144
rect 46750 436132 46756 436144
rect 43680 436104 46756 436132
rect 43680 436092 43686 436104
rect 46750 436092 46756 436104
rect 46808 436092 46814 436144
rect 373626 436092 373632 436144
rect 373684 436132 373690 436144
rect 407206 436132 407212 436144
rect 373684 436104 407212 436132
rect 373684 436092 373690 436104
rect 407206 436092 407212 436104
rect 407264 436092 407270 436144
rect 552658 436092 552664 436144
rect 552716 436132 552722 436144
rect 563514 436132 563520 436144
rect 552716 436104 563520 436132
rect 552716 436092 552722 436104
rect 563514 436092 563520 436104
rect 563572 436092 563578 436144
rect 39850 434732 39856 434784
rect 39908 434772 39914 434784
rect 46750 434772 46756 434784
rect 39908 434744 46756 434772
rect 39908 434732 39914 434744
rect 46750 434732 46756 434744
rect 46808 434732 46814 434784
rect 350442 434732 350448 434784
rect 350500 434772 350506 434784
rect 372706 434772 372712 434784
rect 350500 434744 372712 434772
rect 350500 434732 350506 434744
rect 372706 434732 372712 434744
rect 372764 434732 372770 434784
rect 388806 434732 388812 434784
rect 388864 434772 388870 434784
rect 407206 434772 407212 434784
rect 388864 434744 407212 434772
rect 388864 434732 388870 434744
rect 407206 434732 407212 434744
rect 407264 434732 407270 434784
rect 552658 434732 552664 434784
rect 552716 434772 552722 434784
rect 581362 434772 581368 434784
rect 552716 434744 581368 434772
rect 552716 434732 552722 434744
rect 581362 434732 581368 434744
rect 581420 434732 581426 434784
rect 37918 433304 37924 433356
rect 37976 433344 37982 433356
rect 46750 433344 46756 433356
rect 37976 433316 46756 433344
rect 37976 433304 37982 433316
rect 46750 433304 46756 433316
rect 46808 433304 46814 433356
rect 405274 432488 405280 432540
rect 405332 432528 405338 432540
rect 407206 432528 407212 432540
rect 405332 432500 407212 432528
rect 405332 432488 405338 432500
rect 407206 432488 407212 432500
rect 407264 432488 407270 432540
rect 28902 431944 28908 431996
rect 28960 431984 28966 431996
rect 46382 431984 46388 431996
rect 28960 431956 46388 431984
rect 28960 431944 28966 431956
rect 46382 431944 46388 431956
rect 46440 431944 46446 431996
rect 576302 431876 576308 431928
rect 576360 431916 576366 431928
rect 580166 431916 580172 431928
rect 576360 431888 580172 431916
rect 576360 431876 576366 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 350442 430652 350448 430704
rect 350500 430692 350506 430704
rect 361022 430692 361028 430704
rect 350500 430664 361028 430692
rect 350500 430652 350506 430664
rect 361022 430652 361028 430664
rect 361080 430652 361086 430704
rect 350074 430584 350080 430636
rect 350132 430624 350138 430636
rect 363966 430624 363972 430636
rect 350132 430596 363972 430624
rect 350132 430584 350138 430596
rect 363966 430584 363972 430596
rect 364024 430584 364030 430636
rect 43898 430516 43904 430568
rect 43956 430556 43962 430568
rect 46382 430556 46388 430568
rect 43956 430528 46388 430556
rect 43956 430516 43962 430528
rect 46382 430516 46388 430528
rect 46440 430516 46446 430568
rect 32582 429156 32588 429208
rect 32640 429196 32646 429208
rect 46750 429196 46756 429208
rect 32640 429168 46756 429196
rect 32640 429156 32646 429168
rect 46750 429156 46756 429168
rect 46808 429156 46814 429208
rect 397178 427864 397184 427916
rect 397236 427904 397242 427916
rect 407206 427904 407212 427916
rect 397236 427876 407212 427904
rect 397236 427864 397242 427876
rect 407206 427864 407212 427876
rect 407264 427864 407270 427916
rect 36722 427796 36728 427848
rect 36780 427836 36786 427848
rect 46750 427836 46756 427848
rect 36780 427808 46756 427836
rect 36780 427796 36786 427808
rect 46750 427796 46756 427808
rect 46808 427796 46814 427848
rect 350442 427796 350448 427848
rect 350500 427836 350506 427848
rect 404998 427836 405004 427848
rect 350500 427808 405004 427836
rect 350500 427796 350506 427808
rect 404998 427796 405004 427808
rect 405056 427796 405062 427848
rect 373718 426572 373724 426624
rect 373776 426612 373782 426624
rect 407298 426612 407304 426624
rect 373776 426584 407304 426612
rect 373776 426572 373782 426584
rect 407298 426572 407304 426584
rect 407356 426572 407362 426624
rect 370866 426504 370872 426556
rect 370924 426544 370930 426556
rect 407206 426544 407212 426556
rect 370924 426516 407212 426544
rect 370924 426504 370930 426516
rect 407206 426504 407212 426516
rect 407264 426504 407270 426556
rect 350442 426436 350448 426488
rect 350500 426476 350506 426488
rect 403710 426476 403716 426488
rect 350500 426448 403716 426476
rect 350500 426436 350506 426448
rect 403710 426436 403716 426448
rect 403768 426436 403774 426488
rect 553026 426436 553032 426488
rect 553084 426476 553090 426488
rect 574830 426476 574836 426488
rect 553084 426448 574836 426476
rect 553084 426436 553090 426448
rect 574830 426436 574836 426448
rect 574888 426436 574894 426488
rect 408402 426368 408408 426420
rect 408460 426408 408466 426420
rect 409138 426408 409144 426420
rect 408460 426380 409144 426408
rect 408460 426368 408466 426380
rect 409138 426368 409144 426380
rect 409196 426368 409202 426420
rect 40862 425076 40868 425128
rect 40920 425116 40926 425128
rect 46750 425116 46756 425128
rect 40920 425088 46756 425116
rect 40920 425076 40926 425088
rect 46750 425076 46756 425088
rect 46808 425076 46814 425128
rect 350442 425076 350448 425128
rect 350500 425116 350506 425128
rect 360654 425116 360660 425128
rect 350500 425088 360660 425116
rect 350500 425076 350506 425088
rect 360654 425076 360660 425088
rect 360712 425076 360718 425128
rect 395890 425076 395896 425128
rect 395948 425116 395954 425128
rect 407206 425116 407212 425128
rect 395948 425088 407212 425116
rect 395948 425076 395954 425088
rect 407206 425076 407212 425088
rect 407264 425076 407270 425128
rect 553026 425076 553032 425128
rect 553084 425116 553090 425128
rect 568942 425116 568948 425128
rect 553084 425088 568948 425116
rect 553084 425076 553090 425088
rect 568942 425076 568948 425088
rect 569000 425076 569006 425128
rect 35250 425008 35256 425060
rect 35308 425048 35314 425060
rect 46658 425048 46664 425060
rect 35308 425020 46664 425048
rect 35308 425008 35314 425020
rect 46658 425008 46664 425020
rect 46716 425008 46722 425060
rect 552934 423716 552940 423768
rect 552992 423756 552998 423768
rect 569034 423756 569040 423768
rect 552992 423728 569040 423756
rect 552992 423716 552998 423728
rect 569034 423716 569040 423728
rect 569092 423716 569098 423768
rect 26970 423648 26976 423700
rect 27028 423688 27034 423700
rect 46750 423688 46756 423700
rect 27028 423660 46756 423688
rect 27028 423648 27034 423660
rect 46750 423648 46756 423660
rect 46808 423648 46814 423700
rect 380710 423648 380716 423700
rect 380768 423688 380774 423700
rect 407206 423688 407212 423700
rect 380768 423660 407212 423688
rect 380768 423648 380774 423660
rect 407206 423648 407212 423660
rect 407264 423648 407270 423700
rect 553026 423648 553032 423700
rect 553084 423688 553090 423700
rect 570690 423688 570696 423700
rect 553084 423660 570696 423688
rect 553084 423648 553090 423660
rect 570690 423648 570696 423660
rect 570748 423648 570754 423700
rect 350442 422288 350448 422340
rect 350500 422328 350506 422340
rect 365438 422328 365444 422340
rect 350500 422300 365444 422328
rect 350500 422288 350506 422300
rect 365438 422288 365444 422300
rect 365496 422288 365502 422340
rect 390278 422288 390284 422340
rect 390336 422328 390342 422340
rect 407206 422328 407212 422340
rect 390336 422300 407212 422328
rect 390336 422288 390342 422300
rect 407206 422288 407212 422300
rect 407264 422288 407270 422340
rect 34974 421540 34980 421592
rect 35032 421580 35038 421592
rect 40586 421580 40592 421592
rect 35032 421552 40592 421580
rect 35032 421540 35038 421552
rect 40586 421540 40592 421552
rect 40644 421540 40650 421592
rect 350074 420996 350080 421048
rect 350132 421036 350138 421048
rect 353754 421036 353760 421048
rect 350132 421008 353760 421036
rect 350132 420996 350138 421008
rect 353754 420996 353760 421008
rect 353812 420996 353818 421048
rect 552290 420996 552296 421048
rect 552348 421036 552354 421048
rect 555234 421036 555240 421048
rect 552348 421008 555240 421036
rect 552348 420996 552354 421008
rect 555234 420996 555240 421008
rect 555292 420996 555298 421048
rect 35250 420928 35256 420980
rect 35308 420968 35314 420980
rect 46750 420968 46756 420980
rect 35308 420940 46756 420968
rect 35308 420928 35314 420940
rect 46750 420928 46756 420940
rect 46808 420928 46814 420980
rect 350442 420928 350448 420980
rect 350500 420968 350506 420980
rect 369302 420968 369308 420980
rect 350500 420940 369308 420968
rect 350500 420928 350506 420940
rect 369302 420928 369308 420940
rect 369360 420928 369366 420980
rect 570874 420180 570880 420232
rect 570932 420220 570938 420232
rect 580442 420220 580448 420232
rect 570932 420192 580448 420220
rect 570932 420180 570938 420192
rect 580442 420180 580448 420192
rect 580500 420180 580506 420232
rect 553026 419840 553032 419892
rect 553084 419880 553090 419892
rect 558086 419880 558092 419892
rect 553084 419852 558092 419880
rect 553084 419840 553090 419852
rect 558086 419840 558092 419852
rect 558144 419840 558150 419892
rect 40586 419568 40592 419620
rect 40644 419608 40650 419620
rect 46658 419608 46664 419620
rect 40644 419580 46664 419608
rect 40644 419568 40650 419580
rect 46658 419568 46664 419580
rect 46716 419568 46722 419620
rect 376386 419568 376392 419620
rect 376444 419608 376450 419620
rect 407298 419608 407304 419620
rect 376444 419580 407304 419608
rect 376444 419568 376450 419580
rect 407298 419568 407304 419580
rect 407356 419568 407362 419620
rect 28442 419500 28448 419552
rect 28500 419540 28506 419552
rect 46750 419540 46756 419552
rect 28500 419512 46756 419540
rect 28500 419500 28506 419512
rect 46750 419500 46756 419512
rect 46808 419500 46814 419552
rect 350442 419500 350448 419552
rect 350500 419540 350506 419552
rect 361942 419540 361948 419552
rect 350500 419512 361948 419540
rect 350500 419500 350506 419512
rect 361942 419500 361948 419512
rect 362000 419500 362006 419552
rect 362402 419500 362408 419552
rect 362460 419540 362466 419552
rect 407206 419540 407212 419552
rect 362460 419512 407212 419540
rect 362460 419500 362466 419512
rect 407206 419500 407212 419512
rect 407264 419500 407270 419552
rect 36814 418208 36820 418260
rect 36872 418248 36878 418260
rect 46658 418248 46664 418260
rect 36872 418220 46664 418248
rect 36872 418208 36878 418220
rect 46658 418208 46664 418220
rect 46716 418208 46722 418260
rect 388898 418208 388904 418260
rect 388956 418248 388962 418260
rect 407206 418248 407212 418260
rect 388956 418220 407212 418248
rect 388956 418208 388962 418220
rect 407206 418208 407212 418220
rect 407264 418208 407270 418260
rect 33686 418140 33692 418192
rect 33744 418180 33750 418192
rect 46750 418180 46756 418192
rect 33744 418152 46756 418180
rect 33744 418140 33750 418152
rect 46750 418140 46756 418152
rect 46808 418140 46814 418192
rect 350442 418140 350448 418192
rect 350500 418180 350506 418192
rect 400950 418180 400956 418192
rect 350500 418152 400956 418180
rect 350500 418140 350506 418152
rect 400950 418140 400956 418152
rect 401008 418140 401014 418192
rect 350442 416780 350448 416832
rect 350500 416820 350506 416832
rect 377950 416820 377956 416832
rect 350500 416792 377956 416820
rect 350500 416780 350506 416792
rect 377950 416780 377956 416792
rect 378008 416780 378014 416832
rect 405090 416712 405096 416764
rect 405148 416752 405154 416764
rect 407574 416752 407580 416764
rect 405148 416724 407580 416752
rect 405148 416712 405154 416724
rect 407574 416712 407580 416724
rect 407632 416712 407638 416764
rect 552014 416032 552020 416084
rect 552072 416072 552078 416084
rect 559650 416072 559656 416084
rect 552072 416044 559656 416072
rect 552072 416032 552078 416044
rect 559650 416032 559656 416044
rect 559708 416032 559714 416084
rect 43898 415488 43904 415540
rect 43956 415528 43962 415540
rect 46750 415528 46756 415540
rect 43956 415500 46756 415528
rect 43956 415488 43962 415500
rect 46750 415488 46756 415500
rect 46808 415488 46814 415540
rect 24394 415420 24400 415472
rect 24452 415460 24458 415472
rect 46658 415460 46664 415472
rect 24452 415432 46664 415460
rect 24452 415420 24458 415432
rect 46658 415420 46664 415432
rect 46716 415420 46722 415472
rect 552014 415420 552020 415472
rect 552072 415460 552078 415472
rect 566090 415460 566096 415472
rect 552072 415432 566096 415460
rect 552072 415420 552078 415432
rect 566090 415420 566096 415432
rect 566148 415420 566154 415472
rect 350442 414400 350448 414452
rect 350500 414440 350506 414452
rect 356790 414440 356796 414452
rect 350500 414412 356796 414440
rect 350500 414400 350506 414412
rect 356790 414400 356796 414412
rect 356848 414400 356854 414452
rect 20438 413992 20444 414044
rect 20496 414032 20502 414044
rect 46750 414032 46756 414044
rect 20496 414004 46756 414032
rect 20496 413992 20502 414004
rect 46750 413992 46756 414004
rect 46808 413992 46814 414044
rect 350442 413992 350448 414044
rect 350500 414032 350506 414044
rect 383470 414032 383476 414044
rect 350500 414004 383476 414032
rect 350500 413992 350506 414004
rect 383470 413992 383476 414004
rect 383528 413992 383534 414044
rect 387702 413992 387708 414044
rect 387760 414032 387766 414044
rect 407206 414032 407212 414044
rect 387760 414004 407212 414032
rect 387760 413992 387766 414004
rect 407206 413992 407212 414004
rect 407264 413992 407270 414044
rect 552014 412768 552020 412820
rect 552072 412808 552078 412820
rect 555326 412808 555332 412820
rect 552072 412780 555332 412808
rect 552072 412768 552078 412780
rect 555326 412768 555332 412780
rect 555384 412768 555390 412820
rect 552198 412632 552204 412684
rect 552256 412672 552262 412684
rect 578602 412672 578608 412684
rect 552256 412644 578608 412672
rect 552256 412632 552262 412644
rect 578602 412632 578608 412644
rect 578660 412632 578666 412684
rect 406194 411340 406200 411392
rect 406252 411380 406258 411392
rect 407298 411380 407304 411392
rect 406252 411352 407304 411380
rect 406252 411340 406258 411352
rect 407298 411340 407304 411352
rect 407356 411340 407362 411392
rect 31478 411272 31484 411324
rect 31536 411312 31542 411324
rect 46566 411312 46572 411324
rect 31536 411284 46572 411312
rect 31536 411272 31542 411284
rect 46566 411272 46572 411284
rect 46624 411272 46630 411324
rect 350442 411272 350448 411324
rect 350500 411312 350506 411324
rect 390186 411312 390192 411324
rect 350500 411284 390192 411312
rect 350500 411272 350506 411284
rect 390186 411272 390192 411284
rect 390244 411272 390250 411324
rect 391658 411272 391664 411324
rect 391716 411312 391722 411324
rect 407206 411312 407212 411324
rect 391716 411284 407212 411312
rect 391716 411272 391722 411284
rect 407206 411272 407212 411284
rect 407264 411272 407270 411324
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 31110 411244 31116 411256
rect 3016 411216 31116 411244
rect 3016 411204 3022 411216
rect 31110 411204 31116 411216
rect 31168 411204 31174 411256
rect 387518 409844 387524 409896
rect 387576 409884 387582 409896
rect 407206 409884 407212 409896
rect 387576 409856 407212 409884
rect 387576 409844 387582 409856
rect 407206 409844 407212 409856
rect 407264 409844 407270 409896
rect 406286 408484 406292 408536
rect 406344 408524 406350 408536
rect 408126 408524 408132 408536
rect 406344 408496 408132 408524
rect 406344 408484 406350 408496
rect 408126 408484 408132 408496
rect 408184 408484 408190 408536
rect 350442 407192 350448 407244
rect 350500 407232 350506 407244
rect 375466 407232 375472 407244
rect 350500 407204 375472 407232
rect 350500 407192 350506 407204
rect 375466 407192 375472 407204
rect 375524 407192 375530 407244
rect 21450 407124 21456 407176
rect 21508 407164 21514 407176
rect 46566 407164 46572 407176
rect 21508 407136 46572 407164
rect 21508 407124 21514 407136
rect 46566 407124 46572 407136
rect 46624 407124 46630 407176
rect 370958 407124 370964 407176
rect 371016 407164 371022 407176
rect 407206 407164 407212 407176
rect 371016 407136 407212 407164
rect 371016 407124 371022 407136
rect 407206 407124 407212 407136
rect 407264 407124 407270 407176
rect 391382 405696 391388 405748
rect 391440 405736 391446 405748
rect 407206 405736 407212 405748
rect 391440 405708 407212 405736
rect 391440 405696 391446 405708
rect 407206 405696 407212 405708
rect 407264 405696 407270 405748
rect 402514 405628 402520 405680
rect 402572 405668 402578 405680
rect 407298 405668 407304 405680
rect 402572 405640 407304 405668
rect 402572 405628 402578 405640
rect 407298 405628 407304 405640
rect 407356 405628 407362 405680
rect 552934 405628 552940 405680
rect 552992 405668 552998 405680
rect 579062 405668 579068 405680
rect 552992 405640 579068 405668
rect 552992 405628 552998 405640
rect 579062 405628 579068 405640
rect 579120 405628 579126 405680
rect 350442 404404 350448 404456
rect 350500 404444 350506 404456
rect 358446 404444 358452 404456
rect 350500 404416 358452 404444
rect 350500 404404 350506 404416
rect 358446 404404 358452 404416
rect 358504 404404 358510 404456
rect 350074 404336 350080 404388
rect 350132 404376 350138 404388
rect 367370 404376 367376 404388
rect 350132 404348 367376 404376
rect 350132 404336 350138 404348
rect 367370 404336 367376 404348
rect 367428 404336 367434 404388
rect 552934 403044 552940 403096
rect 552992 403084 552998 403096
rect 562042 403084 562048 403096
rect 552992 403056 562048 403084
rect 552992 403044 552998 403056
rect 562042 403044 562048 403056
rect 562100 403044 562106 403096
rect 35158 402976 35164 403028
rect 35216 403016 35222 403028
rect 45922 403016 45928 403028
rect 35216 402988 45928 403016
rect 35216 402976 35222 402988
rect 45922 402976 45928 402988
rect 45980 402976 45986 403028
rect 552842 402976 552848 403028
rect 552900 403016 552906 403028
rect 575842 403016 575848 403028
rect 552900 402988 575848 403016
rect 552900 402976 552906 402988
rect 575842 402976 575848 402988
rect 575900 402976 575906 403028
rect 42426 401820 42432 401872
rect 42484 401860 42490 401872
rect 43254 401860 43260 401872
rect 42484 401832 43260 401860
rect 42484 401820 42490 401832
rect 43254 401820 43260 401832
rect 43312 401820 43318 401872
rect 391566 401616 391572 401668
rect 391624 401656 391630 401668
rect 407206 401656 407212 401668
rect 391624 401628 407212 401656
rect 391624 401616 391630 401628
rect 407206 401616 407212 401628
rect 407264 401616 407270 401668
rect 41966 400188 41972 400240
rect 42024 400228 42030 400240
rect 46106 400228 46112 400240
rect 42024 400200 46112 400228
rect 42024 400188 42030 400200
rect 46106 400188 46112 400200
rect 46164 400188 46170 400240
rect 350442 400188 350448 400240
rect 350500 400228 350506 400240
rect 365346 400228 365352 400240
rect 350500 400200 365352 400228
rect 350500 400188 350506 400200
rect 365346 400188 365352 400200
rect 365404 400188 365410 400240
rect 33778 398828 33784 398880
rect 33836 398868 33842 398880
rect 46566 398868 46572 398880
rect 33836 398840 46572 398868
rect 33836 398828 33842 398840
rect 46566 398828 46572 398840
rect 46624 398828 46630 398880
rect 350442 398828 350448 398880
rect 350500 398868 350506 398880
rect 359366 398868 359372 398880
rect 350500 398840 359372 398868
rect 350500 398828 350506 398840
rect 359366 398828 359372 398840
rect 359424 398828 359430 398880
rect 387426 397536 387432 397588
rect 387484 397576 387490 397588
rect 407206 397576 407212 397588
rect 387484 397548 407212 397576
rect 387484 397536 387490 397548
rect 407206 397536 407212 397548
rect 407264 397536 407270 397588
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 17310 397508 17316 397520
rect 3568 397480 17316 397508
rect 3568 397468 3574 397480
rect 17310 397468 17316 397480
rect 17368 397468 17374 397520
rect 350442 397468 350448 397520
rect 350500 397508 350506 397520
rect 396994 397508 397000 397520
rect 350500 397480 397000 397508
rect 350500 397468 350506 397480
rect 396994 397468 397000 397480
rect 397052 397468 397058 397520
rect 348510 397264 348516 397316
rect 348568 397304 348574 397316
rect 351178 397304 351184 397316
rect 348568 397276 351184 397304
rect 348568 397264 348574 397276
rect 351178 397264 351184 397276
rect 351236 397264 351242 397316
rect 42426 396448 42432 396500
rect 42484 396488 42490 396500
rect 46474 396488 46480 396500
rect 42484 396460 46480 396488
rect 42484 396448 42490 396460
rect 46474 396448 46480 396460
rect 46532 396448 46538 396500
rect 350442 396040 350448 396092
rect 350500 396080 350506 396092
rect 382826 396080 382832 396092
rect 350500 396052 382832 396080
rect 350500 396040 350506 396052
rect 382826 396040 382832 396052
rect 382884 396040 382890 396092
rect 39574 394748 39580 394800
rect 39632 394788 39638 394800
rect 45830 394788 45836 394800
rect 39632 394760 45836 394788
rect 39632 394748 39638 394760
rect 45830 394748 45836 394760
rect 45888 394748 45894 394800
rect 349798 394748 349804 394800
rect 349856 394788 349862 394800
rect 352006 394788 352012 394800
rect 349856 394760 352012 394788
rect 349856 394748 349862 394760
rect 352006 394748 352012 394760
rect 352064 394748 352070 394800
rect 22738 394680 22744 394732
rect 22796 394720 22802 394732
rect 46566 394720 46572 394732
rect 22796 394692 46572 394720
rect 22796 394680 22802 394692
rect 46566 394680 46572 394692
rect 46624 394680 46630 394732
rect 350074 394680 350080 394732
rect 350132 394720 350138 394732
rect 351454 394720 351460 394732
rect 350132 394692 351460 394720
rect 350132 394680 350138 394692
rect 351454 394680 351460 394692
rect 351512 394680 351518 394732
rect 388346 394680 388352 394732
rect 388404 394720 388410 394732
rect 407206 394720 407212 394732
rect 388404 394692 407212 394720
rect 388404 394680 388410 394692
rect 407206 394680 407212 394692
rect 407264 394680 407270 394732
rect 552934 394680 552940 394732
rect 552992 394720 552998 394732
rect 581822 394720 581828 394732
rect 552992 394692 581828 394720
rect 552992 394680 552998 394692
rect 581822 394680 581828 394692
rect 581880 394680 581886 394732
rect 350442 394612 350448 394664
rect 350500 394652 350506 394664
rect 399754 394652 399760 394664
rect 350500 394624 399760 394652
rect 350500 394612 350506 394624
rect 399754 394612 399760 394624
rect 399812 394612 399818 394664
rect 552014 393456 552020 393508
rect 552072 393496 552078 393508
rect 554314 393496 554320 393508
rect 552072 393468 554320 393496
rect 552072 393456 552078 393468
rect 554314 393456 554320 393468
rect 554372 393456 554378 393508
rect 39574 393320 39580 393372
rect 39632 393360 39638 393372
rect 46566 393360 46572 393372
rect 39632 393332 46572 393360
rect 39632 393320 39638 393332
rect 46566 393320 46572 393332
rect 46624 393320 46630 393372
rect 398374 393320 398380 393372
rect 398432 393360 398438 393372
rect 407206 393360 407212 393372
rect 398432 393332 407212 393360
rect 398432 393320 398438 393332
rect 407206 393320 407212 393332
rect 407264 393320 407270 393372
rect 37826 392028 37832 392080
rect 37884 392068 37890 392080
rect 46566 392068 46572 392080
rect 37884 392040 46572 392068
rect 37884 392028 37890 392040
rect 46566 392028 46572 392040
rect 46624 392028 46630 392080
rect 27338 391960 27344 392012
rect 27396 392000 27402 392012
rect 46474 392000 46480 392012
rect 27396 391972 46480 392000
rect 27396 391960 27402 391972
rect 46474 391960 46480 391972
rect 46532 391960 46538 392012
rect 350442 391960 350448 392012
rect 350500 392000 350506 392012
rect 356882 392000 356888 392012
rect 350500 391972 356888 392000
rect 350500 391960 350506 391972
rect 356882 391960 356888 391972
rect 356940 391960 356946 392012
rect 390094 390600 390100 390652
rect 390152 390640 390158 390652
rect 407206 390640 407212 390652
rect 390152 390612 407212 390640
rect 390152 390600 390158 390612
rect 407206 390600 407212 390612
rect 407264 390600 407270 390652
rect 552842 390600 552848 390652
rect 552900 390640 552906 390652
rect 560846 390640 560852 390652
rect 552900 390612 560852 390640
rect 552900 390600 552906 390612
rect 560846 390600 560852 390612
rect 560904 390600 560910 390652
rect 36262 390532 36268 390584
rect 36320 390572 36326 390584
rect 46474 390572 46480 390584
rect 36320 390544 46480 390572
rect 36320 390532 36326 390544
rect 46474 390532 46480 390544
rect 46532 390532 46538 390584
rect 350074 390532 350080 390584
rect 350132 390572 350138 390584
rect 352742 390572 352748 390584
rect 350132 390544 352748 390572
rect 350132 390532 350138 390544
rect 352742 390532 352748 390544
rect 352800 390532 352806 390584
rect 358354 390532 358360 390584
rect 358412 390572 358418 390584
rect 407298 390572 407304 390584
rect 358412 390544 407304 390572
rect 358412 390532 358418 390544
rect 407298 390532 407304 390544
rect 407356 390532 407362 390584
rect 552934 390532 552940 390584
rect 552992 390572 552998 390584
rect 568850 390572 568856 390584
rect 552992 390544 568856 390572
rect 552992 390532 552998 390544
rect 568850 390532 568856 390544
rect 568908 390532 568914 390584
rect 37182 390464 37188 390516
rect 37240 390504 37246 390516
rect 46566 390504 46572 390516
rect 37240 390476 46572 390504
rect 37240 390464 37246 390476
rect 46566 390464 46572 390476
rect 46624 390464 46630 390516
rect 350442 390464 350448 390516
rect 350500 390504 350506 390516
rect 395430 390504 395436 390516
rect 350500 390476 395436 390504
rect 350500 390464 350506 390476
rect 395430 390464 395436 390476
rect 395488 390464 395494 390516
rect 350074 390056 350080 390108
rect 350132 390096 350138 390108
rect 350350 390096 350356 390108
rect 350132 390068 350356 390096
rect 350132 390056 350138 390068
rect 350350 390056 350356 390068
rect 350408 390056 350414 390108
rect 348878 389376 348884 389428
rect 348936 389416 348942 389428
rect 349522 389416 349528 389428
rect 348936 389388 349528 389416
rect 348936 389376 348942 389388
rect 349522 389376 349528 389388
rect 349580 389376 349586 389428
rect 20530 389172 20536 389224
rect 20588 389212 20594 389224
rect 46566 389212 46572 389224
rect 20588 389184 46572 389212
rect 20588 389172 20594 389184
rect 46566 389172 46572 389184
rect 46624 389172 46630 389224
rect 350350 389172 350356 389224
rect 350408 389212 350414 389224
rect 401134 389212 401140 389224
rect 350408 389184 401140 389212
rect 350408 389172 350414 389184
rect 401134 389172 401140 389184
rect 401192 389172 401198 389224
rect 552290 389172 552296 389224
rect 552348 389212 552354 389224
rect 578786 389212 578792 389224
rect 552348 389184 578792 389212
rect 552348 389172 552354 389184
rect 578786 389172 578792 389184
rect 578844 389172 578850 389224
rect 348878 388424 348884 388476
rect 348936 388464 348942 388476
rect 357710 388464 357716 388476
rect 348936 388436 357716 388464
rect 348936 388424 348942 388436
rect 357710 388424 357716 388436
rect 357768 388424 357774 388476
rect 350442 387812 350448 387864
rect 350500 387852 350506 387864
rect 397086 387852 397092 387864
rect 350500 387824 397092 387852
rect 350500 387812 350506 387824
rect 397086 387812 397092 387824
rect 397144 387812 397150 387864
rect 552934 387812 552940 387864
rect 552992 387852 552998 387864
rect 579798 387852 579804 387864
rect 552992 387824 579804 387852
rect 552992 387812 552998 387824
rect 579798 387812 579804 387824
rect 579856 387812 579862 387864
rect 350350 387744 350356 387796
rect 350408 387784 350414 387796
rect 377858 387784 377864 387796
rect 350408 387756 377864 387784
rect 350408 387744 350414 387756
rect 377858 387744 377864 387756
rect 377916 387744 377922 387796
rect 38010 387064 38016 387116
rect 38068 387104 38074 387116
rect 45554 387104 45560 387116
rect 38068 387076 45560 387104
rect 38068 387064 38074 387076
rect 45554 387064 45560 387076
rect 45612 387064 45618 387116
rect 29914 386384 29920 386436
rect 29972 386424 29978 386436
rect 46566 386424 46572 386436
rect 29972 386396 46572 386424
rect 29972 386384 29978 386396
rect 46566 386384 46572 386396
rect 46624 386384 46630 386436
rect 552934 386384 552940 386436
rect 552992 386424 552998 386436
rect 560938 386424 560944 386436
rect 552992 386396 560944 386424
rect 552992 386384 552998 386396
rect 560938 386384 560944 386396
rect 560996 386384 561002 386436
rect 36446 386316 36452 386368
rect 36504 386356 36510 386368
rect 46474 386356 46480 386368
rect 36504 386328 46480 386356
rect 36504 386316 36510 386328
rect 46474 386316 46480 386328
rect 46532 386316 46538 386368
rect 391474 386316 391480 386368
rect 391532 386356 391538 386368
rect 407206 386356 407212 386368
rect 391532 386328 407212 386356
rect 391532 386316 391538 386328
rect 407206 386316 407212 386328
rect 407264 386316 407270 386368
rect 38010 385024 38016 385076
rect 38068 385064 38074 385076
rect 46566 385064 46572 385076
rect 38068 385036 46572 385064
rect 38068 385024 38074 385036
rect 46566 385024 46572 385036
rect 46624 385024 46630 385076
rect 552934 385024 552940 385076
rect 552992 385064 552998 385076
rect 563238 385064 563244 385076
rect 552992 385036 563244 385064
rect 552992 385024 552998 385036
rect 563238 385024 563244 385036
rect 563296 385024 563302 385076
rect 350074 384956 350080 385008
rect 350132 384996 350138 385008
rect 351178 384996 351184 385008
rect 350132 384968 351184 384996
rect 350132 384956 350138 384968
rect 351178 384956 351184 384968
rect 351236 384956 351242 385008
rect 36446 384276 36452 384328
rect 36504 384316 36510 384328
rect 45646 384316 45652 384328
rect 36504 384288 45652 384316
rect 36504 384276 36510 384288
rect 45646 384276 45652 384288
rect 45704 384276 45710 384328
rect 400674 383664 400680 383716
rect 400732 383704 400738 383716
rect 407206 383704 407212 383716
rect 400732 383676 407212 383704
rect 400732 383664 400738 383676
rect 407206 383664 407212 383676
rect 407264 383664 407270 383716
rect 29638 382236 29644 382288
rect 29696 382276 29702 382288
rect 46566 382276 46572 382288
rect 29696 382248 46572 382276
rect 29696 382236 29702 382248
rect 46566 382236 46572 382248
rect 46624 382236 46630 382288
rect 350442 382236 350448 382288
rect 350500 382276 350506 382288
rect 394326 382276 394332 382288
rect 350500 382248 394332 382276
rect 350500 382236 350506 382248
rect 394326 382236 394332 382248
rect 394384 382236 394390 382288
rect 552934 381080 552940 381132
rect 552992 381120 552998 381132
rect 559742 381120 559748 381132
rect 552992 381092 559748 381120
rect 552992 381080 552998 381092
rect 559742 381080 559748 381092
rect 559800 381080 559806 381132
rect 380066 381012 380072 381064
rect 380124 381052 380130 381064
rect 407206 381052 407212 381064
rect 380124 381024 407212 381052
rect 380124 381012 380130 381024
rect 407206 381012 407212 381024
rect 407264 381012 407270 381064
rect 350350 380944 350356 380996
rect 350408 380984 350414 380996
rect 387794 380984 387800 380996
rect 350408 380956 387800 380984
rect 350408 380944 350414 380956
rect 387794 380944 387800 380956
rect 387852 380944 387858 380996
rect 350442 380876 350448 380928
rect 350500 380916 350506 380928
rect 392946 380916 392952 380928
rect 350500 380888 392952 380916
rect 350500 380876 350506 380888
rect 392946 380876 392952 380888
rect 393004 380876 393010 380928
rect 394418 380128 394424 380180
rect 394476 380168 394482 380180
rect 407850 380168 407856 380180
rect 394476 380140 407856 380168
rect 394476 380128 394482 380140
rect 407850 380128 407856 380140
rect 407908 380128 407914 380180
rect 32490 379516 32496 379568
rect 32548 379556 32554 379568
rect 46566 379556 46572 379568
rect 32548 379528 46572 379556
rect 32548 379516 32554 379528
rect 46566 379516 46572 379528
rect 46624 379516 46630 379568
rect 29546 378156 29552 378208
rect 29604 378196 29610 378208
rect 46566 378196 46572 378208
rect 29604 378168 46572 378196
rect 29604 378156 29610 378168
rect 46566 378156 46572 378168
rect 46624 378156 46630 378208
rect 377858 378156 377864 378208
rect 377916 378196 377922 378208
rect 407206 378196 407212 378208
rect 377916 378168 407212 378196
rect 377916 378156 377922 378168
rect 407206 378156 407212 378168
rect 407264 378156 407270 378208
rect 574922 378156 574928 378208
rect 574980 378196 574986 378208
rect 580166 378196 580172 378208
rect 574980 378168 580172 378196
rect 574980 378156 574986 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 350442 376728 350448 376780
rect 350500 376768 350506 376780
rect 375006 376768 375012 376780
rect 350500 376740 375012 376768
rect 350500 376728 350506 376740
rect 375006 376728 375012 376740
rect 375064 376728 375070 376780
rect 552934 376728 552940 376780
rect 552992 376768 552998 376780
rect 583110 376768 583116 376780
rect 552992 376740 583116 376768
rect 552992 376728 552998 376740
rect 583110 376728 583116 376740
rect 583168 376728 583174 376780
rect 350350 375368 350356 375420
rect 350408 375408 350414 375420
rect 395430 375408 395436 375420
rect 350408 375380 395436 375408
rect 350408 375368 350414 375380
rect 395430 375368 395436 375380
rect 395488 375368 395494 375420
rect 350442 375300 350448 375352
rect 350500 375340 350506 375352
rect 375098 375340 375104 375352
rect 350500 375312 375104 375340
rect 350500 375300 350506 375312
rect 375098 375300 375104 375312
rect 375156 375300 375162 375352
rect 43438 374688 43444 374740
rect 43496 374728 43502 374740
rect 47210 374728 47216 374740
rect 43496 374700 47216 374728
rect 43496 374688 43502 374700
rect 47210 374688 47216 374700
rect 47268 374688 47274 374740
rect 26878 374008 26884 374060
rect 26936 374048 26942 374060
rect 46474 374048 46480 374060
rect 26936 374020 46480 374048
rect 26936 374008 26942 374020
rect 46474 374008 46480 374020
rect 46532 374008 46538 374060
rect 395706 374008 395712 374060
rect 395764 374048 395770 374060
rect 407206 374048 407212 374060
rect 395764 374020 407212 374048
rect 395764 374008 395770 374020
rect 407206 374008 407212 374020
rect 407264 374008 407270 374060
rect 28350 372648 28356 372700
rect 28408 372688 28414 372700
rect 46106 372688 46112 372700
rect 28408 372660 46112 372688
rect 28408 372648 28414 372660
rect 46106 372648 46112 372660
rect 46164 372648 46170 372700
rect 552934 372648 552940 372700
rect 552992 372688 552998 372700
rect 556522 372688 556528 372700
rect 552992 372660 556528 372688
rect 552992 372648 552998 372660
rect 556522 372648 556528 372660
rect 556580 372648 556586 372700
rect 26786 372580 26792 372632
rect 26844 372620 26850 372632
rect 46474 372620 46480 372632
rect 26844 372592 46480 372620
rect 26844 372580 26850 372592
rect 46474 372580 46480 372592
rect 46532 372580 46538 372632
rect 350442 372580 350448 372632
rect 350500 372620 350506 372632
rect 379146 372620 379152 372632
rect 350500 372592 379152 372620
rect 350500 372580 350506 372592
rect 379146 372580 379152 372592
rect 379204 372580 379210 372632
rect 399938 372580 399944 372632
rect 399996 372620 400002 372632
rect 407206 372620 407212 372632
rect 399996 372592 407212 372620
rect 399996 372580 400002 372592
rect 407206 372580 407212 372592
rect 407264 372580 407270 372632
rect 30742 371220 30748 371272
rect 30800 371260 30806 371272
rect 46474 371260 46480 371272
rect 30800 371232 46480 371260
rect 30800 371220 30806 371232
rect 46474 371220 46480 371232
rect 46532 371220 46538 371272
rect 350442 371220 350448 371272
rect 350500 371260 350506 371272
rect 375190 371260 375196 371272
rect 350500 371232 375196 371260
rect 350500 371220 350506 371232
rect 375190 371220 375196 371232
rect 375248 371220 375254 371272
rect 374546 371152 374552 371204
rect 374604 371192 374610 371204
rect 407206 371192 407212 371204
rect 374604 371164 407212 371192
rect 374604 371152 374610 371164
rect 407206 371152 407212 371164
rect 407264 371152 407270 371204
rect 41874 369860 41880 369912
rect 41932 369900 41938 369912
rect 43438 369900 43444 369912
rect 41932 369872 43444 369900
rect 41932 369860 41938 369872
rect 43438 369860 43444 369872
rect 43496 369860 43502 369912
rect 552934 369860 552940 369912
rect 552992 369900 552998 369912
rect 562134 369900 562140 369912
rect 552992 369872 562140 369900
rect 552992 369860 552998 369872
rect 562134 369860 562140 369872
rect 562192 369860 562198 369912
rect 552934 368568 552940 368620
rect 552992 368608 552998 368620
rect 557902 368608 557908 368620
rect 552992 368580 557908 368608
rect 552992 368568 552998 368580
rect 557902 368568 557908 368580
rect 557960 368568 557966 368620
rect 29730 368500 29736 368552
rect 29788 368540 29794 368552
rect 46474 368540 46480 368552
rect 29788 368512 46480 368540
rect 29788 368500 29794 368512
rect 46474 368500 46480 368512
rect 46532 368500 46538 368552
rect 400766 368500 400772 368552
rect 400824 368540 400830 368552
rect 407206 368540 407212 368552
rect 400824 368512 407212 368540
rect 400824 368500 400830 368512
rect 407206 368500 407212 368512
rect 407264 368500 407270 368552
rect 552842 368500 552848 368552
rect 552900 368540 552906 368552
rect 571794 368540 571800 368552
rect 552900 368512 571800 368540
rect 552900 368500 552906 368512
rect 571794 368500 571800 368512
rect 571852 368500 571858 368552
rect 552014 368092 552020 368144
rect 552072 368132 552078 368144
rect 553762 368132 553768 368144
rect 552072 368104 553768 368132
rect 552072 368092 552078 368104
rect 553762 368092 553768 368104
rect 553820 368092 553826 368144
rect 29822 367072 29828 367124
rect 29880 367112 29886 367124
rect 46382 367112 46388 367124
rect 29880 367084 46388 367112
rect 29880 367072 29886 367084
rect 46382 367072 46388 367084
rect 46440 367072 46446 367124
rect 31386 367004 31392 367056
rect 31444 367044 31450 367056
rect 46474 367044 46480 367056
rect 31444 367016 46480 367044
rect 31444 367004 31450 367016
rect 46474 367004 46480 367016
rect 46532 367004 46538 367056
rect 552934 365780 552940 365832
rect 552992 365820 552998 365832
rect 566366 365820 566372 365832
rect 552992 365792 566372 365820
rect 552992 365780 552998 365792
rect 566366 365780 566372 365792
rect 566424 365780 566430 365832
rect 552842 365712 552848 365764
rect 552900 365752 552906 365764
rect 578418 365752 578424 365764
rect 552900 365724 578424 365752
rect 552900 365712 552906 365724
rect 578418 365712 578424 365724
rect 578476 365712 578482 365764
rect 350442 365644 350448 365696
rect 350500 365684 350506 365696
rect 353846 365684 353852 365696
rect 350500 365656 353852 365684
rect 350500 365644 350506 365656
rect 353846 365644 353852 365656
rect 353904 365644 353910 365696
rect 350442 364352 350448 364404
rect 350500 364392 350506 364404
rect 383654 364392 383660 364404
rect 350500 364364 383660 364392
rect 350500 364352 350506 364364
rect 383654 364352 383660 364364
rect 383712 364352 383718 364404
rect 28718 362924 28724 362976
rect 28776 362964 28782 362976
rect 46474 362964 46480 362976
rect 28776 362936 46480 362964
rect 28776 362924 28782 362936
rect 46474 362924 46480 362936
rect 46532 362924 46538 362976
rect 552842 362924 552848 362976
rect 552900 362964 552906 362976
rect 555142 362964 555148 362976
rect 552900 362936 555148 362964
rect 552900 362924 552906 362936
rect 555142 362924 555148 362936
rect 555200 362924 555206 362976
rect 366726 361496 366732 361548
rect 366784 361536 366790 361548
rect 407206 361536 407212 361548
rect 366784 361508 407212 361536
rect 366784 361496 366790 361508
rect 407206 361496 407212 361508
rect 407264 361496 407270 361548
rect 552198 360408 552204 360460
rect 552256 360448 552262 360460
rect 555142 360448 555148 360460
rect 552256 360420 555148 360448
rect 552256 360408 552262 360420
rect 555142 360408 555148 360420
rect 555200 360408 555206 360460
rect 364058 360204 364064 360256
rect 364116 360244 364122 360256
rect 407206 360244 407212 360256
rect 364116 360216 407212 360244
rect 364116 360204 364122 360216
rect 407206 360204 407212 360216
rect 407264 360204 407270 360256
rect 552934 360204 552940 360256
rect 552992 360244 552998 360256
rect 571978 360244 571984 360256
rect 552992 360216 571984 360244
rect 552992 360204 552998 360216
rect 571978 360204 571984 360216
rect 572036 360204 572042 360256
rect 32674 358708 32680 358760
rect 32732 358748 32738 358760
rect 46474 358748 46480 358760
rect 32732 358720 46480 358748
rect 32732 358708 32738 358720
rect 46474 358708 46480 358720
rect 46532 358708 46538 358760
rect 552934 358708 552940 358760
rect 552992 358748 552998 358760
rect 574922 358748 574928 358760
rect 552992 358720 574928 358748
rect 552992 358708 552998 358720
rect 574922 358708 574928 358720
rect 574980 358708 574986 358760
rect 348786 358504 348792 358556
rect 348844 358544 348850 358556
rect 352466 358544 352472 358556
rect 348844 358516 352472 358544
rect 348844 358504 348850 358516
rect 352466 358504 352472 358516
rect 352524 358504 352530 358556
rect 350442 357960 350448 358012
rect 350500 358000 350506 358012
rect 355410 358000 355416 358012
rect 350500 357972 355416 358000
rect 350500 357960 350506 357972
rect 355410 357960 355416 357972
rect 355468 357960 355474 358012
rect 552658 357620 552664 357672
rect 552716 357660 552722 357672
rect 556798 357660 556804 357672
rect 552716 357632 556804 357660
rect 552716 357620 552722 357632
rect 556798 357620 556804 357632
rect 556856 357620 556862 357672
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 24118 357456 24124 357468
rect 3200 357428 24124 357456
rect 3200 357416 3206 357428
rect 24118 357416 24124 357428
rect 24176 357416 24182 357468
rect 386966 357416 386972 357468
rect 387024 357456 387030 357468
rect 407206 357456 407212 357468
rect 387024 357428 407212 357456
rect 387024 357416 387030 357428
rect 407206 357416 407212 357428
rect 407264 357416 407270 357468
rect 349982 356056 349988 356108
rect 350040 356096 350046 356108
rect 352466 356096 352472 356108
rect 350040 356068 352472 356096
rect 350040 356056 350046 356068
rect 352466 356056 352472 356068
rect 352524 356056 352530 356108
rect 395522 356056 395528 356108
rect 395580 356096 395586 356108
rect 407206 356096 407212 356108
rect 395580 356068 407212 356096
rect 395580 356056 395586 356068
rect 407206 356056 407212 356068
rect 407264 356056 407270 356108
rect 350442 355988 350448 356040
rect 350500 356028 350506 356040
rect 388714 356028 388720 356040
rect 350500 356000 388720 356028
rect 350500 355988 350506 356000
rect 388714 355988 388720 356000
rect 388772 355988 388778 356040
rect 25498 354696 25504 354748
rect 25556 354736 25562 354748
rect 46474 354736 46480 354748
rect 25556 354708 46480 354736
rect 25556 354696 25562 354708
rect 46474 354696 46480 354708
rect 46532 354696 46538 354748
rect 350442 354696 350448 354748
rect 350500 354736 350506 354748
rect 375098 354736 375104 354748
rect 350500 354708 375104 354736
rect 350500 354696 350506 354708
rect 375098 354696 375104 354708
rect 375156 354696 375162 354748
rect 552934 354696 552940 354748
rect 552992 354736 552998 354748
rect 571702 354736 571708 354748
rect 552992 354708 571708 354736
rect 552992 354696 552998 354708
rect 571702 354696 571708 354708
rect 571760 354696 571766 354748
rect 552934 354424 552940 354476
rect 552992 354464 552998 354476
rect 553118 354464 553124 354476
rect 552992 354436 553124 354464
rect 552992 354424 552998 354436
rect 553118 354424 553124 354436
rect 553176 354424 553182 354476
rect 553118 353744 553124 353796
rect 553176 353784 553182 353796
rect 558178 353784 558184 353796
rect 553176 353756 558184 353784
rect 553176 353744 553182 353756
rect 558178 353744 558184 353756
rect 558236 353744 558242 353796
rect 378042 353268 378048 353320
rect 378100 353308 378106 353320
rect 407206 353308 407212 353320
rect 378100 353280 407212 353308
rect 378100 353268 378106 353280
rect 407206 353268 407212 353280
rect 407264 353268 407270 353320
rect 553118 353268 553124 353320
rect 553176 353308 553182 353320
rect 574370 353308 574376 353320
rect 553176 353280 574376 353308
rect 553176 353268 553182 353280
rect 574370 353268 574376 353280
rect 574428 353268 574434 353320
rect 35066 353200 35072 353252
rect 35124 353240 35130 353252
rect 46474 353240 46480 353252
rect 35124 353212 46480 353240
rect 35124 353200 35130 353212
rect 46474 353200 46480 353212
rect 46532 353200 46538 353252
rect 402514 351976 402520 352028
rect 402572 352016 402578 352028
rect 407206 352016 407212 352028
rect 402572 351988 407212 352016
rect 402572 351976 402578 351988
rect 407206 351976 407212 351988
rect 407264 351976 407270 352028
rect 350350 351908 350356 351960
rect 350408 351948 350414 351960
rect 352374 351948 352380 351960
rect 350408 351920 352380 351948
rect 350408 351908 350414 351920
rect 352374 351908 352380 351920
rect 352432 351908 352438 351960
rect 379330 351908 379336 351960
rect 379388 351948 379394 351960
rect 407298 351948 407304 351960
rect 379388 351920 407304 351948
rect 379388 351908 379394 351920
rect 407298 351908 407304 351920
rect 407356 351908 407362 351960
rect 35066 351160 35072 351212
rect 35124 351200 35130 351212
rect 39298 351200 39304 351212
rect 35124 351172 39304 351200
rect 35124 351160 35130 351172
rect 39298 351160 39304 351172
rect 39356 351160 39362 351212
rect 552014 350888 552020 350940
rect 552072 350928 552078 350940
rect 554038 350928 554044 350940
rect 552072 350900 554044 350928
rect 552072 350888 552078 350900
rect 554038 350888 554044 350900
rect 554096 350888 554102 350940
rect 350166 350616 350172 350668
rect 350224 350656 350230 350668
rect 352374 350656 352380 350668
rect 350224 350628 352380 350656
rect 350224 350616 350230 350628
rect 352374 350616 352380 350628
rect 352432 350616 352438 350668
rect 350442 350548 350448 350600
rect 350500 350588 350506 350600
rect 362494 350588 362500 350600
rect 350500 350560 362500 350588
rect 350500 350548 350506 350560
rect 362494 350548 362500 350560
rect 362552 350548 362558 350600
rect 391474 350548 391480 350600
rect 391532 350588 391538 350600
rect 407206 350588 407212 350600
rect 391532 350560 407212 350588
rect 391532 350548 391538 350560
rect 407206 350548 407212 350560
rect 407264 350548 407270 350600
rect 552290 350548 552296 350600
rect 552348 350588 552354 350600
rect 583202 350588 583208 350600
rect 552348 350560 583208 350588
rect 552348 350548 552354 350560
rect 583202 350548 583208 350560
rect 583260 350548 583266 350600
rect 348970 349800 348976 349852
rect 349028 349840 349034 349852
rect 349798 349840 349804 349852
rect 349028 349812 349804 349840
rect 349028 349800 349034 349812
rect 349798 349800 349804 349812
rect 349856 349800 349862 349852
rect 350442 349188 350448 349240
rect 350500 349228 350506 349240
rect 368290 349228 368296 349240
rect 350500 349200 368296 349228
rect 350500 349188 350506 349200
rect 368290 349188 368296 349200
rect 368348 349188 368354 349240
rect 379238 349188 379244 349240
rect 379296 349228 379302 349240
rect 407206 349228 407212 349240
rect 379296 349200 407212 349228
rect 379296 349188 379302 349200
rect 407206 349188 407212 349200
rect 407264 349188 407270 349240
rect 17678 349120 17684 349172
rect 17736 349160 17742 349172
rect 46474 349160 46480 349172
rect 17736 349132 46480 349160
rect 17736 349120 17742 349132
rect 46474 349120 46480 349132
rect 46532 349120 46538 349172
rect 350350 349120 350356 349172
rect 350408 349160 350414 349172
rect 388254 349160 388260 349172
rect 350408 349132 388260 349160
rect 350408 349120 350414 349132
rect 388254 349120 388260 349132
rect 388312 349120 388318 349172
rect 553118 349120 553124 349172
rect 553176 349160 553182 349172
rect 583294 349160 583300 349172
rect 553176 349132 583300 349160
rect 553176 349120 553182 349132
rect 583294 349120 583300 349132
rect 583352 349120 583358 349172
rect 36354 348372 36360 348424
rect 36412 348412 36418 348424
rect 47210 348412 47216 348424
rect 36412 348384 47216 348412
rect 36412 348372 36418 348384
rect 47210 348372 47216 348384
rect 47268 348372 47274 348424
rect 553118 346468 553124 346520
rect 553176 346508 553182 346520
rect 573174 346508 573180 346520
rect 553176 346480 573180 346508
rect 553176 346468 553182 346480
rect 573174 346468 573180 346480
rect 573232 346468 573238 346520
rect 25406 346400 25412 346452
rect 25464 346440 25470 346452
rect 46474 346440 46480 346452
rect 25464 346412 46480 346440
rect 25464 346400 25470 346412
rect 46474 346400 46480 346412
rect 46532 346400 46538 346452
rect 552658 346400 552664 346452
rect 552716 346440 552722 346452
rect 578694 346440 578700 346452
rect 552716 346412 578700 346440
rect 552716 346400 552722 346412
rect 578694 346400 578700 346412
rect 578752 346400 578758 346452
rect 402790 346332 402796 346384
rect 402848 346372 402854 346384
rect 407206 346372 407212 346384
rect 402848 346344 407212 346372
rect 402848 346332 402854 346344
rect 407206 346332 407212 346344
rect 407264 346332 407270 346384
rect 350350 345448 350356 345500
rect 350408 345488 350414 345500
rect 353846 345488 353852 345500
rect 350408 345460 353852 345488
rect 350408 345448 350414 345460
rect 353846 345448 353852 345460
rect 353904 345448 353910 345500
rect 22646 345108 22652 345160
rect 22704 345148 22710 345160
rect 45922 345148 45928 345160
rect 22704 345120 45928 345148
rect 22704 345108 22710 345120
rect 45922 345108 45928 345120
rect 45980 345108 45986 345160
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 29454 345080 29460 345092
rect 3384 345052 29460 345080
rect 3384 345040 3390 345052
rect 29454 345040 29460 345052
rect 29512 345040 29518 345092
rect 365438 344972 365444 345024
rect 365496 345012 365502 345024
rect 407206 345012 407212 345024
rect 365496 344984 407212 345012
rect 365496 344972 365502 344984
rect 407206 344972 407212 344984
rect 407264 344972 407270 345024
rect 350350 343680 350356 343732
rect 350408 343720 350414 343732
rect 381446 343720 381452 343732
rect 350408 343692 381452 343720
rect 350408 343680 350414 343692
rect 381446 343680 381452 343692
rect 381504 343680 381510 343732
rect 350166 343612 350172 343664
rect 350224 343652 350230 343664
rect 385494 343652 385500 343664
rect 350224 343624 385500 343652
rect 350224 343612 350230 343624
rect 385494 343612 385500 343624
rect 385552 343612 385558 343664
rect 350350 343544 350356 343596
rect 350408 343584 350414 343596
rect 363138 343584 363144 343596
rect 350408 343556 363144 343584
rect 350408 343544 350414 343556
rect 363138 343544 363144 343556
rect 363196 343544 363202 343596
rect 552014 342796 552020 342848
rect 552072 342836 552078 342848
rect 553670 342836 553676 342848
rect 552072 342808 553676 342836
rect 552072 342796 552078 342808
rect 553670 342796 553676 342808
rect 553728 342796 553734 342848
rect 395246 342252 395252 342304
rect 395304 342292 395310 342304
rect 407206 342292 407212 342304
rect 395304 342264 407212 342292
rect 395304 342252 395310 342264
rect 407206 342252 407212 342264
rect 407264 342252 407270 342304
rect 553118 342252 553124 342304
rect 553176 342292 553182 342304
rect 567470 342292 567476 342304
rect 553176 342264 567476 342292
rect 553176 342252 553182 342264
rect 567470 342252 567476 342264
rect 567528 342252 567534 342304
rect 45186 342184 45192 342236
rect 45244 342224 45250 342236
rect 46290 342224 46296 342236
rect 45244 342196 46296 342224
rect 45244 342184 45250 342196
rect 46290 342184 46296 342196
rect 46348 342184 46354 342236
rect 376662 339464 376668 339516
rect 376720 339504 376726 339516
rect 407206 339504 407212 339516
rect 376720 339476 407212 339504
rect 376720 339464 376726 339476
rect 407206 339464 407212 339476
rect 407264 339464 407270 339516
rect 350350 338104 350356 338156
rect 350408 338144 350414 338156
rect 366082 338144 366088 338156
rect 350408 338116 366088 338144
rect 350408 338104 350414 338116
rect 366082 338104 366088 338116
rect 366140 338104 366146 338156
rect 553118 338104 553124 338156
rect 553176 338144 553182 338156
rect 573450 338144 573456 338156
rect 553176 338116 573456 338144
rect 553176 338104 553182 338116
rect 573450 338104 573456 338116
rect 573508 338104 573514 338156
rect 28258 336744 28264 336796
rect 28316 336784 28322 336796
rect 46474 336784 46480 336796
rect 28316 336756 46480 336784
rect 28316 336744 28322 336756
rect 46474 336744 46480 336756
rect 46532 336744 46538 336796
rect 382182 336676 382188 336728
rect 382240 336716 382246 336728
rect 407206 336716 407212 336728
rect 382240 336688 407212 336716
rect 382240 336676 382246 336688
rect 407206 336676 407212 336688
rect 407264 336676 407270 336728
rect 552934 335316 552940 335368
rect 552992 335356 552998 335368
rect 566458 335356 566464 335368
rect 552992 335328 566464 335356
rect 552992 335316 552998 335328
rect 566458 335316 566464 335328
rect 566516 335316 566522 335368
rect 553118 335248 553124 335300
rect 553176 335288 553182 335300
rect 564710 335288 564716 335300
rect 553176 335260 564716 335288
rect 553176 335248 553182 335260
rect 564710 335248 564716 335260
rect 564768 335248 564774 335300
rect 350350 333956 350356 334008
rect 350408 333996 350414 334008
rect 382182 333996 382188 334008
rect 350408 333968 382188 333996
rect 350408 333956 350414 333968
rect 382182 333956 382188 333968
rect 382240 333956 382246 334008
rect 553118 333956 553124 334008
rect 553176 333996 553182 334008
rect 580074 333996 580080 334008
rect 553176 333968 580080 333996
rect 553176 333956 553182 333968
rect 580074 333956 580080 333968
rect 580132 333956 580138 334008
rect 350350 332596 350356 332648
rect 350408 332636 350414 332648
rect 366818 332636 366824 332648
rect 350408 332608 366824 332636
rect 350408 332596 350414 332608
rect 366818 332596 366824 332608
rect 366876 332596 366882 332648
rect 39298 332528 39304 332580
rect 39356 332568 39362 332580
rect 45646 332568 45652 332580
rect 39356 332540 45652 332568
rect 39356 332528 39362 332540
rect 45646 332528 45652 332540
rect 45704 332528 45710 332580
rect 376570 331236 376576 331288
rect 376628 331276 376634 331288
rect 407206 331276 407212 331288
rect 376628 331248 407212 331276
rect 376628 331236 376634 331248
rect 407206 331236 407212 331248
rect 407264 331236 407270 331288
rect 36630 331168 36636 331220
rect 36688 331208 36694 331220
rect 46842 331208 46848 331220
rect 36688 331180 46848 331208
rect 36688 331168 36694 331180
rect 46842 331168 46848 331180
rect 46900 331168 46906 331220
rect 350350 329808 350356 329860
rect 350408 329848 350414 329860
rect 363138 329848 363144 329860
rect 350408 329820 363144 329848
rect 350408 329808 350414 329820
rect 363138 329808 363144 329820
rect 363196 329808 363202 329860
rect 365530 329808 365536 329860
rect 365588 329848 365594 329860
rect 407206 329848 407212 329860
rect 365588 329820 407212 329848
rect 365588 329808 365594 329820
rect 407206 329808 407212 329820
rect 407264 329808 407270 329860
rect 28166 328448 28172 328500
rect 28224 328488 28230 328500
rect 45830 328488 45836 328500
rect 28224 328460 45836 328488
rect 28224 328448 28230 328460
rect 45830 328448 45836 328460
rect 45888 328448 45894 328500
rect 350350 328448 350356 328500
rect 350408 328488 350414 328500
rect 369394 328488 369400 328500
rect 350408 328460 369400 328488
rect 350408 328448 350414 328460
rect 369394 328448 369400 328460
rect 369452 328448 369458 328500
rect 381354 328448 381360 328500
rect 381412 328488 381418 328500
rect 407206 328488 407212 328500
rect 381412 328460 407212 328488
rect 381412 328448 381418 328460
rect 407206 328448 407212 328460
rect 407264 328448 407270 328500
rect 553118 327088 553124 327140
rect 553176 327128 553182 327140
rect 577590 327128 577596 327140
rect 553176 327100 577596 327128
rect 553176 327088 553182 327100
rect 577590 327088 577596 327100
rect 577648 327088 577654 327140
rect 553118 325728 553124 325780
rect 553176 325768 553182 325780
rect 569126 325768 569132 325780
rect 553176 325740 569132 325768
rect 553176 325728 553182 325740
rect 569126 325728 569132 325740
rect 569184 325728 569190 325780
rect 43714 325660 43720 325712
rect 43772 325700 43778 325712
rect 45738 325700 45744 325712
rect 43772 325672 45744 325700
rect 43772 325660 43778 325672
rect 45738 325660 45744 325672
rect 45796 325660 45802 325712
rect 350350 325660 350356 325712
rect 350408 325700 350414 325712
rect 363230 325700 363236 325712
rect 350408 325672 363236 325700
rect 350408 325660 350414 325672
rect 363230 325660 363236 325672
rect 363288 325660 363294 325712
rect 552934 325660 552940 325712
rect 552992 325700 552998 325712
rect 581638 325700 581644 325712
rect 552992 325672 581644 325700
rect 552992 325660 552998 325672
rect 581638 325660 581644 325672
rect 581696 325660 581702 325712
rect 31294 325592 31300 325644
rect 31352 325632 31358 325644
rect 46842 325632 46848 325644
rect 31352 325604 46848 325632
rect 31352 325592 31358 325604
rect 46842 325592 46848 325604
rect 46900 325592 46906 325644
rect 376478 325592 376484 325644
rect 376536 325632 376542 325644
rect 407206 325632 407212 325644
rect 376536 325604 407212 325632
rect 376536 325592 376542 325604
rect 407206 325592 407212 325604
rect 407264 325592 407270 325644
rect 572070 325592 572076 325644
rect 572128 325632 572134 325644
rect 580166 325632 580172 325644
rect 572128 325604 580172 325632
rect 572128 325592 572134 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 552934 323280 552940 323332
rect 552992 323320 552998 323332
rect 556706 323320 556712 323332
rect 552992 323292 556712 323320
rect 552992 323280 552998 323292
rect 556706 323280 556712 323292
rect 556764 323280 556770 323332
rect 407114 323144 407120 323196
rect 407172 323184 407178 323196
rect 407390 323184 407396 323196
rect 407172 323156 407396 323184
rect 407172 323144 407178 323156
rect 407390 323144 407396 323156
rect 407448 323144 407454 323196
rect 402146 323008 402152 323060
rect 402204 323048 402210 323060
rect 407206 323048 407212 323060
rect 402204 323020 407212 323048
rect 402204 323008 402210 323020
rect 407206 323008 407212 323020
rect 407264 323008 407270 323060
rect 39206 322940 39212 322992
rect 39264 322980 39270 322992
rect 46842 322980 46848 322992
rect 39264 322952 46848 322980
rect 39264 322940 39270 322952
rect 46842 322940 46848 322952
rect 46900 322940 46906 322992
rect 377306 322940 377312 322992
rect 377364 322980 377370 322992
rect 407114 322980 407120 322992
rect 377364 322952 407120 322980
rect 377364 322940 377370 322952
rect 407114 322940 407120 322952
rect 407172 322940 407178 322992
rect 363230 322872 363236 322924
rect 363288 322912 363294 322924
rect 407206 322912 407212 322924
rect 363288 322884 407212 322912
rect 363288 322872 363294 322884
rect 407206 322872 407212 322884
rect 407264 322872 407270 322924
rect 401042 322804 401048 322856
rect 401100 322844 401106 322856
rect 407114 322844 407120 322856
rect 401100 322816 407120 322844
rect 401100 322804 401106 322816
rect 407114 322804 407120 322816
rect 407172 322804 407178 322856
rect 552014 321784 552020 321836
rect 552072 321824 552078 321836
rect 553670 321824 553676 321836
rect 552072 321796 553676 321824
rect 552072 321784 552078 321796
rect 553670 321784 553676 321796
rect 553728 321784 553734 321836
rect 43346 321580 43352 321632
rect 43404 321620 43410 321632
rect 46842 321620 46848 321632
rect 43404 321592 46848 321620
rect 43404 321580 43410 321592
rect 46842 321580 46848 321592
rect 46900 321580 46906 321632
rect 350350 321580 350356 321632
rect 350408 321620 350414 321632
rect 378686 321620 378692 321632
rect 350408 321592 378692 321620
rect 350408 321580 350414 321592
rect 378686 321580 378692 321592
rect 378744 321580 378750 321632
rect 407850 320832 407856 320884
rect 407908 320872 407914 320884
rect 408402 320872 408408 320884
rect 407908 320844 408408 320872
rect 407908 320832 407914 320844
rect 408402 320832 408408 320844
rect 408460 320832 408466 320884
rect 28074 320152 28080 320204
rect 28132 320192 28138 320204
rect 46842 320192 46848 320204
rect 28132 320164 46848 320192
rect 28132 320152 28138 320164
rect 46842 320152 46848 320164
rect 46900 320152 46906 320204
rect 350350 320152 350356 320204
rect 350408 320192 350414 320204
rect 371142 320192 371148 320204
rect 350408 320164 371148 320192
rect 350408 320152 350414 320164
rect 371142 320152 371148 320164
rect 371200 320152 371206 320204
rect 395798 320152 395804 320204
rect 395856 320192 395862 320204
rect 407114 320192 407120 320204
rect 395856 320164 407120 320192
rect 395856 320152 395862 320164
rect 407114 320152 407120 320164
rect 407172 320152 407178 320204
rect 350166 320084 350172 320136
rect 350224 320124 350230 320136
rect 383378 320124 383384 320136
rect 350224 320096 383384 320124
rect 350224 320084 350230 320096
rect 383378 320084 383384 320096
rect 383436 320084 383442 320136
rect 43714 318928 43720 318980
rect 43772 318968 43778 318980
rect 46842 318968 46848 318980
rect 43772 318940 46848 318968
rect 43772 318928 43778 318940
rect 46842 318928 46848 318940
rect 46900 318928 46906 318980
rect 350350 318792 350356 318844
rect 350408 318832 350414 318844
rect 382734 318832 382740 318844
rect 350408 318804 382740 318832
rect 350408 318792 350414 318804
rect 382734 318792 382740 318804
rect 382792 318792 382798 318844
rect 44634 318588 44640 318640
rect 44692 318628 44698 318640
rect 46842 318628 46848 318640
rect 44692 318600 46848 318628
rect 44692 318588 44698 318600
rect 46842 318588 46848 318600
rect 46900 318588 46906 318640
rect 553118 317500 553124 317552
rect 553176 317540 553182 317552
rect 564710 317540 564716 317552
rect 553176 317512 564716 317540
rect 553176 317500 553182 317512
rect 564710 317500 564716 317512
rect 564768 317500 564774 317552
rect 350350 317432 350356 317484
rect 350408 317472 350414 317484
rect 393866 317472 393872 317484
rect 350408 317444 393872 317472
rect 350408 317432 350414 317444
rect 393866 317432 393872 317444
rect 393924 317432 393930 317484
rect 396626 317432 396632 317484
rect 396684 317472 396690 317484
rect 407114 317472 407120 317484
rect 396684 317444 407120 317472
rect 396684 317432 396690 317444
rect 407114 317432 407120 317444
rect 407172 317432 407178 317484
rect 552934 317432 552940 317484
rect 552992 317472 552998 317484
rect 579890 317472 579896 317484
rect 552992 317444 579896 317472
rect 552992 317432 552998 317444
rect 579890 317432 579896 317444
rect 579948 317432 579954 317484
rect 553118 316004 553124 316056
rect 553176 316044 553182 316056
rect 576302 316044 576308 316056
rect 553176 316016 576308 316044
rect 553176 316004 553182 316016
rect 576302 316004 576308 316016
rect 576360 316004 576366 316056
rect 350350 315936 350356 315988
rect 350408 315976 350414 315988
rect 398374 315976 398380 315988
rect 350408 315948 398380 315976
rect 350408 315936 350414 315948
rect 398374 315936 398380 315948
rect 398432 315936 398438 315988
rect 577498 315324 577504 315376
rect 577556 315364 577562 315376
rect 580442 315364 580448 315376
rect 577556 315336 580448 315364
rect 577556 315324 577562 315336
rect 580442 315324 580448 315336
rect 580500 315324 580506 315376
rect 32674 314644 32680 314696
rect 32732 314684 32738 314696
rect 46842 314684 46848 314696
rect 32732 314656 46848 314684
rect 32732 314644 32738 314656
rect 46842 314644 46848 314656
rect 46900 314644 46906 314696
rect 350166 314644 350172 314696
rect 350224 314684 350230 314696
rect 392854 314684 392860 314696
rect 350224 314656 392860 314684
rect 350224 314644 350230 314656
rect 392854 314644 392860 314656
rect 392912 314644 392918 314696
rect 552934 313284 552940 313336
rect 552992 313324 552998 313336
rect 583386 313324 583392 313336
rect 552992 313296 583392 313324
rect 552992 313284 552998 313296
rect 583386 313284 583392 313296
rect 583444 313284 583450 313336
rect 553118 313216 553124 313268
rect 553176 313256 553182 313268
rect 567286 313256 567292 313268
rect 553176 313228 567292 313256
rect 553176 313216 553182 313228
rect 567286 313216 567292 313228
rect 567344 313216 567350 313268
rect 44358 313080 44364 313132
rect 44416 313120 44422 313132
rect 46382 313120 46388 313132
rect 44416 313092 46388 313120
rect 44416 313080 44422 313092
rect 46382 313080 46388 313092
rect 46440 313080 46446 313132
rect 350350 311856 350356 311908
rect 350408 311896 350414 311908
rect 388714 311896 388720 311908
rect 350408 311868 388720 311896
rect 350408 311856 350414 311868
rect 388714 311856 388720 311868
rect 388772 311856 388778 311908
rect 399846 311856 399852 311908
rect 399904 311896 399910 311908
rect 407114 311896 407120 311908
rect 399904 311868 407120 311896
rect 399904 311856 399910 311868
rect 407114 311856 407120 311868
rect 407172 311856 407178 311908
rect 403526 310564 403532 310616
rect 403584 310604 403590 310616
rect 407114 310604 407120 310616
rect 403584 310576 407120 310604
rect 403584 310564 403590 310576
rect 407114 310564 407120 310576
rect 407172 310564 407178 310616
rect 552934 310564 552940 310616
rect 552992 310604 552998 310616
rect 574554 310604 574560 310616
rect 552992 310576 574560 310604
rect 552992 310564 552998 310576
rect 574554 310564 574560 310576
rect 574612 310564 574618 310616
rect 22554 310496 22560 310548
rect 22612 310536 22618 310548
rect 46842 310536 46848 310548
rect 22612 310508 46848 310536
rect 22612 310496 22618 310508
rect 46842 310496 46848 310508
rect 46900 310496 46906 310548
rect 350350 310496 350356 310548
rect 350408 310536 350414 310548
rect 368106 310536 368112 310548
rect 350408 310508 368112 310536
rect 350408 310496 350414 310508
rect 368106 310496 368112 310508
rect 368164 310496 368170 310548
rect 399754 310496 399760 310548
rect 399812 310536 399818 310548
rect 407206 310536 407212 310548
rect 399812 310508 407212 310536
rect 399812 310496 399818 310508
rect 407206 310496 407212 310508
rect 407264 310496 407270 310548
rect 553118 310496 553124 310548
rect 553176 310536 553182 310548
rect 577682 310536 577688 310548
rect 553176 310508 577688 310536
rect 553176 310496 553182 310508
rect 577682 310496 577688 310508
rect 577740 310496 577746 310548
rect 368014 310428 368020 310480
rect 368072 310468 368078 310480
rect 407114 310468 407120 310480
rect 368072 310440 407120 310468
rect 368072 310428 368078 310440
rect 407114 310428 407120 310440
rect 407172 310428 407178 310480
rect 350166 309748 350172 309800
rect 350224 309788 350230 309800
rect 357618 309788 357624 309800
rect 350224 309760 357624 309788
rect 350224 309748 350230 309760
rect 357618 309748 357624 309760
rect 357676 309748 357682 309800
rect 32398 309136 32404 309188
rect 32456 309176 32462 309188
rect 46842 309176 46848 309188
rect 32456 309148 46848 309176
rect 32456 309136 32462 309148
rect 46842 309136 46848 309148
rect 46900 309136 46906 309188
rect 553118 309136 553124 309188
rect 553176 309176 553182 309188
rect 575934 309176 575940 309188
rect 553176 309148 575940 309176
rect 553176 309136 553182 309148
rect 575934 309136 575940 309148
rect 575992 309136 575998 309188
rect 350350 307776 350356 307828
rect 350408 307816 350414 307828
rect 353938 307816 353944 307828
rect 350408 307788 353944 307816
rect 350408 307776 350414 307788
rect 353938 307776 353944 307788
rect 353996 307776 354002 307828
rect 358538 307776 358544 307828
rect 358596 307816 358602 307828
rect 407114 307816 407120 307828
rect 358596 307788 407120 307816
rect 358596 307776 358602 307788
rect 407114 307776 407120 307788
rect 407172 307776 407178 307828
rect 553118 307776 553124 307828
rect 553176 307816 553182 307828
rect 572070 307816 572076 307828
rect 553176 307788 572076 307816
rect 553176 307776 553182 307788
rect 572070 307776 572076 307788
rect 572128 307776 572134 307828
rect 388254 307708 388260 307760
rect 388312 307748 388318 307760
rect 407206 307748 407212 307760
rect 388312 307720 407212 307748
rect 388312 307708 388318 307720
rect 407206 307708 407212 307720
rect 407264 307708 407270 307760
rect 552014 307436 552020 307488
rect 552072 307476 552078 307488
rect 553854 307476 553860 307488
rect 552072 307448 553860 307476
rect 552072 307436 552078 307448
rect 553854 307436 553860 307448
rect 553912 307436 553918 307488
rect 552290 305328 552296 305380
rect 552348 305368 552354 305380
rect 555418 305368 555424 305380
rect 552348 305340 555424 305368
rect 552348 305328 552354 305340
rect 555418 305328 555424 305340
rect 555476 305328 555482 305380
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 26694 305028 26700 305040
rect 3568 305000 26700 305028
rect 3568 304988 3574 305000
rect 26694 304988 26700 305000
rect 26752 304988 26758 305040
rect 349890 304988 349896 305040
rect 349948 305028 349954 305040
rect 350718 305028 350724 305040
rect 349948 305000 350724 305028
rect 349948 304988 349954 305000
rect 350718 304988 350724 305000
rect 350776 304988 350782 305040
rect 398006 304988 398012 305040
rect 398064 305028 398070 305040
rect 407114 305028 407120 305040
rect 398064 305000 407120 305028
rect 398064 304988 398070 305000
rect 407114 304988 407120 305000
rect 407172 304988 407178 305040
rect 553118 304988 553124 305040
rect 553176 305028 553182 305040
rect 583478 305028 583484 305040
rect 553176 305000 583484 305028
rect 553176 304988 553182 305000
rect 583478 304988 583484 305000
rect 583536 304988 583542 305040
rect 351178 304308 351184 304360
rect 351236 304348 351242 304360
rect 352650 304348 352656 304360
rect 351236 304320 352656 304348
rect 351236 304308 351242 304320
rect 352650 304308 352656 304320
rect 352708 304308 352714 304360
rect 350350 303696 350356 303748
rect 350408 303736 350414 303748
rect 374546 303736 374552 303748
rect 350408 303708 374552 303736
rect 350408 303696 350414 303708
rect 374546 303696 374552 303708
rect 374604 303696 374610 303748
rect 31294 303628 31300 303680
rect 31352 303668 31358 303680
rect 46842 303668 46848 303680
rect 31352 303640 46848 303668
rect 31352 303628 31358 303640
rect 46842 303628 46848 303640
rect 46900 303628 46906 303680
rect 359642 303628 359648 303680
rect 359700 303668 359706 303680
rect 407114 303668 407120 303680
rect 359700 303640 407120 303668
rect 359700 303628 359706 303640
rect 407114 303628 407120 303640
rect 407172 303628 407178 303680
rect 372798 302880 372804 302932
rect 372856 302920 372862 302932
rect 379422 302920 379428 302932
rect 372856 302892 379428 302920
rect 372856 302880 372862 302892
rect 379422 302880 379428 302892
rect 379480 302880 379486 302932
rect 350350 302268 350356 302320
rect 350408 302308 350414 302320
rect 354214 302308 354220 302320
rect 350408 302280 354220 302308
rect 350408 302268 350414 302280
rect 354214 302268 354220 302280
rect 354272 302268 354278 302320
rect 25590 302200 25596 302252
rect 25648 302240 25654 302252
rect 46474 302240 46480 302252
rect 25648 302212 46480 302240
rect 25648 302200 25654 302212
rect 46474 302200 46480 302212
rect 46532 302200 46538 302252
rect 349798 302200 349804 302252
rect 349856 302240 349862 302252
rect 350534 302240 350540 302252
rect 349856 302212 350540 302240
rect 349856 302200 349862 302212
rect 350534 302200 350540 302212
rect 350592 302200 350598 302252
rect 405182 302200 405188 302252
rect 405240 302240 405246 302252
rect 407390 302240 407396 302252
rect 405240 302212 407396 302240
rect 405240 302200 405246 302212
rect 407390 302200 407396 302212
rect 407448 302200 407454 302252
rect 43530 302132 43536 302184
rect 43588 302172 43594 302184
rect 46842 302172 46848 302184
rect 43588 302144 46848 302172
rect 43588 302132 43594 302144
rect 46842 302132 46848 302144
rect 46900 302132 46906 302184
rect 401042 300908 401048 300960
rect 401100 300948 401106 300960
rect 407114 300948 407120 300960
rect 401100 300920 407120 300948
rect 401100 300908 401106 300920
rect 407114 300908 407120 300920
rect 407172 300908 407178 300960
rect 21266 300840 21272 300892
rect 21324 300880 21330 300892
rect 46842 300880 46848 300892
rect 21324 300852 46848 300880
rect 21324 300840 21330 300852
rect 46842 300840 46848 300852
rect 46900 300840 46906 300892
rect 350350 300840 350356 300892
rect 350408 300880 350414 300892
rect 365438 300880 365444 300892
rect 350408 300852 365444 300880
rect 350408 300840 350414 300852
rect 365438 300840 365444 300852
rect 365496 300840 365502 300892
rect 366726 300840 366732 300892
rect 366784 300880 366790 300892
rect 407206 300880 407212 300892
rect 366784 300852 407212 300880
rect 366784 300840 366790 300852
rect 407206 300840 407212 300852
rect 407264 300840 407270 300892
rect 553118 300840 553124 300892
rect 553176 300880 553182 300892
rect 570506 300880 570512 300892
rect 553176 300852 570512 300880
rect 553176 300840 553182 300852
rect 570506 300840 570512 300852
rect 570564 300840 570570 300892
rect 350074 300772 350080 300824
rect 350132 300812 350138 300824
rect 353662 300812 353668 300824
rect 350132 300784 353668 300812
rect 350132 300772 350138 300784
rect 353662 300772 353668 300784
rect 353720 300772 353726 300824
rect 350350 299548 350356 299600
rect 350408 299588 350414 299600
rect 379422 299588 379428 299600
rect 350408 299560 379428 299588
rect 350408 299548 350414 299560
rect 379422 299548 379428 299560
rect 379480 299548 379486 299600
rect 368014 299480 368020 299532
rect 368072 299520 368078 299532
rect 407114 299520 407120 299532
rect 368072 299492 407120 299520
rect 368072 299480 368078 299492
rect 407114 299480 407120 299492
rect 407172 299480 407178 299532
rect 553118 299480 553124 299532
rect 553176 299520 553182 299532
rect 571886 299520 571892 299532
rect 553176 299492 571892 299520
rect 553176 299480 553182 299492
rect 571886 299480 571892 299492
rect 571944 299480 571950 299532
rect 18966 298120 18972 298172
rect 19024 298160 19030 298172
rect 46842 298160 46848 298172
rect 19024 298132 46848 298160
rect 19024 298120 19030 298132
rect 46842 298120 46848 298132
rect 46900 298120 46906 298172
rect 350350 298120 350356 298172
rect 350408 298160 350414 298172
rect 354030 298160 354036 298172
rect 350408 298132 354036 298160
rect 350408 298120 350414 298132
rect 354030 298120 354036 298132
rect 354088 298120 354094 298172
rect 350074 297984 350080 298036
rect 350132 298024 350138 298036
rect 350350 298024 350356 298036
rect 350132 297996 350356 298024
rect 350132 297984 350138 297996
rect 350350 297984 350356 297996
rect 350408 297984 350414 298036
rect 553118 297848 553124 297900
rect 553176 297888 553182 297900
rect 556890 297888 556896 297900
rect 553176 297860 556896 297888
rect 553176 297848 553182 297860
rect 556890 297848 556896 297860
rect 556948 297848 556954 297900
rect 18874 296692 18880 296744
rect 18932 296732 18938 296744
rect 46842 296732 46848 296744
rect 18932 296704 46848 296732
rect 18932 296692 18938 296704
rect 46842 296692 46848 296704
rect 46900 296692 46906 296744
rect 553118 296692 553124 296744
rect 553176 296732 553182 296744
rect 572162 296732 572168 296744
rect 553176 296704 572168 296732
rect 553176 296692 553182 296704
rect 572162 296692 572168 296704
rect 572220 296692 572226 296744
rect 350074 295468 350080 295520
rect 350132 295508 350138 295520
rect 350258 295508 350264 295520
rect 350132 295480 350264 295508
rect 350132 295468 350138 295480
rect 350258 295468 350264 295480
rect 350316 295468 350322 295520
rect 348418 295332 348424 295384
rect 348476 295372 348482 295384
rect 349246 295372 349252 295384
rect 348476 295344 349252 295372
rect 348476 295332 348482 295344
rect 349246 295332 349252 295344
rect 349304 295332 349310 295384
rect 350258 295332 350264 295384
rect 350316 295372 350322 295384
rect 379974 295372 379980 295384
rect 350316 295344 379980 295372
rect 350316 295332 350322 295344
rect 379974 295332 379980 295344
rect 380032 295332 380038 295384
rect 399386 295332 399392 295384
rect 399444 295372 399450 295384
rect 407114 295372 407120 295384
rect 399444 295344 407120 295372
rect 399444 295332 399450 295344
rect 407114 295332 407120 295344
rect 407172 295332 407178 295384
rect 365162 294584 365168 294636
rect 365220 294624 365226 294636
rect 384206 294624 384212 294636
rect 365220 294596 384212 294624
rect 365220 294584 365226 294596
rect 384206 294584 384212 294596
rect 384264 294584 384270 294636
rect 348970 294040 348976 294092
rect 349028 294080 349034 294092
rect 350534 294080 350540 294092
rect 349028 294052 350540 294080
rect 349028 294040 349034 294052
rect 350534 294040 350540 294052
rect 350592 294040 350598 294092
rect 350258 293972 350264 294024
rect 350316 294012 350322 294024
rect 368934 294012 368940 294024
rect 350316 293984 368940 294012
rect 350316 293972 350322 293984
rect 368934 293972 368940 293984
rect 368992 293972 368998 294024
rect 32766 293904 32772 293956
rect 32824 293944 32830 293956
rect 46474 293944 46480 293956
rect 32824 293916 46480 293944
rect 32824 293904 32830 293916
rect 46474 293904 46480 293916
rect 46532 293904 46538 293956
rect 552014 293088 552020 293140
rect 552072 293128 552078 293140
rect 553762 293128 553768 293140
rect 552072 293100 553768 293128
rect 552072 293088 552078 293100
rect 553762 293088 553768 293100
rect 553820 293088 553826 293140
rect 371050 292612 371056 292664
rect 371108 292652 371114 292664
rect 407114 292652 407120 292664
rect 371108 292624 407120 292652
rect 371108 292612 371114 292624
rect 407114 292612 407120 292624
rect 407172 292612 407178 292664
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 20162 292584 20168 292596
rect 3568 292556 20168 292584
rect 3568 292544 3574 292556
rect 20162 292544 20168 292556
rect 20220 292544 20226 292596
rect 44634 292544 44640 292596
rect 44692 292584 44698 292596
rect 46842 292584 46848 292596
rect 44692 292556 46848 292584
rect 44692 292544 44698 292556
rect 46842 292544 46848 292556
rect 46900 292544 46906 292596
rect 365162 292544 365168 292596
rect 365220 292584 365226 292596
rect 407206 292584 407212 292596
rect 365220 292556 407212 292584
rect 365220 292544 365226 292556
rect 407206 292544 407212 292556
rect 407264 292544 407270 292596
rect 399662 292476 399668 292528
rect 399720 292516 399726 292528
rect 407114 292516 407120 292528
rect 399720 292488 407120 292516
rect 399720 292476 399726 292488
rect 407114 292476 407120 292488
rect 407172 292476 407178 292528
rect 401226 292408 401232 292460
rect 401284 292448 401290 292460
rect 407206 292448 407212 292460
rect 401284 292420 407212 292448
rect 401284 292408 401290 292420
rect 407206 292408 407212 292420
rect 407264 292408 407270 292460
rect 552198 291728 552204 291780
rect 552256 291768 552262 291780
rect 555510 291768 555516 291780
rect 552256 291740 555516 291768
rect 552256 291728 552262 291740
rect 555510 291728 555516 291740
rect 555568 291728 555574 291780
rect 43530 291184 43536 291236
rect 43588 291224 43594 291236
rect 46842 291224 46848 291236
rect 43588 291196 46848 291224
rect 43588 291184 43594 291196
rect 46842 291184 46848 291196
rect 46900 291184 46906 291236
rect 553118 291184 553124 291236
rect 553176 291224 553182 291236
rect 562318 291224 562324 291236
rect 553176 291196 562324 291224
rect 553176 291184 553182 291196
rect 562318 291184 562324 291196
rect 562376 291184 562382 291236
rect 552014 290096 552020 290148
rect 552072 290136 552078 290148
rect 553854 290136 553860 290148
rect 552072 290108 553860 290136
rect 552072 290096 552078 290108
rect 553854 290096 553860 290108
rect 553912 290096 553918 290148
rect 351178 288464 351184 288516
rect 351236 288504 351242 288516
rect 356514 288504 356520 288516
rect 351236 288476 356520 288504
rect 351236 288464 351242 288476
rect 356514 288464 356520 288476
rect 356572 288464 356578 288516
rect 395614 288464 395620 288516
rect 395672 288504 395678 288516
rect 407114 288504 407120 288516
rect 395672 288476 407120 288504
rect 395672 288464 395678 288476
rect 407114 288464 407120 288476
rect 407172 288464 407178 288516
rect 552934 288464 552940 288516
rect 552992 288504 552998 288516
rect 563882 288504 563888 288516
rect 552992 288476 563888 288504
rect 552992 288464 552998 288476
rect 563882 288464 563888 288476
rect 563940 288464 563946 288516
rect 28534 288396 28540 288448
rect 28592 288436 28598 288448
rect 46842 288436 46848 288448
rect 28592 288408 46848 288436
rect 28592 288396 28598 288408
rect 46842 288396 46848 288408
rect 46900 288396 46906 288448
rect 350258 288396 350264 288448
rect 350316 288436 350322 288448
rect 386874 288436 386880 288448
rect 350316 288408 386880 288436
rect 350316 288396 350322 288408
rect 386874 288396 386880 288408
rect 386932 288396 386938 288448
rect 553118 288396 553124 288448
rect 553176 288436 553182 288448
rect 578510 288436 578516 288448
rect 553176 288408 578516 288436
rect 553176 288396 553182 288408
rect 578510 288396 578516 288408
rect 578568 288396 578574 288448
rect 404906 287376 404912 287428
rect 404964 287416 404970 287428
rect 407206 287416 407212 287428
rect 404964 287388 407212 287416
rect 404964 287376 404970 287388
rect 407206 287376 407212 287388
rect 407264 287376 407270 287428
rect 391106 287172 391112 287224
rect 391164 287212 391170 287224
rect 407114 287212 407120 287224
rect 391164 287184 407120 287212
rect 391164 287172 391170 287184
rect 407114 287172 407120 287184
rect 407172 287172 407178 287224
rect 350258 287104 350264 287156
rect 350316 287144 350322 287156
rect 357066 287144 357072 287156
rect 350316 287116 357072 287144
rect 350316 287104 350322 287116
rect 357066 287104 357072 287116
rect 357124 287104 357130 287156
rect 350258 286968 350264 287020
rect 350316 287008 350322 287020
rect 356422 287008 356428 287020
rect 350316 286980 356428 287008
rect 350316 286968 350322 286980
rect 356422 286968 356428 286980
rect 356480 286968 356486 287020
rect 349338 286220 349344 286272
rect 349396 286260 349402 286272
rect 350626 286260 350632 286272
rect 349396 286232 350632 286260
rect 349396 286220 349402 286232
rect 350626 286220 350632 286232
rect 350684 286220 350690 286272
rect 355502 285744 355508 285796
rect 355560 285784 355566 285796
rect 399294 285784 399300 285796
rect 355560 285756 399300 285784
rect 355560 285744 355566 285756
rect 399294 285744 399300 285756
rect 399352 285744 399358 285796
rect 30926 285676 30932 285728
rect 30984 285716 30990 285728
rect 46842 285716 46848 285728
rect 30984 285688 46848 285716
rect 30984 285676 30990 285688
rect 46842 285676 46848 285688
rect 46900 285676 46906 285728
rect 349798 285676 349804 285728
rect 349856 285716 349862 285728
rect 407114 285716 407120 285728
rect 349856 285688 407120 285716
rect 349856 285676 349862 285688
rect 407114 285676 407120 285688
rect 407172 285676 407178 285728
rect 553118 285676 553124 285728
rect 553176 285716 553182 285728
rect 569586 285716 569592 285728
rect 553176 285688 569592 285716
rect 553176 285676 553182 285688
rect 569586 285676 569592 285688
rect 569644 285676 569650 285728
rect 350258 285608 350264 285660
rect 350316 285648 350322 285660
rect 365530 285648 365536 285660
rect 350316 285620 365536 285648
rect 350316 285608 350322 285620
rect 365530 285608 365536 285620
rect 365588 285608 365594 285660
rect 403894 285608 403900 285660
rect 403952 285648 403958 285660
rect 407206 285648 407212 285660
rect 403952 285620 407212 285648
rect 403952 285608 403958 285620
rect 407206 285608 407212 285620
rect 407264 285608 407270 285660
rect 43438 284316 43444 284368
rect 43496 284356 43502 284368
rect 44818 284356 44824 284368
rect 43496 284328 44824 284356
rect 43496 284316 43502 284328
rect 44818 284316 44824 284328
rect 44876 284316 44882 284368
rect 392486 284316 392492 284368
rect 392544 284356 392550 284368
rect 407114 284356 407120 284368
rect 392544 284328 407120 284356
rect 392544 284316 392550 284328
rect 407114 284316 407120 284328
rect 407172 284316 407178 284368
rect 368290 284248 368296 284300
rect 368348 284288 368354 284300
rect 407206 284288 407212 284300
rect 368348 284260 407212 284288
rect 368348 284248 368354 284260
rect 407206 284248 407212 284260
rect 407264 284248 407270 284300
rect 553118 283568 553124 283620
rect 553176 283608 553182 283620
rect 564710 283608 564716 283620
rect 553176 283580 564716 283608
rect 553176 283568 553182 283580
rect 564710 283568 564716 283580
rect 564768 283568 564774 283620
rect 368198 282888 368204 282940
rect 368256 282928 368262 282940
rect 407114 282928 407120 282940
rect 368256 282900 407120 282928
rect 368256 282888 368262 282900
rect 407114 282888 407120 282900
rect 407172 282888 407178 282940
rect 553118 282820 553124 282872
rect 553176 282860 553182 282872
rect 568758 282860 568764 282872
rect 553176 282832 568764 282860
rect 553176 282820 553182 282832
rect 568758 282820 568764 282832
rect 568816 282820 568822 282872
rect 348418 282004 348424 282056
rect 348476 282044 348482 282056
rect 349154 282044 349160 282056
rect 348476 282016 349160 282044
rect 348476 282004 348482 282016
rect 349154 282004 349160 282016
rect 349212 282004 349218 282056
rect 25314 281528 25320 281580
rect 25372 281568 25378 281580
rect 46842 281568 46848 281580
rect 25372 281540 46848 281568
rect 25372 281528 25378 281540
rect 46842 281528 46848 281540
rect 46900 281528 46906 281580
rect 405090 281392 405096 281444
rect 405148 281432 405154 281444
rect 409230 281432 409236 281444
rect 405148 281404 409236 281432
rect 405148 281392 405154 281404
rect 409230 281392 409236 281404
rect 409288 281392 409294 281444
rect 553118 280848 553124 280900
rect 553176 280888 553182 280900
rect 558270 280888 558276 280900
rect 553176 280860 558276 280888
rect 553176 280848 553182 280860
rect 558270 280848 558276 280860
rect 558328 280848 558334 280900
rect 553118 280168 553124 280220
rect 553176 280208 553182 280220
rect 564986 280208 564992 280220
rect 553176 280180 564992 280208
rect 553176 280168 553182 280180
rect 564986 280168 564992 280180
rect 565044 280168 565050 280220
rect 552934 280100 552940 280152
rect 552992 280140 552998 280152
rect 564802 280140 564808 280152
rect 552992 280112 564808 280140
rect 552992 280100 552998 280112
rect 564802 280100 564808 280112
rect 564860 280100 564866 280152
rect 395154 278740 395160 278792
rect 395212 278780 395218 278792
rect 407114 278780 407120 278792
rect 395212 278752 407120 278780
rect 395212 278740 395218 278752
rect 407114 278740 407120 278752
rect 407172 278740 407178 278792
rect 553118 278740 553124 278792
rect 553176 278780 553182 278792
rect 570874 278780 570880 278792
rect 553176 278752 570880 278780
rect 553176 278740 553182 278752
rect 570874 278740 570880 278752
rect 570932 278740 570938 278792
rect 402054 277992 402060 278044
rect 402112 278032 402118 278044
rect 408034 278032 408040 278044
rect 402112 278004 408040 278032
rect 402112 277992 402118 278004
rect 408034 277992 408040 278004
rect 408092 277992 408098 278044
rect 20346 277380 20352 277432
rect 20404 277420 20410 277432
rect 46842 277420 46848 277432
rect 20404 277392 46848 277420
rect 20404 277380 20410 277392
rect 46842 277380 46848 277392
rect 46900 277380 46906 277432
rect 350258 277380 350264 277432
rect 350316 277420 350322 277432
rect 403434 277420 403440 277432
rect 350316 277392 403440 277420
rect 350316 277380 350322 277392
rect 403434 277380 403440 277392
rect 403492 277380 403498 277432
rect 553118 277380 553124 277432
rect 553176 277420 553182 277432
rect 563790 277420 563796 277432
rect 553176 277392 563796 277420
rect 553176 277380 553182 277392
rect 563790 277380 563796 277392
rect 563848 277380 563854 277432
rect 391290 277312 391296 277364
rect 391348 277352 391354 277364
rect 407114 277352 407120 277364
rect 391348 277324 407120 277352
rect 391348 277312 391354 277324
rect 407114 277312 407120 277324
rect 407172 277312 407178 277364
rect 348878 276020 348884 276072
rect 348936 276060 348942 276072
rect 350534 276060 350540 276072
rect 348936 276032 350540 276060
rect 348936 276020 348942 276032
rect 350534 276020 350540 276032
rect 350592 276020 350598 276072
rect 553118 276020 553124 276072
rect 553176 276060 553182 276072
rect 576026 276060 576032 276072
rect 553176 276032 576032 276060
rect 553176 276020 553182 276032
rect 576026 276020 576032 276032
rect 576084 276020 576090 276072
rect 365070 275952 365076 276004
rect 365128 275992 365134 276004
rect 407114 275992 407120 276004
rect 365128 275964 407120 275992
rect 365128 275952 365134 275964
rect 407114 275952 407120 275964
rect 407172 275952 407178 276004
rect 350258 275884 350264 275936
rect 350316 275924 350322 275936
rect 387242 275924 387248 275936
rect 350316 275896 387248 275924
rect 350316 275884 350322 275896
rect 387242 275884 387248 275896
rect 387300 275884 387306 275936
rect 352558 275272 352564 275324
rect 352616 275312 352622 275324
rect 357618 275312 357624 275324
rect 352616 275284 357624 275312
rect 352616 275272 352622 275284
rect 357618 275272 357624 275284
rect 357676 275272 357682 275324
rect 40770 274864 40776 274916
rect 40828 274904 40834 274916
rect 46934 274904 46940 274916
rect 40828 274876 46940 274904
rect 40828 274864 40834 274876
rect 46934 274864 46940 274876
rect 46992 274864 46998 274916
rect 552290 274728 552296 274780
rect 552348 274768 552354 274780
rect 555234 274768 555240 274780
rect 552348 274740 555240 274768
rect 552348 274728 552354 274740
rect 555234 274728 555240 274740
rect 555292 274728 555298 274780
rect 350258 273368 350264 273420
rect 350316 273408 350322 273420
rect 355502 273408 355508 273420
rect 350316 273380 355508 273408
rect 350316 273368 350322 273380
rect 355502 273368 355508 273380
rect 355560 273368 355566 273420
rect 349982 273300 349988 273352
rect 350040 273340 350046 273352
rect 353570 273340 353576 273352
rect 350040 273312 353576 273340
rect 350040 273300 350046 273312
rect 353570 273300 353576 273312
rect 353628 273300 353634 273352
rect 350166 273232 350172 273284
rect 350224 273272 350230 273284
rect 391014 273272 391020 273284
rect 350224 273244 391020 273272
rect 350224 273232 350230 273244
rect 391014 273232 391020 273244
rect 391072 273232 391078 273284
rect 553118 273232 553124 273284
rect 553176 273272 553182 273284
rect 579982 273272 579988 273284
rect 553176 273244 579988 273272
rect 553176 273232 553182 273244
rect 579982 273232 579988 273244
rect 580040 273232 580046 273284
rect 572070 273164 572076 273216
rect 572128 273204 572134 273216
rect 580166 273204 580172 273216
rect 572128 273176 580172 273204
rect 572128 273164 572134 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 407482 272552 407488 272604
rect 407540 272592 407546 272604
rect 407758 272592 407764 272604
rect 407540 272564 407764 272592
rect 407540 272552 407546 272564
rect 407758 272552 407764 272564
rect 407816 272552 407822 272604
rect 350258 271872 350264 271924
rect 350316 271912 350322 271924
rect 353570 271912 353576 271924
rect 350316 271884 353576 271912
rect 350316 271872 350322 271884
rect 353570 271872 353576 271884
rect 353628 271872 353634 271924
rect 398374 271872 398380 271924
rect 398432 271912 398438 271924
rect 407114 271912 407120 271924
rect 398432 271884 407120 271912
rect 398432 271872 398438 271884
rect 407114 271872 407120 271884
rect 407172 271872 407178 271924
rect 403986 271804 403992 271856
rect 404044 271844 404050 271856
rect 407206 271844 407212 271856
rect 404044 271816 407212 271844
rect 404044 271804 404050 271816
rect 407206 271804 407212 271816
rect 407264 271804 407270 271856
rect 553118 270512 553124 270564
rect 553176 270552 553182 270564
rect 577498 270552 577504 270564
rect 553176 270524 577504 270552
rect 553176 270512 553182 270524
rect 577498 270512 577504 270524
rect 577556 270512 577562 270564
rect 350258 270444 350264 270496
rect 350316 270484 350322 270496
rect 395338 270484 395344 270496
rect 350316 270456 395344 270484
rect 350316 270444 350322 270456
rect 395338 270444 395344 270456
rect 395396 270444 395402 270496
rect 350074 270376 350080 270428
rect 350132 270416 350138 270428
rect 350810 270416 350816 270428
rect 350132 270388 350816 270416
rect 350132 270376 350138 270388
rect 350810 270376 350816 270388
rect 350868 270376 350874 270428
rect 40494 270240 40500 270292
rect 40552 270280 40558 270292
rect 43438 270280 43444 270292
rect 40552 270252 43444 270280
rect 40552 270240 40558 270252
rect 43438 270240 43444 270252
rect 43496 270240 43502 270292
rect 551922 270036 551928 270088
rect 551980 270076 551986 270088
rect 552842 270076 552848 270088
rect 551980 270048 552848 270076
rect 551980 270036 551986 270048
rect 552842 270036 552848 270048
rect 552900 270036 552906 270088
rect 376478 269084 376484 269136
rect 376536 269124 376542 269136
rect 407114 269124 407120 269136
rect 376536 269096 407120 269124
rect 376536 269084 376542 269096
rect 407114 269084 407120 269096
rect 407172 269084 407178 269136
rect 348878 269016 348884 269068
rect 348936 269056 348942 269068
rect 350534 269056 350540 269068
rect 348936 269028 350540 269056
rect 348936 269016 348942 269028
rect 350534 269016 350540 269028
rect 350592 269016 350598 269068
rect 348970 268948 348976 269000
rect 349028 268988 349034 269000
rect 349154 268988 349160 269000
rect 349028 268960 349160 268988
rect 349028 268948 349034 268960
rect 349154 268948 349160 268960
rect 349212 268948 349218 269000
rect 350258 268948 350264 269000
rect 350316 268988 350322 269000
rect 355134 268988 355140 269000
rect 350316 268960 355140 268988
rect 350316 268948 350322 268960
rect 355134 268948 355140 268960
rect 355192 268948 355198 269000
rect 348970 268812 348976 268864
rect 349028 268852 349034 268864
rect 349522 268852 349528 268864
rect 349028 268824 349528 268852
rect 349028 268812 349034 268824
rect 349522 268812 349528 268824
rect 349580 268812 349586 268864
rect 553118 268608 553124 268660
rect 553176 268648 553182 268660
rect 556982 268648 556988 268660
rect 553176 268620 556988 268648
rect 553176 268608 553182 268620
rect 556982 268608 556988 268620
rect 557040 268608 557046 268660
rect 36630 268064 36636 268116
rect 36688 268104 36694 268116
rect 39298 268104 39304 268116
rect 36688 268076 39304 268104
rect 36688 268064 36694 268076
rect 39298 268064 39304 268076
rect 39356 268064 39362 268116
rect 43438 267792 43444 267844
rect 43496 267832 43502 267844
rect 46842 267832 46848 267844
rect 43496 267804 46848 267832
rect 43496 267792 43502 267804
rect 46842 267792 46848 267804
rect 46900 267792 46906 267844
rect 43254 267724 43260 267776
rect 43312 267764 43318 267776
rect 44174 267764 44180 267776
rect 43312 267736 44180 267764
rect 43312 267724 43318 267736
rect 44174 267724 44180 267736
rect 44232 267724 44238 267776
rect 402790 267724 402796 267776
rect 402848 267764 402854 267776
rect 407114 267764 407120 267776
rect 402848 267736 407120 267764
rect 402848 267724 402854 267736
rect 407114 267724 407120 267736
rect 407172 267724 407178 267776
rect 35066 266976 35072 267028
rect 35124 267016 35130 267028
rect 39114 267016 39120 267028
rect 35124 266988 39120 267016
rect 35124 266976 35130 266988
rect 39114 266976 39120 266988
rect 39172 266976 39178 267028
rect 350258 266364 350264 266416
rect 350316 266404 350322 266416
rect 389726 266404 389732 266416
rect 350316 266376 389732 266404
rect 350316 266364 350322 266376
rect 389726 266364 389732 266376
rect 389784 266364 389790 266416
rect 405642 266364 405648 266416
rect 405700 266404 405706 266416
rect 407758 266404 407764 266416
rect 405700 266376 407764 266404
rect 405700 266364 405706 266376
rect 407758 266364 407764 266376
rect 407816 266364 407822 266416
rect 367922 265616 367928 265668
rect 367980 265656 367986 265668
rect 396442 265656 396448 265668
rect 367980 265628 396448 265656
rect 367980 265616 367986 265628
rect 396442 265616 396448 265628
rect 396500 265616 396506 265668
rect 553118 264936 553124 264988
rect 553176 264976 553182 264988
rect 570322 264976 570328 264988
rect 553176 264948 570328 264976
rect 553176 264936 553182 264948
rect 570322 264936 570328 264948
rect 570380 264936 570386 264988
rect 350258 263644 350264 263696
rect 350316 263684 350322 263696
rect 367462 263684 367468 263696
rect 350316 263656 367468 263684
rect 350316 263644 350322 263656
rect 367462 263644 367468 263656
rect 367520 263644 367526 263696
rect 553118 263644 553124 263696
rect 553176 263684 553182 263696
rect 567746 263684 567752 263696
rect 553176 263656 567752 263684
rect 553176 263644 553182 263656
rect 567746 263644 567752 263656
rect 567804 263644 567810 263696
rect 46290 263576 46296 263628
rect 46348 263616 46354 263628
rect 46934 263616 46940 263628
rect 46348 263588 46940 263616
rect 46348 263576 46354 263588
rect 46934 263576 46940 263588
rect 46992 263576 46998 263628
rect 365622 263576 365628 263628
rect 365680 263616 365686 263628
rect 407114 263616 407120 263628
rect 365680 263588 407120 263616
rect 365680 263576 365686 263588
rect 407114 263576 407120 263588
rect 407172 263576 407178 263628
rect 552934 263576 552940 263628
rect 552992 263616 552998 263628
rect 568574 263616 568580 263628
rect 552992 263588 568580 263616
rect 552992 263576 552998 263588
rect 568574 263576 568580 263588
rect 568632 263576 568638 263628
rect 365530 262896 365536 262948
rect 365588 262936 365594 262948
rect 367186 262936 367192 262948
rect 365588 262908 367192 262936
rect 365588 262896 365594 262908
rect 367186 262896 367192 262908
rect 367244 262896 367250 262948
rect 552014 262352 552020 262404
rect 552072 262392 552078 262404
rect 554774 262392 554780 262404
rect 552072 262364 554780 262392
rect 552072 262352 552078 262364
rect 554774 262352 554780 262364
rect 554832 262352 554838 262404
rect 349430 262216 349436 262268
rect 349488 262256 349494 262268
rect 351270 262256 351276 262268
rect 349488 262228 351276 262256
rect 349488 262216 349494 262228
rect 351270 262216 351276 262228
rect 351328 262216 351334 262268
rect 403894 262216 403900 262268
rect 403952 262256 403958 262268
rect 407114 262256 407120 262268
rect 403952 262228 407120 262256
rect 403952 262216 403958 262228
rect 407114 262216 407120 262228
rect 407172 262216 407178 262268
rect 36354 262148 36360 262200
rect 36412 262188 36418 262200
rect 43254 262188 43260 262200
rect 36412 262160 43260 262188
rect 36412 262148 36418 262160
rect 43254 262148 43260 262160
rect 43312 262148 43318 262200
rect 348970 262148 348976 262200
rect 349028 262188 349034 262200
rect 349246 262188 349252 262200
rect 349028 262160 349252 262188
rect 349028 262148 349034 262160
rect 349246 262148 349252 262160
rect 349304 262148 349310 262200
rect 350258 262148 350264 262200
rect 350316 262188 350322 262200
rect 365622 262188 365628 262200
rect 350316 262160 365628 262188
rect 350316 262148 350322 262160
rect 365622 262148 365628 262160
rect 365680 262148 365686 262200
rect 404998 262148 405004 262200
rect 405056 262188 405062 262200
rect 406562 262188 406568 262200
rect 405056 262160 406568 262188
rect 405056 262148 405062 262160
rect 406562 262148 406568 262160
rect 406620 262148 406626 262200
rect 395062 261060 395068 261112
rect 395120 261100 395126 261112
rect 396718 261100 396724 261112
rect 395120 261072 396724 261100
rect 395120 261060 395126 261072
rect 396718 261060 396724 261072
rect 396776 261060 396782 261112
rect 401226 260856 401232 260908
rect 401284 260896 401290 260908
rect 407114 260896 407120 260908
rect 401284 260868 407120 260896
rect 401284 260856 401290 260868
rect 407114 260856 407120 260868
rect 407172 260856 407178 260908
rect 553118 260856 553124 260908
rect 553176 260896 553182 260908
rect 564802 260896 564808 260908
rect 553176 260868 564808 260896
rect 553176 260856 553182 260868
rect 564802 260856 564808 260868
rect 564860 260856 564866 260908
rect 348970 260788 348976 260840
rect 349028 260828 349034 260840
rect 349154 260828 349160 260840
rect 349028 260800 349160 260828
rect 349028 260788 349034 260800
rect 349154 260788 349160 260800
rect 349212 260788 349218 260840
rect 385494 260788 385500 260840
rect 385552 260828 385558 260840
rect 387242 260828 387248 260840
rect 385552 260800 387248 260828
rect 385552 260788 385558 260800
rect 387242 260788 387248 260800
rect 387300 260788 387306 260840
rect 552934 259496 552940 259548
rect 552992 259536 552998 259548
rect 567286 259536 567292 259548
rect 552992 259508 567292 259536
rect 552992 259496 552998 259508
rect 567286 259496 567292 259508
rect 567344 259496 567350 259548
rect 45462 259428 45468 259480
rect 45520 259468 45526 259480
rect 46934 259468 46940 259480
rect 45520 259440 46940 259468
rect 45520 259428 45526 259440
rect 46934 259428 46940 259440
rect 46992 259428 46998 259480
rect 396534 259428 396540 259480
rect 396592 259468 396598 259480
rect 407114 259468 407120 259480
rect 396592 259440 407120 259468
rect 396592 259428 396598 259440
rect 407114 259428 407120 259440
rect 407172 259428 407178 259480
rect 553118 259428 553124 259480
rect 553176 259468 553182 259480
rect 583570 259468 583576 259480
rect 553176 259440 583576 259468
rect 553176 259428 553182 259440
rect 583570 259428 583576 259440
rect 583628 259428 583634 259480
rect 376294 259360 376300 259412
rect 376352 259400 376358 259412
rect 377214 259400 377220 259412
rect 376352 259372 377220 259400
rect 376352 259360 376358 259372
rect 377214 259360 377220 259372
rect 377272 259360 377278 259412
rect 570598 259360 570604 259412
rect 570656 259400 570662 259412
rect 580166 259400 580172 259412
rect 570656 259372 580172 259400
rect 570656 259360 570662 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 349522 258068 349528 258120
rect 349580 258108 349586 258120
rect 385494 258108 385500 258120
rect 349580 258080 385500 258108
rect 349580 258068 349586 258080
rect 385494 258068 385500 258080
rect 385552 258068 385558 258120
rect 553118 258068 553124 258120
rect 553176 258108 553182 258120
rect 560294 258108 560300 258120
rect 553176 258080 560300 258108
rect 553176 258068 553182 258080
rect 560294 258068 560300 258080
rect 560352 258068 560358 258120
rect 376294 256776 376300 256828
rect 376352 256816 376358 256828
rect 407114 256816 407120 256828
rect 376352 256788 407120 256816
rect 376352 256776 376358 256788
rect 407114 256776 407120 256788
rect 407172 256776 407178 256828
rect 356974 256708 356980 256760
rect 357032 256748 357038 256760
rect 407206 256748 407212 256760
rect 357032 256720 407212 256748
rect 357032 256708 357038 256720
rect 407206 256708 407212 256720
rect 407264 256708 407270 256760
rect 553118 256708 553124 256760
rect 553176 256748 553182 256760
rect 564434 256748 564440 256760
rect 553176 256720 564440 256748
rect 553176 256708 553182 256720
rect 564434 256708 564440 256720
rect 564492 256708 564498 256760
rect 45278 255688 45284 255740
rect 45336 255728 45342 255740
rect 45738 255728 45744 255740
rect 45336 255700 45744 255728
rect 45336 255688 45342 255700
rect 45738 255688 45744 255700
rect 45796 255688 45802 255740
rect 350166 255416 350172 255468
rect 350224 255456 350230 255468
rect 350442 255456 350448 255468
rect 350224 255428 350448 255456
rect 350224 255416 350230 255428
rect 350442 255416 350448 255428
rect 350500 255416 350506 255468
rect 350442 255280 350448 255332
rect 350500 255320 350506 255332
rect 393774 255320 393780 255332
rect 350500 255292 393780 255320
rect 350500 255280 350506 255292
rect 393774 255280 393780 255292
rect 393832 255280 393838 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 31018 255252 31024 255264
rect 3200 255224 31024 255252
rect 3200 255212 3206 255224
rect 31018 255212 31024 255224
rect 31076 255212 31082 255264
rect 405366 255212 405372 255264
rect 405424 255252 405430 255264
rect 407390 255252 407396 255264
rect 405424 255224 407396 255252
rect 405424 255212 405430 255224
rect 407390 255212 407396 255224
rect 407448 255212 407454 255264
rect 46382 254328 46388 254380
rect 46440 254368 46446 254380
rect 46566 254368 46572 254380
rect 46440 254340 46572 254368
rect 46440 254328 46446 254340
rect 46566 254328 46572 254340
rect 46624 254328 46630 254380
rect 552934 253988 552940 254040
rect 552992 254028 552998 254040
rect 564710 254028 564716 254040
rect 552992 254000 564716 254028
rect 552992 253988 552998 254000
rect 564710 253988 564716 254000
rect 564768 253988 564774 254040
rect 35066 253920 35072 253972
rect 35124 253960 35130 253972
rect 46566 253960 46572 253972
rect 35124 253932 46572 253960
rect 35124 253920 35130 253932
rect 46566 253920 46572 253932
rect 46624 253920 46630 253972
rect 350442 253920 350448 253972
rect 350500 253960 350506 253972
rect 355134 253960 355140 253972
rect 350500 253932 355140 253960
rect 350500 253920 350506 253932
rect 355134 253920 355140 253932
rect 355192 253920 355198 253972
rect 391290 253920 391296 253972
rect 391348 253960 391354 253972
rect 407114 253960 407120 253972
rect 391348 253932 407120 253960
rect 391348 253920 391354 253932
rect 407114 253920 407120 253932
rect 407172 253920 407178 253972
rect 553118 253920 553124 253972
rect 553176 253960 553182 253972
rect 570414 253960 570420 253972
rect 553176 253932 570420 253960
rect 553176 253920 553182 253932
rect 570414 253920 570420 253932
rect 570472 253920 570478 253972
rect 553118 252560 553124 252612
rect 553176 252600 553182 252612
rect 569310 252600 569316 252612
rect 553176 252572 569316 252600
rect 553176 252560 553182 252572
rect 569310 252560 569316 252572
rect 569368 252560 569374 252612
rect 403986 251200 403992 251252
rect 404044 251240 404050 251252
rect 407206 251240 407212 251252
rect 404044 251212 407212 251240
rect 404044 251200 404050 251212
rect 407206 251200 407212 251212
rect 407264 251200 407270 251252
rect 553118 251200 553124 251252
rect 553176 251240 553182 251252
rect 573542 251240 573548 251252
rect 553176 251212 573548 251240
rect 553176 251200 553182 251212
rect 573542 251200 573548 251212
rect 573600 251200 573606 251252
rect 400122 251132 400128 251184
rect 400180 251172 400186 251184
rect 407114 251172 407120 251184
rect 400180 251144 407120 251172
rect 400180 251132 400186 251144
rect 407114 251132 407120 251144
rect 407172 251132 407178 251184
rect 405366 251064 405372 251116
rect 405424 251104 405430 251116
rect 408494 251104 408500 251116
rect 405424 251076 408500 251104
rect 405424 251064 405430 251076
rect 408494 251064 408500 251076
rect 408552 251064 408558 251116
rect 361114 249840 361120 249892
rect 361172 249880 361178 249892
rect 407206 249880 407212 249892
rect 361172 249852 407212 249880
rect 361172 249840 361178 249852
rect 407206 249840 407212 249852
rect 407264 249840 407270 249892
rect 350442 249772 350448 249824
rect 350500 249812 350506 249824
rect 397914 249812 397920 249824
rect 350500 249784 397920 249812
rect 350500 249772 350506 249784
rect 397914 249772 397920 249784
rect 397972 249772 397978 249824
rect 552934 249772 552940 249824
rect 552992 249812 552998 249824
rect 568022 249812 568028 249824
rect 552992 249784 568028 249812
rect 552992 249772 552998 249784
rect 568022 249772 568028 249784
rect 568080 249772 568086 249824
rect 348786 249704 348792 249756
rect 348844 249744 348850 249756
rect 349338 249744 349344 249756
rect 348844 249716 349344 249744
rect 348844 249704 348850 249716
rect 349338 249704 349344 249716
rect 349396 249704 349402 249756
rect 553118 249704 553124 249756
rect 553176 249744 553182 249756
rect 567194 249744 567200 249756
rect 553176 249716 567200 249744
rect 553176 249704 553182 249716
rect 567194 249704 567200 249716
rect 567252 249704 567258 249756
rect 34974 249024 34980 249076
rect 35032 249064 35038 249076
rect 46290 249064 46296 249076
rect 35032 249036 46296 249064
rect 35032 249024 35038 249036
rect 46290 249024 46296 249036
rect 46348 249024 46354 249076
rect 350442 248412 350448 248464
rect 350500 248452 350506 248464
rect 400122 248452 400128 248464
rect 350500 248424 400128 248452
rect 350500 248412 350506 248424
rect 400122 248412 400128 248424
rect 400180 248412 400186 248464
rect 350074 248344 350080 248396
rect 350132 248384 350138 248396
rect 355042 248384 355048 248396
rect 350132 248356 355048 248384
rect 350132 248344 350138 248356
rect 355042 248344 355048 248356
rect 355100 248344 355106 248396
rect 563698 247664 563704 247716
rect 563756 247704 563762 247716
rect 575014 247704 575020 247716
rect 563756 247676 575020 247704
rect 563756 247664 563762 247676
rect 575014 247664 575020 247676
rect 575072 247664 575078 247716
rect 45370 247256 45376 247308
rect 45428 247296 45434 247308
rect 46566 247296 46572 247308
rect 45428 247268 46572 247296
rect 45428 247256 45434 247268
rect 46566 247256 46572 247268
rect 46624 247256 46630 247308
rect 45094 247120 45100 247172
rect 45152 247160 45158 247172
rect 45830 247160 45836 247172
rect 45152 247132 45836 247160
rect 45152 247120 45158 247132
rect 45830 247120 45836 247132
rect 45888 247120 45894 247172
rect 553118 247120 553124 247172
rect 553176 247160 553182 247172
rect 562410 247160 562416 247172
rect 553176 247132 562416 247160
rect 553176 247120 553182 247132
rect 562410 247120 562416 247132
rect 562468 247120 562474 247172
rect 36354 247052 36360 247104
rect 36412 247092 36418 247104
rect 46750 247092 46756 247104
rect 36412 247064 46756 247092
rect 36412 247052 36418 247064
rect 46750 247052 46756 247064
rect 46808 247052 46814 247104
rect 348602 247052 348608 247104
rect 348660 247092 348666 247104
rect 352190 247092 352196 247104
rect 348660 247064 352196 247092
rect 348660 247052 348666 247064
rect 352190 247052 352196 247064
rect 352248 247052 352254 247104
rect 352558 247052 352564 247104
rect 352616 247092 352622 247104
rect 353386 247092 353392 247104
rect 352616 247064 353392 247092
rect 352616 247052 352622 247064
rect 353386 247052 353392 247064
rect 353444 247052 353450 247104
rect 395890 246304 395896 246356
rect 395948 246344 395954 246356
rect 406838 246344 406844 246356
rect 395948 246316 406844 246344
rect 395948 246304 395954 246316
rect 406838 246304 406844 246316
rect 406896 246304 406902 246356
rect 357710 245800 357716 245812
rect 355704 245772 357716 245800
rect 350442 245692 350448 245744
rect 350500 245732 350506 245744
rect 355704 245732 355732 245772
rect 357710 245760 357716 245772
rect 357768 245760 357774 245812
rect 404998 245760 405004 245812
rect 405056 245800 405062 245812
rect 406378 245800 406384 245812
rect 405056 245772 406384 245800
rect 405056 245760 405062 245772
rect 406378 245760 406384 245772
rect 406436 245760 406442 245812
rect 363230 245732 363236 245744
rect 350500 245704 355732 245732
rect 355796 245704 363236 245732
rect 350500 245692 350506 245704
rect 350350 245624 350356 245676
rect 350408 245664 350414 245676
rect 355796 245664 355824 245704
rect 363230 245692 363236 245704
rect 363288 245692 363294 245744
rect 399662 245692 399668 245744
rect 399720 245732 399726 245744
rect 407206 245732 407212 245744
rect 399720 245704 407212 245732
rect 399720 245692 399726 245704
rect 407206 245692 407212 245704
rect 407264 245692 407270 245744
rect 350408 245636 355824 245664
rect 350408 245624 350414 245636
rect 355870 245624 355876 245676
rect 355928 245664 355934 245676
rect 359274 245664 359280 245676
rect 355928 245636 359280 245664
rect 355928 245624 355934 245636
rect 359274 245624 359280 245636
rect 359332 245624 359338 245676
rect 395338 245624 395344 245676
rect 395396 245664 395402 245676
rect 407114 245664 407120 245676
rect 395396 245636 407120 245664
rect 395396 245624 395402 245636
rect 407114 245624 407120 245636
rect 407172 245624 407178 245676
rect 553118 245624 553124 245676
rect 553176 245664 553182 245676
rect 563698 245664 563704 245676
rect 553176 245636 563704 245664
rect 553176 245624 553182 245636
rect 563698 245624 563704 245636
rect 563756 245624 563762 245676
rect 348878 244876 348884 244928
rect 348936 244916 348942 244928
rect 359274 244916 359280 244928
rect 348936 244888 359280 244916
rect 348936 244876 348942 244888
rect 359274 244876 359280 244888
rect 359332 244876 359338 244928
rect 402606 244876 402612 244928
rect 402664 244916 402670 244928
rect 407206 244916 407212 244928
rect 402664 244888 407212 244916
rect 402664 244876 402670 244888
rect 407206 244876 407212 244888
rect 407264 244876 407270 244928
rect 350166 244604 350172 244656
rect 350224 244644 350230 244656
rect 352190 244644 352196 244656
rect 350224 244616 352196 244644
rect 350224 244604 350230 244616
rect 352190 244604 352196 244616
rect 352248 244604 352254 244656
rect 392394 244264 392400 244316
rect 392452 244304 392458 244316
rect 407114 244304 407120 244316
rect 392452 244276 407120 244304
rect 392452 244264 392458 244276
rect 407114 244264 407120 244276
rect 407172 244264 407178 244316
rect 553118 244264 553124 244316
rect 553176 244304 553182 244316
rect 583662 244304 583668 244316
rect 553176 244276 583668 244304
rect 553176 244264 553182 244276
rect 583662 244264 583668 244276
rect 583720 244264 583726 244316
rect 550174 243924 550180 243976
rect 550232 243964 550238 243976
rect 550542 243964 550548 243976
rect 550232 243936 550548 243964
rect 550232 243924 550238 243936
rect 550542 243924 550548 243936
rect 550600 243924 550606 243976
rect 31018 242904 31024 242956
rect 31076 242944 31082 242956
rect 45830 242944 45836 242956
rect 31076 242916 45836 242944
rect 31076 242904 31082 242916
rect 45830 242904 45836 242916
rect 45888 242904 45894 242956
rect 350442 242904 350448 242956
rect 350500 242944 350506 242956
rect 396718 242944 396724 242956
rect 350500 242916 396724 242944
rect 350500 242904 350506 242916
rect 396718 242904 396724 242916
rect 396776 242904 396782 242956
rect 390186 242836 390192 242888
rect 390244 242876 390250 242888
rect 407114 242876 407120 242888
rect 390244 242848 407120 242876
rect 390244 242836 390250 242848
rect 407114 242836 407120 242848
rect 407172 242836 407178 242888
rect 36630 242156 36636 242208
rect 36688 242196 36694 242208
rect 47118 242196 47124 242208
rect 36688 242168 47124 242196
rect 36688 242156 36694 242168
rect 47118 242156 47124 242168
rect 47176 242156 47182 242208
rect 387242 241272 387248 241324
rect 387300 241312 387306 241324
rect 581546 241312 581552 241324
rect 387300 241284 581552 241312
rect 387300 241272 387306 241284
rect 581546 241272 581552 241284
rect 581604 241272 581610 241324
rect 390002 241204 390008 241256
rect 390060 241244 390066 241256
rect 563882 241244 563888 241256
rect 390060 241216 563888 241244
rect 390060 241204 390066 241216
rect 563882 241204 563888 241216
rect 563940 241204 563946 241256
rect 409506 241136 409512 241188
rect 409564 241176 409570 241188
rect 571610 241176 571616 241188
rect 409564 241148 571616 241176
rect 409564 241136 409570 241148
rect 571610 241136 571616 241148
rect 571668 241136 571674 241188
rect 562318 240836 562324 240848
rect 547846 240808 562324 240836
rect 384942 240728 384948 240780
rect 385000 240768 385006 240780
rect 385000 240740 410288 240768
rect 385000 240728 385006 240740
rect 410260 240644 410288 240740
rect 409506 240592 409512 240644
rect 409564 240632 409570 240644
rect 410150 240632 410156 240644
rect 409564 240604 410156 240632
rect 409564 240592 409570 240604
rect 410150 240592 410156 240604
rect 410208 240592 410214 240644
rect 410242 240592 410248 240644
rect 410300 240592 410306 240644
rect 547322 240592 547328 240644
rect 547380 240632 547386 240644
rect 547846 240632 547874 240808
rect 562318 240796 562324 240808
rect 562376 240796 562382 240848
rect 574646 240768 574652 240780
rect 557506 240740 574652 240768
rect 547380 240604 547874 240632
rect 547380 240592 547386 240604
rect 548702 240592 548708 240644
rect 548760 240632 548766 240644
rect 557506 240632 557534 240740
rect 574646 240728 574652 240740
rect 574704 240728 574710 240780
rect 548760 240604 557534 240632
rect 548760 240592 548766 240604
rect 409230 240524 409236 240576
rect 409288 240564 409294 240576
rect 412266 240564 412272 240576
rect 409288 240536 412272 240564
rect 409288 240524 409294 240536
rect 412266 240524 412272 240536
rect 412324 240524 412330 240576
rect 404078 240456 404084 240508
rect 404136 240496 404142 240508
rect 410794 240496 410800 240508
rect 404136 240468 410800 240496
rect 404136 240456 404142 240468
rect 410794 240456 410800 240468
rect 410852 240456 410858 240508
rect 549990 240320 549996 240372
rect 550048 240360 550054 240372
rect 552382 240360 552388 240372
rect 550048 240332 552388 240360
rect 550048 240320 550054 240332
rect 552382 240320 552388 240332
rect 552440 240320 552446 240372
rect 544286 240184 544292 240236
rect 544344 240224 544350 240236
rect 544746 240224 544752 240236
rect 544344 240196 544752 240224
rect 544344 240184 544350 240196
rect 544746 240184 544752 240196
rect 544804 240184 544810 240236
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 30834 240156 30840 240168
rect 3108 240128 30840 240156
rect 3108 240116 3114 240128
rect 30834 240116 30840 240128
rect 30892 240116 30898 240168
rect 549530 240116 549536 240168
rect 549588 240156 549594 240168
rect 550082 240156 550088 240168
rect 549588 240128 550088 240156
rect 549588 240116 549594 240128
rect 550082 240116 550088 240128
rect 550140 240116 550146 240168
rect 365622 240048 365628 240100
rect 365680 240088 365686 240100
rect 577590 240088 577596 240100
rect 365680 240060 577596 240088
rect 365680 240048 365686 240060
rect 577590 240048 577596 240060
rect 577648 240048 577654 240100
rect 373810 239980 373816 240032
rect 373868 240020 373874 240032
rect 567746 240020 567752 240032
rect 373868 239992 567752 240020
rect 373868 239980 373874 239992
rect 567746 239980 567752 239992
rect 567804 239980 567810 240032
rect 406746 239912 406752 239964
rect 406804 239952 406810 239964
rect 580534 239952 580540 239964
rect 406804 239924 580540 239952
rect 406804 239912 406810 239924
rect 580534 239912 580540 239924
rect 580592 239912 580598 239964
rect 394510 239844 394516 239896
rect 394568 239884 394574 239896
rect 564802 239884 564808 239896
rect 394568 239856 564808 239884
rect 394568 239844 394574 239856
rect 564802 239844 564808 239856
rect 564860 239844 564866 239896
rect 405642 239776 405648 239828
rect 405700 239816 405706 239828
rect 573358 239816 573364 239828
rect 405700 239788 573364 239816
rect 405700 239776 405706 239788
rect 573358 239776 573364 239788
rect 573416 239776 573422 239828
rect 400122 239708 400128 239760
rect 400180 239748 400186 239760
rect 567654 239748 567660 239760
rect 400180 239720 567660 239748
rect 400180 239708 400186 239720
rect 567654 239708 567660 239720
rect 567712 239708 567718 239760
rect 402606 239640 402612 239692
rect 402664 239680 402670 239692
rect 564894 239680 564900 239692
rect 402664 239652 564900 239680
rect 402664 239640 402670 239652
rect 564894 239640 564900 239652
rect 564952 239640 564958 239692
rect 392946 239572 392952 239624
rect 393004 239612 393010 239624
rect 548702 239612 548708 239624
rect 393004 239584 548708 239612
rect 393004 239572 393010 239584
rect 548702 239572 548708 239584
rect 548760 239572 548766 239624
rect 549898 239504 549904 239556
rect 549956 239544 549962 239556
rect 564434 239544 564440 239556
rect 549956 239516 564440 239544
rect 549956 239504 549962 239516
rect 564434 239504 564440 239516
rect 564492 239504 564498 239556
rect 406194 239436 406200 239488
rect 406252 239476 406258 239488
rect 551094 239476 551100 239488
rect 406252 239448 551100 239476
rect 406252 239436 406258 239448
rect 551094 239436 551100 239448
rect 551152 239436 551158 239488
rect 35802 239368 35808 239420
rect 35860 239408 35866 239420
rect 45646 239408 45652 239420
rect 35860 239380 45652 239408
rect 35860 239368 35866 239380
rect 45646 239368 45652 239380
rect 45704 239368 45710 239420
rect 406838 239368 406844 239420
rect 406896 239408 406902 239420
rect 549990 239408 549996 239420
rect 406896 239380 549996 239408
rect 406896 239368 406902 239380
rect 549990 239368 549996 239380
rect 550048 239368 550054 239420
rect 551462 239368 551468 239420
rect 551520 239408 551526 239420
rect 560294 239408 560300 239420
rect 551520 239380 560300 239408
rect 551520 239368 551526 239380
rect 560294 239368 560300 239380
rect 560352 239368 560358 239420
rect 532050 239300 532056 239352
rect 532108 239340 532114 239352
rect 554038 239340 554044 239352
rect 532108 239312 554044 239340
rect 532108 239300 532114 239312
rect 554038 239300 554044 239312
rect 554096 239300 554102 239352
rect 396626 239232 396632 239284
rect 396684 239272 396690 239284
rect 550174 239272 550180 239284
rect 396684 239244 550180 239272
rect 396684 239232 396690 239244
rect 550174 239232 550180 239244
rect 550232 239232 550238 239284
rect 350350 238892 350356 238944
rect 350408 238932 350414 238944
rect 499850 238932 499856 238944
rect 350408 238904 499856 238932
rect 350408 238892 350414 238904
rect 499850 238892 499856 238904
rect 499908 238892 499914 238944
rect 505646 238892 505652 238944
rect 505704 238932 505710 238944
rect 570782 238932 570788 238944
rect 505704 238904 570788 238932
rect 505704 238892 505710 238904
rect 570782 238892 570788 238904
rect 570840 238892 570846 238944
rect 350442 238824 350448 238876
rect 350500 238864 350506 238876
rect 392302 238864 392308 238876
rect 350500 238836 392308 238864
rect 350500 238824 350506 238836
rect 392302 238824 392308 238836
rect 392360 238824 392366 238876
rect 447042 238824 447048 238876
rect 447100 238864 447106 238876
rect 551186 238864 551192 238876
rect 447100 238836 551192 238864
rect 447100 238824 447106 238836
rect 551186 238824 551192 238836
rect 551244 238824 551250 238876
rect 381538 238756 381544 238808
rect 381596 238796 381602 238808
rect 509234 238796 509240 238808
rect 381596 238768 509240 238796
rect 381596 238756 381602 238768
rect 509234 238756 509240 238768
rect 509292 238756 509298 238808
rect 35342 238688 35348 238740
rect 35400 238728 35406 238740
rect 46842 238728 46848 238740
rect 35400 238700 46848 238728
rect 35400 238688 35406 238700
rect 46842 238688 46848 238700
rect 46900 238688 46906 238740
rect 400858 238688 400864 238740
rect 400916 238728 400922 238740
rect 427814 238728 427820 238740
rect 400916 238700 427820 238728
rect 400916 238688 400922 238700
rect 427814 238688 427820 238700
rect 427872 238688 427878 238740
rect 403710 238620 403716 238672
rect 403768 238660 403774 238672
rect 440234 238660 440240 238672
rect 403768 238632 440240 238660
rect 403768 238620 403774 238632
rect 440234 238620 440240 238632
rect 440292 238620 440298 238672
rect 445110 238620 445116 238672
rect 445168 238660 445174 238672
rect 570322 238660 570328 238672
rect 445168 238632 570328 238660
rect 445168 238620 445174 238632
rect 570322 238620 570328 238632
rect 570380 238620 570386 238672
rect 399294 238552 399300 238604
rect 399352 238592 399358 238604
rect 428366 238592 428372 238604
rect 399352 238564 428372 238592
rect 399352 238552 399358 238564
rect 428366 238552 428372 238564
rect 428424 238552 428430 238604
rect 436738 238552 436744 238604
rect 436796 238592 436802 238604
rect 559558 238592 559564 238604
rect 436796 238564 559564 238592
rect 436796 238552 436802 238564
rect 559558 238552 559564 238564
rect 559616 238552 559622 238604
rect 408954 238484 408960 238536
rect 409012 238524 409018 238536
rect 504358 238524 504364 238536
rect 409012 238496 504364 238524
rect 409012 238484 409018 238496
rect 504358 238484 504364 238496
rect 504416 238484 504422 238536
rect 506658 238484 506664 238536
rect 506716 238524 506722 238536
rect 555326 238524 555332 238536
rect 506716 238496 555332 238524
rect 506716 238484 506722 238496
rect 555326 238484 555332 238496
rect 555384 238484 555390 238536
rect 405550 238416 405556 238468
rect 405608 238456 405614 238468
rect 514754 238456 514760 238468
rect 405608 238428 514760 238456
rect 405608 238416 405614 238428
rect 514754 238416 514760 238428
rect 514812 238416 514818 238468
rect 535270 238416 535276 238468
rect 535328 238456 535334 238468
rect 550634 238456 550640 238468
rect 535328 238428 550640 238456
rect 535328 238416 535334 238428
rect 550634 238416 550640 238428
rect 550692 238416 550698 238468
rect 497918 238348 497924 238400
rect 497976 238388 497982 238400
rect 557994 238388 558000 238400
rect 497976 238360 558000 238388
rect 497976 238348 497982 238360
rect 557994 238348 558000 238360
rect 558052 238348 558058 238400
rect 403434 238280 403440 238332
rect 403492 238320 403498 238332
rect 463142 238320 463148 238332
rect 403492 238292 463148 238320
rect 403492 238280 403498 238292
rect 463142 238280 463148 238292
rect 463200 238280 463206 238332
rect 472618 238280 472624 238332
rect 472676 238320 472682 238332
rect 551370 238320 551376 238332
rect 472676 238292 551376 238320
rect 472676 238280 472682 238292
rect 551370 238280 551376 238292
rect 551428 238280 551434 238332
rect 409138 238212 409144 238264
rect 409196 238252 409202 238264
rect 442534 238252 442540 238264
rect 409196 238224 442540 238252
rect 409196 238212 409202 238224
rect 442534 238212 442540 238224
rect 442592 238212 442598 238264
rect 476390 238212 476396 238264
rect 476448 238252 476454 238264
rect 554774 238252 554780 238264
rect 476448 238224 554780 238252
rect 476448 238212 476454 238224
rect 554774 238212 554780 238224
rect 554832 238212 554838 238264
rect 569218 238212 569224 238264
rect 569276 238252 569282 238264
rect 570322 238252 570328 238264
rect 569276 238224 570328 238252
rect 569276 238212 569282 238224
rect 570322 238212 570328 238224
rect 570380 238212 570386 238264
rect 400030 238144 400036 238196
rect 400088 238184 400094 238196
rect 432230 238184 432236 238196
rect 400088 238156 432236 238184
rect 400088 238144 400094 238156
rect 432230 238144 432236 238156
rect 432288 238144 432294 238196
rect 475378 238144 475384 238196
rect 475436 238184 475442 238196
rect 571610 238184 571616 238196
rect 475436 238156 571616 238184
rect 475436 238144 475442 238156
rect 571610 238144 571616 238156
rect 571668 238144 571674 238196
rect 355318 238076 355324 238128
rect 355376 238116 355382 238128
rect 416682 238116 416688 238128
rect 355376 238088 416688 238116
rect 355376 238076 355382 238088
rect 416682 238076 416688 238088
rect 416740 238076 416746 238128
rect 421282 238076 421288 238128
rect 421340 238116 421346 238128
rect 547506 238116 547512 238128
rect 421340 238088 547512 238116
rect 421340 238076 421346 238088
rect 547506 238076 547512 238088
rect 547564 238076 547570 238128
rect 554038 238076 554044 238128
rect 554096 238116 554102 238128
rect 561030 238116 561036 238128
rect 554096 238088 561036 238116
rect 554096 238076 554102 238088
rect 561030 238076 561036 238088
rect 561088 238076 561094 238128
rect 349890 238008 349896 238060
rect 349948 238048 349954 238060
rect 540422 238048 540428 238060
rect 349948 238020 540428 238048
rect 349948 238008 349954 238020
rect 540422 238008 540428 238020
rect 540480 238008 540486 238060
rect 548058 238008 548064 238060
rect 548116 238048 548122 238060
rect 557994 238048 558000 238060
rect 548116 238020 558000 238048
rect 548116 238008 548122 238020
rect 557994 238008 558000 238020
rect 558052 238008 558058 238060
rect 416682 237940 416688 237992
rect 416740 237980 416746 237992
rect 490558 237980 490564 237992
rect 416740 237952 490564 237980
rect 416740 237940 416746 237952
rect 490558 237940 490564 237952
rect 490616 237980 490622 237992
rect 491110 237980 491116 237992
rect 490616 237952 491116 237980
rect 490616 237940 490622 237952
rect 491110 237940 491116 237952
rect 491168 237940 491174 237992
rect 501782 237940 501788 237992
rect 501840 237980 501846 237992
rect 547598 237980 547604 237992
rect 501840 237952 547604 237980
rect 501840 237940 501846 237952
rect 547598 237940 547604 237952
rect 547656 237940 547662 237992
rect 372062 237872 372068 237924
rect 372120 237912 372126 237924
rect 422846 237912 422852 237924
rect 372120 237884 422852 237912
rect 372120 237872 372126 237884
rect 422846 237872 422852 237884
rect 422904 237912 422910 237924
rect 482922 237912 482928 237924
rect 422904 237884 482928 237912
rect 422904 237872 422910 237884
rect 482922 237872 482928 237884
rect 482980 237872 482986 237924
rect 528186 237872 528192 237924
rect 528244 237912 528250 237924
rect 544838 237912 544844 237924
rect 528244 237884 544844 237912
rect 528244 237872 528250 237884
rect 544838 237872 544844 237884
rect 544896 237872 544902 237924
rect 545850 237872 545856 237924
rect 545908 237912 545914 237924
rect 552106 237912 552112 237924
rect 545908 237884 552112 237912
rect 545908 237872 545914 237884
rect 552106 237872 552112 237884
rect 552164 237872 552170 237924
rect 396810 237804 396816 237856
rect 396868 237844 396874 237856
rect 515306 237844 515312 237856
rect 396868 237816 515312 237844
rect 396868 237804 396874 237816
rect 515306 237804 515312 237816
rect 515364 237804 515370 237856
rect 529842 237804 529848 237856
rect 529900 237844 529906 237856
rect 545666 237844 545672 237856
rect 529900 237816 545672 237844
rect 529900 237804 529906 237816
rect 545666 237804 545672 237816
rect 545724 237804 545730 237856
rect 382826 237668 382832 237720
rect 382884 237708 382890 237720
rect 567562 237708 567568 237720
rect 382884 237680 567568 237708
rect 382884 237668 382890 237680
rect 567562 237668 567568 237680
rect 567620 237668 567626 237720
rect 542078 237464 542084 237516
rect 542136 237504 542142 237516
rect 549622 237504 549628 237516
rect 542136 237476 549628 237504
rect 542136 237464 542142 237476
rect 549622 237464 549628 237476
rect 549680 237464 549686 237516
rect 32766 237396 32772 237448
rect 32824 237436 32830 237448
rect 46842 237436 46848 237448
rect 32824 237408 46848 237436
rect 32824 237396 32830 237408
rect 46842 237396 46848 237408
rect 46900 237396 46906 237448
rect 482922 237396 482928 237448
rect 482980 237436 482986 237448
rect 483750 237436 483756 237448
rect 482980 237408 483756 237436
rect 482980 237396 482986 237408
rect 483750 237396 483756 237408
rect 483808 237396 483814 237448
rect 545758 237396 545764 237448
rect 545816 237436 545822 237448
rect 548794 237436 548800 237448
rect 545816 237408 548800 237436
rect 545816 237396 545822 237408
rect 548794 237396 548800 237408
rect 548852 237396 548858 237448
rect 363782 237328 363788 237380
rect 363840 237368 363846 237380
rect 552014 237368 552020 237380
rect 363840 237340 552020 237368
rect 363840 237328 363846 237340
rect 552014 237328 552020 237340
rect 552072 237328 552078 237380
rect 350442 237260 350448 237312
rect 350500 237300 350506 237312
rect 376662 237300 376668 237312
rect 350500 237272 376668 237300
rect 350500 237260 350506 237272
rect 376662 237260 376668 237272
rect 376720 237260 376726 237312
rect 391750 237260 391756 237312
rect 391808 237300 391814 237312
rect 578694 237300 578700 237312
rect 391808 237272 578700 237300
rect 391808 237260 391814 237272
rect 578694 237260 578700 237272
rect 578752 237260 578758 237312
rect 394326 237192 394332 237244
rect 394384 237232 394390 237244
rect 574554 237232 574560 237244
rect 394384 237204 574560 237232
rect 394384 237192 394390 237204
rect 574554 237192 574560 237204
rect 574612 237192 574618 237244
rect 406562 237124 406568 237176
rect 406620 237164 406626 237176
rect 580074 237164 580080 237176
rect 406620 237136 580080 237164
rect 406620 237124 406626 237136
rect 580074 237124 580080 237136
rect 580132 237124 580138 237176
rect 391566 237056 391572 237108
rect 391624 237096 391630 237108
rect 563606 237096 563612 237108
rect 391624 237068 563612 237096
rect 391624 237056 391630 237068
rect 563606 237056 563612 237068
rect 563664 237056 563670 237108
rect 402054 236988 402060 237040
rect 402112 237028 402118 237040
rect 573450 237028 573456 237040
rect 402112 237000 573456 237028
rect 402112 236988 402118 237000
rect 573450 236988 573456 237000
rect 573508 236988 573514 237040
rect 395706 236920 395712 236972
rect 395764 236960 395770 236972
rect 566274 236960 566280 236972
rect 395764 236932 566280 236960
rect 395764 236920 395770 236932
rect 566274 236920 566280 236932
rect 566332 236920 566338 236972
rect 381998 236852 382004 236904
rect 382056 236892 382062 236904
rect 550910 236892 550916 236904
rect 382056 236864 550916 236892
rect 382056 236852 382062 236864
rect 550910 236852 550916 236864
rect 550968 236852 550974 236904
rect 386874 236784 386880 236836
rect 386932 236824 386938 236836
rect 545574 236824 545580 236836
rect 386932 236796 545580 236824
rect 386932 236784 386938 236796
rect 545574 236784 545580 236796
rect 545632 236784 545638 236836
rect 386138 236716 386144 236768
rect 386196 236756 386202 236768
rect 532694 236756 532700 236768
rect 386196 236728 532700 236756
rect 386196 236716 386202 236728
rect 532694 236716 532700 236728
rect 532752 236716 532758 236768
rect 45370 236648 45376 236700
rect 45428 236688 45434 236700
rect 46934 236688 46940 236700
rect 45428 236660 46940 236688
rect 45428 236648 45434 236660
rect 46934 236648 46940 236660
rect 46992 236648 46998 236700
rect 417418 236648 417424 236700
rect 417476 236688 417482 236700
rect 553486 236688 553492 236700
rect 417476 236660 553492 236688
rect 417476 236648 417482 236660
rect 553486 236648 553492 236660
rect 553544 236648 553550 236700
rect 409322 236580 409328 236632
rect 409380 236620 409386 236632
rect 419350 236620 419356 236632
rect 409380 236592 419356 236620
rect 409380 236580 409386 236592
rect 419350 236580 419356 236592
rect 419408 236580 419414 236632
rect 430298 236580 430304 236632
rect 430356 236620 430362 236632
rect 556798 236620 556804 236632
rect 430356 236592 556804 236620
rect 430356 236580 430362 236592
rect 556798 236580 556804 236592
rect 556856 236580 556862 236632
rect 374822 236512 374828 236564
rect 374880 236552 374886 236564
rect 454126 236552 454132 236564
rect 374880 236524 454132 236552
rect 374880 236512 374886 236524
rect 454126 236512 454132 236524
rect 454184 236512 454190 236564
rect 478598 236512 478604 236564
rect 478656 236552 478662 236564
rect 556614 236552 556620 236564
rect 478656 236524 556620 236552
rect 478656 236512 478662 236524
rect 556614 236512 556620 236524
rect 556672 236512 556678 236564
rect 499206 236444 499212 236496
rect 499264 236484 499270 236496
rect 571794 236484 571800 236496
rect 499264 236456 571800 236484
rect 499264 236444 499270 236456
rect 571794 236444 571800 236456
rect 571852 236444 571858 236496
rect 349890 235968 349896 236020
rect 349948 236008 349954 236020
rect 350810 236008 350816 236020
rect 349948 235980 350816 236008
rect 349948 235968 349954 235980
rect 350810 235968 350816 235980
rect 350868 235968 350874 236020
rect 481542 235900 481548 235952
rect 481600 235940 481606 235952
rect 564894 235940 564900 235952
rect 481600 235912 564900 235940
rect 481600 235900 481606 235912
rect 564894 235900 564900 235912
rect 564952 235900 564958 235952
rect 461210 235832 461216 235884
rect 461268 235872 461274 235884
rect 550542 235872 550548 235884
rect 461268 235844 550548 235872
rect 461268 235832 461274 235844
rect 550542 235832 550548 235844
rect 550600 235832 550606 235884
rect 474642 235764 474648 235816
rect 474700 235804 474706 235816
rect 568758 235804 568764 235816
rect 474700 235776 568764 235804
rect 474700 235764 474706 235776
rect 568758 235764 568764 235776
rect 568816 235764 568822 235816
rect 460934 235696 460940 235748
rect 460992 235736 460998 235748
rect 564802 235736 564808 235748
rect 460992 235708 564808 235736
rect 460992 235696 460998 235708
rect 564802 235696 564808 235708
rect 564860 235696 564866 235748
rect 452562 235628 452568 235680
rect 452620 235668 452626 235680
rect 563606 235668 563612 235680
rect 452620 235640 563612 235668
rect 452620 235628 452626 235640
rect 563606 235628 563612 235640
rect 563664 235628 563670 235680
rect 393866 235560 393872 235612
rect 393924 235600 393930 235612
rect 511442 235600 511448 235612
rect 393924 235572 511448 235600
rect 393924 235560 393930 235572
rect 511442 235560 511448 235572
rect 511500 235560 511506 235612
rect 456702 235492 456708 235544
rect 456760 235532 456766 235544
rect 573358 235532 573364 235544
rect 456760 235504 573364 235532
rect 456760 235492 456766 235504
rect 573358 235492 573364 235504
rect 573416 235492 573422 235544
rect 385586 235424 385592 235476
rect 385644 235464 385650 235476
rect 551370 235464 551376 235476
rect 385644 235436 551376 235464
rect 385644 235424 385650 235436
rect 551370 235424 551376 235436
rect 551428 235424 551434 235476
rect 385034 235356 385040 235408
rect 385092 235396 385098 235408
rect 554222 235396 554228 235408
rect 385092 235368 554228 235396
rect 385092 235356 385098 235368
rect 554222 235356 554228 235368
rect 554280 235356 554286 235408
rect 378134 235288 378140 235340
rect 378192 235328 378198 235340
rect 558086 235328 558092 235340
rect 378192 235300 558092 235328
rect 378192 235288 378198 235300
rect 558086 235288 558092 235300
rect 558144 235288 558150 235340
rect 567654 235288 567660 235340
rect 567712 235328 567718 235340
rect 569034 235328 569040 235340
rect 567712 235300 569040 235328
rect 567712 235288 567718 235300
rect 569034 235288 569040 235300
rect 569092 235288 569098 235340
rect 350166 235220 350172 235272
rect 350224 235260 350230 235272
rect 541066 235260 541072 235272
rect 350224 235232 541072 235260
rect 350224 235220 350230 235232
rect 541066 235220 541072 235232
rect 541124 235220 541130 235272
rect 409414 235152 409420 235204
rect 409472 235192 409478 235204
rect 491294 235192 491300 235204
rect 409472 235164 491300 235192
rect 409472 235152 409478 235164
rect 491294 235152 491300 235164
rect 491352 235152 491358 235204
rect 491110 235084 491116 235136
rect 491168 235124 491174 235136
rect 562318 235124 562324 235136
rect 491168 235096 562324 235124
rect 491168 235084 491174 235096
rect 562318 235084 562324 235096
rect 562376 235084 562382 235136
rect 491202 235016 491208 235068
rect 491260 235056 491266 235068
rect 552750 235056 552756 235068
rect 491260 235028 552756 235056
rect 491260 235016 491266 235028
rect 552750 235016 552756 235028
rect 552808 235016 552814 235068
rect 350442 234880 350448 234932
rect 350500 234920 350506 234932
rect 356146 234920 356152 234932
rect 350500 234892 356152 234920
rect 350500 234880 350506 234892
rect 356146 234880 356152 234892
rect 356204 234880 356210 234932
rect 355502 234676 355508 234728
rect 355560 234716 355566 234728
rect 363414 234716 363420 234728
rect 355560 234688 363420 234716
rect 355560 234676 355566 234688
rect 363414 234676 363420 234688
rect 363472 234676 363478 234728
rect 44450 234608 44456 234660
rect 44508 234648 44514 234660
rect 45646 234648 45652 234660
rect 44508 234620 45652 234648
rect 44508 234608 44514 234620
rect 45646 234608 45652 234620
rect 45704 234608 45710 234660
rect 384758 234540 384764 234592
rect 384816 234580 384822 234592
rect 580350 234580 580356 234592
rect 384816 234552 580356 234580
rect 384816 234540 384822 234552
rect 580350 234540 580356 234552
rect 580408 234540 580414 234592
rect 395154 234472 395160 234524
rect 395212 234512 395218 234524
rect 545942 234512 545948 234524
rect 395212 234484 545948 234512
rect 395212 234472 395218 234484
rect 545942 234472 545948 234484
rect 546000 234472 546006 234524
rect 398466 234404 398472 234456
rect 398524 234444 398530 234456
rect 555602 234444 555608 234456
rect 398524 234416 555608 234444
rect 398524 234404 398530 234416
rect 555602 234404 555608 234416
rect 555660 234404 555666 234456
rect 380618 234336 380624 234388
rect 380676 234376 380682 234388
rect 540330 234376 540336 234388
rect 380676 234348 540336 234376
rect 380676 234336 380682 234348
rect 540330 234336 540336 234348
rect 540388 234336 540394 234388
rect 387702 234268 387708 234320
rect 387760 234308 387766 234320
rect 548058 234308 548064 234320
rect 387760 234280 548064 234308
rect 387760 234268 387766 234280
rect 548058 234268 548064 234280
rect 548116 234268 548122 234320
rect 395246 234200 395252 234252
rect 395304 234240 395310 234252
rect 566642 234240 566648 234252
rect 395304 234212 566648 234240
rect 395304 234200 395310 234212
rect 566642 234200 566648 234212
rect 566700 234200 566706 234252
rect 386230 234132 386236 234184
rect 386288 234172 386294 234184
rect 561030 234172 561036 234184
rect 386288 234144 561036 234172
rect 386288 234132 386294 234144
rect 561030 234132 561036 234144
rect 561088 234132 561094 234184
rect 363966 234064 363972 234116
rect 364024 234104 364030 234116
rect 544378 234104 544384 234116
rect 364024 234076 544384 234104
rect 364024 234064 364030 234076
rect 544378 234064 544384 234076
rect 544436 234064 544442 234116
rect 376754 233996 376760 234048
rect 376812 234036 376818 234048
rect 559466 234036 559472 234048
rect 376812 234008 559472 234036
rect 376812 233996 376818 234008
rect 559466 233996 559472 234008
rect 559524 233996 559530 234048
rect 355594 233928 355600 233980
rect 355652 233968 355658 233980
rect 555510 233968 555516 233980
rect 355652 233940 555516 233968
rect 355652 233928 355658 233940
rect 555510 233928 555516 233940
rect 555568 233928 555574 233980
rect 349062 233860 349068 233912
rect 349120 233900 349126 233912
rect 349430 233900 349436 233912
rect 349120 233872 349436 233900
rect 349120 233860 349126 233872
rect 349430 233860 349436 233872
rect 349488 233860 349494 233912
rect 349982 233860 349988 233912
rect 350040 233900 350046 233912
rect 580074 233900 580080 233912
rect 350040 233872 580080 233900
rect 350040 233860 350046 233872
rect 580074 233860 580080 233872
rect 580132 233860 580138 233912
rect 398006 233792 398012 233844
rect 398064 233832 398070 233844
rect 547046 233832 547052 233844
rect 398064 233804 547052 233832
rect 398064 233792 398070 233804
rect 547046 233792 547052 233804
rect 547104 233792 547110 233844
rect 349062 233724 349068 233776
rect 349120 233764 349126 233776
rect 352558 233764 352564 233776
rect 349120 233736 352564 233764
rect 349120 233724 349126 233736
rect 352558 233724 352564 233736
rect 352616 233724 352622 233776
rect 393130 233724 393136 233776
rect 393188 233764 393194 233776
rect 541618 233764 541624 233776
rect 393188 233736 541624 233764
rect 393188 233724 393194 233736
rect 541618 233724 541624 233736
rect 541676 233724 541682 233776
rect 409966 233656 409972 233708
rect 410024 233696 410030 233708
rect 410334 233696 410340 233708
rect 410024 233668 410340 233696
rect 410024 233656 410030 233668
rect 410334 233656 410340 233668
rect 410392 233656 410398 233708
rect 412634 233656 412640 233708
rect 412692 233696 412698 233708
rect 412910 233696 412916 233708
rect 412692 233668 412916 233696
rect 412692 233656 412698 233668
rect 412910 233656 412916 233668
rect 412968 233656 412974 233708
rect 418798 233656 418804 233708
rect 418856 233696 418862 233708
rect 419994 233696 420000 233708
rect 418856 233668 420000 233696
rect 418856 233656 418862 233668
rect 419994 233656 420000 233668
rect 420052 233656 420058 233708
rect 486970 233656 486976 233708
rect 487028 233696 487034 233708
rect 496814 233696 496820 233708
rect 487028 233668 496820 233696
rect 487028 233656 487034 233668
rect 496814 233656 496820 233668
rect 496872 233656 496878 233708
rect 46658 233180 46664 233232
rect 46716 233220 46722 233232
rect 47118 233220 47124 233232
rect 46716 233192 47124 233220
rect 46716 233180 46722 233192
rect 47118 233180 47124 233192
rect 47176 233180 47182 233232
rect 355870 233180 355876 233232
rect 355928 233220 355934 233232
rect 356054 233220 356060 233232
rect 355928 233192 356060 233220
rect 355928 233180 355934 233192
rect 356054 233180 356060 233192
rect 356112 233180 356118 233232
rect 406930 233180 406936 233232
rect 406988 233220 406994 233232
rect 580166 233220 580172 233232
rect 406988 233192 580172 233220
rect 406988 233180 406994 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 372430 233112 372436 233164
rect 372488 233152 372494 233164
rect 540054 233152 540060 233164
rect 372488 233124 540060 233152
rect 372488 233112 372494 233124
rect 540054 233112 540060 233124
rect 540112 233112 540118 233164
rect 378686 233044 378692 233096
rect 378744 233084 378750 233096
rect 547138 233084 547144 233096
rect 378744 233056 547144 233084
rect 378744 233044 378750 233056
rect 547138 233044 547144 233056
rect 547196 233044 547202 233096
rect 371142 232976 371148 233028
rect 371200 233016 371206 233028
rect 541710 233016 541716 233028
rect 371200 232988 541716 233016
rect 371200 232976 371206 232988
rect 541710 232976 541716 232988
rect 541768 232976 541774 233028
rect 406286 232908 406292 232960
rect 406344 232948 406350 232960
rect 578694 232948 578700 232960
rect 406344 232920 578700 232948
rect 406344 232908 406350 232920
rect 578694 232908 578700 232920
rect 578752 232908 578758 232960
rect 369210 232840 369216 232892
rect 369268 232880 369274 232892
rect 542446 232880 542452 232892
rect 369268 232852 542452 232880
rect 369268 232840 369274 232852
rect 542446 232840 542452 232852
rect 542504 232840 542510 232892
rect 374546 232772 374552 232824
rect 374604 232812 374610 232824
rect 547966 232812 547972 232824
rect 374604 232784 547972 232812
rect 374604 232772 374610 232784
rect 547966 232772 547972 232784
rect 548024 232772 548030 232824
rect 403802 232704 403808 232756
rect 403860 232744 403866 232756
rect 577682 232744 577688 232756
rect 403860 232716 577688 232744
rect 403860 232704 403866 232716
rect 577682 232704 577688 232716
rect 577740 232704 577746 232756
rect 362494 232636 362500 232688
rect 362552 232676 362558 232688
rect 540238 232676 540244 232688
rect 362552 232648 540244 232676
rect 362552 232636 362558 232648
rect 540238 232636 540244 232648
rect 540296 232636 540302 232688
rect 46842 232568 46848 232620
rect 46900 232608 46906 232620
rect 47670 232608 47676 232620
rect 46900 232580 47676 232608
rect 46900 232568 46906 232580
rect 47670 232568 47676 232580
rect 47728 232568 47734 232620
rect 365438 232568 365444 232620
rect 365496 232608 365502 232620
rect 548150 232608 548156 232620
rect 365496 232580 548156 232608
rect 365496 232568 365502 232580
rect 548150 232568 548156 232580
rect 548208 232568 548214 232620
rect 358446 232500 358452 232552
rect 358504 232540 358510 232552
rect 541894 232540 541900 232552
rect 358504 232512 541900 232540
rect 358504 232500 358510 232512
rect 541894 232500 541900 232512
rect 541952 232500 541958 232552
rect 379422 232432 379428 232484
rect 379480 232472 379486 232484
rect 471974 232472 471980 232484
rect 379480 232444 471980 232472
rect 379480 232432 379486 232444
rect 471974 232432 471980 232444
rect 472032 232432 472038 232484
rect 493410 232432 493416 232484
rect 493468 232472 493474 232484
rect 563422 232472 563428 232484
rect 493468 232444 563428 232472
rect 493468 232432 493474 232444
rect 563422 232432 563428 232444
rect 563480 232432 563486 232484
rect 408862 232364 408868 232416
rect 408920 232404 408926 232416
rect 470226 232404 470232 232416
rect 408920 232376 470232 232404
rect 408920 232364 408926 232376
rect 470226 232364 470232 232376
rect 470284 232364 470290 232416
rect 525610 232364 525616 232416
rect 525668 232404 525674 232416
rect 554958 232404 554964 232416
rect 525668 232376 554964 232404
rect 525668 232364 525674 232376
rect 554958 232364 554964 232376
rect 555016 232364 555022 232416
rect 402882 232296 402888 232348
rect 402940 232336 402946 232348
rect 416774 232336 416780 232348
rect 402940 232308 416780 232336
rect 402940 232296 402946 232308
rect 416774 232296 416780 232308
rect 416832 232296 416838 232348
rect 33594 231820 33600 231872
rect 33652 231860 33658 231872
rect 46842 231860 46848 231872
rect 33652 231832 46848 231860
rect 33652 231820 33658 231832
rect 46842 231820 46848 231832
rect 46900 231820 46906 231872
rect 350442 231820 350448 231872
rect 350500 231860 350506 231872
rect 353386 231860 353392 231872
rect 350500 231832 353392 231860
rect 350500 231820 350506 231832
rect 353386 231820 353392 231832
rect 353444 231820 353450 231872
rect 36446 231752 36452 231804
rect 36504 231792 36510 231804
rect 45462 231792 45468 231804
rect 36504 231764 45468 231792
rect 36504 231752 36510 231764
rect 45462 231752 45468 231764
rect 45520 231752 45526 231804
rect 410794 231752 410800 231804
rect 410852 231792 410858 231804
rect 538950 231792 538956 231804
rect 410852 231764 538956 231792
rect 410852 231752 410858 231764
rect 538950 231752 538956 231764
rect 539008 231752 539014 231804
rect 408218 231684 408224 231736
rect 408276 231724 408282 231736
rect 544010 231724 544016 231736
rect 408276 231696 544016 231724
rect 408276 231684 408282 231696
rect 544010 231684 544016 231696
rect 544068 231684 544074 231736
rect 407758 231616 407764 231668
rect 407816 231656 407822 231668
rect 546034 231656 546040 231668
rect 407816 231628 546040 231656
rect 407816 231616 407822 231628
rect 546034 231616 546040 231628
rect 546092 231616 546098 231668
rect 414014 231548 414020 231600
rect 414072 231588 414078 231600
rect 558362 231588 558368 231600
rect 414072 231560 558368 231588
rect 414072 231548 414078 231560
rect 558362 231548 558368 231560
rect 558420 231548 558426 231600
rect 404998 231480 405004 231532
rect 405056 231520 405062 231532
rect 549990 231520 549996 231532
rect 405056 231492 549996 231520
rect 405056 231480 405062 231492
rect 549990 231480 549996 231492
rect 550048 231480 550054 231532
rect 399386 231412 399392 231464
rect 399444 231452 399450 231464
rect 548242 231452 548248 231464
rect 399444 231424 548248 231452
rect 399444 231412 399450 231424
rect 548242 231412 548248 231424
rect 548300 231412 548306 231464
rect 402146 231344 402152 231396
rect 402204 231384 402210 231396
rect 562502 231384 562508 231396
rect 402204 231356 562508 231384
rect 402204 231344 402210 231356
rect 562502 231344 562508 231356
rect 562560 231344 562566 231396
rect 388346 231276 388352 231328
rect 388404 231316 388410 231328
rect 552842 231316 552848 231328
rect 388404 231288 552848 231316
rect 388404 231276 388410 231288
rect 552842 231276 552848 231288
rect 552900 231276 552906 231328
rect 390370 231208 390376 231260
rect 390428 231248 390434 231260
rect 563882 231248 563888 231260
rect 390428 231220 563888 231248
rect 390428 231208 390434 231220
rect 563882 231208 563888 231220
rect 563940 231208 563946 231260
rect 401318 231140 401324 231192
rect 401376 231180 401382 231192
rect 583754 231180 583760 231192
rect 401376 231152 583760 231180
rect 401376 231140 401382 231152
rect 583754 231140 583760 231152
rect 583812 231140 583818 231192
rect 398558 231072 398564 231124
rect 398616 231112 398622 231124
rect 581730 231112 581736 231124
rect 398616 231084 581736 231112
rect 398616 231072 398622 231084
rect 581730 231072 581736 231084
rect 581788 231072 581794 231124
rect 452654 231004 452660 231056
rect 452712 231044 452718 231056
rect 574646 231044 574652 231056
rect 452712 231016 574652 231044
rect 452712 231004 452718 231016
rect 574646 231004 574652 231016
rect 574704 231004 574710 231056
rect 534718 230936 534724 230988
rect 534776 230976 534782 230988
rect 536834 230976 536840 230988
rect 534776 230948 536840 230976
rect 534776 230936 534782 230948
rect 536834 230936 536840 230948
rect 536892 230936 536898 230988
rect 45278 230528 45284 230580
rect 45336 230568 45342 230580
rect 45738 230568 45744 230580
rect 45336 230540 45744 230568
rect 45336 230528 45342 230540
rect 45738 230528 45744 230540
rect 45796 230528 45802 230580
rect 36630 230460 36636 230512
rect 36688 230500 36694 230512
rect 46842 230500 46848 230512
rect 36688 230472 46848 230500
rect 36688 230460 36694 230472
rect 46842 230460 46848 230472
rect 46900 230460 46906 230512
rect 350442 230460 350448 230512
rect 350500 230500 350506 230512
rect 542998 230500 543004 230512
rect 350500 230472 543004 230500
rect 350500 230460 350506 230472
rect 542998 230460 543004 230472
rect 543056 230460 543062 230512
rect 388714 229916 388720 229968
rect 388772 229956 388778 229968
rect 448330 229956 448336 229968
rect 388772 229928 448336 229956
rect 388772 229916 388778 229928
rect 448330 229916 448336 229928
rect 448388 229916 448394 229968
rect 409046 229848 409052 229900
rect 409104 229888 409110 229900
rect 503714 229888 503720 229900
rect 409104 229860 503720 229888
rect 409104 229848 409110 229860
rect 503714 229848 503720 229860
rect 503772 229848 503778 229900
rect 518158 229848 518164 229900
rect 518216 229888 518222 229900
rect 543918 229888 543924 229900
rect 518216 229860 543924 229888
rect 518216 229848 518222 229860
rect 543918 229848 543924 229860
rect 543976 229848 543982 229900
rect 377766 229780 377772 229832
rect 377824 229820 377830 229832
rect 497918 229820 497924 229832
rect 377824 229792 497924 229820
rect 377824 229780 377830 229792
rect 497918 229780 497924 229792
rect 497976 229780 497982 229832
rect 378962 229712 378968 229764
rect 379020 229752 379026 229764
rect 401318 229752 401324 229764
rect 379020 229724 401324 229752
rect 379020 229712 379026 229724
rect 401318 229712 401324 229724
rect 401376 229712 401382 229764
rect 407942 229712 407948 229764
rect 408000 229752 408006 229764
rect 543918 229752 543924 229764
rect 408000 229724 543924 229752
rect 408000 229712 408006 229724
rect 543918 229712 543924 229724
rect 543976 229712 543982 229764
rect 350442 229100 350448 229152
rect 350500 229140 350506 229152
rect 366174 229140 366180 229152
rect 350500 229112 366180 229140
rect 350500 229100 350506 229112
rect 366174 229100 366180 229112
rect 366232 229100 366238 229152
rect 356790 228896 356796 228948
rect 356848 228936 356854 228948
rect 411622 228936 411628 228948
rect 356848 228908 411628 228936
rect 356848 228896 356854 228908
rect 411622 228896 411628 228908
rect 411680 228896 411686 228948
rect 509326 228896 509332 228948
rect 509384 228936 509390 228948
rect 572070 228936 572076 228948
rect 509384 228908 572076 228936
rect 509384 228896 509390 228908
rect 572070 228896 572076 228908
rect 572128 228896 572134 228948
rect 380526 228828 380532 228880
rect 380584 228868 380590 228880
rect 543182 228868 543188 228880
rect 380584 228840 543188 228868
rect 380584 228828 380590 228840
rect 543182 228828 543188 228840
rect 543240 228828 543246 228880
rect 375190 228760 375196 228812
rect 375248 228800 375254 228812
rect 541802 228800 541808 228812
rect 375248 228772 541808 228800
rect 375248 228760 375254 228772
rect 541802 228760 541808 228772
rect 541860 228760 541866 228812
rect 379974 228692 379980 228744
rect 380032 228732 380038 228744
rect 549714 228732 549720 228744
rect 380032 228704 549720 228732
rect 380032 228692 380038 228704
rect 549714 228692 549720 228704
rect 549772 228692 549778 228744
rect 404906 228624 404912 228676
rect 404964 228664 404970 228676
rect 576302 228664 576308 228676
rect 404964 228636 576308 228664
rect 404964 228624 404970 228636
rect 576302 228624 576308 228636
rect 576360 228624 576366 228676
rect 386966 228556 386972 228608
rect 387024 228596 387030 228608
rect 559558 228596 559564 228608
rect 387024 228568 559564 228596
rect 387024 228556 387030 228568
rect 559558 228556 559564 228568
rect 559616 228556 559622 228608
rect 390278 228488 390284 228540
rect 390336 228528 390342 228540
rect 563422 228528 563428 228540
rect 390336 228500 563428 228528
rect 390336 228488 390342 228500
rect 563422 228488 563428 228500
rect 563480 228488 563486 228540
rect 369394 228420 369400 228472
rect 369452 228460 369458 228472
rect 546770 228460 546776 228472
rect 369452 228432 546776 228460
rect 369452 228420 369458 228432
rect 546770 228420 546776 228432
rect 546828 228420 546834 228472
rect 384850 228352 384856 228404
rect 384908 228392 384914 228404
rect 577590 228392 577596 228404
rect 384908 228364 577596 228392
rect 384908 228352 384914 228364
rect 577590 228352 577596 228364
rect 577648 228352 577654 228404
rect 43254 227808 43260 227860
rect 43312 227848 43318 227860
rect 47118 227848 47124 227860
rect 43312 227820 47124 227848
rect 43312 227808 43318 227820
rect 47118 227808 47124 227820
rect 47176 227808 47182 227860
rect 44082 227740 44088 227792
rect 44140 227780 44146 227792
rect 46842 227780 46848 227792
rect 44140 227752 46848 227780
rect 44140 227740 44146 227752
rect 46842 227740 46848 227752
rect 46900 227740 46906 227792
rect 357066 227196 357072 227248
rect 357124 227236 357130 227248
rect 418062 227236 418068 227248
rect 357124 227208 418068 227236
rect 357124 227196 357130 227208
rect 418062 227196 418068 227208
rect 418120 227196 418126 227248
rect 380802 227128 380808 227180
rect 380860 227168 380866 227180
rect 512086 227168 512092 227180
rect 380860 227140 512092 227168
rect 380860 227128 380866 227140
rect 512086 227128 512092 227140
rect 512144 227128 512150 227180
rect 391014 227060 391020 227112
rect 391072 227100 391078 227112
rect 527542 227100 527548 227112
rect 391072 227072 527548 227100
rect 391072 227060 391078 227072
rect 527542 227060 527548 227072
rect 527600 227060 527606 227112
rect 45370 226992 45376 227044
rect 45428 227032 45434 227044
rect 46934 227032 46940 227044
rect 45428 227004 46940 227032
rect 45428 226992 45434 227004
rect 46934 226992 46940 227004
rect 46992 226992 46998 227044
rect 369302 226992 369308 227044
rect 369360 227032 369366 227044
rect 525794 227032 525800 227044
rect 369360 227004 525800 227032
rect 369360 226992 369366 227004
rect 525794 226992 525800 227004
rect 525852 226992 525858 227044
rect 355318 226312 355324 226364
rect 355376 226352 355382 226364
rect 360562 226352 360568 226364
rect 355376 226324 360568 226352
rect 355376 226312 355382 226324
rect 360562 226312 360568 226324
rect 360620 226312 360626 226364
rect 367830 225564 367836 225616
rect 367888 225604 367894 225616
rect 481174 225604 481180 225616
rect 367888 225576 481180 225604
rect 367888 225564 367894 225576
rect 481174 225564 481180 225576
rect 481232 225564 481238 225616
rect 39298 225496 39304 225548
rect 39356 225536 39362 225548
rect 46658 225536 46664 225548
rect 39356 225508 46664 225536
rect 39356 225496 39362 225508
rect 46658 225496 46664 225508
rect 46716 225496 46722 225548
rect 350442 224952 350448 225004
rect 350500 224992 350506 225004
rect 360562 224992 360568 225004
rect 350500 224964 360568 224992
rect 350500 224952 350506 224964
rect 360562 224952 360568 224964
rect 360620 224952 360626 225004
rect 39114 224680 39120 224732
rect 39172 224720 39178 224732
rect 44266 224720 44272 224732
rect 39172 224692 44272 224720
rect 39172 224680 39178 224692
rect 44266 224680 44272 224692
rect 44324 224680 44330 224732
rect 404170 224408 404176 224460
rect 404228 224448 404234 224460
rect 444466 224448 444472 224460
rect 404228 224420 444472 224448
rect 404228 224408 404234 224420
rect 444466 224408 444472 224420
rect 444524 224408 444530 224460
rect 380250 224340 380256 224392
rect 380308 224380 380314 224392
rect 459922 224380 459928 224392
rect 380308 224352 459928 224380
rect 380308 224340 380314 224352
rect 459922 224340 459928 224352
rect 459980 224340 459986 224392
rect 361022 224272 361028 224324
rect 361080 224312 361086 224324
rect 429194 224312 429200 224324
rect 361080 224284 429200 224312
rect 361080 224272 361086 224284
rect 429194 224272 429200 224284
rect 429252 224272 429258 224324
rect 436738 224272 436744 224324
rect 436796 224312 436802 224324
rect 563330 224312 563336 224324
rect 436796 224284 563336 224312
rect 436796 224272 436802 224284
rect 563330 224272 563336 224284
rect 563388 224272 563394 224324
rect 387610 224204 387616 224256
rect 387668 224244 387674 224256
rect 521654 224244 521660 224256
rect 387668 224216 521660 224244
rect 387668 224204 387674 224216
rect 521654 224204 521660 224216
rect 521712 224204 521718 224256
rect 348786 223864 348792 223916
rect 348844 223904 348850 223916
rect 349154 223904 349160 223916
rect 348844 223876 349160 223904
rect 348844 223864 348850 223876
rect 349154 223864 349160 223876
rect 349212 223864 349218 223916
rect 31110 223592 31116 223644
rect 31168 223632 31174 223644
rect 46842 223632 46848 223644
rect 31168 223604 46848 223632
rect 31168 223592 31174 223604
rect 46842 223592 46848 223604
rect 46900 223592 46906 223644
rect 350442 223524 350448 223576
rect 350500 223564 350506 223576
rect 388898 223564 388904 223576
rect 350500 223536 388904 223564
rect 350500 223524 350506 223536
rect 388898 223524 388904 223536
rect 388956 223524 388962 223576
rect 392302 222912 392308 222964
rect 392360 222952 392366 222964
rect 413554 222952 413560 222964
rect 392360 222924 413560 222952
rect 392360 222912 392366 222924
rect 413554 222912 413560 222924
rect 413612 222912 413618 222964
rect 409874 222844 409880 222896
rect 409932 222884 409938 222896
rect 472802 222884 472808 222896
rect 409932 222856 472808 222884
rect 409932 222844 409938 222856
rect 472802 222844 472808 222856
rect 472860 222844 472866 222896
rect 350166 222572 350172 222624
rect 350224 222612 350230 222624
rect 352650 222612 352656 222624
rect 350224 222584 352656 222612
rect 350224 222572 350230 222584
rect 352650 222572 352656 222584
rect 352708 222572 352714 222624
rect 35342 222164 35348 222216
rect 35400 222204 35406 222216
rect 46842 222204 46848 222216
rect 35400 222176 46848 222204
rect 35400 222164 35406 222176
rect 46842 222164 46848 222176
rect 46900 222164 46906 222216
rect 350258 222096 350264 222148
rect 350316 222136 350322 222148
rect 351914 222136 351920 222148
rect 350316 222108 351920 222136
rect 350316 222096 350322 222108
rect 351914 222096 351920 222108
rect 351972 222096 351978 222148
rect 39942 221416 39948 221468
rect 40000 221456 40006 221468
rect 40678 221456 40684 221468
rect 40000 221428 40684 221456
rect 40000 221416 40006 221428
rect 40678 221416 40684 221428
rect 40736 221416 40742 221468
rect 397914 221416 397920 221468
rect 397972 221456 397978 221468
rect 477954 221456 477960 221468
rect 397972 221428 477960 221456
rect 397972 221416 397978 221428
rect 477954 221416 477960 221428
rect 478012 221416 478018 221468
rect 350442 221144 350448 221196
rect 350500 221184 350506 221196
rect 356422 221184 356428 221196
rect 350500 221156 356428 221184
rect 350500 221144 350506 221156
rect 356422 221144 356428 221156
rect 356480 221144 356486 221196
rect 31202 220804 31208 220856
rect 31260 220844 31266 220856
rect 46842 220844 46848 220856
rect 31260 220816 46848 220844
rect 31260 220804 31266 220816
rect 46842 220804 46848 220816
rect 46900 220804 46906 220856
rect 355962 220736 355968 220788
rect 356020 220776 356026 220788
rect 356606 220776 356612 220788
rect 356020 220748 356612 220776
rect 356020 220736 356026 220748
rect 356606 220736 356612 220748
rect 356664 220736 356670 220788
rect 41046 220396 41052 220448
rect 41104 220436 41110 220448
rect 46014 220436 46020 220448
rect 41104 220408 46020 220436
rect 41104 220396 41110 220408
rect 46014 220396 46020 220408
rect 46072 220396 46078 220448
rect 44266 220260 44272 220312
rect 44324 220300 44330 220312
rect 46014 220300 46020 220312
rect 44324 220272 46020 220300
rect 44324 220260 44330 220272
rect 46014 220260 46020 220272
rect 46072 220260 46078 220312
rect 377950 220124 377956 220176
rect 378008 220164 378014 220176
rect 435450 220164 435456 220176
rect 378008 220136 435456 220164
rect 378008 220124 378014 220136
rect 435450 220124 435456 220136
rect 435508 220124 435514 220176
rect 354030 220056 354036 220108
rect 354088 220096 354094 220108
rect 494054 220096 494060 220108
rect 354088 220068 494060 220096
rect 354088 220056 354094 220068
rect 494054 220056 494060 220068
rect 494112 220056 494118 220108
rect 354582 219444 354588 219496
rect 354640 219484 354646 219496
rect 356054 219484 356060 219496
rect 354640 219456 356060 219484
rect 354640 219444 354646 219456
rect 356054 219444 356060 219456
rect 356112 219444 356118 219496
rect 36906 218696 36912 218748
rect 36964 218736 36970 218748
rect 46106 218736 46112 218748
rect 36964 218708 46112 218736
rect 36964 218696 36970 218708
rect 46106 218696 46112 218708
rect 46164 218696 46170 218748
rect 369118 218696 369124 218748
rect 369176 218736 369182 218748
rect 476666 218736 476672 218748
rect 369176 218708 476672 218736
rect 369176 218696 369182 218708
rect 476666 218696 476672 218708
rect 476724 218696 476730 218748
rect 35802 218084 35808 218136
rect 35860 218124 35866 218136
rect 46566 218124 46572 218136
rect 35860 218096 46572 218124
rect 35860 218084 35866 218096
rect 46566 218084 46572 218096
rect 46624 218084 46630 218136
rect 348970 218084 348976 218136
rect 349028 218124 349034 218136
rect 349154 218124 349160 218136
rect 349028 218096 349160 218124
rect 349028 218084 349034 218096
rect 349154 218084 349160 218096
rect 349212 218084 349218 218136
rect 32306 218016 32312 218068
rect 32364 218056 32370 218068
rect 46842 218056 46848 218068
rect 32364 218028 46848 218056
rect 32364 218016 32370 218028
rect 46842 218016 46848 218028
rect 46900 218016 46906 218068
rect 348694 218016 348700 218068
rect 348752 218056 348758 218068
rect 349430 218056 349436 218068
rect 348752 218028 349436 218056
rect 348752 218016 348758 218028
rect 349430 218016 349436 218028
rect 349488 218016 349494 218068
rect 350442 218016 350448 218068
rect 350500 218056 350506 218068
rect 355502 218056 355508 218068
rect 350500 218028 355508 218056
rect 350500 218016 350506 218028
rect 355502 218016 355508 218028
rect 355560 218016 355566 218068
rect 350258 217948 350264 218000
rect 350316 217988 350322 218000
rect 354950 217988 354956 218000
rect 350316 217960 354956 217988
rect 350316 217948 350322 217960
rect 354950 217948 354956 217960
rect 355008 217948 355014 218000
rect 45922 217472 45928 217524
rect 45980 217472 45986 217524
rect 45940 217320 45968 217472
rect 45922 217268 45928 217320
rect 45980 217268 45986 217320
rect 356698 217268 356704 217320
rect 356756 217308 356762 217320
rect 445754 217308 445760 217320
rect 356756 217280 445760 217308
rect 356756 217268 356762 217280
rect 445754 217268 445760 217280
rect 445812 217268 445818 217320
rect 350442 217200 350448 217252
rect 350500 217240 350506 217252
rect 355042 217240 355048 217252
rect 350500 217212 355048 217240
rect 350500 217200 350506 217212
rect 355042 217200 355048 217212
rect 355100 217200 355106 217252
rect 36906 216656 36912 216708
rect 36964 216696 36970 216708
rect 46014 216696 46020 216708
rect 36964 216668 46020 216696
rect 36964 216656 36970 216668
rect 46014 216656 46020 216668
rect 46072 216656 46078 216708
rect 388622 215908 388628 215960
rect 388680 215948 388686 215960
rect 535914 215948 535920 215960
rect 388680 215920 535920 215948
rect 388680 215908 388686 215920
rect 535914 215908 535920 215920
rect 535972 215908 535978 215960
rect 46382 215364 46388 215416
rect 46440 215404 46446 215416
rect 47118 215404 47124 215416
rect 46440 215376 47124 215404
rect 46440 215364 46446 215376
rect 47118 215364 47124 215376
rect 47176 215364 47182 215416
rect 32214 215296 32220 215348
rect 32272 215336 32278 215348
rect 46842 215336 46848 215348
rect 32272 215308 46848 215336
rect 32272 215296 32278 215308
rect 46842 215296 46848 215308
rect 46900 215296 46906 215348
rect 350442 215296 350448 215348
rect 350500 215336 350506 215348
rect 353294 215336 353300 215348
rect 350500 215308 353300 215336
rect 350500 215296 350506 215308
rect 353294 215296 353300 215308
rect 353352 215296 353358 215348
rect 354582 215228 354588 215280
rect 354640 215268 354646 215280
rect 356514 215268 356520 215280
rect 354640 215240 356520 215268
rect 354640 215228 354646 215240
rect 356514 215228 356520 215240
rect 356572 215228 356578 215280
rect 41782 214548 41788 214600
rect 41840 214588 41846 214600
rect 44174 214588 44180 214600
rect 41840 214560 44180 214588
rect 41840 214548 41846 214560
rect 44174 214548 44180 214560
rect 44232 214548 44238 214600
rect 45094 214548 45100 214600
rect 45152 214588 45158 214600
rect 45370 214588 45376 214600
rect 45152 214560 45376 214588
rect 45152 214548 45158 214560
rect 45370 214548 45376 214560
rect 45428 214548 45434 214600
rect 45830 214548 45836 214600
rect 45888 214588 45894 214600
rect 47118 214588 47124 214600
rect 45888 214560 47124 214588
rect 45888 214548 45894 214560
rect 47118 214548 47124 214560
rect 47176 214548 47182 214600
rect 433334 214548 433340 214600
rect 433392 214588 433398 214600
rect 581546 214588 581552 214600
rect 433392 214560 581552 214588
rect 433392 214548 433398 214560
rect 581546 214548 581552 214560
rect 581604 214548 581610 214600
rect 38102 213936 38108 213988
rect 38160 213976 38166 213988
rect 46842 213976 46848 213988
rect 38160 213948 46848 213976
rect 38160 213936 38166 213948
rect 46842 213936 46848 213948
rect 46900 213936 46906 213988
rect 45370 213868 45376 213920
rect 45428 213908 45434 213920
rect 45738 213908 45744 213920
rect 45428 213880 45744 213908
rect 45428 213868 45434 213880
rect 45738 213868 45744 213880
rect 45796 213868 45802 213920
rect 407022 213256 407028 213308
rect 407080 213296 407086 213308
rect 485038 213296 485044 213308
rect 407080 213268 485044 213296
rect 407080 213256 407086 213268
rect 485038 213256 485044 213268
rect 485096 213256 485102 213308
rect 356882 213188 356888 213240
rect 356940 213228 356946 213240
rect 542538 213228 542544 213240
rect 356940 213200 542544 213228
rect 356940 213188 356946 213200
rect 542538 213188 542544 213200
rect 542596 213188 542602 213240
rect 46566 213120 46572 213172
rect 46624 213160 46630 213172
rect 47578 213160 47584 213172
rect 46624 213132 47584 213160
rect 46624 213120 46630 213132
rect 47578 213120 47584 213132
rect 47636 213120 47642 213172
rect 350442 212508 350448 212560
rect 350500 212548 350506 212560
rect 508498 212548 508504 212560
rect 350500 212520 508504 212548
rect 350500 212508 350506 212520
rect 508498 212508 508504 212520
rect 508556 212508 508562 212560
rect 348970 212440 348976 212492
rect 349028 212480 349034 212492
rect 349338 212480 349344 212492
rect 349028 212452 349344 212480
rect 349028 212440 349034 212452
rect 349338 212440 349344 212452
rect 349396 212440 349402 212492
rect 349062 212372 349068 212424
rect 349120 212412 349126 212424
rect 349706 212412 349712 212424
rect 349120 212384 349712 212412
rect 349120 212372 349126 212384
rect 349706 212372 349712 212384
rect 349764 212372 349770 212424
rect 438670 211964 438676 212016
rect 438728 212004 438734 212016
rect 477586 212004 477592 212016
rect 438728 211976 477592 212004
rect 438728 211964 438734 211976
rect 477586 211964 477592 211976
rect 477644 211964 477650 212016
rect 388530 211896 388536 211948
rect 388588 211936 388594 211948
rect 441614 211936 441620 211948
rect 388588 211908 441620 211936
rect 388588 211896 388594 211908
rect 441614 211896 441620 211908
rect 441672 211896 441678 211948
rect 382734 211828 382740 211880
rect 382792 211868 382798 211880
rect 524966 211868 524972 211880
rect 382792 211840 524972 211868
rect 382792 211828 382798 211840
rect 524966 211828 524972 211840
rect 525024 211828 525030 211880
rect 33870 211760 33876 211812
rect 33928 211800 33934 211812
rect 47578 211800 47584 211812
rect 33928 211772 47584 211800
rect 33928 211760 33934 211772
rect 47578 211760 47584 211772
rect 47636 211760 47642 211812
rect 416958 211760 416964 211812
rect 417016 211800 417022 211812
rect 583294 211800 583300 211812
rect 417016 211772 583300 211800
rect 417016 211760 417022 211772
rect 583294 211760 583300 211772
rect 583352 211760 583358 211812
rect 33870 211148 33876 211200
rect 33928 211188 33934 211200
rect 46842 211188 46848 211200
rect 33928 211160 46848 211188
rect 33928 211148 33934 211160
rect 46842 211148 46848 211160
rect 46900 211148 46906 211200
rect 350442 208360 350448 208412
rect 350500 208400 350506 208412
rect 539042 208400 539048 208412
rect 350500 208372 539048 208400
rect 350500 208360 350506 208372
rect 539042 208360 539048 208372
rect 539100 208360 539106 208412
rect 43806 208292 43812 208344
rect 43864 208332 43870 208344
rect 46842 208332 46848 208344
rect 43864 208304 46848 208332
rect 43864 208292 43870 208304
rect 46842 208292 46848 208304
rect 46900 208292 46906 208344
rect 350442 207068 350448 207120
rect 350500 207108 350506 207120
rect 541986 207108 541992 207120
rect 350500 207080 541992 207108
rect 350500 207068 350506 207080
rect 541986 207068 541992 207080
rect 542044 207068 542050 207120
rect 350258 207000 350264 207052
rect 350316 207040 350322 207052
rect 566550 207040 566556 207052
rect 350316 207012 566556 207040
rect 350316 207000 350322 207012
rect 566550 207000 566556 207012
rect 566608 207000 566614 207052
rect 41230 206932 41236 206984
rect 41288 206972 41294 206984
rect 46842 206972 46848 206984
rect 41288 206944 46848 206972
rect 41288 206932 41294 206944
rect 46842 206932 46848 206944
rect 46900 206932 46906 206984
rect 350442 206932 350448 206984
rect 350500 206972 350506 206984
rect 376294 206972 376300 206984
rect 350500 206944 376300 206972
rect 350500 206932 350506 206944
rect 376294 206932 376300 206944
rect 376352 206932 376358 206984
rect 410058 206252 410064 206304
rect 410116 206292 410122 206304
rect 507578 206292 507584 206304
rect 410116 206264 507584 206292
rect 410116 206252 410122 206264
rect 507578 206252 507584 206264
rect 507636 206252 507642 206304
rect 348970 206116 348976 206168
rect 349028 206156 349034 206168
rect 352558 206156 352564 206168
rect 349028 206128 352564 206156
rect 349028 206116 349034 206128
rect 352558 206116 352564 206128
rect 352616 206116 352622 206168
rect 37182 205640 37188 205692
rect 37240 205680 37246 205692
rect 46842 205680 46848 205692
rect 37240 205652 46848 205680
rect 37240 205640 37246 205652
rect 46842 205640 46848 205652
rect 46900 205640 46906 205692
rect 36998 205164 37004 205216
rect 37056 205204 37062 205216
rect 37734 205204 37740 205216
rect 37056 205176 37740 205204
rect 37056 205164 37062 205176
rect 37734 205164 37740 205176
rect 37792 205164 37798 205216
rect 442994 204892 443000 204944
rect 443052 204932 443058 204944
rect 508222 204932 508228 204944
rect 443052 204904 508228 204932
rect 443052 204892 443058 204904
rect 508222 204892 508228 204904
rect 508280 204892 508286 204944
rect 349982 204416 349988 204468
rect 350040 204456 350046 204468
rect 351914 204456 351920 204468
rect 350040 204428 351920 204456
rect 350040 204416 350046 204428
rect 351914 204416 351920 204428
rect 351972 204416 351978 204468
rect 46842 204280 46848 204332
rect 46900 204320 46906 204332
rect 47118 204320 47124 204332
rect 46900 204292 47124 204320
rect 46900 204280 46906 204292
rect 47118 204280 47124 204292
rect 47176 204280 47182 204332
rect 350258 204280 350264 204332
rect 350316 204320 350322 204332
rect 389082 204320 389088 204332
rect 350316 204292 389088 204320
rect 350316 204280 350322 204292
rect 389082 204280 389088 204292
rect 389140 204280 389146 204332
rect 350442 204212 350448 204264
rect 350500 204252 350506 204264
rect 418798 204252 418804 204264
rect 350500 204224 418804 204252
rect 350500 204212 350506 204224
rect 418798 204212 418804 204224
rect 418856 204212 418862 204264
rect 406470 203600 406476 203652
rect 406528 203640 406534 203652
rect 519170 203640 519176 203652
rect 406528 203612 519176 203640
rect 406528 203600 406534 203612
rect 519170 203600 519176 203612
rect 519228 203600 519234 203652
rect 350074 203532 350080 203584
rect 350132 203572 350138 203584
rect 545298 203572 545304 203584
rect 350132 203544 545304 203572
rect 350132 203532 350138 203544
rect 545298 203532 545304 203544
rect 545356 203532 545362 203584
rect 36998 202852 37004 202904
rect 37056 202892 37062 202904
rect 45646 202892 45652 202904
rect 37056 202864 45652 202892
rect 37056 202852 37062 202864
rect 45646 202852 45652 202864
rect 45704 202852 45710 202904
rect 350442 202852 350448 202904
rect 350500 202892 350506 202904
rect 414658 202892 414664 202904
rect 350500 202864 414664 202892
rect 350500 202852 350506 202864
rect 414658 202852 414664 202864
rect 414716 202852 414722 202904
rect 34882 202784 34888 202836
rect 34940 202824 34946 202836
rect 45554 202824 45560 202836
rect 34940 202796 45560 202824
rect 34940 202784 34946 202796
rect 45554 202784 45560 202796
rect 45612 202784 45618 202836
rect 46382 202308 46388 202360
rect 46440 202348 46446 202360
rect 47854 202348 47860 202360
rect 46440 202320 47860 202348
rect 46440 202308 46446 202320
rect 47854 202308 47860 202320
rect 47912 202308 47918 202360
rect 411346 202104 411352 202156
rect 411404 202144 411410 202156
rect 476022 202144 476028 202156
rect 411404 202116 476028 202144
rect 411404 202104 411410 202116
rect 476022 202104 476028 202116
rect 476080 202104 476086 202156
rect 350442 201492 350448 201544
rect 350500 201532 350506 201544
rect 383378 201532 383384 201544
rect 350500 201504 383384 201532
rect 350500 201492 350506 201504
rect 383378 201492 383384 201504
rect 383436 201492 383442 201544
rect 349062 200744 349068 200796
rect 349120 200784 349126 200796
rect 359182 200784 359188 200796
rect 349120 200756 359188 200784
rect 349120 200744 349126 200756
rect 359182 200744 359188 200756
rect 359240 200744 359246 200796
rect 363322 200744 363328 200796
rect 363380 200784 363386 200796
rect 507946 200784 507952 200796
rect 363380 200756 507952 200784
rect 363380 200744 363386 200756
rect 507946 200744 507952 200756
rect 508004 200744 508010 200796
rect 347682 200336 347688 200388
rect 347740 200336 347746 200388
rect 42334 200064 42340 200116
rect 42392 200104 42398 200116
rect 44266 200104 44272 200116
rect 42392 200076 44272 200104
rect 42392 200064 42398 200076
rect 44266 200064 44272 200076
rect 44324 200064 44330 200116
rect 46658 199928 46664 199980
rect 46716 199968 46722 199980
rect 50338 199968 50344 199980
rect 46716 199940 50344 199968
rect 46716 199928 46722 199940
rect 50338 199928 50344 199940
rect 50396 199928 50402 199980
rect 347700 199912 347728 200336
rect 347682 199860 347688 199912
rect 347740 199860 347746 199912
rect 41046 199656 41052 199708
rect 41104 199696 41110 199708
rect 75454 199696 75460 199708
rect 41104 199668 75460 199696
rect 41104 199656 41110 199668
rect 75454 199656 75460 199668
rect 75512 199656 75518 199708
rect 44542 199588 44548 199640
rect 44600 199628 44606 199640
rect 90910 199628 90916 199640
rect 44600 199600 90916 199628
rect 44600 199588 44606 199600
rect 90910 199588 90916 199600
rect 90968 199588 90974 199640
rect 104066 199588 104072 199640
rect 104124 199628 104130 199640
rect 104710 199628 104716 199640
rect 104124 199600 104716 199628
rect 104124 199588 104130 199600
rect 104710 199588 104716 199600
rect 104768 199588 104774 199640
rect 346302 199588 346308 199640
rect 346360 199628 346366 199640
rect 348786 199628 348792 199640
rect 346360 199600 348792 199628
rect 346360 199588 346366 199600
rect 348786 199588 348792 199600
rect 348844 199588 348850 199640
rect 43438 199520 43444 199572
rect 43496 199560 43502 199572
rect 92658 199560 92664 199572
rect 43496 199532 92664 199560
rect 43496 199520 43502 199532
rect 92658 199520 92664 199532
rect 92716 199520 92722 199572
rect 275830 199520 275836 199572
rect 275888 199560 275894 199572
rect 340874 199560 340880 199572
rect 275888 199532 340880 199560
rect 275888 199520 275894 199532
rect 340874 199520 340880 199532
rect 340932 199520 340938 199572
rect 347498 199520 347504 199572
rect 347556 199560 347562 199572
rect 350166 199560 350172 199572
rect 347556 199532 350172 199560
rect 347556 199520 347562 199532
rect 350166 199520 350172 199532
rect 350224 199520 350230 199572
rect 47026 199452 47032 199504
rect 47084 199492 47090 199504
rect 108942 199492 108948 199504
rect 47084 199464 108948 199492
rect 47084 199452 47090 199464
rect 108942 199452 108948 199464
rect 109000 199452 109006 199504
rect 328178 199452 328184 199504
rect 328236 199492 328242 199504
rect 348602 199492 348608 199504
rect 328236 199464 348608 199492
rect 328236 199452 328242 199464
rect 348602 199452 348608 199464
rect 348660 199452 348666 199504
rect 44818 199384 44824 199436
rect 44876 199424 44882 199436
rect 158530 199424 158536 199436
rect 44876 199396 158536 199424
rect 44876 199384 44882 199396
rect 158530 199384 158536 199396
rect 158588 199384 158594 199436
rect 317230 199384 317236 199436
rect 317288 199424 317294 199436
rect 348510 199424 348516 199436
rect 317288 199396 348516 199424
rect 317288 199384 317294 199396
rect 348510 199384 348516 199396
rect 348568 199384 348574 199436
rect 348970 199384 348976 199436
rect 349028 199424 349034 199436
rect 354858 199424 354864 199436
rect 349028 199396 354864 199424
rect 349028 199384 349034 199396
rect 354858 199384 354864 199396
rect 354916 199384 354922 199436
rect 319806 199316 319812 199368
rect 319864 199356 319870 199368
rect 360838 199356 360844 199368
rect 319864 199328 360844 199356
rect 319864 199316 319870 199328
rect 360838 199316 360844 199328
rect 360896 199316 360902 199368
rect 35434 199248 35440 199300
rect 35492 199288 35498 199300
rect 105998 199288 106004 199300
rect 35492 199260 106004 199288
rect 35492 199248 35498 199260
rect 105998 199248 106004 199260
rect 106056 199248 106062 199300
rect 271506 199248 271512 199300
rect 271564 199288 271570 199300
rect 358262 199288 358268 199300
rect 271564 199260 358268 199288
rect 271564 199248 271570 199260
rect 358262 199248 358268 199260
rect 358320 199248 358326 199300
rect 38194 199180 38200 199232
rect 38252 199220 38258 199232
rect 118786 199220 118792 199232
rect 38252 199192 118792 199220
rect 38252 199180 38258 199192
rect 118786 199180 118792 199192
rect 118844 199180 118850 199232
rect 208394 199180 208400 199232
rect 208452 199220 208458 199232
rect 366450 199220 366456 199232
rect 208452 199192 366456 199220
rect 208452 199180 208458 199192
rect 366450 199180 366456 199192
rect 366508 199180 366514 199232
rect 27154 199112 27160 199164
rect 27212 199152 27218 199164
rect 127250 199152 127256 199164
rect 27212 199124 127256 199152
rect 27212 199112 27218 199124
rect 127250 199112 127256 199124
rect 127308 199112 127314 199164
rect 300486 199112 300492 199164
rect 300544 199152 300550 199164
rect 560938 199152 560944 199164
rect 300544 199124 560944 199152
rect 300544 199112 300550 199124
rect 560938 199112 560944 199124
rect 560996 199112 561002 199164
rect 39482 199044 39488 199096
rect 39540 199084 39546 199096
rect 104618 199084 104624 199096
rect 39540 199056 104624 199084
rect 39540 199044 39546 199056
rect 104618 199044 104624 199056
rect 104676 199044 104682 199096
rect 104710 199044 104716 199096
rect 104768 199084 104774 199096
rect 370866 199084 370872 199096
rect 104768 199056 370872 199084
rect 104768 199044 104774 199056
rect 370866 199044 370872 199056
rect 370924 199044 370930 199096
rect 84102 198976 84108 199028
rect 84160 199016 84166 199028
rect 371878 199016 371884 199028
rect 84160 198988 371884 199016
rect 84160 198976 84166 198988
rect 371878 198976 371884 198988
rect 371936 198976 371942 199028
rect 37090 198908 37096 198960
rect 37148 198948 37154 198960
rect 167822 198948 167828 198960
rect 37148 198920 167828 198948
rect 37148 198908 37154 198920
rect 167822 198908 167828 198920
rect 167880 198908 167886 198960
rect 233510 198908 233516 198960
rect 233568 198948 233574 198960
rect 542078 198948 542084 198960
rect 233568 198920 542084 198948
rect 233568 198908 233574 198920
rect 542078 198908 542084 198920
rect 542136 198908 542142 198960
rect 40494 198840 40500 198892
rect 40552 198880 40558 198892
rect 221918 198880 221924 198892
rect 40552 198852 221924 198880
rect 40552 198840 40558 198852
rect 221918 198840 221924 198852
rect 221976 198840 221982 198892
rect 247034 198840 247040 198892
rect 247092 198880 247098 198892
rect 559374 198880 559380 198892
rect 247092 198852 559380 198880
rect 247092 198840 247098 198852
rect 559374 198840 559380 198852
rect 559432 198840 559438 198892
rect 30006 198772 30012 198824
rect 30064 198812 30070 198824
rect 160094 198812 160100 198824
rect 30064 198784 160100 198812
rect 30064 198772 30070 198784
rect 160094 198772 160100 198784
rect 160152 198772 160158 198824
rect 194226 198772 194232 198824
rect 194284 198812 194290 198824
rect 559650 198812 559656 198824
rect 194284 198784 559656 198812
rect 194284 198772 194290 198784
rect 559650 198772 559656 198784
rect 559708 198772 559714 198824
rect 100846 198704 100852 198756
rect 100904 198744 100910 198756
rect 467926 198744 467932 198756
rect 100904 198716 467932 198744
rect 100904 198704 100910 198716
rect 467926 198704 467932 198716
rect 467984 198704 467990 198756
rect 22922 198636 22928 198688
rect 22980 198676 22986 198688
rect 48682 198676 48688 198688
rect 22980 198648 48688 198676
rect 22980 198636 22986 198648
rect 48682 198636 48688 198648
rect 48740 198636 48746 198688
rect 346210 198636 346216 198688
rect 346268 198676 346274 198688
rect 360378 198676 360384 198688
rect 346268 198648 360384 198676
rect 346268 198636 346274 198648
rect 360378 198636 360384 198648
rect 360436 198636 360442 198688
rect 25682 198568 25688 198620
rect 25740 198608 25746 198620
rect 101490 198608 101496 198620
rect 25740 198580 101496 198608
rect 25740 198568 25746 198580
rect 101490 198568 101496 198580
rect 101548 198568 101554 198620
rect 123386 198568 123392 198620
rect 123444 198608 123450 198620
rect 570874 198608 570880 198620
rect 123444 198580 570880 198608
rect 123444 198568 123450 198580
rect 570874 198568 570880 198580
rect 570932 198568 570938 198620
rect 46566 198500 46572 198552
rect 46624 198540 46630 198552
rect 168466 198540 168472 198552
rect 46624 198512 168472 198540
rect 46624 198500 46630 198512
rect 168466 198500 168472 198512
rect 168524 198500 168530 198552
rect 223850 198500 223856 198552
rect 223908 198540 223914 198552
rect 553946 198540 553952 198552
rect 223908 198512 553952 198540
rect 223908 198500 223914 198512
rect 553946 198500 553952 198512
rect 554004 198500 554010 198552
rect 33042 198432 33048 198484
rect 33100 198472 33106 198484
rect 67358 198472 67364 198484
rect 33100 198444 67364 198472
rect 33100 198432 33106 198444
rect 67358 198432 67364 198444
rect 67416 198432 67422 198484
rect 244458 198432 244464 198484
rect 244516 198472 244522 198484
rect 558270 198472 558276 198484
rect 244516 198444 558276 198472
rect 244516 198432 244522 198444
rect 558270 198432 558276 198444
rect 558328 198432 558334 198484
rect 22830 198364 22836 198416
rect 22888 198404 22894 198416
rect 55766 198404 55772 198416
rect 22888 198376 55772 198404
rect 22888 198364 22894 198376
rect 55766 198364 55772 198376
rect 55824 198364 55830 198416
rect 58618 198364 58624 198416
rect 58676 198404 58682 198416
rect 77662 198404 77668 198416
rect 58676 198376 77668 198404
rect 58676 198364 58682 198376
rect 77662 198364 77668 198376
rect 77720 198364 77726 198416
rect 201954 198364 201960 198416
rect 202012 198404 202018 198416
rect 491386 198404 491392 198416
rect 202012 198376 491392 198404
rect 202012 198364 202018 198376
rect 491386 198364 491392 198376
rect 491444 198364 491450 198416
rect 44726 198296 44732 198348
rect 44784 198336 44790 198348
rect 88610 198336 88616 198348
rect 44784 198308 88616 198336
rect 44784 198296 44790 198308
rect 88610 198296 88616 198308
rect 88668 198296 88674 198348
rect 147858 198296 147864 198348
rect 147916 198336 147922 198348
rect 254854 198336 254860 198348
rect 147916 198308 254860 198336
rect 147916 198296 147922 198308
rect 254854 198296 254860 198308
rect 254912 198296 254918 198348
rect 287606 198296 287612 198348
rect 287664 198336 287670 198348
rect 551002 198336 551008 198348
rect 287664 198308 551008 198336
rect 287664 198296 287670 198308
rect 551002 198296 551008 198308
rect 551060 198296 551066 198348
rect 31570 198228 31576 198280
rect 31628 198268 31634 198280
rect 64138 198268 64144 198280
rect 31628 198240 64144 198268
rect 31628 198228 31634 198240
rect 64138 198228 64144 198240
rect 64196 198228 64202 198280
rect 342990 198228 342996 198280
rect 343048 198268 343054 198280
rect 365254 198268 365260 198280
rect 343048 198240 365260 198268
rect 343048 198228 343054 198240
rect 365254 198228 365260 198240
rect 365312 198228 365318 198280
rect 40402 198160 40408 198212
rect 40460 198200 40466 198212
rect 145650 198200 145656 198212
rect 40460 198172 145656 198200
rect 40460 198160 40466 198172
rect 145650 198160 145656 198172
rect 145708 198160 145714 198212
rect 160738 198160 160744 198212
rect 160796 198200 160802 198212
rect 166258 198200 166264 198212
rect 160796 198172 166264 198200
rect 160796 198160 160802 198172
rect 166258 198160 166264 198172
rect 166316 198160 166322 198212
rect 190362 198160 190368 198212
rect 190420 198200 190426 198212
rect 383010 198200 383016 198212
rect 190420 198172 383016 198200
rect 190420 198160 190426 198172
rect 383010 198160 383016 198172
rect 383068 198160 383074 198212
rect 17770 198092 17776 198144
rect 17828 198132 17834 198144
rect 49970 198132 49976 198144
rect 17828 198104 49976 198132
rect 17828 198092 17834 198104
rect 49970 198092 49976 198104
rect 50028 198092 50034 198144
rect 51902 198092 51908 198144
rect 51960 198132 51966 198144
rect 165246 198132 165252 198144
rect 51960 198104 165252 198132
rect 51960 198092 51966 198104
rect 165246 198092 165252 198104
rect 165304 198092 165310 198144
rect 201310 198092 201316 198144
rect 201368 198132 201374 198144
rect 268378 198132 268384 198144
rect 201368 198104 268384 198132
rect 201368 198092 201374 198104
rect 268378 198092 268384 198104
rect 268436 198092 268442 198144
rect 275370 198092 275376 198144
rect 275428 198132 275434 198144
rect 364334 198132 364340 198144
rect 275428 198104 364340 198132
rect 275428 198092 275434 198104
rect 364334 198092 364340 198104
rect 364392 198092 364398 198144
rect 44082 198024 44088 198076
rect 44140 198064 44146 198076
rect 208762 198064 208768 198076
rect 44140 198036 208768 198064
rect 44140 198024 44146 198036
rect 208762 198024 208768 198036
rect 208820 198024 208826 198076
rect 272150 198024 272156 198076
rect 272208 198064 272214 198076
rect 307018 198064 307024 198076
rect 272208 198036 307024 198064
rect 272208 198024 272214 198036
rect 307018 198024 307024 198036
rect 307076 198024 307082 198076
rect 332042 198024 332048 198076
rect 332100 198064 332106 198076
rect 401042 198064 401048 198076
rect 332100 198036 401048 198064
rect 332100 198024 332106 198036
rect 401042 198024 401048 198036
rect 401100 198024 401106 198076
rect 25774 197956 25780 198008
rect 25832 197996 25838 198008
rect 48038 197996 48044 198008
rect 25832 197968 48044 197996
rect 25832 197956 25838 197968
rect 48038 197956 48044 197968
rect 48096 197956 48102 198008
rect 50062 197956 50068 198008
rect 50120 197996 50126 198008
rect 50614 197996 50620 198008
rect 50120 197968 50620 197996
rect 50120 197956 50126 197968
rect 50614 197956 50620 197968
rect 50672 197956 50678 198008
rect 53006 197956 53012 198008
rect 53064 197996 53070 198008
rect 395338 197996 395344 198008
rect 53064 197968 395344 197996
rect 53064 197956 53070 197968
rect 395338 197956 395344 197968
rect 395396 197956 395402 198008
rect 32858 197888 32864 197940
rect 32916 197928 32922 197940
rect 63494 197928 63500 197940
rect 32916 197900 63500 197928
rect 32916 197888 32922 197900
rect 63494 197888 63500 197900
rect 63552 197888 63558 197940
rect 317874 197888 317880 197940
rect 317932 197928 317938 197940
rect 385678 197928 385684 197940
rect 317932 197900 385684 197928
rect 317932 197888 317938 197900
rect 385678 197888 385684 197900
rect 385736 197888 385742 197940
rect 49510 197820 49516 197872
rect 49568 197860 49574 197872
rect 72510 197860 72516 197872
rect 49568 197832 72516 197860
rect 49568 197820 49574 197832
rect 72510 197820 72516 197832
rect 72568 197820 72574 197872
rect 315298 197820 315304 197872
rect 315356 197860 315362 197872
rect 349062 197860 349068 197872
rect 315356 197832 349068 197860
rect 315356 197820 315362 197832
rect 349062 197820 349068 197832
rect 349120 197820 349126 197872
rect 86678 197752 86684 197804
rect 86736 197792 86742 197804
rect 346118 197792 346124 197804
rect 86736 197764 346124 197792
rect 86736 197752 86742 197764
rect 346118 197752 346124 197764
rect 346176 197752 346182 197804
rect 36906 197684 36912 197736
rect 36964 197724 36970 197736
rect 487154 197724 487160 197736
rect 36964 197696 487160 197724
rect 36964 197684 36970 197696
rect 487154 197684 487160 197696
rect 487212 197684 487218 197736
rect 49326 197412 49332 197464
rect 49384 197452 49390 197464
rect 54478 197452 54484 197464
rect 49384 197424 54484 197452
rect 49384 197412 49390 197424
rect 54478 197412 54484 197424
rect 54536 197412 54542 197464
rect 51258 197344 51264 197396
rect 51316 197384 51322 197396
rect 53190 197384 53196 197396
rect 51316 197356 53196 197384
rect 51316 197344 51322 197356
rect 53190 197344 53196 197356
rect 53248 197344 53254 197396
rect 68278 197344 68284 197396
rect 68336 197384 68342 197396
rect 71130 197384 71136 197396
rect 68336 197356 71136 197384
rect 68336 197344 68342 197356
rect 71130 197344 71136 197356
rect 71188 197344 71194 197396
rect 108574 197344 108580 197396
rect 108632 197384 108638 197396
rect 109678 197384 109684 197396
rect 108632 197356 109684 197384
rect 108632 197344 108638 197356
rect 109678 197344 109684 197356
rect 109736 197344 109742 197396
rect 262490 197344 262496 197396
rect 262548 197384 262554 197396
rect 264238 197384 264244 197396
rect 262548 197356 264244 197384
rect 262548 197344 262554 197356
rect 264238 197344 264244 197356
rect 264296 197344 264302 197396
rect 41322 197276 41328 197328
rect 41380 197316 41386 197328
rect 73798 197316 73804 197328
rect 41380 197288 73804 197316
rect 41380 197276 41386 197288
rect 73798 197276 73804 197288
rect 73856 197276 73862 197328
rect 340414 197276 340420 197328
rect 340472 197316 340478 197328
rect 369946 197316 369952 197328
rect 340472 197288 369952 197316
rect 340472 197276 340478 197288
rect 369946 197276 369952 197288
rect 370004 197276 370010 197328
rect 45370 197208 45376 197260
rect 45428 197248 45434 197260
rect 89254 197248 89260 197260
rect 45428 197220 89260 197248
rect 45428 197208 45434 197220
rect 89254 197208 89260 197220
rect 89312 197208 89318 197260
rect 340874 197208 340880 197260
rect 340932 197248 340938 197260
rect 349798 197248 349804 197260
rect 340932 197220 349804 197248
rect 340932 197208 340938 197220
rect 349798 197208 349804 197220
rect 349856 197208 349862 197260
rect 24118 197140 24124 197192
rect 24176 197180 24182 197192
rect 422294 197180 422300 197192
rect 24176 197152 422300 197180
rect 24176 197140 24182 197152
rect 422294 197140 422300 197152
rect 422352 197140 422358 197192
rect 29454 197072 29460 197124
rect 29512 197112 29518 197124
rect 412818 197112 412824 197124
rect 29512 197084 412824 197112
rect 29512 197072 29518 197084
rect 412818 197072 412824 197084
rect 412876 197072 412882 197124
rect 20070 197004 20076 197056
rect 20128 197044 20134 197056
rect 392486 197044 392492 197056
rect 20128 197016 392492 197044
rect 20128 197004 20134 197016
rect 392486 197004 392492 197016
rect 392544 197004 392550 197056
rect 82170 196936 82176 196988
rect 82228 196976 82234 196988
rect 379054 196976 379060 196988
rect 82228 196948 379060 196976
rect 82228 196936 82234 196948
rect 379054 196936 379060 196948
rect 379112 196936 379118 196988
rect 32950 196868 32956 196920
rect 33008 196908 33014 196920
rect 295334 196908 295340 196920
rect 33008 196880 295340 196908
rect 33008 196868 33014 196880
rect 295334 196868 295340 196880
rect 295392 196868 295398 196920
rect 304350 196868 304356 196920
rect 304408 196908 304414 196920
rect 371234 196908 371240 196920
rect 304408 196880 371240 196908
rect 304408 196868 304414 196880
rect 371234 196868 371240 196880
rect 371292 196868 371298 196920
rect 21450 196800 21456 196852
rect 21508 196840 21514 196852
rect 275830 196840 275836 196852
rect 21508 196812 275836 196840
rect 21508 196800 21514 196812
rect 275830 196800 275836 196812
rect 275888 196800 275894 196852
rect 276658 196800 276664 196852
rect 276716 196840 276722 196852
rect 352558 196840 352564 196852
rect 276716 196812 352564 196840
rect 276716 196800 276722 196812
rect 352558 196800 352564 196812
rect 352616 196800 352622 196852
rect 24302 196732 24308 196784
rect 24360 196772 24366 196784
rect 246390 196772 246396 196784
rect 24360 196744 246396 196772
rect 24360 196732 24366 196744
rect 246390 196732 246396 196744
rect 246448 196732 246454 196784
rect 266078 196732 266084 196784
rect 266136 196772 266142 196784
rect 351270 196772 351276 196784
rect 266136 196744 351276 196772
rect 266136 196732 266142 196744
rect 351270 196732 351276 196744
rect 351328 196732 351334 196784
rect 42242 196664 42248 196716
rect 42300 196704 42306 196716
rect 220354 196704 220360 196716
rect 42300 196676 220360 196704
rect 42300 196664 42306 196676
rect 220354 196664 220360 196676
rect 220412 196664 220418 196716
rect 227714 196664 227720 196716
rect 227772 196704 227778 196716
rect 361574 196704 361580 196716
rect 227772 196676 361580 196704
rect 227772 196664 227778 196676
rect 361574 196664 361580 196676
rect 361632 196664 361638 196716
rect 34238 196596 34244 196648
rect 34296 196636 34302 196648
rect 75638 196636 75644 196648
rect 34296 196608 75644 196636
rect 34296 196596 34302 196608
rect 75638 196596 75644 196608
rect 75696 196596 75702 196648
rect 80146 196596 80152 196648
rect 80204 196636 80210 196648
rect 556982 196636 556988 196648
rect 80204 196608 556988 196636
rect 80204 196596 80210 196608
rect 556982 196596 556988 196608
rect 557040 196596 557046 196648
rect 36722 196528 36728 196580
rect 36780 196568 36786 196580
rect 135254 196568 135260 196580
rect 36780 196540 135260 196568
rect 36780 196528 36786 196540
rect 135254 196528 135260 196540
rect 135312 196528 135318 196580
rect 182634 196528 182640 196580
rect 182692 196568 182698 196580
rect 354766 196568 354772 196580
rect 182692 196540 354772 196568
rect 182692 196528 182698 196540
rect 354766 196528 354772 196540
rect 354824 196528 354830 196580
rect 40586 196460 40592 196512
rect 40644 196500 40650 196512
rect 125042 196500 125048 196512
rect 40644 196472 125048 196500
rect 40644 196460 40650 196472
rect 125042 196460 125048 196472
rect 125100 196460 125106 196512
rect 28442 196392 28448 196444
rect 28500 196432 28506 196444
rect 551462 196432 551468 196444
rect 28500 196404 551468 196432
rect 28500 196392 28506 196404
rect 551462 196392 551468 196404
rect 551520 196392 551526 196444
rect 36630 196324 36636 196376
rect 36688 196364 36694 196376
rect 463694 196364 463700 196376
rect 36688 196336 463700 196364
rect 36688 196324 36694 196336
rect 463694 196324 463700 196336
rect 463752 196324 463758 196376
rect 32398 195916 32404 195968
rect 32456 195956 32462 195968
rect 519078 195956 519084 195968
rect 32456 195928 519084 195956
rect 32456 195916 32462 195928
rect 519078 195916 519084 195928
rect 519136 195916 519142 195968
rect 30834 195848 30840 195900
rect 30892 195888 30898 195900
rect 465074 195888 465080 195900
rect 30892 195860 465080 195888
rect 30892 195848 30898 195860
rect 465074 195848 465080 195860
rect 465132 195848 465138 195900
rect 39942 195780 39948 195832
rect 40000 195820 40006 195832
rect 121454 195820 121460 195832
rect 40000 195792 121460 195820
rect 40000 195780 40006 195792
rect 121454 195780 121460 195792
rect 121512 195780 121518 195832
rect 138198 195780 138204 195832
rect 138256 195820 138262 195832
rect 569310 195820 569316 195832
rect 138256 195792 569316 195820
rect 138256 195780 138262 195792
rect 569310 195780 569316 195792
rect 569368 195780 569374 195832
rect 52270 195712 52276 195764
rect 52328 195752 52334 195764
rect 128446 195752 128452 195764
rect 52328 195724 128452 195752
rect 52328 195712 52334 195724
rect 128446 195712 128452 195724
rect 128504 195712 128510 195764
rect 174262 195712 174268 195764
rect 174320 195752 174326 195764
rect 549530 195752 549536 195764
rect 174320 195724 549536 195752
rect 174320 195712 174326 195724
rect 549530 195712 549536 195724
rect 549588 195712 549594 195764
rect 28074 195644 28080 195696
rect 28132 195684 28138 195696
rect 395522 195684 395528 195696
rect 28132 195656 395528 195684
rect 28132 195644 28138 195656
rect 395522 195644 395528 195656
rect 395580 195644 395586 195696
rect 40770 195576 40776 195628
rect 40828 195616 40834 195628
rect 228358 195616 228364 195628
rect 40828 195588 228364 195616
rect 40828 195576 40834 195588
rect 228358 195576 228364 195588
rect 228416 195576 228422 195628
rect 312722 195576 312728 195628
rect 312780 195616 312786 195628
rect 573266 195616 573272 195628
rect 312780 195588 573272 195616
rect 312780 195576 312786 195588
rect 573266 195576 573272 195588
rect 573324 195576 573330 195628
rect 38378 195508 38384 195560
rect 38436 195548 38442 195560
rect 86402 195548 86408 195560
rect 38436 195520 86408 195548
rect 38436 195508 38442 195520
rect 86402 195508 86408 195520
rect 86460 195508 86466 195560
rect 116946 195508 116952 195560
rect 117004 195548 117010 195560
rect 363874 195548 363880 195560
rect 117004 195520 363880 195548
rect 117004 195508 117010 195520
rect 363874 195508 363880 195520
rect 363932 195508 363938 195560
rect 54754 195440 54760 195492
rect 54812 195480 54818 195492
rect 247678 195480 247684 195492
rect 54812 195452 247684 195480
rect 54812 195440 54818 195452
rect 247678 195440 247684 195452
rect 247736 195440 247742 195492
rect 266906 195480 266912 195492
rect 258046 195452 266912 195480
rect 50890 195372 50896 195424
rect 50948 195412 50954 195424
rect 258046 195412 258074 195452
rect 266906 195440 266912 195452
rect 266964 195440 266970 195492
rect 281166 195440 281172 195492
rect 281224 195480 281230 195492
rect 348970 195480 348976 195492
rect 281224 195452 348976 195480
rect 281224 195440 281230 195452
rect 348970 195440 348976 195452
rect 349028 195440 349034 195492
rect 50948 195384 258074 195412
rect 50948 195372 50954 195384
rect 259454 195372 259460 195424
rect 259512 195412 259518 195424
rect 260558 195412 260564 195424
rect 259512 195384 260564 195412
rect 259512 195372 259518 195384
rect 260558 195372 260564 195384
rect 260616 195372 260622 195424
rect 293954 195372 293960 195424
rect 294012 195412 294018 195424
rect 294690 195412 294696 195424
rect 294012 195384 294696 195412
rect 294012 195372 294018 195384
rect 294690 195372 294696 195384
rect 294748 195372 294754 195424
rect 297910 195372 297916 195424
rect 297968 195412 297974 195424
rect 356606 195412 356612 195424
rect 297968 195384 356612 195412
rect 297968 195372 297974 195384
rect 356606 195372 356612 195384
rect 356664 195372 356670 195424
rect 55582 195304 55588 195356
rect 55640 195344 55646 195356
rect 350350 195344 350356 195356
rect 55640 195316 350356 195344
rect 55640 195304 55646 195316
rect 350350 195304 350356 195316
rect 350408 195304 350414 195356
rect 46750 195236 46756 195288
rect 46808 195276 46814 195288
rect 452838 195276 452844 195288
rect 46808 195248 452844 195276
rect 46808 195236 46814 195248
rect 452838 195236 452844 195248
rect 452896 195236 452902 195288
rect 551922 195236 551928 195288
rect 551980 195276 551986 195288
rect 556798 195276 556804 195288
rect 551980 195248 556804 195276
rect 551980 195236 551986 195248
rect 556798 195236 556804 195248
rect 556856 195236 556862 195288
rect 42150 195168 42156 195220
rect 42208 195208 42214 195220
rect 175918 195208 175924 195220
rect 42208 195180 175924 195208
rect 42208 195168 42214 195180
rect 175918 195168 175924 195180
rect 175976 195168 175982 195220
rect 204530 195168 204536 195220
rect 204588 195208 204594 195220
rect 361850 195208 361856 195220
rect 204588 195180 361856 195208
rect 204588 195168 204594 195180
rect 361850 195168 361856 195180
rect 361908 195168 361914 195220
rect 35526 195100 35532 195152
rect 35584 195140 35590 195152
rect 69014 195140 69020 195152
rect 35584 195112 69020 195140
rect 35584 195100 35590 195112
rect 69014 195100 69020 195112
rect 69072 195100 69078 195152
rect 78674 195100 78680 195152
rect 78732 195140 78738 195152
rect 79594 195140 79600 195152
rect 78732 195112 79600 195140
rect 78732 195100 78738 195112
rect 79594 195100 79600 195112
rect 79652 195100 79658 195152
rect 80054 195100 80060 195152
rect 80112 195140 80118 195152
rect 80790 195140 80796 195152
rect 80112 195112 80796 195140
rect 80112 195100 80118 195112
rect 80790 195100 80796 195112
rect 80848 195100 80854 195152
rect 111794 195100 111800 195152
rect 111852 195140 111858 195152
rect 113082 195140 113088 195152
rect 111852 195112 113088 195140
rect 111852 195100 111858 195112
rect 113082 195100 113088 195112
rect 113140 195100 113146 195152
rect 113174 195100 113180 195152
rect 113232 195140 113238 195152
rect 114278 195140 114284 195152
rect 113232 195112 114284 195140
rect 113232 195100 113238 195112
rect 114278 195100 114284 195112
rect 114336 195100 114342 195152
rect 150526 195100 150532 195152
rect 150584 195140 150590 195152
rect 151722 195140 151728 195152
rect 150584 195112 151728 195140
rect 150584 195100 150590 195112
rect 151722 195100 151728 195112
rect 151780 195100 151786 195152
rect 160094 195100 160100 195152
rect 160152 195140 160158 195152
rect 161382 195140 161388 195152
rect 160152 195112 161388 195140
rect 160152 195100 160158 195112
rect 161382 195100 161388 195112
rect 161440 195100 161446 195152
rect 179506 195100 179512 195152
rect 179564 195140 179570 195152
rect 180702 195140 180708 195152
rect 179564 195112 180708 195140
rect 179564 195100 179570 195112
rect 180702 195100 180708 195112
rect 180760 195100 180766 195152
rect 209774 195100 209780 195152
rect 209832 195140 209838 195152
rect 210970 195140 210976 195152
rect 209832 195112 210976 195140
rect 209832 195100 209838 195112
rect 210970 195100 210976 195112
rect 211028 195100 211034 195152
rect 238754 195100 238760 195152
rect 238812 195140 238818 195152
rect 239950 195140 239956 195152
rect 238812 195112 239956 195140
rect 238812 195100 238818 195112
rect 239950 195100 239956 195112
rect 240008 195100 240014 195152
rect 324314 195100 324320 195152
rect 324372 195140 324378 195152
rect 324866 195140 324872 195152
rect 324372 195112 324872 195140
rect 324372 195100 324378 195112
rect 324866 195100 324872 195112
rect 324924 195100 324930 195152
rect 325694 195100 325700 195152
rect 325752 195140 325758 195152
rect 326890 195140 326896 195152
rect 325752 195112 326896 195140
rect 325752 195100 325758 195112
rect 326890 195100 326896 195112
rect 326948 195100 326954 195152
rect 333974 195100 333980 195152
rect 334032 195140 334038 195152
rect 335262 195140 335268 195152
rect 334032 195112 335268 195140
rect 334032 195100 334038 195112
rect 335262 195100 335268 195112
rect 335320 195100 335326 195152
rect 342714 195100 342720 195152
rect 342772 195140 342778 195152
rect 355226 195140 355232 195152
rect 342772 195112 355232 195140
rect 342772 195100 342778 195112
rect 355226 195100 355232 195112
rect 355284 195100 355290 195152
rect 39758 195032 39764 195084
rect 39816 195072 39822 195084
rect 73522 195072 73528 195084
rect 39816 195044 73528 195072
rect 39816 195032 39822 195044
rect 73522 195032 73528 195044
rect 73580 195032 73586 195084
rect 237374 194896 237380 194948
rect 237432 194936 237438 194948
rect 238570 194936 238576 194948
rect 237432 194908 238576 194936
rect 237432 194896 237438 194908
rect 238570 194896 238576 194908
rect 238628 194896 238634 194948
rect 20438 194488 20444 194540
rect 20496 194528 20502 194540
rect 572162 194528 572168 194540
rect 20496 194500 572168 194528
rect 20496 194488 20502 194500
rect 572162 194488 572168 194500
rect 572220 194488 572226 194540
rect 25314 194420 25320 194472
rect 25372 194460 25378 194472
rect 566458 194460 566464 194472
rect 25372 194432 566464 194460
rect 25372 194420 25378 194432
rect 566458 194420 566464 194432
rect 566516 194420 566522 194472
rect 25406 194352 25412 194404
rect 25464 194392 25470 194404
rect 566366 194392 566372 194404
rect 25464 194364 566372 194392
rect 25464 194352 25470 194364
rect 566366 194352 566372 194364
rect 566424 194352 566430 194404
rect 142062 194284 142068 194336
rect 142120 194324 142126 194336
rect 529934 194324 529940 194336
rect 142120 194296 529940 194324
rect 142120 194284 142126 194296
rect 529934 194284 529940 194296
rect 529992 194284 529998 194336
rect 181346 194216 181352 194268
rect 181404 194256 181410 194268
rect 449894 194256 449900 194268
rect 181404 194228 449900 194256
rect 181404 194216 181410 194228
rect 449894 194216 449900 194228
rect 449952 194216 449958 194268
rect 17218 194148 17224 194200
rect 17276 194188 17282 194200
rect 281718 194188 281724 194200
rect 17276 194160 281724 194188
rect 17276 194148 17282 194160
rect 281718 194148 281724 194160
rect 281776 194148 281782 194200
rect 284754 194148 284760 194200
rect 284812 194188 284818 194200
rect 364426 194188 364432 194200
rect 284812 194160 364432 194188
rect 284812 194148 284818 194160
rect 364426 194148 364432 194160
rect 364484 194148 364490 194200
rect 102134 194080 102140 194132
rect 102192 194120 102198 194132
rect 364058 194120 364064 194132
rect 102192 194092 364064 194120
rect 102192 194080 102198 194092
rect 364058 194080 364064 194092
rect 364116 194080 364122 194132
rect 249610 194012 249616 194064
rect 249668 194052 249674 194064
rect 390094 194052 390100 194064
rect 249668 194024 390100 194052
rect 249668 194012 249674 194024
rect 390094 194012 390100 194024
rect 390152 194012 390158 194064
rect 241238 193944 241244 193996
rect 241296 193984 241302 193996
rect 370774 193984 370780 193996
rect 241296 193956 370780 193984
rect 241296 193944 241302 193956
rect 370774 193944 370780 193956
rect 370832 193944 370838 193996
rect 242986 193876 242992 193928
rect 243044 193916 243050 193928
rect 365806 193916 365812 193928
rect 243044 193888 365812 193916
rect 243044 193876 243050 193888
rect 365806 193876 365812 193888
rect 365864 193876 365870 193928
rect 41138 193808 41144 193860
rect 41196 193848 41202 193860
rect 141786 193848 141792 193860
rect 41196 193820 141792 193848
rect 41196 193808 41202 193820
rect 141786 193808 141792 193820
rect 141844 193808 141850 193860
rect 318886 193808 318892 193860
rect 318944 193848 318950 193860
rect 562226 193848 562232 193860
rect 318944 193820 562232 193848
rect 318944 193808 318950 193820
rect 562226 193808 562232 193820
rect 562284 193808 562290 193860
rect 276014 193740 276020 193792
rect 276072 193780 276078 193792
rect 352190 193780 352196 193792
rect 276072 193752 352196 193780
rect 276072 193740 276078 193752
rect 352190 193740 352196 193752
rect 352248 193740 352254 193792
rect 280522 193672 280528 193724
rect 280580 193712 280586 193724
rect 351178 193712 351184 193724
rect 280580 193684 351184 193712
rect 280580 193672 280586 193684
rect 351178 193672 351184 193684
rect 351236 193672 351242 193724
rect 287974 193604 287980 193656
rect 288032 193644 288038 193656
rect 358354 193644 358360 193656
rect 288032 193616 358360 193644
rect 288032 193604 288038 193616
rect 358354 193604 358360 193616
rect 358412 193604 358418 193656
rect 26694 193128 26700 193180
rect 26752 193168 26758 193180
rect 478874 193168 478880 193180
rect 26752 193140 478880 193168
rect 26752 193128 26758 193140
rect 478874 193128 478880 193140
rect 478932 193128 478938 193180
rect 49602 193060 49608 193112
rect 49660 193100 49666 193112
rect 189074 193100 189080 193112
rect 49660 193072 189080 193100
rect 49660 193060 49666 193072
rect 189074 193060 189080 193072
rect 189132 193060 189138 193112
rect 205174 193060 205180 193112
rect 205232 193100 205238 193112
rect 575658 193100 575664 193112
rect 205232 193072 575664 193100
rect 205232 193060 205238 193072
rect 575658 193060 575664 193072
rect 575716 193060 575722 193112
rect 34146 192992 34152 193044
rect 34204 193032 34210 193044
rect 337838 193032 337844 193044
rect 34204 193004 337844 193032
rect 34204 192992 34210 193004
rect 337838 192992 337844 193004
rect 337896 192992 337902 193044
rect 39666 192924 39672 192976
rect 39724 192964 39730 192976
rect 87690 192964 87696 192976
rect 39724 192936 87696 192964
rect 39724 192924 39730 192936
rect 87690 192924 87696 192936
rect 87748 192924 87754 192976
rect 134334 192924 134340 192976
rect 134392 192964 134398 192976
rect 346302 192964 346308 192976
rect 134392 192936 346308 192964
rect 134392 192924 134398 192936
rect 346302 192924 346308 192936
rect 346360 192924 346366 192976
rect 36906 192856 36912 192908
rect 36964 192896 36970 192908
rect 154298 192896 154304 192908
rect 36964 192868 154304 192896
rect 36964 192856 36970 192868
rect 154298 192856 154304 192868
rect 154356 192856 154362 192908
rect 173618 192856 173624 192908
rect 173676 192896 173682 192908
rect 361758 192896 361764 192908
rect 173676 192868 361764 192896
rect 173676 192856 173682 192868
rect 361758 192856 361764 192868
rect 361816 192856 361822 192908
rect 51442 192788 51448 192840
rect 51500 192828 51506 192840
rect 194870 192828 194876 192840
rect 51500 192800 194876 192828
rect 51500 192788 51506 192800
rect 194870 192788 194876 192800
rect 194928 192788 194934 192840
rect 217778 192788 217784 192840
rect 217836 192828 217842 192840
rect 349246 192828 349252 192840
rect 217836 192800 349252 192828
rect 217836 192788 217842 192800
rect 349246 192788 349252 192800
rect 349304 192788 349310 192840
rect 45462 192720 45468 192772
rect 45520 192760 45526 192772
rect 243078 192760 243084 192772
rect 45520 192732 243084 192760
rect 45520 192720 45526 192732
rect 243078 192720 243084 192732
rect 243136 192720 243142 192772
rect 48958 192652 48964 192704
rect 49016 192692 49022 192704
rect 263778 192692 263784 192704
rect 49016 192664 263784 192692
rect 49016 192652 49022 192664
rect 263778 192652 263784 192664
rect 263836 192652 263842 192704
rect 54202 192584 54208 192636
rect 54260 192624 54266 192636
rect 355134 192624 355140 192636
rect 54260 192596 355140 192624
rect 54260 192584 54266 192596
rect 355134 192584 355140 192596
rect 355192 192584 355198 192636
rect 50798 192516 50804 192568
rect 50856 192556 50862 192568
rect 356146 192556 356152 192568
rect 50856 192528 356152 192556
rect 50856 192516 50862 192528
rect 356146 192516 356152 192528
rect 356204 192516 356210 192568
rect 4798 192448 4804 192500
rect 4856 192488 4862 192500
rect 506566 192488 506572 192500
rect 4856 192460 506572 192488
rect 4856 192448 4862 192460
rect 506566 192448 506572 192460
rect 506624 192448 506630 192500
rect 49970 192380 49976 192432
rect 50028 192420 50034 192432
rect 172974 192420 172980 192432
rect 50028 192392 172980 192420
rect 50028 192380 50034 192392
rect 172974 192380 172980 192392
rect 173032 192380 173038 192432
rect 46842 192312 46848 192364
rect 46900 192352 46906 192364
rect 151814 192352 151820 192364
rect 46900 192324 151820 192352
rect 46900 192312 46906 192324
rect 151814 192312 151820 192324
rect 151872 192312 151878 192364
rect 40586 192244 40592 192296
rect 40644 192284 40650 192296
rect 85298 192284 85304 192296
rect 40644 192256 85304 192284
rect 40644 192244 40650 192256
rect 85298 192244 85304 192256
rect 85356 192244 85362 192296
rect 20162 191768 20168 191820
rect 20220 191808 20226 191820
rect 574462 191808 574468 191820
rect 20220 191780 574468 191808
rect 20220 191768 20226 191780
rect 574462 191768 574468 191780
rect 574520 191768 574526 191820
rect 17310 191700 17316 191752
rect 17368 191740 17374 191752
rect 391106 191740 391112 191752
rect 17368 191712 391112 191740
rect 17368 191700 17374 191712
rect 391106 191700 391112 191712
rect 391164 191700 391170 191752
rect 184566 191632 184572 191684
rect 184624 191672 184630 191684
rect 359274 191672 359280 191684
rect 184624 191644 359280 191672
rect 184624 191632 184630 191644
rect 359274 191632 359280 191644
rect 359332 191632 359338 191684
rect 300854 191428 300860 191480
rect 300912 191468 300918 191480
rect 348050 191468 348056 191480
rect 300912 191440 348056 191468
rect 300912 191428 300918 191440
rect 348050 191428 348056 191440
rect 348108 191428 348114 191480
rect 44634 191360 44640 191412
rect 44692 191400 44698 191412
rect 202966 191400 202972 191412
rect 44692 191372 202972 191400
rect 44692 191360 44698 191372
rect 202966 191360 202972 191372
rect 203024 191360 203030 191412
rect 285398 191360 285404 191412
rect 285456 191400 285462 191412
rect 353478 191400 353484 191412
rect 285456 191372 353484 191400
rect 285456 191360 285462 191372
rect 353478 191360 353484 191372
rect 353536 191360 353542 191412
rect 61562 191292 61568 191344
rect 61620 191332 61626 191344
rect 307938 191332 307944 191344
rect 61620 191304 307944 191332
rect 61620 191292 61626 191304
rect 307938 191292 307944 191304
rect 307996 191292 308002 191344
rect 98638 191224 98644 191276
rect 98696 191264 98702 191276
rect 366082 191264 366088 191276
rect 98696 191236 366088 191264
rect 98696 191224 98702 191236
rect 366082 191224 366088 191236
rect 366140 191224 366146 191276
rect 46842 191156 46848 191208
rect 46900 191196 46906 191208
rect 333330 191196 333336 191208
rect 46900 191168 333336 191196
rect 46900 191156 46906 191168
rect 333330 191156 333336 191168
rect 333388 191156 333394 191208
rect 339494 191156 339500 191208
rect 339552 191196 339558 191208
rect 350994 191196 351000 191208
rect 339552 191168 351000 191196
rect 339552 191156 339558 191168
rect 350994 191156 351000 191168
rect 351052 191156 351058 191208
rect 49418 191088 49424 191140
rect 49476 191128 49482 191140
rect 472158 191128 472164 191140
rect 49476 191100 472164 191128
rect 49476 191088 49482 191100
rect 472158 191088 472164 191100
rect 472216 191088 472222 191140
rect 20346 190408 20352 190460
rect 20404 190448 20410 190460
rect 578786 190448 578792 190460
rect 20404 190420 578792 190448
rect 20404 190408 20410 190420
rect 578786 190408 578792 190420
rect 578844 190408 578850 190460
rect 42058 190340 42064 190392
rect 42116 190380 42122 190392
rect 275738 190380 275744 190392
rect 42116 190352 275744 190380
rect 42116 190340 42122 190352
rect 275738 190340 275744 190352
rect 275796 190340 275802 190392
rect 58802 190272 58808 190324
rect 58860 190312 58866 190324
rect 341058 190312 341064 190324
rect 58860 190284 341064 190312
rect 58860 190272 58866 190284
rect 341058 190272 341064 190284
rect 341116 190272 341122 190324
rect 55950 190204 55956 190256
rect 56008 190244 56014 190256
rect 349614 190244 349620 190256
rect 56008 190216 349620 190244
rect 56008 190204 56014 190216
rect 349614 190204 349620 190216
rect 349672 190204 349678 190256
rect 42242 190136 42248 190188
rect 42300 190176 42306 190188
rect 380710 190176 380716 190188
rect 42300 190148 380716 190176
rect 42300 190136 42306 190148
rect 380710 190136 380716 190148
rect 380768 190136 380774 190188
rect 41322 190068 41328 190120
rect 41380 190108 41386 190120
rect 392394 190108 392400 190120
rect 41380 190080 392400 190108
rect 41380 190068 41386 190080
rect 392394 190068 392400 190080
rect 392452 190068 392458 190120
rect 55030 190000 55036 190052
rect 55088 190040 55094 190052
rect 409966 190040 409972 190052
rect 55088 190012 409972 190040
rect 55088 190000 55094 190012
rect 409966 190000 409972 190012
rect 410024 190000 410030 190052
rect 34146 189932 34152 189984
rect 34204 189972 34210 189984
rect 169110 189972 169116 189984
rect 34204 189944 169116 189972
rect 34204 189932 34210 189944
rect 169110 189932 169116 189944
rect 169168 189932 169174 189984
rect 174630 189932 174636 189984
rect 174688 189972 174694 189984
rect 560846 189972 560852 189984
rect 174688 189944 560852 189972
rect 174688 189932 174694 189944
rect 560846 189932 560852 189944
rect 560904 189932 560910 189984
rect 85758 189864 85764 189916
rect 85816 189904 85822 189916
rect 556890 189904 556896 189916
rect 85816 189876 556896 189904
rect 85816 189864 85822 189876
rect 556890 189864 556896 189876
rect 556948 189864 556954 189916
rect 19334 189796 19340 189848
rect 19392 189836 19398 189848
rect 556430 189836 556436 189848
rect 19392 189808 556436 189836
rect 19392 189796 19398 189808
rect 556430 189796 556436 189808
rect 556488 189796 556494 189848
rect 3510 189728 3516 189780
rect 3568 189768 3574 189780
rect 567378 189768 567384 189780
rect 3568 189740 567384 189768
rect 3568 189728 3574 189740
rect 567378 189728 567384 189740
rect 567436 189728 567442 189780
rect 43806 189660 43812 189712
rect 43864 189700 43870 189712
rect 216122 189700 216128 189712
rect 43864 189672 216128 189700
rect 43864 189660 43870 189672
rect 216122 189660 216128 189672
rect 216180 189660 216186 189712
rect 59446 189592 59452 189644
rect 59504 189632 59510 189644
rect 226426 189632 226432 189644
rect 59504 189604 226432 189632
rect 59504 189592 59510 189604
rect 226426 189592 226432 189604
rect 226484 189592 226490 189644
rect 183922 188980 183928 189032
rect 183980 189020 183986 189032
rect 582834 189020 582840 189032
rect 183980 188992 582840 189020
rect 183980 188980 183986 188992
rect 582834 188980 582840 188992
rect 582892 188980 582898 189032
rect 3418 188912 3424 188964
rect 3476 188952 3482 188964
rect 396902 188952 396908 188964
rect 3476 188924 396908 188952
rect 3476 188912 3482 188924
rect 396902 188912 396908 188924
rect 396960 188912 396966 188964
rect 169754 188844 169760 188896
rect 169812 188884 169818 188896
rect 356514 188884 356520 188896
rect 169812 188856 356520 188884
rect 169812 188844 169818 188856
rect 356514 188844 356520 188856
rect 356572 188844 356578 188896
rect 293126 188368 293132 188420
rect 293184 188408 293190 188420
rect 352742 188408 352748 188420
rect 293184 188380 352748 188408
rect 293184 188368 293190 188380
rect 352742 188368 352748 188380
rect 352800 188368 352806 188420
rect 221274 188300 221280 188352
rect 221332 188340 221338 188352
rect 252646 188340 252652 188352
rect 221332 188312 252652 188340
rect 221332 188300 221338 188312
rect 252646 188300 252652 188312
rect 252704 188300 252710 188352
rect 296346 188300 296352 188352
rect 296404 188340 296410 188352
rect 379330 188340 379336 188352
rect 296404 188312 379336 188340
rect 296404 188300 296410 188312
rect 379330 188300 379336 188312
rect 379388 188300 379394 188352
rect 38194 187620 38200 187672
rect 38252 187660 38258 187672
rect 179506 187660 179512 187672
rect 38252 187632 179512 187660
rect 38252 187620 38258 187632
rect 179506 187620 179512 187632
rect 179564 187620 179570 187672
rect 192018 187620 192024 187672
rect 192076 187660 192082 187672
rect 360654 187660 360660 187672
rect 192076 187632 360660 187660
rect 192076 187620 192082 187632
rect 360654 187620 360660 187632
rect 360712 187620 360718 187672
rect 53466 187552 53472 187604
rect 53524 187592 53530 187604
rect 236730 187592 236736 187604
rect 53524 187564 236736 187592
rect 53524 187552 53530 187564
rect 236730 187552 236736 187564
rect 236788 187552 236794 187604
rect 322106 187552 322112 187604
rect 322164 187592 322170 187604
rect 559742 187592 559748 187604
rect 322164 187564 559748 187592
rect 322164 187552 322170 187564
rect 559742 187552 559748 187564
rect 559800 187552 559806 187604
rect 99926 187484 99932 187536
rect 99984 187524 99990 187536
rect 370682 187524 370688 187536
rect 99984 187496 370688 187524
rect 99984 187484 99990 187496
rect 370682 187484 370688 187496
rect 370740 187484 370746 187536
rect 58710 187416 58716 187468
rect 58768 187456 58774 187468
rect 357710 187456 357716 187468
rect 58768 187428 357716 187456
rect 58768 187416 58774 187428
rect 357710 187416 357716 187428
rect 357768 187416 357774 187468
rect 53558 187348 53564 187400
rect 53616 187388 53622 187400
rect 354214 187388 354220 187400
rect 53616 187360 354220 187388
rect 53616 187348 53622 187360
rect 354214 187348 354220 187360
rect 354272 187348 354278 187400
rect 59722 187280 59728 187332
rect 59780 187320 59786 187332
rect 363046 187320 363052 187332
rect 59780 187292 363052 187320
rect 59780 187280 59786 187292
rect 363046 187280 363052 187292
rect 363104 187280 363110 187332
rect 35526 187212 35532 187264
rect 35584 187252 35590 187264
rect 349522 187252 349528 187264
rect 35584 187224 349528 187252
rect 35584 187212 35590 187224
rect 349522 187212 349528 187224
rect 349580 187212 349586 187264
rect 38286 187144 38292 187196
rect 38344 187184 38350 187196
rect 370590 187184 370596 187196
rect 38344 187156 370596 187184
rect 38344 187144 38350 187156
rect 370590 187144 370596 187156
rect 370648 187144 370654 187196
rect 36538 187076 36544 187128
rect 36596 187116 36602 187128
rect 371326 187116 371332 187128
rect 36596 187088 371332 187116
rect 36596 187076 36602 187088
rect 371326 187076 371332 187088
rect 371384 187076 371390 187128
rect 34330 187008 34336 187060
rect 34388 187048 34394 187060
rect 377674 187048 377680 187060
rect 34388 187020 377680 187048
rect 34388 187008 34394 187020
rect 377674 187008 377680 187020
rect 377732 187008 377738 187060
rect 33686 186940 33692 186992
rect 33744 186980 33750 186992
rect 490190 186980 490196 186992
rect 33744 186952 490196 186980
rect 33744 186940 33750 186952
rect 490190 186940 490196 186952
rect 490248 186940 490254 186992
rect 239030 186872 239036 186924
rect 239088 186912 239094 186924
rect 353754 186912 353760 186924
rect 239088 186884 353760 186912
rect 239088 186872 239094 186884
rect 353754 186872 353760 186884
rect 353812 186872 353818 186924
rect 278958 186124 278964 186176
rect 279016 186164 279022 186176
rect 366726 186164 366732 186176
rect 279016 186136 366732 186164
rect 279016 186124 279022 186136
rect 366726 186124 366732 186136
rect 366784 186124 366790 186176
rect 187510 186056 187516 186108
rect 187568 186096 187574 186108
rect 354122 186096 354128 186108
rect 187568 186068 354128 186096
rect 187568 186056 187574 186068
rect 354122 186056 354128 186068
rect 354180 186056 354186 186108
rect 116670 185988 116676 186040
rect 116728 186028 116734 186040
rect 351454 186028 351460 186040
rect 116728 186000 351460 186028
rect 116728 185988 116734 186000
rect 351454 185988 351460 186000
rect 351512 185988 351518 186040
rect 58250 185920 58256 185972
rect 58308 185960 58314 185972
rect 303706 185960 303712 185972
rect 58308 185932 303712 185960
rect 58308 185920 58314 185932
rect 303706 185920 303712 185932
rect 303764 185920 303770 185972
rect 53374 185852 53380 185904
rect 53432 185892 53438 185904
rect 356422 185892 356428 185904
rect 53432 185864 356428 185892
rect 53432 185852 53438 185864
rect 356422 185852 356428 185864
rect 356480 185852 356486 185904
rect 40770 185784 40776 185836
rect 40828 185824 40834 185836
rect 359366 185824 359372 185836
rect 40828 185796 359372 185824
rect 40828 185784 40834 185796
rect 359366 185784 359372 185796
rect 359424 185784 359430 185836
rect 42150 185716 42156 185768
rect 42208 185756 42214 185768
rect 381630 185756 381636 185768
rect 42208 185728 381636 185756
rect 42208 185716 42214 185728
rect 381630 185716 381636 185728
rect 381688 185716 381694 185768
rect 407114 185716 407120 185768
rect 407172 185756 407178 185768
rect 438854 185756 438860 185768
rect 407172 185728 438860 185756
rect 407172 185716 407178 185728
rect 438854 185716 438860 185728
rect 438912 185716 438918 185768
rect 222286 185648 222292 185700
rect 222344 185688 222350 185700
rect 561858 185688 561864 185700
rect 222344 185660 561864 185688
rect 222344 185648 222350 185660
rect 561858 185648 561864 185660
rect 561916 185648 561922 185700
rect 55858 185580 55864 185632
rect 55916 185620 55922 185632
rect 408034 185620 408040 185632
rect 55916 185592 408040 185620
rect 55916 185580 55922 185592
rect 408034 185580 408040 185592
rect 408092 185580 408098 185632
rect 194962 184832 194968 184884
rect 195020 184872 195026 184884
rect 201494 184872 201500 184884
rect 195020 184844 201500 184872
rect 195020 184832 195026 184844
rect 201494 184832 201500 184844
rect 201552 184832 201558 184884
rect 216490 184832 216496 184884
rect 216548 184872 216554 184884
rect 347774 184872 347780 184884
rect 216548 184844 347780 184872
rect 216548 184832 216554 184844
rect 347774 184832 347780 184844
rect 347832 184832 347838 184884
rect 209866 184764 209872 184816
rect 209924 184804 209930 184816
rect 352834 184804 352840 184816
rect 209924 184776 352840 184804
rect 209924 184764 209930 184776
rect 352834 184764 352840 184776
rect 352892 184764 352898 184816
rect 159174 184696 159180 184748
rect 159232 184736 159238 184748
rect 352374 184736 352380 184748
rect 159232 184708 352380 184736
rect 159232 184696 159238 184708
rect 352374 184696 352380 184708
rect 352432 184696 352438 184748
rect 146938 184628 146944 184680
rect 146996 184668 147002 184680
rect 351086 184668 351092 184680
rect 146996 184640 351092 184668
rect 146996 184628 147002 184640
rect 351086 184628 351092 184640
rect 351144 184628 351150 184680
rect 37826 184560 37832 184612
rect 37884 184600 37890 184612
rect 245470 184600 245476 184612
rect 37884 184572 245476 184600
rect 37884 184560 37890 184572
rect 245470 184560 245476 184572
rect 245528 184560 245534 184612
rect 272518 184560 272524 184612
rect 272576 184600 272582 184612
rect 383654 184600 383660 184612
rect 272576 184572 383660 184600
rect 272576 184560 272582 184572
rect 383654 184560 383660 184572
rect 383712 184560 383718 184612
rect 59814 184492 59820 184544
rect 59872 184532 59878 184544
rect 355042 184532 355048 184544
rect 59872 184504 355048 184532
rect 59872 184492 59878 184504
rect 355042 184492 355048 184504
rect 355100 184492 355106 184544
rect 59630 184424 59636 184476
rect 59688 184464 59694 184476
rect 357434 184464 357440 184476
rect 59688 184436 357440 184464
rect 59688 184424 59694 184436
rect 357434 184424 357440 184436
rect 357492 184424 357498 184476
rect 59078 184356 59084 184408
rect 59136 184396 59142 184408
rect 363414 184396 363420 184408
rect 59136 184368 363420 184396
rect 59136 184356 59142 184368
rect 363414 184356 363420 184368
rect 363472 184356 363478 184408
rect 40954 184288 40960 184340
rect 41012 184328 41018 184340
rect 183002 184328 183008 184340
rect 41012 184300 183008 184328
rect 41012 184288 41018 184300
rect 183002 184288 183008 184300
rect 183060 184288 183066 184340
rect 234522 184288 234528 184340
rect 234580 184328 234586 184340
rect 560570 184328 560576 184340
rect 234580 184300 560576 184328
rect 234580 184288 234586 184300
rect 560570 184288 560576 184300
rect 560628 184288 560634 184340
rect 35710 184220 35716 184272
rect 35768 184260 35774 184272
rect 367278 184260 367284 184272
rect 35768 184232 367284 184260
rect 35768 184220 35774 184232
rect 367278 184220 367284 184232
rect 367336 184220 367342 184272
rect 36630 184152 36636 184204
rect 36688 184192 36694 184204
rect 371418 184192 371424 184204
rect 36688 184164 371424 184192
rect 36688 184152 36694 184164
rect 371418 184152 371424 184164
rect 371476 184152 371482 184204
rect 249978 184084 249984 184136
rect 250036 184124 250042 184136
rect 352282 184124 352288 184136
rect 250036 184096 352288 184124
rect 250036 184084 250042 184096
rect 352282 184084 352288 184096
rect 352340 184084 352346 184136
rect 283466 184016 283472 184068
rect 283524 184056 283530 184068
rect 347498 184056 347504 184068
rect 283524 184028 347504 184056
rect 283524 184016 283530 184028
rect 347498 184016 347504 184028
rect 347556 184016 347562 184068
rect 163038 183472 163044 183524
rect 163096 183512 163102 183524
rect 348878 183512 348884 183524
rect 163096 183484 348884 183512
rect 163096 183472 163102 183484
rect 348878 183472 348884 183484
rect 348936 183472 348942 183524
rect 52178 183404 52184 183456
rect 52236 183444 52242 183456
rect 358998 183444 359004 183456
rect 52236 183416 359004 183444
rect 52236 183404 52242 183416
rect 358998 183404 359004 183416
rect 359056 183404 359062 183456
rect 398834 183404 398840 183456
rect 398892 183444 398898 183456
rect 402514 183444 402520 183456
rect 398892 183416 402520 183444
rect 398892 183404 398898 183416
rect 402514 183404 402520 183416
rect 402572 183404 402578 183456
rect 44082 183336 44088 183388
rect 44140 183376 44146 183388
rect 353386 183376 353392 183388
rect 44140 183348 353392 183376
rect 44140 183336 44146 183348
rect 353386 183336 353392 183348
rect 353444 183336 353450 183388
rect 46014 183268 46020 183320
rect 46072 183308 46078 183320
rect 360562 183308 360568 183320
rect 46072 183280 360568 183308
rect 46072 183268 46078 183280
rect 360562 183268 360568 183280
rect 360620 183268 360626 183320
rect 393774 183268 393780 183320
rect 393832 183308 393838 183320
rect 407206 183308 407212 183320
rect 393832 183280 407212 183308
rect 393832 183268 393838 183280
rect 407206 183268 407212 183280
rect 407264 183268 407270 183320
rect 224218 183200 224224 183252
rect 224276 183240 224282 183252
rect 552474 183240 552480 183252
rect 224276 183212 552480 183240
rect 224276 183200 224282 183212
rect 552474 183200 552480 183212
rect 552532 183200 552538 183252
rect 54662 183132 54668 183184
rect 54720 183172 54726 183184
rect 399754 183172 399760 183184
rect 54720 183144 399760 183172
rect 54720 183132 54726 183144
rect 399754 183132 399760 183144
rect 399812 183132 399818 183184
rect 44726 183064 44732 183116
rect 44784 183104 44790 183116
rect 407850 183104 407856 183116
rect 44784 183076 407856 183104
rect 44784 183064 44790 183076
rect 407850 183064 407856 183076
rect 407908 183064 407914 183116
rect 39666 182996 39672 183048
rect 39724 183036 39730 183048
rect 459646 183036 459652 183048
rect 39724 183008 459652 183036
rect 39724 182996 39730 183008
rect 459646 182996 459652 183008
rect 459704 182996 459710 183048
rect 116026 182928 116032 182980
rect 116084 182968 116090 182980
rect 558178 182968 558184 182980
rect 116084 182940 558184 182968
rect 116084 182928 116090 182940
rect 558178 182928 558184 182940
rect 558236 182928 558242 182980
rect 37918 182860 37924 182912
rect 37976 182900 37982 182912
rect 529934 182900 529940 182912
rect 37976 182872 529940 182900
rect 37976 182860 37982 182872
rect 529934 182860 529940 182872
rect 529992 182860 529998 182912
rect 47854 182792 47860 182844
rect 47912 182832 47918 182844
rect 573542 182832 573548 182844
rect 47912 182804 573548 182832
rect 47912 182792 47918 182804
rect 573542 182792 573548 182804
rect 573600 182792 573606 182844
rect 246114 182724 246120 182776
rect 246172 182764 246178 182776
rect 351362 182764 351368 182776
rect 246172 182736 351368 182764
rect 246172 182724 246178 182736
rect 351362 182724 351368 182736
rect 351420 182724 351426 182776
rect 198090 182112 198096 182164
rect 198148 182152 198154 182164
rect 302142 182152 302148 182164
rect 198148 182124 302148 182152
rect 198148 182112 198154 182124
rect 302142 182112 302148 182124
rect 302200 182112 302206 182164
rect 58894 182044 58900 182096
rect 58952 182084 58958 182096
rect 364518 182084 364524 182096
rect 58952 182056 364524 182084
rect 58952 182044 58958 182056
rect 364518 182044 364524 182056
rect 364576 182044 364582 182096
rect 255774 181976 255780 182028
rect 255832 182016 255838 182028
rect 561950 182016 561956 182028
rect 255832 181988 561956 182016
rect 255832 181976 255838 181988
rect 561950 181976 561956 181988
rect 562008 181976 562014 182028
rect 54938 181908 54944 181960
rect 54996 181948 55002 181960
rect 376570 181948 376576 181960
rect 54996 181920 376576 181948
rect 54996 181908 55002 181920
rect 376570 181908 376576 181920
rect 376628 181908 376634 181960
rect 42058 181840 42064 181892
rect 42116 181880 42122 181892
rect 368934 181880 368940 181892
rect 42116 181852 368940 181880
rect 42116 181840 42122 181852
rect 368934 181840 368940 181852
rect 368992 181840 368998 181892
rect 34238 181772 34244 181824
rect 34296 181812 34302 181824
rect 373626 181812 373632 181824
rect 34296 181784 373632 181812
rect 34296 181772 34302 181784
rect 373626 181772 373632 181784
rect 373684 181772 373690 181824
rect 35618 181704 35624 181756
rect 35676 181744 35682 181756
rect 381354 181744 381360 181756
rect 35676 181716 381360 181744
rect 35676 181704 35682 181716
rect 381354 181704 381360 181716
rect 381412 181704 381418 181756
rect 37090 181636 37096 181688
rect 37148 181676 37154 181688
rect 387334 181676 387340 181688
rect 37148 181648 387340 181676
rect 37148 181636 37154 181648
rect 387334 181636 387340 181648
rect 387392 181636 387398 181688
rect 33962 181568 33968 181620
rect 34020 181608 34026 181620
rect 391290 181608 391296 181620
rect 34020 181580 391296 181608
rect 34020 181568 34026 181580
rect 391290 181568 391296 181580
rect 391348 181568 391354 181620
rect 43530 181500 43536 181552
rect 43588 181540 43594 181552
rect 412818 181540 412824 181552
rect 43588 181512 412824 181540
rect 43588 181500 43594 181512
rect 412818 181500 412824 181512
rect 412876 181500 412882 181552
rect 48866 181432 48872 181484
rect 48924 181472 48930 181484
rect 426526 181472 426532 181484
rect 48924 181444 426532 181472
rect 48924 181432 48930 181444
rect 426526 181432 426532 181444
rect 426584 181432 426590 181484
rect 576118 181432 576124 181484
rect 576176 181472 576182 181484
rect 580718 181472 580724 181484
rect 576176 181444 580724 181472
rect 576176 181432 576182 181444
rect 580718 181432 580724 181444
rect 580776 181432 580782 181484
rect 191834 180412 191840 180464
rect 191892 180452 191898 180464
rect 274450 180452 274456 180464
rect 191892 180424 274456 180452
rect 191892 180412 191898 180424
rect 274450 180412 274456 180424
rect 274508 180412 274514 180464
rect 279602 180412 279608 180464
rect 279660 180452 279666 180464
rect 357526 180452 357532 180464
rect 279660 180424 357532 180452
rect 279660 180412 279666 180424
rect 357526 180412 357532 180424
rect 357584 180412 357590 180464
rect 226794 180344 226800 180396
rect 226852 180384 226858 180396
rect 358078 180384 358084 180396
rect 226852 180356 358084 180384
rect 226852 180344 226858 180356
rect 358078 180344 358084 180356
rect 358136 180344 358142 180396
rect 69658 180276 69664 180328
rect 69716 180316 69722 180328
rect 197354 180316 197360 180328
rect 69716 180288 197360 180316
rect 69716 180276 69722 180288
rect 197354 180276 197360 180288
rect 197412 180276 197418 180328
rect 330478 180276 330484 180328
rect 330536 180316 330542 180328
rect 552566 180316 552572 180328
rect 330536 180288 552572 180316
rect 330536 180276 330542 180288
rect 552566 180276 552572 180288
rect 552624 180276 552630 180328
rect 53098 180208 53104 180260
rect 53156 180248 53162 180260
rect 65794 180248 65800 180260
rect 53156 180220 65800 180248
rect 53156 180208 53162 180220
rect 65794 180208 65800 180220
rect 65852 180208 65858 180260
rect 103790 180208 103796 180260
rect 103848 180248 103854 180260
rect 347866 180248 347872 180260
rect 103848 180220 347872 180248
rect 103848 180208 103854 180220
rect 347866 180208 347872 180220
rect 347924 180208 347930 180260
rect 59906 180140 59912 180192
rect 59964 180180 59970 180192
rect 372706 180180 372712 180192
rect 59964 180152 372712 180180
rect 59964 180140 59970 180152
rect 372706 180140 372712 180152
rect 372764 180140 372770 180192
rect 50246 180072 50252 180124
rect 50304 180112 50310 180124
rect 400766 180112 400772 180124
rect 50304 180084 400772 180112
rect 50304 180072 50310 180084
rect 400766 180072 400772 180084
rect 400824 180072 400830 180124
rect 111978 179052 111984 179104
rect 112036 179092 112042 179104
rect 130194 179092 130200 179104
rect 112036 179064 130200 179092
rect 112036 179052 112042 179064
rect 130194 179052 130200 179064
rect 130252 179052 130258 179104
rect 213914 179052 213920 179104
rect 213972 179092 213978 179104
rect 346578 179092 346584 179104
rect 213972 179064 346584 179092
rect 213972 179052 213978 179064
rect 346578 179052 346584 179064
rect 346636 179052 346642 179104
rect 41966 178984 41972 179036
rect 42024 179024 42030 179036
rect 345014 179024 345020 179036
rect 42024 178996 345020 179024
rect 42024 178984 42030 178996
rect 345014 178984 345020 178996
rect 345072 178984 345078 179036
rect 49326 178916 49332 178968
rect 49384 178956 49390 178968
rect 367370 178956 367376 178968
rect 49384 178928 367376 178956
rect 49384 178916 49390 178928
rect 367370 178916 367376 178928
rect 367428 178916 367434 178968
rect 34054 178848 34060 178900
rect 34112 178888 34118 178900
rect 401962 178888 401968 178900
rect 34112 178860 401968 178888
rect 34112 178848 34118 178860
rect 401962 178848 401968 178860
rect 402020 178848 402026 178900
rect 13814 178780 13820 178832
rect 13872 178820 13878 178832
rect 432046 178820 432052 178832
rect 13872 178792 432052 178820
rect 13872 178780 13878 178792
rect 432046 178780 432052 178792
rect 432104 178780 432110 178832
rect 40494 178712 40500 178764
rect 40552 178752 40558 178764
rect 460934 178752 460940 178764
rect 40552 178724 460940 178752
rect 40552 178712 40558 178724
rect 460934 178712 460940 178724
rect 460992 178712 460998 178764
rect 43254 178644 43260 178696
rect 43312 178684 43318 178696
rect 488626 178684 488632 178696
rect 43312 178656 488632 178684
rect 43312 178644 43318 178656
rect 488626 178644 488632 178656
rect 488684 178644 488690 178696
rect 241606 177828 241612 177880
rect 241664 177868 241670 177880
rect 375374 177868 375380 177880
rect 241664 177840 375380 177868
rect 241664 177828 241670 177840
rect 375374 177828 375380 177840
rect 375432 177828 375438 177880
rect 227714 177760 227720 177812
rect 227772 177800 227778 177812
rect 469306 177800 469312 177812
rect 227772 177772 469312 177800
rect 227772 177760 227778 177772
rect 469306 177760 469312 177772
rect 469364 177760 469370 177812
rect 74810 177692 74816 177744
rect 74868 177732 74874 177744
rect 378042 177732 378048 177744
rect 74868 177704 378048 177732
rect 74868 177692 74874 177704
rect 378042 177692 378048 177704
rect 378100 177692 378106 177744
rect 268654 177624 268660 177676
rect 268712 177664 268718 177676
rect 578602 177664 578608 177676
rect 268712 177636 578608 177664
rect 268712 177624 268718 177636
rect 578602 177624 578608 177636
rect 578660 177624 578666 177676
rect 54570 177556 54576 177608
rect 54628 177596 54634 177608
rect 368842 177596 368848 177608
rect 54628 177568 368848 177596
rect 54628 177556 54634 177568
rect 368842 177556 368848 177568
rect 368900 177556 368906 177608
rect 89806 177488 89812 177540
rect 89864 177528 89870 177540
rect 99282 177528 99288 177540
rect 89864 177500 99288 177528
rect 89864 177488 89870 177500
rect 99282 177488 99288 177500
rect 99340 177488 99346 177540
rect 250622 177488 250628 177540
rect 250680 177528 250686 177540
rect 571886 177528 571892 177540
rect 250680 177500 571892 177528
rect 250680 177488 250686 177500
rect 571886 177488 571892 177500
rect 571944 177488 571950 177540
rect 49050 177420 49056 177472
rect 49108 177460 49114 177472
rect 391474 177460 391480 177472
rect 49108 177432 391480 177460
rect 49108 177420 49114 177432
rect 391474 177420 391480 177432
rect 391532 177420 391538 177472
rect 52638 177352 52644 177404
rect 52696 177392 52702 177404
rect 398374 177392 398380 177404
rect 52696 177364 398380 177392
rect 52696 177352 52702 177364
rect 398374 177352 398380 177364
rect 398432 177352 398438 177404
rect 48222 177284 48228 177336
rect 48280 177324 48286 177336
rect 399662 177324 399668 177336
rect 48280 177296 399668 177324
rect 48280 177284 48286 177296
rect 399662 177284 399668 177296
rect 399720 177284 399726 177336
rect 213270 176332 213276 176384
rect 213328 176372 213334 176384
rect 273346 176372 273352 176384
rect 213328 176344 273352 176372
rect 213328 176332 213334 176344
rect 273346 176332 273352 176344
rect 273404 176332 273410 176384
rect 313090 176332 313096 176384
rect 313148 176372 313154 176384
rect 380158 176372 380164 176384
rect 313148 176344 380164 176372
rect 313148 176332 313154 176344
rect 380158 176332 380164 176344
rect 380216 176332 380222 176384
rect 188154 176264 188160 176316
rect 188212 176304 188218 176316
rect 362310 176304 362316 176316
rect 188212 176276 362316 176304
rect 188212 176264 188218 176276
rect 362310 176264 362316 176276
rect 362368 176264 362374 176316
rect 113358 176196 113364 176248
rect 113416 176236 113422 176248
rect 379238 176236 379244 176248
rect 113416 176208 379244 176236
rect 113416 176196 113422 176208
rect 379238 176196 379244 176208
rect 379296 176196 379302 176248
rect 48130 176128 48136 176180
rect 48188 176168 48194 176180
rect 353846 176168 353852 176180
rect 48188 176140 353852 176168
rect 48188 176128 48194 176140
rect 353846 176128 353852 176140
rect 353904 176128 353910 176180
rect 44450 176060 44456 176112
rect 44508 176100 44514 176112
rect 360102 176100 360108 176112
rect 44508 176072 360108 176100
rect 44508 176060 44514 176072
rect 360102 176060 360108 176072
rect 360160 176060 360166 176112
rect 95234 175992 95240 176044
rect 95292 176032 95298 176044
rect 443178 176032 443184 176044
rect 95292 176004 443184 176032
rect 95292 175992 95298 176004
rect 443178 175992 443184 176004
rect 443236 175992 443242 176044
rect 49786 175924 49792 175976
rect 49844 175964 49850 175976
rect 526438 175964 526444 175976
rect 49844 175936 526444 175964
rect 49844 175924 49850 175936
rect 526438 175924 526444 175936
rect 526496 175924 526502 175976
rect 312446 175040 312452 175092
rect 312504 175080 312510 175092
rect 352098 175080 352104 175092
rect 312504 175052 352104 175080
rect 312504 175040 312510 175052
rect 352098 175040 352104 175052
rect 352156 175040 352162 175092
rect 53282 174972 53288 175024
rect 53340 175012 53346 175024
rect 349338 175012 349344 175024
rect 53340 174984 349344 175012
rect 53340 174972 53346 174984
rect 349338 174972 349344 174984
rect 349396 174972 349402 175024
rect 354306 174972 354312 175024
rect 354364 175012 354370 175024
rect 467834 175012 467840 175024
rect 354364 174984 467840 175012
rect 354364 174972 354370 174984
rect 467834 174972 467840 174984
rect 467892 174972 467898 175024
rect 59538 174904 59544 174956
rect 59596 174944 59602 174956
rect 380066 174944 380072 174956
rect 59596 174916 380072 174944
rect 59596 174904 59602 174916
rect 380066 174904 380072 174916
rect 380124 174904 380130 174956
rect 46750 174836 46756 174888
rect 46808 174876 46814 174888
rect 385862 174876 385868 174888
rect 46808 174848 385868 174876
rect 46808 174836 46814 174848
rect 385862 174836 385868 174848
rect 385920 174836 385926 174888
rect 55674 174768 55680 174820
rect 55732 174808 55738 174820
rect 401226 174808 401232 174820
rect 55732 174780 401232 174808
rect 55732 174768 55738 174780
rect 401226 174768 401232 174780
rect 401284 174768 401290 174820
rect 39758 174700 39764 174752
rect 39816 174740 39822 174752
rect 391382 174740 391388 174752
rect 39816 174712 391388 174740
rect 39816 174700 39822 174712
rect 391382 174700 391388 174712
rect 391440 174700 391446 174752
rect 40402 174632 40408 174684
rect 40460 174672 40466 174684
rect 483106 174672 483112 174684
rect 40460 174644 483112 174672
rect 40460 174632 40466 174644
rect 483106 174632 483112 174644
rect 483164 174632 483170 174684
rect 36722 174564 36728 174616
rect 36780 174604 36786 174616
rect 552658 174604 552664 174616
rect 36780 174576 552664 174604
rect 36780 174564 36786 174576
rect 552658 174564 552664 174576
rect 552716 174564 552722 174616
rect 50062 174496 50068 174548
rect 50120 174536 50126 174548
rect 574278 174536 574284 174548
rect 50120 174508 574284 174536
rect 50120 174496 50126 174508
rect 574278 174496 574284 174508
rect 574336 174496 574342 174548
rect 249334 173340 249340 173392
rect 249392 173380 249398 173392
rect 352466 173380 352472 173392
rect 249392 173352 352472 173380
rect 249392 173340 249398 173352
rect 352466 173340 352472 173352
rect 352524 173340 352530 173392
rect 268378 173272 268384 173324
rect 268436 173312 268442 173324
rect 506290 173312 506296 173324
rect 268436 173284 506296 173312
rect 268436 173272 268442 173284
rect 506290 173272 506296 173284
rect 506348 173272 506354 173324
rect 38654 173204 38660 173256
rect 38712 173244 38718 173256
rect 368014 173244 368020 173256
rect 38712 173216 368020 173244
rect 38712 173204 38718 173216
rect 368014 173204 368020 173216
rect 368072 173204 368078 173256
rect 88426 173136 88432 173188
rect 88484 173176 88490 173188
rect 480530 173176 480536 173188
rect 88484 173148 480536 173176
rect 88484 173136 88490 173148
rect 480530 173136 480536 173148
rect 480588 173136 480594 173188
rect 264146 172116 264152 172168
rect 264204 172156 264210 172168
rect 353570 172156 353576 172168
rect 264204 172128 353576 172156
rect 264204 172116 264210 172128
rect 353570 172116 353576 172128
rect 353628 172116 353634 172168
rect 112162 172048 112168 172100
rect 112220 172088 112226 172100
rect 129826 172088 129832 172100
rect 112220 172060 129832 172088
rect 112220 172048 112226 172060
rect 129826 172048 129832 172060
rect 129884 172048 129890 172100
rect 180794 172048 180800 172100
rect 180852 172088 180858 172100
rect 327074 172088 327080 172100
rect 180852 172060 327080 172088
rect 180852 172048 180858 172060
rect 327074 172048 327080 172060
rect 327132 172048 327138 172100
rect 96706 171980 96712 172032
rect 96764 172020 96770 172032
rect 242250 172020 242256 172032
rect 96764 171992 242256 172020
rect 96764 171980 96770 171992
rect 242250 171980 242256 171992
rect 242308 171980 242314 172032
rect 301038 171980 301044 172032
rect 301096 172020 301102 172032
rect 468294 172020 468300 172032
rect 301096 171992 468300 172020
rect 301096 171980 301102 171992
rect 468294 171980 468300 171992
rect 468352 171980 468358 172032
rect 115934 171912 115940 171964
rect 115992 171952 115998 171964
rect 343358 171952 343364 171964
rect 115992 171924 343364 171952
rect 115992 171912 115998 171924
rect 343358 171912 343364 171924
rect 343416 171912 343422 171964
rect 79318 171844 79324 171896
rect 79376 171884 79382 171896
rect 355502 171884 355508 171896
rect 79376 171856 355508 171884
rect 79376 171844 79382 171856
rect 355502 171844 355508 171856
rect 355560 171844 355566 171896
rect 50706 171776 50712 171828
rect 50764 171816 50770 171828
rect 375466 171816 375472 171828
rect 50764 171788 375472 171816
rect 50764 171776 50770 171788
rect 375466 171776 375472 171788
rect 375524 171776 375530 171828
rect 383378 171776 383384 171828
rect 383436 171816 383442 171828
rect 386414 171816 386420 171828
rect 383436 171788 386420 171816
rect 383436 171776 383442 171788
rect 386414 171776 386420 171788
rect 386472 171776 386478 171828
rect 35250 170552 35256 170604
rect 35308 170592 35314 170604
rect 193214 170592 193220 170604
rect 35308 170564 193220 170592
rect 35308 170552 35314 170564
rect 193214 170552 193220 170564
rect 193272 170552 193278 170604
rect 56410 170484 56416 170536
rect 56468 170524 56474 170536
rect 230474 170524 230480 170536
rect 56468 170496 230480 170524
rect 56468 170484 56474 170496
rect 230474 170484 230480 170496
rect 230532 170484 230538 170536
rect 233878 170484 233884 170536
rect 233936 170524 233942 170536
rect 389818 170524 389824 170536
rect 233936 170496 389824 170524
rect 233936 170484 233942 170496
rect 389818 170484 389824 170496
rect 389876 170484 389882 170536
rect 66438 170416 66444 170468
rect 66496 170456 66502 170468
rect 347958 170456 347964 170468
rect 66496 170428 347964 170456
rect 66496 170416 66502 170428
rect 347958 170416 347964 170428
rect 348016 170416 348022 170468
rect 57882 170348 57888 170400
rect 57940 170388 57946 170400
rect 387518 170388 387524 170400
rect 57940 170360 387524 170388
rect 57940 170348 57946 170360
rect 387518 170348 387524 170360
rect 387576 170348 387582 170400
rect 306466 169668 306472 169720
rect 306524 169708 306530 169720
rect 367738 169708 367744 169720
rect 306524 169680 367744 169708
rect 306524 169668 306530 169680
rect 367738 169668 367744 169680
rect 367796 169668 367802 169720
rect 225506 169600 225512 169652
rect 225564 169640 225570 169652
rect 365162 169640 365168 169652
rect 225564 169612 365168 169640
rect 225564 169600 225570 169612
rect 365162 169600 365168 169612
rect 365220 169600 365226 169652
rect 176654 169532 176660 169584
rect 176712 169572 176718 169584
rect 294046 169572 294052 169584
rect 176712 169544 294052 169572
rect 176712 169532 176718 169544
rect 294046 169532 294052 169544
rect 294104 169532 294110 169584
rect 315298 169532 315304 169584
rect 315356 169572 315362 169584
rect 484394 169572 484400 169584
rect 315356 169544 484400 169572
rect 315356 169532 315362 169544
rect 484394 169532 484400 169544
rect 484452 169532 484458 169584
rect 170766 169464 170772 169516
rect 170824 169504 170830 169516
rect 355410 169504 355416 169516
rect 170824 169476 355416 169504
rect 170824 169464 170830 169476
rect 355410 169464 355416 169476
rect 355468 169464 355474 169516
rect 124398 169396 124404 169448
rect 124456 169436 124462 169448
rect 363138 169436 363144 169448
rect 124456 169408 363144 169436
rect 124456 169396 124462 169408
rect 363138 169396 363144 169408
rect 363196 169396 363202 169448
rect 46566 169328 46572 169380
rect 46624 169368 46630 169380
rect 325694 169368 325700 169380
rect 46624 169340 325700 169368
rect 46624 169328 46630 169340
rect 325694 169328 325700 169340
rect 325752 169328 325758 169380
rect 328730 169328 328736 169380
rect 328788 169368 328794 169380
rect 394142 169368 394148 169380
rect 328788 169340 394148 169368
rect 328788 169328 328794 169340
rect 394142 169328 394148 169340
rect 394200 169328 394206 169380
rect 30098 169260 30104 169312
rect 30156 169300 30162 169312
rect 335630 169300 335636 169312
rect 30156 169272 335636 169300
rect 30156 169260 30162 169272
rect 335630 169260 335636 169272
rect 335688 169260 335694 169312
rect 78030 169192 78036 169244
rect 78088 169232 78094 169244
rect 388806 169232 388812 169244
rect 78088 169204 388812 169232
rect 78088 169192 78094 169204
rect 388806 169192 388812 169204
rect 388864 169192 388870 169244
rect 52822 169124 52828 169176
rect 52880 169164 52886 169176
rect 371050 169164 371056 169176
rect 52880 169136 371056 169164
rect 52880 169124 52886 169136
rect 371050 169124 371056 169136
rect 371108 169124 371114 169176
rect 64506 169056 64512 169108
rect 64564 169096 64570 169108
rect 563514 169096 563520 169108
rect 64564 169068 563520 169096
rect 64564 169056 64570 169068
rect 563514 169056 563520 169068
rect 563572 169056 563578 169108
rect 26786 168988 26792 169040
rect 26844 169028 26850 169040
rect 552566 169028 552572 169040
rect 26844 169000 552572 169028
rect 26844 168988 26850 169000
rect 552566 168988 552572 169000
rect 552624 168988 552630 169040
rect 207474 167696 207480 167748
rect 207532 167736 207538 167748
rect 402238 167736 402244 167748
rect 207532 167708 402244 167736
rect 207532 167696 207538 167708
rect 402238 167696 402244 167708
rect 402296 167696 402302 167748
rect 40862 167628 40868 167680
rect 40920 167668 40926 167680
rect 314378 167668 314384 167680
rect 40920 167640 314384 167668
rect 40920 167628 40926 167640
rect 314378 167628 314384 167640
rect 314436 167628 314442 167680
rect 405274 167628 405280 167680
rect 405332 167668 405338 167680
rect 565906 167668 565912 167680
rect 405332 167640 565912 167668
rect 405332 167628 405338 167640
rect 565906 167628 565912 167640
rect 565964 167628 565970 167680
rect 277394 166812 277400 166864
rect 277452 166852 277458 166864
rect 356974 166852 356980 166864
rect 277452 166824 356980 166852
rect 277452 166812 277458 166824
rect 356974 166812 356980 166824
rect 357032 166812 357038 166864
rect 258994 166744 259000 166796
rect 259052 166784 259058 166796
rect 350626 166784 350632 166796
rect 259052 166756 350632 166784
rect 259052 166744 259058 166756
rect 350626 166744 350632 166756
rect 350684 166744 350690 166796
rect 392854 166744 392860 166796
rect 392912 166784 392918 166796
rect 549530 166784 549536 166796
rect 392912 166756 549536 166784
rect 392912 166744 392918 166756
rect 549530 166744 549536 166756
rect 549588 166744 549594 166796
rect 199746 166676 199752 166728
rect 199804 166716 199810 166728
rect 372246 166716 372252 166728
rect 199804 166688 372252 166716
rect 199804 166676 199810 166688
rect 372246 166676 372252 166688
rect 372304 166676 372310 166728
rect 395062 166676 395068 166728
rect 395120 166716 395126 166728
rect 561214 166716 561220 166728
rect 395120 166688 561220 166716
rect 395120 166676 395126 166688
rect 561214 166676 561220 166688
rect 561272 166676 561278 166728
rect 324406 166608 324412 166660
rect 324464 166648 324470 166660
rect 563514 166648 563520 166660
rect 324464 166620 563520 166648
rect 324464 166608 324470 166620
rect 563514 166608 563520 166620
rect 563572 166608 563578 166660
rect 84194 166540 84200 166592
rect 84252 166580 84258 166592
rect 367462 166580 367468 166592
rect 84252 166552 367468 166580
rect 84252 166540 84258 166552
rect 367462 166540 367468 166552
rect 367520 166540 367526 166592
rect 391198 166540 391204 166592
rect 391256 166580 391262 166592
rect 560478 166580 560484 166592
rect 391256 166552 560484 166580
rect 391256 166540 391262 166552
rect 560478 166540 560484 166552
rect 560536 166540 560542 166592
rect 41138 166472 41144 166524
rect 41196 166512 41202 166524
rect 377582 166512 377588 166524
rect 41196 166484 377588 166512
rect 41196 166472 41202 166484
rect 377582 166472 377588 166484
rect 377640 166472 377646 166524
rect 391842 166472 391848 166524
rect 391900 166512 391906 166524
rect 566274 166512 566280 166524
rect 391900 166484 566280 166512
rect 391900 166472 391906 166484
rect 566274 166472 566280 166484
rect 566332 166472 566338 166524
rect 150526 166404 150532 166456
rect 150584 166444 150590 166456
rect 539226 166444 539232 166456
rect 150584 166416 539232 166444
rect 150584 166404 150590 166416
rect 539226 166404 539232 166416
rect 539284 166404 539290 166456
rect 54846 166336 54852 166388
rect 54904 166376 54910 166388
rect 470594 166376 470600 166388
rect 54904 166348 470600 166376
rect 54904 166336 54910 166348
rect 470594 166336 470600 166348
rect 470652 166336 470658 166388
rect 508498 166336 508504 166388
rect 508556 166376 508562 166388
rect 514018 166376 514024 166388
rect 508556 166348 514024 166376
rect 508556 166336 508562 166348
rect 514018 166336 514024 166348
rect 514076 166336 514082 166388
rect 150434 166268 150440 166320
rect 150492 166308 150498 166320
rect 567746 166308 567752 166320
rect 150492 166280 567752 166308
rect 150492 166268 150498 166280
rect 567746 166268 567752 166280
rect 567804 166268 567810 166320
rect 228726 165112 228732 165164
rect 228784 165152 228790 165164
rect 374638 165152 374644 165164
rect 228784 165124 374644 165152
rect 228784 165112 228790 165124
rect 374638 165112 374644 165124
rect 374696 165112 374702 165164
rect 81894 165044 81900 165096
rect 81952 165084 81958 165096
rect 231946 165084 231952 165096
rect 81952 165056 231952 165084
rect 81952 165044 81958 165056
rect 231946 165044 231952 165056
rect 232004 165044 232010 165096
rect 237374 165044 237380 165096
rect 237432 165084 237438 165096
rect 506934 165084 506940 165096
rect 237432 165056 506940 165084
rect 237432 165044 237438 165056
rect 506934 165044 506940 165056
rect 506992 165044 506998 165096
rect 43346 164976 43352 165028
rect 43404 165016 43410 165028
rect 350442 165016 350448 165028
rect 43404 164988 350448 165016
rect 43404 164976 43410 164988
rect 350442 164976 350448 164988
rect 350500 164976 350506 165028
rect 29546 164908 29552 164960
rect 29604 164948 29610 164960
rect 376846 164948 376852 164960
rect 29604 164920 376852 164948
rect 29604 164908 29610 164920
rect 376846 164908 376852 164920
rect 376904 164908 376910 164960
rect 197170 164840 197176 164892
rect 197228 164880 197234 164892
rect 560386 164880 560392 164892
rect 197228 164852 560392 164880
rect 197228 164840 197234 164852
rect 560386 164840 560392 164852
rect 560444 164840 560450 164892
rect 307018 164160 307024 164212
rect 307076 164200 307082 164212
rect 309870 164200 309876 164212
rect 307076 164172 309876 164200
rect 307076 164160 307082 164172
rect 309870 164160 309876 164172
rect 309928 164160 309934 164212
rect 397270 164160 397276 164212
rect 397328 164200 397334 164212
rect 548334 164200 548340 164212
rect 397328 164172 548340 164200
rect 397328 164160 397334 164172
rect 548334 164160 548340 164172
rect 548392 164160 548398 164212
rect 408126 164092 408132 164144
rect 408184 164132 408190 164144
rect 560570 164132 560576 164144
rect 408184 164104 560576 164132
rect 408184 164092 408190 164104
rect 560570 164092 560576 164104
rect 560628 164092 560634 164144
rect 237742 164024 237748 164076
rect 237800 164064 237806 164076
rect 384390 164064 384396 164076
rect 237800 164036 384396 164064
rect 237800 164024 237806 164036
rect 384390 164024 384396 164036
rect 384448 164024 384454 164076
rect 404722 164024 404728 164076
rect 404780 164064 404786 164076
rect 570598 164064 570604 164076
rect 404780 164036 570604 164064
rect 404780 164024 404786 164036
rect 570598 164024 570604 164036
rect 570656 164024 570662 164076
rect 226150 163956 226156 164008
rect 226208 163996 226214 164008
rect 324314 163996 324320 164008
rect 226208 163968 324320 163996
rect 226208 163956 226214 163968
rect 324314 163956 324320 163968
rect 324372 163956 324378 164008
rect 346394 163956 346400 164008
rect 346452 163996 346458 164008
rect 560938 163996 560944 164008
rect 346452 163968 560944 163996
rect 346452 163956 346458 163968
rect 560938 163956 560944 163968
rect 560996 163956 561002 164008
rect 137278 163888 137284 163940
rect 137336 163928 137342 163940
rect 360470 163928 360476 163940
rect 137336 163900 360476 163928
rect 137336 163888 137342 163900
rect 360470 163888 360476 163900
rect 360528 163888 360534 163940
rect 384482 163888 384488 163940
rect 384540 163928 384546 163940
rect 552106 163928 552112 163940
rect 384540 163900 552112 163928
rect 384540 163888 384546 163900
rect 552106 163888 552112 163900
rect 552164 163888 552170 163940
rect 110874 163820 110880 163872
rect 110932 163860 110938 163872
rect 278774 163860 278780 163872
rect 110932 163832 278780 163860
rect 110932 163820 110938 163832
rect 278774 163820 278780 163832
rect 278832 163820 278838 163872
rect 305086 163820 305092 163872
rect 305144 163860 305150 163872
rect 550910 163860 550916 163872
rect 305144 163832 550916 163860
rect 305144 163820 305150 163832
rect 550910 163820 550916 163832
rect 550968 163820 550974 163872
rect 43622 163752 43628 163804
rect 43680 163792 43686 163804
rect 260834 163792 260840 163804
rect 43680 163764 260840 163792
rect 43680 163752 43686 163764
rect 260834 163752 260840 163764
rect 260892 163752 260898 163804
rect 302234 163752 302240 163804
rect 302292 163792 302298 163804
rect 551094 163792 551100 163804
rect 302292 163764 551100 163792
rect 302292 163752 302298 163764
rect 551094 163752 551100 163764
rect 551152 163752 551158 163804
rect 35158 163684 35164 163736
rect 35216 163724 35222 163736
rect 214098 163724 214104 163736
rect 35216 163696 214104 163724
rect 35216 163684 35222 163696
rect 214098 163684 214104 163696
rect 214156 163684 214162 163736
rect 222194 163684 222200 163736
rect 222252 163724 222258 163736
rect 546862 163724 546868 163736
rect 222252 163696 546868 163724
rect 222252 163684 222258 163696
rect 546862 163684 546868 163696
rect 546920 163684 546926 163736
rect 212534 163616 212540 163668
rect 212592 163656 212598 163668
rect 541250 163656 541256 163668
rect 212592 163628 541256 163656
rect 212592 163616 212598 163628
rect 541250 163616 541256 163628
rect 541308 163616 541314 163668
rect 184934 163548 184940 163600
rect 184992 163588 184998 163600
rect 540698 163588 540704 163600
rect 184992 163560 540704 163588
rect 184992 163548 184998 163560
rect 540698 163548 540704 163560
rect 540756 163548 540762 163600
rect 29638 163480 29644 163532
rect 29696 163520 29702 163532
rect 460566 163520 460572 163532
rect 29696 163492 460572 163520
rect 29696 163480 29702 163492
rect 460566 163480 460572 163492
rect 460624 163480 460630 163532
rect 395614 163412 395620 163464
rect 395672 163452 395678 163464
rect 510154 163452 510160 163464
rect 395672 163424 510160 163452
rect 395672 163412 395678 163424
rect 510154 163412 510160 163424
rect 510212 163412 510218 163464
rect 414658 162800 414664 162852
rect 414716 162840 414722 162852
rect 419994 162840 420000 162852
rect 414716 162812 420000 162840
rect 414716 162800 414722 162812
rect 419994 162800 420000 162812
rect 420052 162800 420058 162852
rect 351086 162324 351092 162376
rect 351144 162364 351150 162376
rect 377858 162364 377864 162376
rect 351144 162336 377864 162364
rect 351144 162324 351150 162336
rect 377858 162324 377864 162336
rect 377916 162324 377922 162376
rect 266354 162256 266360 162308
rect 266412 162296 266418 162308
rect 356054 162296 356060 162308
rect 266412 162268 356060 162296
rect 266412 162256 266418 162268
rect 356054 162256 356060 162268
rect 356112 162256 356118 162308
rect 382182 162256 382188 162308
rect 382240 162296 382246 162308
rect 400674 162296 400680 162308
rect 382240 162268 400680 162296
rect 382240 162256 382246 162268
rect 400674 162256 400680 162268
rect 400732 162256 400738 162308
rect 285674 162188 285680 162240
rect 285732 162228 285738 162240
rect 403894 162228 403900 162240
rect 285732 162200 403900 162228
rect 285732 162188 285738 162200
rect 403894 162188 403900 162200
rect 403952 162188 403958 162240
rect 127066 162120 127072 162172
rect 127124 162160 127130 162172
rect 383286 162160 383292 162172
rect 127124 162132 383292 162160
rect 127124 162120 127130 162132
rect 383286 162120 383292 162132
rect 383344 162120 383350 162172
rect 406654 162120 406660 162172
rect 406712 162160 406718 162172
rect 551462 162160 551468 162172
rect 406712 162132 551468 162160
rect 406712 162120 406718 162132
rect 551462 162120 551468 162132
rect 551520 162120 551526 162172
rect 389726 161372 389732 161424
rect 389784 161412 389790 161424
rect 549622 161412 549628 161424
rect 389784 161384 549628 161412
rect 389784 161372 389790 161384
rect 549622 161372 549628 161384
rect 549680 161372 549686 161424
rect 378870 161304 378876 161356
rect 378928 161344 378934 161356
rect 545390 161344 545396 161356
rect 378928 161316 545396 161344
rect 378928 161304 378934 161316
rect 545390 161304 545396 161316
rect 545448 161304 545454 161356
rect 371970 161236 371976 161288
rect 372028 161276 372034 161288
rect 552474 161276 552480 161288
rect 372028 161248 552480 161276
rect 372028 161236 372034 161248
rect 552474 161236 552480 161248
rect 552532 161236 552538 161288
rect 248414 161168 248420 161220
rect 248472 161208 248478 161220
rect 376478 161208 376484 161220
rect 248472 161180 376484 161208
rect 248472 161168 248478 161180
rect 376478 161168 376484 161180
rect 376536 161168 376542 161220
rect 396718 161168 396724 161220
rect 396776 161208 396782 161220
rect 580258 161208 580264 161220
rect 396776 161180 580264 161208
rect 396776 161168 396782 161180
rect 580258 161168 580264 161180
rect 580316 161168 580322 161220
rect 221642 161100 221648 161152
rect 221700 161140 221706 161152
rect 356238 161140 356244 161152
rect 221700 161112 356244 161140
rect 221700 161100 221706 161112
rect 356238 161100 356244 161112
rect 356296 161100 356302 161152
rect 391658 161100 391664 161152
rect 391716 161140 391722 161152
rect 578602 161140 578608 161152
rect 391716 161112 578608 161140
rect 391716 161100 391722 161112
rect 578602 161100 578608 161112
rect 578660 161100 578666 161152
rect 142430 161032 142436 161084
rect 142488 161072 142494 161084
rect 361114 161072 361120 161084
rect 142488 161044 361120 161072
rect 142488 161032 142494 161044
rect 361114 161032 361120 161044
rect 361172 161032 361178 161084
rect 365346 161032 365352 161084
rect 365404 161072 365410 161084
rect 560662 161072 560668 161084
rect 365404 161044 560668 161072
rect 365404 161032 365410 161044
rect 560662 161032 560668 161044
rect 560720 161032 560726 161084
rect 320174 160964 320180 161016
rect 320232 161004 320238 161016
rect 578234 161004 578240 161016
rect 320232 160976 578240 161004
rect 320232 160964 320238 160976
rect 578234 160964 578240 160976
rect 578292 160964 578298 161016
rect 56778 160896 56784 160948
rect 56836 160936 56842 160948
rect 358538 160936 358544 160948
rect 56836 160908 358544 160936
rect 56836 160896 56842 160908
rect 358538 160896 358544 160908
rect 358596 160896 358602 160948
rect 375098 160896 375104 160948
rect 375156 160936 375162 160948
rect 578786 160936 578792 160948
rect 375156 160908 578792 160936
rect 375156 160896 375162 160908
rect 578786 160896 578792 160908
rect 578844 160896 578850 160948
rect 39390 160828 39396 160880
rect 39448 160868 39454 160880
rect 240134 160868 240140 160880
rect 39448 160840 240140 160868
rect 39448 160828 39454 160840
rect 240134 160828 240140 160840
rect 240192 160828 240198 160880
rect 253934 160828 253940 160880
rect 253992 160868 253998 160880
rect 581822 160868 581828 160880
rect 253992 160840 581828 160868
rect 253992 160828 253998 160840
rect 581822 160828 581828 160840
rect 581880 160828 581886 160880
rect 219710 160760 219716 160812
rect 219768 160800 219774 160812
rect 566182 160800 566188 160812
rect 219768 160772 566188 160800
rect 219768 160760 219774 160772
rect 566182 160760 566188 160772
rect 566240 160760 566246 160812
rect 178126 160692 178132 160744
rect 178184 160732 178190 160744
rect 553302 160732 553308 160744
rect 178184 160704 553308 160732
rect 178184 160692 178190 160704
rect 553302 160692 553308 160704
rect 553360 160692 553366 160744
rect 282822 160624 282828 160676
rect 282880 160664 282886 160676
rect 426434 160664 426440 160676
rect 282880 160636 426440 160664
rect 282880 160624 282886 160636
rect 426434 160624 426440 160636
rect 426492 160624 426498 160676
rect 405090 160556 405096 160608
rect 405148 160596 405154 160608
rect 548518 160596 548524 160608
rect 405148 160568 548524 160596
rect 405148 160556 405154 160568
rect 548518 160556 548524 160568
rect 548576 160556 548582 160608
rect 155310 159740 155316 159792
rect 155368 159780 155374 159792
rect 388438 159780 388444 159792
rect 155368 159752 388444 159780
rect 155368 159740 155374 159752
rect 388438 159740 388444 159752
rect 388496 159740 388502 159792
rect 96706 159672 96712 159724
rect 96764 159712 96770 159724
rect 366358 159712 366364 159724
rect 96764 159684 366364 159712
rect 96764 159672 96770 159684
rect 366358 159672 366364 159684
rect 366416 159672 366422 159724
rect 402790 159672 402796 159724
rect 402848 159712 402854 159724
rect 549070 159712 549076 159724
rect 402848 159684 549076 159712
rect 402848 159672 402854 159684
rect 549070 159672 549076 159684
rect 549128 159672 549134 159724
rect 252554 159604 252560 159656
rect 252612 159644 252618 159656
rect 546218 159644 546224 159656
rect 252612 159616 546224 159644
rect 252612 159604 252618 159616
rect 546218 159604 546224 159616
rect 546276 159604 546282 159656
rect 168374 159536 168380 159588
rect 168432 159576 168438 159588
rect 480254 159576 480260 159588
rect 168432 159548 480260 159576
rect 168432 159536 168438 159548
rect 480254 159536 480260 159548
rect 480312 159536 480318 159588
rect 121454 159468 121460 159520
rect 121512 159508 121518 159520
rect 454126 159508 454132 159520
rect 121512 159480 454132 159508
rect 121512 159468 121518 159480
rect 454126 159468 454132 159480
rect 454184 159468 454190 159520
rect 216766 159400 216772 159452
rect 216824 159440 216830 159452
rect 553026 159440 553032 159452
rect 216824 159412 553032 159440
rect 216824 159400 216830 159412
rect 553026 159400 553032 159412
rect 553084 159400 553090 159452
rect 3418 159332 3424 159384
rect 3476 159372 3482 159384
rect 359642 159372 359648 159384
rect 3476 159344 359648 159372
rect 3476 159332 3482 159344
rect 359642 159332 359648 159344
rect 359700 159332 359706 159384
rect 379146 159332 379152 159384
rect 379204 159372 379210 159384
rect 539962 159372 539968 159384
rect 379204 159344 539968 159372
rect 379204 159332 379210 159344
rect 539962 159332 539968 159344
rect 540020 159332 540026 159384
rect 292574 158652 292580 158704
rect 292632 158692 292638 158704
rect 439314 158692 439320 158704
rect 292632 158664 439320 158692
rect 292632 158652 292638 158664
rect 439314 158652 439320 158664
rect 439372 158652 439378 158704
rect 268010 158584 268016 158636
rect 268068 158624 268074 158636
rect 349890 158624 349896 158636
rect 268068 158596 349896 158624
rect 268068 158584 268074 158596
rect 349890 158584 349896 158596
rect 349948 158584 349954 158636
rect 383102 158584 383108 158636
rect 383160 158624 383166 158636
rect 540514 158624 540520 158636
rect 383160 158596 540520 158624
rect 383160 158584 383166 158596
rect 540514 158584 540520 158596
rect 540572 158584 540578 158636
rect 150158 158516 150164 158568
rect 150216 158556 150222 158568
rect 359090 158556 359096 158568
rect 150216 158528 359096 158556
rect 150216 158516 150222 158528
rect 359090 158516 359096 158528
rect 359148 158516 359154 158568
rect 368106 158516 368112 158568
rect 368164 158556 368170 158568
rect 539318 158556 539324 158568
rect 368164 158528 539324 158556
rect 368164 158516 368170 158528
rect 539318 158516 539324 158528
rect 539376 158516 539382 158568
rect 92566 158448 92572 158500
rect 92624 158488 92630 158500
rect 320818 158488 320824 158500
rect 92624 158460 320824 158488
rect 92624 158448 92630 158460
rect 320818 158448 320824 158460
rect 320876 158448 320882 158500
rect 386046 158448 386052 158500
rect 386104 158488 386110 158500
rect 559466 158488 559472 158500
rect 386104 158460 559472 158488
rect 386104 158448 386110 158460
rect 559466 158448 559472 158460
rect 559524 158448 559530 158500
rect 282914 158380 282920 158432
rect 282972 158420 282978 158432
rect 540606 158420 540612 158432
rect 282972 158392 540612 158420
rect 282972 158380 282978 158392
rect 540606 158380 540612 158392
rect 540664 158380 540670 158432
rect 304994 158312 305000 158364
rect 305052 158352 305058 158364
rect 571794 158352 571800 158364
rect 305052 158324 571800 158352
rect 305052 158312 305058 158324
rect 571794 158312 571800 158324
rect 571852 158312 571858 158364
rect 259546 158244 259552 158296
rect 259604 158284 259610 158296
rect 552014 158284 552020 158296
rect 259604 158256 552020 158284
rect 259604 158244 259610 158256
rect 552014 158244 552020 158256
rect 552072 158244 552078 158296
rect 231854 158176 231860 158228
rect 231912 158216 231918 158228
rect 539410 158216 539416 158228
rect 231912 158188 539416 158216
rect 231912 158176 231918 158188
rect 539410 158176 539416 158188
rect 539468 158176 539474 158228
rect 155954 158108 155960 158160
rect 156012 158148 156018 158160
rect 481818 158148 481824 158160
rect 156012 158120 481824 158148
rect 156012 158108 156018 158120
rect 481818 158108 481824 158120
rect 481876 158108 481882 158160
rect 158714 158040 158720 158092
rect 158772 158080 158778 158092
rect 551002 158080 551008 158092
rect 158772 158052 551008 158080
rect 158772 158040 158778 158052
rect 551002 158040 551008 158052
rect 551060 158040 551066 158092
rect 28166 157972 28172 158024
rect 28224 158012 28230 158024
rect 559374 158012 559380 158024
rect 28224 157984 559380 158012
rect 28224 157972 28230 157984
rect 559374 157972 559380 157984
rect 559432 157972 559438 158024
rect 394602 157904 394608 157956
rect 394660 157944 394666 157956
rect 537478 157944 537484 157956
rect 394660 157916 537484 157944
rect 394660 157904 394666 157916
rect 537478 157904 537484 157916
rect 537536 157904 537542 157956
rect 264238 157836 264244 157888
rect 264296 157876 264302 157888
rect 406470 157876 406476 157888
rect 264296 157848 406476 157876
rect 264296 157836 264302 157848
rect 406470 157836 406476 157848
rect 406528 157836 406534 157888
rect 398650 157768 398656 157820
rect 398708 157808 398714 157820
rect 537570 157808 537576 157820
rect 398708 157780 537576 157808
rect 398708 157768 398714 157780
rect 537570 157768 537576 157780
rect 537628 157768 537634 157820
rect 400950 157020 400956 157072
rect 401008 157060 401014 157072
rect 551554 157060 551560 157072
rect 401008 157032 551560 157060
rect 401008 157020 401014 157032
rect 551554 157020 551560 157032
rect 551612 157020 551618 157072
rect 166258 156952 166264 157004
rect 166316 156992 166322 157004
rect 188798 156992 188804 157004
rect 166316 156964 188804 156992
rect 166316 156952 166322 156964
rect 188798 156952 188804 156964
rect 188856 156952 188862 157004
rect 259638 156952 259644 157004
rect 259696 156992 259702 157004
rect 309134 156992 309140 157004
rect 259696 156964 309140 156992
rect 259696 156952 259702 156964
rect 309134 156952 309140 156964
rect 309192 156952 309198 157004
rect 398742 156952 398748 157004
rect 398800 156992 398806 157004
rect 556614 156992 556620 157004
rect 398800 156964 556620 156992
rect 398800 156952 398806 156964
rect 556614 156952 556620 156964
rect 556672 156952 556678 157004
rect 47578 156884 47584 156936
rect 47636 156924 47642 156936
rect 204254 156924 204260 156936
rect 47636 156896 204260 156924
rect 47636 156884 47642 156896
rect 204254 156884 204260 156896
rect 204312 156884 204318 156936
rect 271874 156884 271880 156936
rect 271932 156924 271938 156936
rect 368198 156924 368204 156936
rect 271932 156896 368204 156924
rect 271932 156884 271938 156896
rect 368198 156884 368204 156896
rect 368256 156884 368262 156936
rect 381446 156884 381452 156936
rect 381504 156924 381510 156936
rect 571886 156924 571892 156936
rect 381504 156896 571892 156924
rect 381504 156884 381510 156896
rect 571886 156884 571892 156896
rect 571944 156884 571950 156936
rect 45922 156816 45928 156868
rect 45980 156856 45986 156868
rect 361942 156856 361948 156868
rect 45980 156828 361948 156856
rect 45980 156816 45986 156828
rect 361942 156816 361948 156828
rect 362000 156816 362006 156868
rect 375006 156816 375012 156868
rect 375064 156856 375070 156868
rect 574278 156856 574284 156868
rect 375064 156828 574284 156856
rect 375064 156816 375070 156828
rect 574278 156816 574284 156828
rect 574336 156816 574342 156868
rect 80238 156748 80244 156800
rect 80296 156788 80302 156800
rect 281534 156788 281540 156800
rect 80296 156760 281540 156788
rect 80296 156748 80302 156760
rect 281534 156748 281540 156760
rect 281592 156748 281598 156800
rect 318242 156748 318248 156800
rect 318300 156788 318306 156800
rect 328454 156788 328460 156800
rect 318300 156760 328460 156788
rect 318300 156748 318306 156760
rect 328454 156748 328460 156760
rect 328512 156748 328518 156800
rect 333974 156748 333980 156800
rect 334032 156788 334038 156800
rect 541158 156788 541164 156800
rect 334032 156760 541164 156788
rect 334032 156748 334038 156760
rect 541158 156748 541164 156760
rect 541216 156748 541222 156800
rect 78766 156680 78772 156732
rect 78824 156720 78830 156732
rect 323394 156720 323400 156732
rect 78824 156692 323400 156720
rect 78824 156680 78830 156692
rect 323394 156680 323400 156692
rect 323452 156680 323458 156732
rect 328546 156680 328552 156732
rect 328604 156720 328610 156732
rect 558086 156720 558092 156732
rect 328604 156692 558092 156720
rect 328604 156680 328610 156692
rect 558086 156680 558092 156692
rect 558144 156680 558150 156732
rect 59354 156612 59360 156664
rect 59412 156652 59418 156664
rect 59630 156652 59636 156664
rect 59412 156624 59636 156652
rect 59412 156612 59418 156624
rect 59630 156612 59636 156624
rect 59688 156612 59694 156664
rect 124306 156612 124312 156664
rect 124364 156652 124370 156664
rect 574462 156652 574468 156664
rect 124364 156624 574468 156652
rect 124364 156612 124370 156624
rect 574462 156612 574468 156624
rect 574520 156612 574526 156664
rect 376754 156544 376760 156596
rect 376812 156584 376818 156596
rect 377214 156584 377220 156596
rect 376812 156556 377220 156584
rect 376812 156544 376818 156556
rect 377214 156544 377220 156556
rect 377272 156544 377278 156596
rect 254578 155864 254584 155916
rect 254636 155904 254642 155916
rect 369118 155904 369124 155916
rect 254636 155876 369124 155904
rect 254636 155864 254642 155876
rect 369118 155864 369124 155876
rect 369176 155864 369182 155916
rect 383470 155864 383476 155916
rect 383528 155904 383534 155916
rect 537110 155904 537116 155916
rect 383528 155876 537116 155904
rect 383528 155864 383534 155876
rect 537110 155864 537116 155876
rect 537168 155864 537174 155916
rect 538950 155864 538956 155916
rect 539008 155904 539014 155916
rect 539502 155904 539508 155916
rect 539008 155876 539508 155904
rect 539008 155864 539014 155876
rect 539502 155864 539508 155876
rect 539560 155864 539566 155916
rect 109678 155796 109684 155848
rect 109736 155836 109742 155848
rect 161750 155836 161756 155848
rect 109736 155808 161756 155836
rect 109736 155796 109742 155808
rect 161750 155796 161756 155808
rect 161808 155796 161814 155848
rect 232590 155796 232596 155848
rect 232648 155836 232654 155848
rect 348418 155836 348424 155848
rect 232648 155808 348424 155836
rect 232648 155796 232654 155808
rect 348418 155796 348424 155808
rect 348476 155796 348482 155848
rect 409782 155796 409788 155848
rect 409840 155836 409846 155848
rect 565078 155836 565084 155848
rect 409840 155808 565084 155836
rect 409840 155796 409846 155808
rect 565078 155796 565084 155808
rect 565136 155796 565142 155848
rect 47946 155728 47952 155780
rect 48004 155768 48010 155780
rect 136634 155768 136640 155780
rect 48004 155740 136640 155768
rect 48004 155728 48010 155740
rect 136634 155728 136640 155740
rect 136692 155728 136698 155780
rect 179414 155728 179420 155780
rect 179472 155768 179478 155780
rect 229370 155768 229376 155780
rect 179472 155740 229376 155768
rect 179472 155728 179478 155740
rect 229370 155728 229376 155740
rect 229428 155728 229434 155780
rect 230014 155728 230020 155780
rect 230072 155768 230078 155780
rect 355318 155768 355324 155780
rect 230072 155740 355324 155768
rect 230072 155728 230078 155740
rect 355318 155728 355324 155740
rect 355376 155728 355382 155780
rect 401410 155728 401416 155780
rect 401468 155768 401474 155780
rect 557810 155768 557816 155780
rect 401468 155740 557816 155768
rect 401468 155728 401474 155740
rect 557810 155728 557816 155740
rect 557868 155728 557874 155780
rect 56042 155660 56048 155712
rect 56100 155700 56106 155712
rect 154574 155700 154580 155712
rect 56100 155672 154580 155700
rect 56100 155660 56106 155672
rect 154574 155660 154580 155672
rect 154632 155660 154638 155712
rect 205634 155660 205640 155712
rect 205692 155700 205698 155712
rect 360930 155700 360936 155712
rect 205692 155672 360936 155700
rect 205692 155660 205698 155672
rect 360930 155660 360936 155672
rect 360988 155660 360994 155712
rect 409598 155660 409604 155712
rect 409656 155700 409662 155712
rect 567378 155700 567384 155712
rect 409656 155672 567384 155700
rect 409656 155660 409662 155672
rect 567378 155660 567384 155672
rect 567436 155660 567442 155712
rect 40954 155592 40960 155644
rect 41012 155632 41018 155644
rect 238754 155632 238760 155644
rect 41012 155604 238760 155632
rect 41012 155592 41018 155604
rect 238754 155592 238760 155604
rect 238812 155592 238818 155644
rect 292482 155592 292488 155644
rect 292540 155632 292546 155644
rect 349982 155632 349988 155644
rect 292540 155604 349988 155632
rect 292540 155592 292546 155604
rect 349982 155592 349988 155604
rect 350040 155592 350046 155644
rect 353938 155592 353944 155644
rect 353996 155632 354002 155644
rect 554130 155632 554136 155644
rect 353996 155604 554136 155632
rect 353996 155592 354002 155604
rect 554130 155592 554136 155604
rect 554188 155592 554194 155644
rect 57606 155524 57612 155576
rect 57664 155564 57670 155576
rect 361666 155564 361672 155576
rect 57664 155536 361672 155564
rect 57664 155524 57670 155536
rect 361666 155524 361672 155536
rect 361724 155524 361730 155576
rect 394418 155524 394424 155576
rect 394476 155564 394482 155576
rect 555050 155564 555056 155576
rect 394476 155536 555056 155564
rect 394476 155524 394482 155536
rect 555050 155524 555056 155536
rect 555108 155524 555114 155576
rect 32214 155456 32220 155508
rect 32272 155496 32278 155508
rect 284110 155496 284116 155508
rect 32272 155468 284116 155496
rect 32272 155456 32278 155468
rect 284110 155456 284116 155468
rect 284168 155456 284174 155508
rect 338114 155456 338120 155508
rect 338172 155496 338178 155508
rect 562226 155496 562232 155508
rect 338172 155468 562232 155496
rect 338172 155456 338178 155468
rect 562226 155456 562232 155468
rect 562284 155456 562290 155508
rect 57698 155388 57704 155440
rect 57756 155428 57762 155440
rect 372338 155428 372344 155440
rect 57756 155400 372344 155428
rect 57756 155388 57762 155400
rect 372338 155388 372344 155400
rect 372396 155388 372402 155440
rect 390462 155388 390468 155440
rect 390520 155428 390526 155440
rect 565354 155428 565360 155440
rect 390520 155400 565360 155428
rect 390520 155388 390526 155400
rect 565354 155388 565360 155400
rect 565412 155388 565418 155440
rect 43622 155320 43628 155372
rect 43680 155360 43686 155372
rect 368566 155360 368572 155372
rect 43680 155332 368572 155360
rect 43680 155320 43686 155332
rect 368566 155320 368572 155332
rect 368624 155320 368630 155372
rect 370498 155320 370504 155372
rect 370556 155360 370562 155372
rect 576118 155360 576124 155372
rect 370556 155332 576124 155360
rect 370556 155320 370562 155332
rect 576118 155320 576124 155332
rect 576176 155320 576182 155372
rect 46382 155252 46388 155304
rect 46440 155292 46446 155304
rect 162854 155292 162860 155304
rect 46440 155264 162860 155292
rect 46440 155252 46446 155264
rect 162854 155252 162860 155264
rect 162912 155252 162918 155304
rect 216674 155252 216680 155304
rect 216732 155292 216738 155304
rect 547782 155292 547788 155304
rect 216732 155264 547788 155292
rect 216732 155252 216738 155264
rect 547782 155252 547788 155264
rect 547840 155252 547846 155304
rect 32582 155184 32588 155236
rect 32640 155224 32646 155236
rect 396166 155224 396172 155236
rect 32640 155196 396172 155224
rect 32640 155184 32646 155196
rect 396166 155184 396172 155196
rect 396224 155184 396230 155236
rect 408310 155184 408316 155236
rect 408368 155224 408374 155236
rect 570506 155224 570512 155236
rect 408368 155196 570512 155224
rect 408368 155184 408374 155196
rect 570506 155184 570512 155196
rect 570564 155184 570570 155236
rect 295702 155116 295708 155168
rect 295760 155156 295766 155168
rect 350534 155156 350540 155168
rect 295760 155128 350540 155156
rect 295760 155116 295766 155128
rect 350534 155116 350540 155128
rect 350592 155116 350598 155168
rect 405366 155116 405372 155168
rect 405424 155156 405430 155168
rect 556430 155156 556436 155168
rect 405424 155128 556436 155156
rect 405424 155116 405430 155128
rect 556430 155116 556436 155128
rect 556488 155116 556494 155168
rect 269114 155048 269120 155100
rect 269172 155088 269178 155100
rect 322750 155088 322756 155100
rect 269172 155060 322756 155088
rect 269172 155048 269178 155060
rect 322750 155048 322756 155060
rect 322808 155048 322814 155100
rect 403986 155048 403992 155100
rect 404044 155088 404050 155100
rect 553946 155088 553952 155100
rect 404044 155060 553952 155088
rect 404044 155048 404050 155060
rect 553946 155048 553952 155060
rect 554004 155048 554010 155100
rect 309226 154980 309232 155032
rect 309284 155020 309290 155032
rect 357158 155020 357164 155032
rect 309284 154992 357164 155020
rect 309284 154980 309290 154992
rect 357158 154980 357164 154992
rect 357216 154980 357222 155032
rect 410150 154980 410156 155032
rect 410208 155020 410214 155032
rect 538950 155020 538956 155032
rect 410208 154992 538956 155020
rect 410208 154980 410214 154992
rect 538950 154980 538956 154992
rect 539008 154980 539014 155032
rect 405182 154504 405188 154556
rect 405240 154544 405246 154556
rect 542722 154544 542728 154556
rect 405240 154516 542728 154544
rect 405240 154504 405246 154516
rect 542722 154504 542728 154516
rect 542780 154504 542786 154556
rect 396994 154436 397000 154488
rect 397052 154476 397058 154488
rect 542630 154476 542636 154488
rect 397052 154448 542636 154476
rect 397052 154436 397058 154448
rect 542630 154436 542636 154448
rect 542688 154436 542694 154488
rect 382090 154368 382096 154420
rect 382148 154408 382154 154420
rect 539594 154408 539600 154420
rect 382148 154380 539600 154408
rect 382148 154368 382154 154380
rect 539594 154368 539600 154380
rect 539652 154368 539658 154420
rect 409690 154300 409696 154352
rect 409748 154340 409754 154352
rect 569310 154340 569316 154352
rect 409748 154312 569316 154340
rect 409748 154300 409754 154312
rect 569310 154300 569316 154312
rect 569368 154300 569374 154352
rect 260282 154232 260288 154284
rect 260340 154272 260346 154284
rect 299474 154272 299480 154284
rect 260340 154244 299480 154272
rect 260340 154232 260346 154244
rect 299474 154232 299480 154244
rect 299532 154232 299538 154284
rect 373258 154232 373264 154284
rect 373316 154272 373322 154284
rect 542446 154272 542452 154284
rect 373316 154244 542452 154272
rect 373316 154232 373322 154244
rect 542446 154232 542452 154244
rect 542504 154232 542510 154284
rect 175274 154164 175280 154216
rect 175332 154204 175338 154216
rect 289814 154204 289820 154216
rect 175332 154176 289820 154204
rect 175332 154164 175338 154176
rect 289814 154164 289820 154176
rect 289872 154164 289878 154216
rect 291194 154164 291200 154216
rect 291252 154204 291258 154216
rect 340138 154204 340144 154216
rect 291252 154176 340144 154204
rect 291252 154164 291258 154176
rect 340138 154164 340144 154176
rect 340196 154164 340202 154216
rect 397086 154164 397092 154216
rect 397144 154204 397150 154216
rect 573450 154204 573456 154216
rect 397144 154176 573456 154204
rect 397144 154164 397150 154176
rect 573450 154164 573456 154176
rect 573508 154164 573514 154216
rect 106274 154096 106280 154148
rect 106332 154136 106338 154148
rect 308582 154136 308588 154148
rect 106332 154108 308588 154136
rect 106332 154096 106338 154108
rect 308582 154096 308588 154108
rect 308640 154096 308646 154148
rect 313734 154096 313740 154148
rect 313792 154136 313798 154148
rect 377306 154136 377312 154148
rect 313792 154108 377312 154136
rect 313792 154096 313798 154108
rect 377306 154096 377312 154108
rect 377364 154096 377370 154148
rect 387058 154096 387064 154148
rect 387116 154136 387122 154148
rect 572162 154136 572168 154148
rect 387116 154108 572168 154136
rect 387116 154096 387122 154108
rect 572162 154096 572168 154108
rect 572220 154096 572226 154148
rect 73246 154028 73252 154080
rect 73304 154068 73310 154080
rect 223942 154068 223948 154080
rect 73304 154040 223948 154068
rect 73304 154028 73310 154040
rect 223942 154028 223948 154040
rect 224000 154028 224006 154080
rect 224862 154028 224868 154080
rect 224920 154068 224926 154080
rect 581454 154068 581460 154080
rect 224920 154040 581460 154068
rect 224920 154028 224926 154040
rect 581454 154028 581460 154040
rect 581512 154028 581518 154080
rect 91094 153960 91100 154012
rect 91152 154000 91158 154012
rect 166902 154000 166908 154012
rect 91152 153972 166908 154000
rect 91152 153960 91158 153972
rect 166902 153960 166908 153972
rect 166960 153960 166966 154012
rect 178034 153960 178040 154012
rect 178092 154000 178098 154012
rect 544194 154000 544200 154012
rect 178092 153972 544200 154000
rect 178092 153960 178098 153972
rect 544194 153960 544200 153972
rect 544252 153960 544258 154012
rect 31018 153892 31024 153944
rect 31076 153932 31082 153944
rect 519814 153932 519820 153944
rect 31076 153904 519820 153932
rect 31076 153892 31082 153904
rect 519814 153892 519820 153904
rect 519872 153892 519878 153944
rect 33870 153824 33876 153876
rect 33928 153864 33934 153876
rect 548426 153864 548432 153876
rect 33928 153836 548432 153864
rect 33928 153824 33934 153836
rect 548426 153824 548432 153836
rect 548484 153824 548490 153876
rect 251910 153212 251916 153264
rect 251968 153252 251974 153264
rect 259454 153252 259460 153264
rect 251968 153224 259460 153252
rect 251968 153212 251974 153224
rect 259454 153212 259460 153224
rect 259512 153212 259518 153264
rect 37734 153144 37740 153196
rect 37792 153184 37798 153196
rect 129550 153184 129556 153196
rect 37792 153156 129556 153184
rect 37792 153144 37798 153156
rect 129550 153144 129556 153156
rect 129608 153144 129614 153196
rect 135990 153144 135996 153196
rect 136048 153184 136054 153196
rect 224218 153184 224224 153196
rect 136048 153156 224224 153184
rect 136048 153144 136054 153156
rect 224218 153144 224224 153156
rect 224276 153144 224282 153196
rect 291194 153144 291200 153196
rect 291252 153184 291258 153196
rect 348694 153184 348700 153196
rect 291252 153156 348700 153184
rect 291252 153144 291258 153156
rect 348694 153144 348700 153156
rect 348752 153144 348758 153196
rect 385770 153144 385776 153196
rect 385828 153184 385834 153196
rect 391658 153184 391664 153196
rect 385828 153156 391664 153184
rect 385828 153144 385834 153156
rect 391658 153144 391664 153156
rect 391716 153144 391722 153196
rect 402698 153144 402704 153196
rect 402756 153184 402762 153196
rect 580166 153184 580172 153196
rect 402756 153156 580172 153184
rect 402756 153144 402762 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 46106 153076 46112 153128
rect 46164 153116 46170 153128
rect 141142 153116 141148 153128
rect 46164 153088 141148 153116
rect 46164 153076 46170 153088
rect 141142 153076 141148 153088
rect 141200 153076 141206 153128
rect 145006 153076 145012 153128
rect 145064 153116 145070 153128
rect 178126 153116 178132 153128
rect 145064 153088 178132 153116
rect 145064 153076 145070 153088
rect 178126 153076 178132 153088
rect 178184 153076 178190 153128
rect 179782 153076 179788 153128
rect 179840 153116 179846 153128
rect 216766 153116 216772 153128
rect 179840 153088 216772 153116
rect 179840 153076 179846 153088
rect 216766 153076 216772 153088
rect 216824 153076 216830 153128
rect 254486 153076 254492 153128
rect 254544 153116 254550 153128
rect 373442 153116 373448 153128
rect 254544 153088 373448 153116
rect 254544 153076 254550 153088
rect 373442 153076 373448 153088
rect 373500 153076 373506 153128
rect 378778 153076 378784 153128
rect 378836 153116 378842 153128
rect 414842 153116 414848 153128
rect 378836 153088 414848 153116
rect 378836 153076 378842 153088
rect 414842 153076 414848 153088
rect 414900 153076 414906 153128
rect 482922 153076 482928 153128
rect 482980 153116 482986 153128
rect 555418 153116 555424 153128
rect 482980 153088 555424 153116
rect 482980 153076 482986 153088
rect 555418 153076 555424 153088
rect 555476 153076 555482 153128
rect 56594 153008 56600 153060
rect 56652 153048 56658 153060
rect 208486 153048 208492 153060
rect 56652 153020 208492 153048
rect 56652 153008 56658 153020
rect 208486 153008 208492 153020
rect 208544 153008 208550 153060
rect 209406 153008 209412 153060
rect 209464 153048 209470 153060
rect 354674 153048 354680 153060
rect 209464 153020 354680 153048
rect 209464 153008 209470 153020
rect 354674 153008 354680 153020
rect 354732 153008 354738 153060
rect 354766 153008 354772 153060
rect 354824 153048 354830 153060
rect 363598 153048 363604 153060
rect 354824 153020 363604 153048
rect 354824 153008 354830 153020
rect 363598 153008 363604 153020
rect 363656 153008 363662 153060
rect 403618 153008 403624 153060
rect 403676 153048 403682 153060
rect 448974 153048 448980 153060
rect 403676 153020 448980 153048
rect 403676 153008 403682 153020
rect 448974 153008 448980 153020
rect 449032 153008 449038 153060
rect 499666 153008 499672 153060
rect 499724 153048 499730 153060
rect 580350 153048 580356 153060
rect 499724 153020 580356 153048
rect 499724 153008 499730 153020
rect 580350 153008 580356 153020
rect 580408 153008 580414 153060
rect 38378 152940 38384 152992
rect 38436 152980 38442 152992
rect 209774 152980 209780 152992
rect 38436 152952 209780 152980
rect 38436 152940 38442 152952
rect 209774 152940 209780 152952
rect 209832 152940 209838 152992
rect 213914 152940 213920 152992
rect 213972 152980 213978 152992
rect 384298 152980 384304 152992
rect 213972 152952 384304 152980
rect 213972 152940 213978 152952
rect 384298 152940 384304 152952
rect 384356 152940 384362 152992
rect 394050 152940 394056 152992
rect 394108 152980 394114 152992
rect 447686 152980 447692 152992
rect 394108 152952 447692 152980
rect 394108 152940 394114 152952
rect 447686 152940 447692 152952
rect 447744 152940 447750 152992
rect 462406 152940 462412 152992
rect 462464 152980 462470 152992
rect 563330 152980 563336 152992
rect 462464 152952 563336 152980
rect 462464 152940 462470 152952
rect 563330 152940 563336 152952
rect 563388 152940 563394 152992
rect 51350 152872 51356 152924
rect 51408 152912 51414 152924
rect 126974 152912 126980 152924
rect 51408 152884 126980 152912
rect 51408 152872 51414 152884
rect 126974 152872 126980 152884
rect 127032 152872 127038 152924
rect 127618 152872 127624 152924
rect 127676 152912 127682 152924
rect 315298 152912 315304 152924
rect 127676 152884 315304 152912
rect 127676 152872 127682 152884
rect 315298 152872 315304 152884
rect 315356 152872 315362 152924
rect 316586 152872 316592 152924
rect 316644 152912 316650 152924
rect 360286 152912 360292 152924
rect 316644 152884 360292 152912
rect 316644 152872 316650 152884
rect 360286 152872 360292 152884
rect 360344 152872 360350 152924
rect 364978 152872 364984 152924
rect 365036 152912 365042 152924
rect 421926 152912 421932 152924
rect 365036 152884 421932 152912
rect 365036 152872 365042 152884
rect 421926 152872 421932 152884
rect 421984 152872 421990 152924
rect 451274 152872 451280 152924
rect 451332 152912 451338 152924
rect 561858 152912 561864 152924
rect 451332 152884 561864 152912
rect 451332 152872 451338 152884
rect 561858 152872 561864 152884
rect 561916 152872 561922 152924
rect 44910 152804 44916 152856
rect 44968 152844 44974 152856
rect 160094 152844 160100 152856
rect 44968 152816 160100 152844
rect 44968 152804 44974 152816
rect 160094 152804 160100 152816
rect 160152 152804 160158 152856
rect 200390 152804 200396 152856
rect 200448 152844 200454 152856
rect 392578 152844 392584 152856
rect 200448 152816 392584 152844
rect 200448 152804 200454 152816
rect 392578 152804 392584 152816
rect 392636 152804 392642 152856
rect 398190 152804 398196 152856
rect 398248 152844 398254 152856
rect 529198 152844 529204 152856
rect 398248 152816 529204 152844
rect 398248 152804 398254 152816
rect 529198 152804 529204 152816
rect 529256 152804 529262 152856
rect 531406 152804 531412 152856
rect 531464 152844 531470 152856
rect 534718 152844 534724 152856
rect 531464 152816 534724 152844
rect 531464 152804 531470 152816
rect 534718 152804 534724 152816
rect 534776 152804 534782 152856
rect 536098 152804 536104 152856
rect 536156 152844 536162 152856
rect 539778 152844 539784 152856
rect 536156 152816 539784 152844
rect 536156 152804 536162 152816
rect 539778 152804 539784 152816
rect 539836 152804 539842 152856
rect 543090 152804 543096 152856
rect 543148 152844 543154 152856
rect 561674 152844 561680 152856
rect 543148 152816 561680 152844
rect 543148 152804 543154 152816
rect 561674 152804 561680 152816
rect 561732 152804 561738 152856
rect 26970 152736 26976 152788
rect 27028 152776 27034 152788
rect 107654 152776 107660 152788
rect 27028 152748 107660 152776
rect 27028 152736 27034 152748
rect 107654 152736 107660 152748
rect 107712 152736 107718 152788
rect 122742 152736 122748 152788
rect 122800 152776 122806 152788
rect 330478 152776 330484 152788
rect 122800 152748 330484 152776
rect 122800 152736 122806 152748
rect 330478 152736 330484 152748
rect 330536 152736 330542 152788
rect 334986 152736 334992 152788
rect 335044 152776 335050 152788
rect 354766 152776 354772 152788
rect 335044 152748 354772 152776
rect 335044 152736 335050 152748
rect 354766 152736 354772 152748
rect 354824 152736 354830 152788
rect 354858 152736 354864 152788
rect 354916 152776 354922 152788
rect 358906 152776 358912 152788
rect 354916 152748 358912 152776
rect 354916 152736 354922 152748
rect 358906 152736 358912 152748
rect 358964 152736 358970 152788
rect 395430 152736 395436 152788
rect 395488 152776 395494 152788
rect 543826 152776 543832 152788
rect 395488 152748 543832 152776
rect 395488 152736 395494 152748
rect 543826 152736 543832 152748
rect 543884 152736 543890 152788
rect 547230 152736 547236 152788
rect 547288 152776 547294 152788
rect 566366 152776 566372 152788
rect 547288 152748 566372 152776
rect 547288 152736 547294 152748
rect 566366 152736 566372 152748
rect 566424 152736 566430 152788
rect 50338 152668 50344 152720
rect 50396 152708 50402 152720
rect 82538 152708 82544 152720
rect 50396 152680 82544 152708
rect 50396 152668 50402 152680
rect 82538 152668 82544 152680
rect 82596 152668 82602 152720
rect 106366 152668 106372 152720
rect 106424 152708 106430 152720
rect 358170 152708 358176 152720
rect 106424 152680 358176 152708
rect 106424 152668 106430 152680
rect 358170 152668 358176 152680
rect 358228 152668 358234 152720
rect 406010 152668 406016 152720
rect 406068 152708 406074 152720
rect 555326 152708 555332 152720
rect 406068 152680 555332 152708
rect 406068 152668 406074 152680
rect 555326 152668 555332 152680
rect 555384 152668 555390 152720
rect 35066 152600 35072 152652
rect 35124 152640 35130 152652
rect 297634 152640 297640 152652
rect 35124 152612 297640 152640
rect 35124 152600 35130 152612
rect 297634 152600 297640 152612
rect 297692 152600 297698 152652
rect 310514 152600 310520 152652
rect 310572 152640 310578 152652
rect 354858 152640 354864 152652
rect 310572 152612 354864 152640
rect 310572 152600 310578 152612
rect 354858 152600 354864 152612
rect 354916 152600 354922 152652
rect 354950 152600 354956 152652
rect 355008 152640 355014 152652
rect 362218 152640 362224 152652
rect 355008 152612 362224 152640
rect 355008 152600 355014 152612
rect 362218 152600 362224 152612
rect 362276 152600 362282 152652
rect 405458 152600 405464 152652
rect 405516 152640 405522 152652
rect 560754 152640 560760 152652
rect 405516 152612 560760 152640
rect 405516 152600 405522 152612
rect 560754 152600 560760 152612
rect 560812 152600 560818 152652
rect 36354 152532 36360 152584
rect 36412 152572 36418 152584
rect 326614 152572 326620 152584
rect 36412 152544 326620 152572
rect 36412 152532 36418 152544
rect 326614 152532 326620 152544
rect 326672 152532 326678 152584
rect 327258 152532 327264 152584
rect 327316 152572 327322 152584
rect 357618 152572 357624 152584
rect 327316 152544 357624 152572
rect 327316 152532 327322 152544
rect 357618 152532 357624 152544
rect 357676 152532 357682 152584
rect 401502 152532 401508 152584
rect 401560 152572 401566 152584
rect 561306 152572 561312 152584
rect 401560 152544 561312 152572
rect 401560 152532 401566 152544
rect 561306 152532 561312 152544
rect 561364 152532 561370 152584
rect 28350 152464 28356 152516
rect 28408 152504 28414 152516
rect 67082 152504 67088 152516
rect 28408 152476 67088 152504
rect 28408 152464 28414 152476
rect 67082 152464 67088 152476
rect 67140 152464 67146 152516
rect 81250 152464 81256 152516
rect 81308 152504 81314 152516
rect 377490 152504 377496 152516
rect 81308 152476 377496 152504
rect 81308 152464 81314 152476
rect 377490 152464 377496 152476
rect 377548 152464 377554 152516
rect 403526 152464 403532 152516
rect 403584 152504 403590 152516
rect 580442 152504 580448 152516
rect 403584 152476 580448 152504
rect 403584 152464 403590 152476
rect 580442 152464 580448 152476
rect 580500 152464 580506 152516
rect 51994 152396 52000 152448
rect 52052 152436 52058 152448
rect 57974 152436 57980 152448
rect 52052 152408 57980 152436
rect 52052 152396 52058 152408
rect 57974 152396 57980 152408
rect 58032 152396 58038 152448
rect 58158 152396 58164 152448
rect 58216 152436 58222 152448
rect 111794 152436 111800 152448
rect 58216 152408 111800 152436
rect 58216 152396 58222 152408
rect 111794 152396 111800 152408
rect 111852 152396 111858 152448
rect 315022 152396 315028 152448
rect 315080 152436 315086 152448
rect 359458 152436 359464 152448
rect 315080 152408 359464 152436
rect 315080 152396 315086 152408
rect 359458 152396 359464 152408
rect 359516 152396 359522 152448
rect 389910 152396 389916 152448
rect 389968 152436 389974 152448
rect 425146 152436 425152 152448
rect 389968 152408 425152 152436
rect 389968 152396 389974 152408
rect 425146 152396 425152 152408
rect 425204 152396 425210 152448
rect 498194 152396 498200 152448
rect 498252 152436 498258 152448
rect 557534 152436 557540 152448
rect 498252 152408 557540 152436
rect 498252 152396 498258 152408
rect 557534 152396 557540 152408
rect 557592 152396 557598 152448
rect 44358 152328 44364 152380
rect 44416 152368 44422 152380
rect 76742 152368 76748 152380
rect 44416 152340 76748 152368
rect 44416 152328 44422 152340
rect 76742 152328 76748 152340
rect 76800 152328 76806 152380
rect 94774 152328 94780 152380
rect 94832 152368 94838 152380
rect 121454 152368 121460 152380
rect 94832 152340 121460 152368
rect 94832 152328 94838 152340
rect 121454 152328 121460 152340
rect 121512 152328 121518 152380
rect 344002 152328 344008 152380
rect 344060 152368 344066 152380
rect 360194 152368 360200 152380
rect 344060 152340 360200 152368
rect 344060 152328 344066 152340
rect 360194 152328 360200 152340
rect 360252 152328 360258 152380
rect 399478 152328 399484 152380
rect 399536 152368 399542 152380
rect 434162 152368 434168 152380
rect 399536 152340 434168 152368
rect 399536 152328 399542 152340
rect 434162 152328 434168 152340
rect 434220 152328 434226 152380
rect 503070 152328 503076 152380
rect 503128 152368 503134 152380
rect 538858 152368 538864 152380
rect 503128 152340 538864 152368
rect 503128 152328 503134 152340
rect 538858 152328 538864 152340
rect 538916 152328 538922 152380
rect 540422 152328 540428 152380
rect 540480 152368 540486 152380
rect 543366 152368 543372 152380
rect 540480 152340 543372 152368
rect 540480 152328 540486 152340
rect 543366 152328 543372 152340
rect 543424 152328 543430 152380
rect 61286 152260 61292 152312
rect 61344 152300 61350 152312
rect 68278 152300 68284 152312
rect 61344 152272 68284 152300
rect 61344 152260 61350 152272
rect 68278 152260 68284 152272
rect 68336 152260 68342 152312
rect 347866 152260 347872 152312
rect 347924 152300 347930 152312
rect 358814 152300 358820 152312
rect 347924 152272 358820 152300
rect 347924 152260 347930 152272
rect 358814 152260 358820 152272
rect 358872 152260 358878 152312
rect 392762 152260 392768 152312
rect 392820 152300 392826 152312
rect 410334 152300 410340 152312
rect 392820 152272 410340 152300
rect 392820 152260 392826 152272
rect 410334 152260 410340 152272
rect 410392 152260 410398 152312
rect 505646 152260 505652 152312
rect 505704 152300 505710 152312
rect 518158 152300 518164 152312
rect 505704 152272 518164 152300
rect 505704 152260 505710 152272
rect 518158 152260 518164 152272
rect 518216 152260 518222 152312
rect 529198 152260 529204 152312
rect 529256 152300 529262 152312
rect 534626 152300 534632 152312
rect 529256 152272 534632 152300
rect 529256 152260 529262 152272
rect 534626 152260 534632 152272
rect 534684 152260 534690 152312
rect 68738 152192 68744 152244
rect 68796 152232 68802 152244
rect 69658 152232 69664 152244
rect 68796 152204 69664 152232
rect 68796 152192 68802 152204
rect 69658 152192 69664 152204
rect 69716 152192 69722 152244
rect 342070 152192 342076 152244
rect 342128 152232 342134 152244
rect 350718 152232 350724 152244
rect 342128 152204 350724 152232
rect 342128 152192 342134 152204
rect 350718 152192 350724 152204
rect 350776 152192 350782 152244
rect 526438 151920 526444 151972
rect 526496 151960 526502 151972
rect 528830 151960 528836 151972
rect 526496 151932 528836 151960
rect 526496 151920 526502 151932
rect 528830 151920 528836 151932
rect 528888 151920 528894 151972
rect 402330 151852 402336 151904
rect 402388 151892 402394 151904
rect 403250 151892 403256 151904
rect 402388 151864 403256 151892
rect 402388 151852 402394 151864
rect 403250 151852 403256 151864
rect 403308 151852 403314 151904
rect 50614 151716 50620 151768
rect 50672 151756 50678 151768
rect 96614 151756 96620 151768
rect 50672 151728 96620 151756
rect 50672 151716 50678 151728
rect 96614 151716 96620 151728
rect 96672 151716 96678 151768
rect 385494 151716 385500 151768
rect 385552 151756 385558 151768
rect 549162 151756 549168 151768
rect 385552 151728 549168 151756
rect 385552 151716 385558 151728
rect 549162 151716 549168 151728
rect 549220 151716 549226 151768
rect 52730 151648 52736 151700
rect 52788 151688 52794 151700
rect 113174 151688 113180 151700
rect 52788 151660 113180 151688
rect 52788 151648 52794 151660
rect 113174 151648 113180 151660
rect 113232 151648 113238 151700
rect 381906 151648 381912 151700
rect 381964 151688 381970 151700
rect 540974 151688 540980 151700
rect 381964 151660 540980 151688
rect 381964 151648 381970 151660
rect 540974 151648 540980 151660
rect 541032 151648 541038 151700
rect 59446 151580 59452 151632
rect 59504 151620 59510 151632
rect 198734 151620 198740 151632
rect 59504 151592 198740 151620
rect 59504 151580 59510 151592
rect 198734 151580 198740 151592
rect 198792 151580 198798 151632
rect 306374 151580 306380 151632
rect 306432 151620 306438 151632
rect 543734 151620 543740 151632
rect 306432 151592 543740 151620
rect 306432 151580 306438 151592
rect 543734 151580 543740 151592
rect 543792 151580 543798 151632
rect 52086 151512 52092 151564
rect 52144 151552 52150 151564
rect 113266 151552 113272 151564
rect 52144 151524 113272 151552
rect 52144 151512 52150 151524
rect 113266 151512 113272 151524
rect 113324 151512 113330 151564
rect 119890 151512 119896 151564
rect 119948 151552 119954 151564
rect 366174 151552 366180 151564
rect 119948 151524 366180 151552
rect 119948 151512 119954 151524
rect 366174 151512 366180 151524
rect 366232 151512 366238 151564
rect 399846 151512 399852 151564
rect 399904 151552 399910 151564
rect 564986 151552 564992 151564
rect 399904 151524 564992 151552
rect 399904 151512 399910 151524
rect 564986 151512 564992 151524
rect 565044 151512 565050 151564
rect 45278 151444 45284 151496
rect 45336 151484 45342 151496
rect 356330 151484 356336 151496
rect 45336 151456 356336 151484
rect 45336 151444 45342 151456
rect 356330 151444 356336 151456
rect 356388 151444 356394 151496
rect 381814 151444 381820 151496
rect 381872 151484 381878 151496
rect 549346 151484 549352 151496
rect 381872 151456 549352 151484
rect 381872 151444 381878 151456
rect 549346 151444 549352 151456
rect 549404 151444 549410 151496
rect 43990 151376 43996 151428
rect 44048 151416 44054 151428
rect 368750 151416 368756 151428
rect 44048 151388 368756 151416
rect 44048 151376 44054 151388
rect 368750 151376 368756 151388
rect 368808 151376 368814 151428
rect 392670 151376 392676 151428
rect 392728 151416 392734 151428
rect 569218 151416 569224 151428
rect 392728 151388 569224 151416
rect 392728 151376 392734 151388
rect 569218 151376 569224 151388
rect 569276 151376 569282 151428
rect 48038 151308 48044 151360
rect 48096 151348 48102 151360
rect 387794 151348 387800 151360
rect 48096 151320 387800 151348
rect 48096 151308 48102 151320
rect 387794 151308 387800 151320
rect 387852 151308 387858 151360
rect 395798 151308 395804 151360
rect 395856 151348 395862 151360
rect 573266 151348 573272 151360
rect 395856 151320 573272 151348
rect 395856 151308 395862 151320
rect 573266 151308 573272 151320
rect 573324 151308 573330 151360
rect 380342 151240 380348 151292
rect 380400 151280 380406 151292
rect 559834 151280 559840 151292
rect 380400 151252 559840 151280
rect 380400 151240 380406 151252
rect 559834 151240 559840 151252
rect 559892 151240 559898 151292
rect 46106 151172 46112 151224
rect 46164 151212 46170 151224
rect 412634 151212 412640 151224
rect 46164 151184 412640 151212
rect 46164 151172 46170 151184
rect 412634 151172 412640 151184
rect 412692 151172 412698 151224
rect 518894 151172 518900 151224
rect 518952 151212 518958 151224
rect 556890 151212 556896 151224
rect 518952 151184 556896 151212
rect 518952 151172 518958 151184
rect 556890 151172 556896 151184
rect 556948 151172 556954 151224
rect 50522 151104 50528 151156
rect 50580 151144 50586 151156
rect 75914 151144 75920 151156
rect 50580 151116 75920 151144
rect 50580 151104 50586 151116
rect 75914 151104 75920 151116
rect 75972 151104 75978 151156
rect 80054 151104 80060 151156
rect 80112 151144 80118 151156
rect 552382 151144 552388 151156
rect 80112 151116 552388 151144
rect 80112 151104 80118 151116
rect 552382 151104 552388 151116
rect 552440 151104 552446 151156
rect 28258 151036 28264 151088
rect 28316 151076 28322 151088
rect 572714 151076 572720 151088
rect 28316 151048 572720 151076
rect 28316 151036 28322 151048
rect 572714 151036 572720 151048
rect 572772 151036 572778 151088
rect 49142 150968 49148 151020
rect 49200 151008 49206 151020
rect 70486 151008 70492 151020
rect 49200 150980 70492 151008
rect 49200 150968 49206 150980
rect 70486 150968 70492 150980
rect 70544 150968 70550 151020
rect 407298 150968 407304 151020
rect 407356 151008 407362 151020
rect 567194 151008 567200 151020
rect 407356 150980 567200 151008
rect 407356 150968 407362 150980
rect 567194 150968 567200 150980
rect 567252 150968 567258 151020
rect 58986 150900 58992 150952
rect 59044 150940 59050 150952
rect 78674 150940 78680 150952
rect 59044 150912 78680 150940
rect 59044 150900 59050 150912
rect 78674 150900 78680 150912
rect 78732 150900 78738 150952
rect 383194 150900 383200 150952
rect 383252 150940 383258 150952
rect 537386 150940 537392 150952
rect 383252 150912 537392 150940
rect 383252 150900 383258 150912
rect 537386 150900 537392 150912
rect 537444 150900 537450 150952
rect 49234 150832 49240 150884
rect 49292 150872 49298 150884
rect 60734 150872 60740 150884
rect 49292 150844 60740 150872
rect 49292 150832 49298 150844
rect 60734 150832 60740 150844
rect 60792 150832 60798 150884
rect 537110 150832 537116 150884
rect 537168 150872 537174 150884
rect 540882 150872 540888 150884
rect 537168 150844 540888 150872
rect 537168 150832 537174 150844
rect 540882 150832 540888 150844
rect 540940 150832 540946 150884
rect 25498 150764 25504 150816
rect 25556 150804 25562 150816
rect 380710 150804 380716 150816
rect 25556 150776 380716 150804
rect 25556 150764 25562 150776
rect 380710 150764 380716 150776
rect 380768 150764 380774 150816
rect 539042 150424 539048 150476
rect 539100 150464 539106 150476
rect 540146 150464 540152 150476
rect 539100 150436 540152 150464
rect 539100 150424 539106 150436
rect 540146 150424 540152 150436
rect 540204 150424 540210 150476
rect 397178 150356 397184 150408
rect 397236 150396 397242 150408
rect 538858 150396 538864 150408
rect 397236 150368 538864 150396
rect 397236 150356 397242 150368
rect 538858 150356 538864 150368
rect 538916 150356 538922 150408
rect 539502 150356 539508 150408
rect 539560 150396 539566 150408
rect 539870 150396 539876 150408
rect 539560 150368 539876 150396
rect 539560 150356 539566 150368
rect 539870 150356 539876 150368
rect 539928 150356 539934 150408
rect 540698 150356 540704 150408
rect 540756 150396 540762 150408
rect 542170 150396 542176 150408
rect 540756 150368 542176 150396
rect 540756 150356 540762 150368
rect 542170 150356 542176 150368
rect 542228 150356 542234 150408
rect 545298 150396 545304 150408
rect 542372 150368 545304 150396
rect 537478 150288 537484 150340
rect 537536 150328 537542 150340
rect 540422 150328 540428 150340
rect 537536 150300 540428 150328
rect 537536 150288 537542 150300
rect 540422 150288 540428 150300
rect 540480 150288 540486 150340
rect 539410 150220 539416 150272
rect 539468 150260 539474 150272
rect 542372 150260 542400 150368
rect 545298 150356 545304 150368
rect 545356 150356 545362 150408
rect 539468 150232 542400 150260
rect 539468 150220 539474 150232
rect 54386 150152 54392 150204
rect 54444 150192 54450 150204
rect 59538 150192 59544 150204
rect 54444 150164 59544 150192
rect 54444 150152 54450 150164
rect 59538 150152 59544 150164
rect 59596 150152 59602 150204
rect 538950 150152 538956 150204
rect 539008 150192 539014 150204
rect 545574 150192 545580 150204
rect 539008 150164 545580 150192
rect 539008 150152 539014 150164
rect 545574 150152 545580 150164
rect 545632 150152 545638 150204
rect 48774 150084 48780 150136
rect 48832 150124 48838 150136
rect 59906 150124 59912 150136
rect 48832 150096 59912 150124
rect 48832 150084 48838 150096
rect 59906 150084 59912 150096
rect 59964 150084 59970 150136
rect 539594 150084 539600 150136
rect 539652 150124 539658 150136
rect 551186 150124 551192 150136
rect 539652 150096 551192 150124
rect 539652 150084 539658 150096
rect 551186 150084 551192 150096
rect 551244 150084 551250 150136
rect 57330 150016 57336 150068
rect 57388 150056 57394 150068
rect 255314 150056 255320 150068
rect 57388 150028 255320 150056
rect 57388 150016 57394 150028
rect 255314 150016 255320 150028
rect 255372 150016 255378 150068
rect 523586 150056 523592 150068
rect 518866 150028 523592 150056
rect 59262 149948 59268 150000
rect 59320 149988 59326 150000
rect 293954 149988 293960 150000
rect 59320 149960 293960 149988
rect 59320 149948 59326 149960
rect 293954 149948 293960 149960
rect 294012 149948 294018 150000
rect 52914 149880 52920 149932
rect 52972 149920 52978 149932
rect 313274 149920 313280 149932
rect 52972 149892 313280 149920
rect 52972 149880 52978 149892
rect 313274 149880 313280 149892
rect 313332 149880 313338 149932
rect 366818 149920 366824 149932
rect 354646 149892 366824 149920
rect 51258 149812 51264 149864
rect 51316 149852 51322 149864
rect 354646 149852 354674 149892
rect 366818 149880 366824 149892
rect 366876 149880 366882 149932
rect 387426 149920 387432 149932
rect 373966 149892 387432 149920
rect 51316 149824 354674 149852
rect 51316 149812 51322 149824
rect 50154 149744 50160 149796
rect 50212 149784 50218 149796
rect 373966 149784 373994 149892
rect 387426 149880 387432 149892
rect 387484 149880 387490 149932
rect 488534 149880 488540 149932
rect 488592 149880 488598 149932
rect 50212 149756 373994 149784
rect 488552 149784 488580 149880
rect 518866 149784 518894 150028
rect 523586 150016 523592 150028
rect 523644 150016 523650 150068
rect 488552 149756 518894 149784
rect 523512 149960 529934 149988
rect 50212 149744 50218 149756
rect 3326 149676 3332 149728
rect 3384 149716 3390 149728
rect 3384 149688 518894 149716
rect 3384 149676 3390 149688
rect 518866 149648 518894 149688
rect 523512 149648 523540 149960
rect 523586 149880 523592 149932
rect 523644 149920 523650 149932
rect 529906 149920 529934 149960
rect 537386 149948 537392 150000
rect 537444 149988 537450 150000
rect 543182 149988 543188 150000
rect 537444 149960 543188 149988
rect 537444 149948 537450 149960
rect 543182 149948 543188 149960
rect 543240 149948 543246 150000
rect 538766 149920 538772 149932
rect 523644 149892 528554 149920
rect 529906 149892 531314 149920
rect 523644 149880 523650 149892
rect 528526 149852 528554 149892
rect 531286 149852 531314 149892
rect 534046 149892 538772 149920
rect 534046 149852 534074 149892
rect 538766 149880 538772 149892
rect 538824 149880 538830 149932
rect 539042 149880 539048 149932
rect 539100 149920 539106 149932
rect 539100 149892 539180 149920
rect 539100 149880 539106 149892
rect 528526 149824 529796 149852
rect 531286 149824 534074 149852
rect 539152 149852 539180 149892
rect 539410 149880 539416 149932
rect 539468 149920 539474 149932
rect 550634 149920 550640 149932
rect 539468 149892 550640 149920
rect 539468 149880 539474 149892
rect 550634 149880 550640 149892
rect 550692 149880 550698 149932
rect 540698 149852 540704 149864
rect 539152 149824 540704 149852
rect 529768 149716 529796 149824
rect 540698 149812 540704 149824
rect 540756 149812 540762 149864
rect 546034 149812 546040 149864
rect 546092 149852 546098 149864
rect 560386 149852 560392 149864
rect 546092 149824 560392 149852
rect 546092 149812 546098 149824
rect 560386 149812 560392 149824
rect 560444 149812 560450 149864
rect 549806 149784 549812 149796
rect 531286 149756 549812 149784
rect 531286 149716 531314 149756
rect 549806 149744 549812 149756
rect 549864 149744 549870 149796
rect 551370 149744 551376 149796
rect 551428 149784 551434 149796
rect 565446 149784 565452 149796
rect 551428 149756 565452 149784
rect 551428 149744 551434 149756
rect 565446 149744 565452 149756
rect 565504 149744 565510 149796
rect 529768 149688 531314 149716
rect 543550 149676 543556 149728
rect 543608 149716 543614 149728
rect 565814 149716 565820 149728
rect 543608 149688 565820 149716
rect 543608 149676 543614 149688
rect 565814 149676 565820 149688
rect 565872 149676 565878 149728
rect 518866 149620 523540 149648
rect 546126 148996 546132 149048
rect 546184 149036 546190 149048
rect 548702 149036 548708 149048
rect 546184 149008 548708 149036
rect 546184 148996 546190 149008
rect 548702 148996 548708 149008
rect 548760 148996 548766 149048
rect 547782 148316 547788 148368
rect 547840 148356 547846 148368
rect 568574 148356 568580 148368
rect 547840 148328 568580 148356
rect 547840 148316 547846 148328
rect 568574 148316 568580 148328
rect 568632 148316 568638 148368
rect 541894 148248 541900 148300
rect 541952 148288 541958 148300
rect 545482 148288 545488 148300
rect 541952 148260 545488 148288
rect 541952 148248 541958 148260
rect 545482 148248 545488 148260
rect 545540 148248 545546 148300
rect 547138 147636 547144 147688
rect 547196 147676 547202 147688
rect 547966 147676 547972 147688
rect 547196 147648 547972 147676
rect 547196 147636 547202 147648
rect 547966 147636 547972 147648
rect 548024 147636 548030 147688
rect 540698 147568 540704 147620
rect 540756 147608 540762 147620
rect 542262 147608 542268 147620
rect 540756 147580 542268 147608
rect 540756 147568 540762 147580
rect 542262 147568 542268 147580
rect 542320 147568 542326 147620
rect 543458 147568 543464 147620
rect 543516 147608 543522 147620
rect 564526 147608 564532 147620
rect 543516 147580 564532 147608
rect 543516 147568 543522 147580
rect 564526 147568 564532 147580
rect 564584 147568 564590 147620
rect 552842 147500 552848 147552
rect 552900 147540 552906 147552
rect 559742 147540 559748 147552
rect 552900 147512 559748 147540
rect 552900 147500 552906 147512
rect 559742 147500 559748 147512
rect 559800 147500 559806 147552
rect 542170 146956 542176 147008
rect 542228 146996 542234 147008
rect 542906 146996 542912 147008
rect 542228 146968 542912 146996
rect 542228 146956 542234 146968
rect 542906 146956 542912 146968
rect 542964 146956 542970 147008
rect 540882 146888 540888 146940
rect 540940 146928 540946 146940
rect 545022 146928 545028 146940
rect 540940 146900 545028 146928
rect 540940 146888 540946 146900
rect 545022 146888 545028 146900
rect 545080 146888 545086 146940
rect 555602 146888 555608 146940
rect 555660 146928 555666 146940
rect 564526 146928 564532 146940
rect 555660 146900 564532 146928
rect 555660 146888 555666 146900
rect 564526 146888 564532 146900
rect 564584 146888 564590 146940
rect 55122 146344 55128 146396
rect 55180 146384 55186 146396
rect 59538 146384 59544 146396
rect 55180 146356 59544 146384
rect 55180 146344 55186 146356
rect 59538 146344 59544 146356
rect 59596 146344 59602 146396
rect 58526 146276 58532 146328
rect 58584 146316 58590 146328
rect 59446 146316 59452 146328
rect 58584 146288 59452 146316
rect 58584 146276 58590 146288
rect 59446 146276 59452 146288
rect 59504 146276 59510 146328
rect 542814 146208 542820 146260
rect 542872 146248 542878 146260
rect 543826 146248 543832 146260
rect 542872 146220 543832 146248
rect 542872 146208 542878 146220
rect 543826 146208 543832 146220
rect 543884 146208 543890 146260
rect 546494 146140 546500 146192
rect 546552 146180 546558 146192
rect 548242 146180 548248 146192
rect 546552 146152 548248 146180
rect 546552 146140 546558 146152
rect 548242 146140 548248 146152
rect 548300 146140 548306 146192
rect 53466 146072 53472 146124
rect 53524 146112 53530 146124
rect 58434 146112 58440 146124
rect 53524 146084 58440 146112
rect 53524 146072 53530 146084
rect 58434 146072 58440 146084
rect 58492 146072 58498 146124
rect 543274 146072 543280 146124
rect 543332 146112 543338 146124
rect 547966 146112 547972 146124
rect 543332 146084 547972 146112
rect 543332 146072 543338 146084
rect 547966 146072 547972 146084
rect 548024 146072 548030 146124
rect 547230 146004 547236 146056
rect 547288 146044 547294 146056
rect 548242 146044 548248 146056
rect 547288 146016 548248 146044
rect 547288 146004 547294 146016
rect 548242 146004 548248 146016
rect 548300 146004 548306 146056
rect 546954 145868 546960 145920
rect 547012 145908 547018 145920
rect 547230 145908 547236 145920
rect 547012 145880 547236 145908
rect 547012 145868 547018 145880
rect 547230 145868 547236 145880
rect 547288 145868 547294 145920
rect 57422 144984 57428 145036
rect 57480 145024 57486 145036
rect 59354 145024 59360 145036
rect 57480 144996 59360 145024
rect 57480 144984 57486 144996
rect 59354 144984 59360 144996
rect 59412 144984 59418 145036
rect 541342 144848 541348 144900
rect 541400 144888 541406 144900
rect 542354 144888 542360 144900
rect 541400 144860 542360 144888
rect 541400 144848 541406 144860
rect 542354 144848 542360 144860
rect 542412 144848 542418 144900
rect 544378 144848 544384 144900
rect 544436 144888 544442 144900
rect 546954 144888 546960 144900
rect 544436 144860 546960 144888
rect 544436 144848 544442 144860
rect 546954 144848 546960 144860
rect 547012 144848 547018 144900
rect 542262 144508 542268 144560
rect 542320 144548 542326 144560
rect 546770 144548 546776 144560
rect 542320 144520 546776 144548
rect 542320 144508 542326 144520
rect 546770 144508 546776 144520
rect 546828 144508 546834 144560
rect 541710 144372 541716 144424
rect 541768 144412 541774 144424
rect 546770 144412 546776 144424
rect 541768 144384 546776 144412
rect 541768 144372 541774 144384
rect 546770 144372 546776 144384
rect 546828 144372 546834 144424
rect 544562 144236 544568 144288
rect 544620 144276 544626 144288
rect 560386 144276 560392 144288
rect 544620 144248 560392 144276
rect 544620 144236 544626 144248
rect 560386 144236 560392 144248
rect 560444 144236 560450 144288
rect 542998 144168 543004 144220
rect 543056 144208 543062 144220
rect 560846 144208 560852 144220
rect 543056 144180 560852 144208
rect 543056 144168 543062 144180
rect 560846 144168 560852 144180
rect 560904 144168 560910 144220
rect 545022 144100 545028 144152
rect 545080 144140 545086 144152
rect 547782 144140 547788 144152
rect 545080 144112 547788 144140
rect 545080 144100 545086 144112
rect 547782 144100 547788 144112
rect 547840 144100 547846 144152
rect 543090 144032 543096 144084
rect 543148 144072 543154 144084
rect 546494 144072 546500 144084
rect 543148 144044 546500 144072
rect 543148 144032 543154 144044
rect 546494 144032 546500 144044
rect 546552 144032 546558 144084
rect 55122 143596 55128 143608
rect 52472 143568 55128 143596
rect 51626 143488 51632 143540
rect 51684 143528 51690 143540
rect 52472 143528 52500 143568
rect 55122 143556 55128 143568
rect 55180 143556 55186 143608
rect 51684 143500 52500 143528
rect 51684 143488 51690 143500
rect 543274 143488 543280 143540
rect 543332 143528 543338 143540
rect 558914 143528 558920 143540
rect 543332 143500 558920 143528
rect 543332 143488 543338 143500
rect 558914 143488 558920 143500
rect 558972 143488 558978 143540
rect 542538 143420 542544 143472
rect 542596 143460 542602 143472
rect 543734 143460 543740 143472
rect 542596 143432 543740 143460
rect 542596 143420 542602 143432
rect 543734 143420 543740 143432
rect 543792 143420 543798 143472
rect 542906 143352 542912 143404
rect 542964 143392 542970 143404
rect 545114 143392 545120 143404
rect 542964 143364 545120 143392
rect 542964 143352 542970 143364
rect 545114 143352 545120 143364
rect 545172 143352 545178 143404
rect 543366 142536 543372 142588
rect 543424 142576 543430 142588
rect 548610 142576 548616 142588
rect 543424 142548 548616 142576
rect 543424 142536 543430 142548
rect 548610 142536 548616 142548
rect 548668 142536 548674 142588
rect 543458 142332 543464 142384
rect 543516 142372 543522 142384
rect 548150 142372 548156 142384
rect 543516 142344 548156 142372
rect 543516 142332 543522 142344
rect 548150 142332 548156 142344
rect 548208 142332 548214 142384
rect 53834 142128 53840 142180
rect 53892 142168 53898 142180
rect 55674 142168 55680 142180
rect 53892 142140 55680 142168
rect 53892 142128 53898 142140
rect 55674 142128 55680 142140
rect 55732 142128 55738 142180
rect 47854 142060 47860 142112
rect 47912 142100 47918 142112
rect 56686 142100 56692 142112
rect 47912 142072 56692 142100
rect 47912 142060 47918 142072
rect 56686 142060 56692 142072
rect 56744 142060 56750 142112
rect 57790 142060 57796 142112
rect 57848 142100 57854 142112
rect 59078 142100 59084 142112
rect 57848 142072 59084 142100
rect 57848 142060 57854 142072
rect 59078 142060 59084 142072
rect 59136 142060 59142 142112
rect 543550 142060 543556 142112
rect 543608 142100 543614 142112
rect 569126 142100 569132 142112
rect 543608 142072 569132 142100
rect 543608 142060 543614 142072
rect 569126 142060 569132 142072
rect 569184 142060 569190 142112
rect 542906 141652 542912 141704
rect 542964 141692 542970 141704
rect 545390 141692 545396 141704
rect 542964 141664 545396 141692
rect 542964 141652 542970 141664
rect 545390 141652 545396 141664
rect 545448 141652 545454 141704
rect 547414 141380 547420 141432
rect 547472 141420 547478 141432
rect 550726 141420 550732 141432
rect 547472 141392 550732 141420
rect 547472 141380 547478 141392
rect 550726 141380 550732 141392
rect 550784 141380 550790 141432
rect 546586 140904 546592 140956
rect 546644 140944 546650 140956
rect 547046 140944 547052 140956
rect 546644 140916 547052 140944
rect 546644 140904 546650 140916
rect 547046 140904 547052 140916
rect 547104 140904 547110 140956
rect 559558 140904 559564 140956
rect 559616 140944 559622 140956
rect 561122 140944 561128 140956
rect 559616 140916 561128 140944
rect 559616 140904 559622 140916
rect 561122 140904 561128 140916
rect 561180 140904 561186 140956
rect 547230 140836 547236 140888
rect 547288 140876 547294 140888
rect 547874 140876 547880 140888
rect 547288 140848 547880 140876
rect 547288 140836 547294 140848
rect 547874 140836 547880 140848
rect 547932 140836 547938 140888
rect 558270 140836 558276 140888
rect 558328 140876 558334 140888
rect 560294 140876 560300 140888
rect 558328 140848 560300 140876
rect 558328 140836 558334 140848
rect 560294 140836 560300 140848
rect 560352 140836 560358 140888
rect 51258 140768 51264 140820
rect 51316 140808 51322 140820
rect 55214 140808 55220 140820
rect 51316 140780 55220 140808
rect 51316 140768 51322 140780
rect 55214 140768 55220 140780
rect 55272 140768 55278 140820
rect 541802 140768 541808 140820
rect 541860 140808 541866 140820
rect 547046 140808 547052 140820
rect 541860 140780 547052 140808
rect 541860 140768 541866 140780
rect 547046 140768 547052 140780
rect 547104 140768 547110 140820
rect 547782 140768 547788 140820
rect 547840 140808 547846 140820
rect 548702 140808 548708 140820
rect 547840 140780 548708 140808
rect 547840 140768 547846 140780
rect 548702 140768 548708 140780
rect 548760 140768 548766 140820
rect 558362 140768 558368 140820
rect 558420 140808 558426 140820
rect 558914 140808 558920 140820
rect 558420 140780 558920 140808
rect 558420 140768 558426 140780
rect 558914 140768 558920 140780
rect 558972 140768 558978 140820
rect 32490 140700 32496 140752
rect 32548 140740 32554 140752
rect 56686 140740 56692 140752
rect 32548 140712 56692 140740
rect 32548 140700 32554 140712
rect 56686 140700 56692 140712
rect 56744 140700 56750 140752
rect 54570 140632 54576 140684
rect 54628 140672 54634 140684
rect 57238 140672 57244 140684
rect 54628 140644 57244 140672
rect 54628 140632 54634 140644
rect 57238 140632 57244 140644
rect 57296 140632 57302 140684
rect 545942 140428 545948 140480
rect 546000 140468 546006 140480
rect 548150 140468 548156 140480
rect 546000 140440 548156 140468
rect 546000 140428 546006 140440
rect 548150 140428 548156 140440
rect 548208 140428 548214 140480
rect 542814 140020 542820 140072
rect 542872 140060 542878 140072
rect 544102 140060 544108 140072
rect 542872 140032 544108 140060
rect 542872 140020 542878 140032
rect 544102 140020 544108 140032
rect 544160 140020 544166 140072
rect 47854 139408 47860 139460
rect 47912 139448 47918 139460
rect 48774 139448 48780 139460
rect 47912 139420 48780 139448
rect 47912 139408 47918 139420
rect 48774 139408 48780 139420
rect 48832 139408 48838 139460
rect 543366 139408 543372 139460
rect 543424 139448 543430 139460
rect 544562 139448 544568 139460
rect 543424 139420 544568 139448
rect 543424 139408 543430 139420
rect 544562 139408 544568 139420
rect 544620 139408 544626 139460
rect 544930 139408 544936 139460
rect 544988 139448 544994 139460
rect 545574 139448 545580 139460
rect 544988 139420 545580 139448
rect 544988 139408 544994 139420
rect 545574 139408 545580 139420
rect 545632 139408 545638 139460
rect 551922 139408 551928 139460
rect 551980 139448 551986 139460
rect 555510 139448 555516 139460
rect 551980 139420 555516 139448
rect 551980 139408 551986 139420
rect 555510 139408 555516 139420
rect 555568 139408 555574 139460
rect 543550 139340 543556 139392
rect 543608 139380 543614 139392
rect 559374 139380 559380 139392
rect 543608 139352 559380 139380
rect 543608 139340 543614 139352
rect 559374 139340 559380 139352
rect 559432 139340 559438 139392
rect 567930 139340 567936 139392
rect 567988 139380 567994 139392
rect 580534 139380 580540 139392
rect 567988 139352 580540 139380
rect 567988 139340 567994 139352
rect 580534 139340 580540 139352
rect 580592 139340 580598 139392
rect 549714 139272 549720 139324
rect 549772 139312 549778 139324
rect 555510 139312 555516 139324
rect 549772 139284 555516 139312
rect 549772 139272 549778 139284
rect 555510 139272 555516 139284
rect 555568 139272 555574 139324
rect 544654 139204 544660 139256
rect 544712 139244 544718 139256
rect 547966 139244 547972 139256
rect 544712 139216 547972 139244
rect 544712 139204 544718 139216
rect 547966 139204 547972 139216
rect 548024 139204 548030 139256
rect 51718 138728 51724 138780
rect 51776 138768 51782 138780
rect 52454 138768 52460 138780
rect 51776 138740 52460 138768
rect 51776 138728 51782 138740
rect 52454 138728 52460 138740
rect 52512 138728 52518 138780
rect 545022 137980 545028 138032
rect 545080 138020 545086 138032
rect 545390 138020 545396 138032
rect 545080 137992 545396 138020
rect 545080 137980 545086 137992
rect 545390 137980 545396 137992
rect 545448 137980 545454 138032
rect 17678 137912 17684 137964
rect 17736 137952 17742 137964
rect 57606 137952 57612 137964
rect 17736 137924 57612 137952
rect 17736 137912 17742 137924
rect 57606 137912 57612 137924
rect 57664 137912 57670 137964
rect 559742 137708 559748 137760
rect 559800 137748 559806 137760
rect 566458 137748 566464 137760
rect 559800 137720 566464 137748
rect 559800 137708 559806 137720
rect 566458 137708 566464 137720
rect 566516 137708 566522 137760
rect 559558 137300 559564 137352
rect 559616 137340 559622 137352
rect 566642 137340 566648 137352
rect 559616 137312 566648 137340
rect 559616 137300 559622 137312
rect 566642 137300 566648 137312
rect 566700 137300 566706 137352
rect 54570 137232 54576 137284
rect 54628 137272 54634 137284
rect 55214 137272 55220 137284
rect 54628 137244 55220 137272
rect 54628 137232 54634 137244
rect 55214 137232 55220 137244
rect 55272 137232 55278 137284
rect 542446 136620 542452 136672
rect 542504 136660 542510 136672
rect 542906 136660 542912 136672
rect 542504 136632 542912 136660
rect 542504 136620 542510 136632
rect 542906 136620 542912 136632
rect 542964 136620 542970 136672
rect 542814 136552 542820 136604
rect 542872 136592 542878 136604
rect 564618 136592 564624 136604
rect 542872 136564 564624 136592
rect 542872 136552 542878 136564
rect 564618 136552 564624 136564
rect 564676 136552 564682 136604
rect 58710 136484 58716 136536
rect 58768 136524 58774 136536
rect 58894 136524 58900 136536
rect 58768 136496 58900 136524
rect 58768 136484 58774 136496
rect 58894 136484 58900 136496
rect 58952 136484 58958 136536
rect 542446 136484 542452 136536
rect 542504 136524 542510 136536
rect 557534 136524 557540 136536
rect 542504 136496 557540 136524
rect 542504 136484 542510 136496
rect 557534 136484 557540 136496
rect 557592 136484 557598 136536
rect 544378 136416 544384 136468
rect 544436 136456 544442 136468
rect 547874 136456 547880 136468
rect 544436 136428 547880 136456
rect 544436 136416 544442 136428
rect 547874 136416 547880 136428
rect 547932 136416 547938 136468
rect 544930 136348 544936 136400
rect 544988 136388 544994 136400
rect 549254 136388 549260 136400
rect 544988 136360 549260 136388
rect 544988 136348 544994 136360
rect 549254 136348 549260 136360
rect 549312 136348 549318 136400
rect 53558 135872 53564 135924
rect 53616 135912 53622 135924
rect 57974 135912 57980 135924
rect 53616 135884 57980 135912
rect 53616 135872 53622 135884
rect 57974 135872 57980 135884
rect 58032 135872 58038 135924
rect 542262 135260 542268 135312
rect 542320 135300 542326 135312
rect 544654 135300 544660 135312
rect 542320 135272 544660 135300
rect 542320 135260 542326 135272
rect 544654 135260 544660 135272
rect 544712 135260 544718 135312
rect 26142 135192 26148 135244
rect 26200 135232 26206 135244
rect 57606 135232 57612 135244
rect 26200 135204 57612 135232
rect 26200 135192 26206 135204
rect 57606 135192 57612 135204
rect 57664 135192 57670 135244
rect 58434 135192 58440 135244
rect 58492 135232 58498 135244
rect 59354 135232 59360 135244
rect 58492 135204 59360 135232
rect 58492 135192 58498 135204
rect 59354 135192 59360 135204
rect 59412 135192 59418 135244
rect 542446 135192 542452 135244
rect 542504 135232 542510 135244
rect 572714 135232 572720 135244
rect 542504 135204 572720 135232
rect 542504 135192 542510 135204
rect 572714 135192 572720 135204
rect 572772 135192 572778 135244
rect 541986 135124 541992 135176
rect 542044 135164 542050 135176
rect 546678 135164 546684 135176
rect 542044 135136 546684 135164
rect 542044 135124 542050 135136
rect 546678 135124 546684 135136
rect 546736 135124 546742 135176
rect 548610 135124 548616 135176
rect 548668 135164 548674 135176
rect 549346 135164 549352 135176
rect 548668 135136 549352 135164
rect 548668 135124 548674 135136
rect 549346 135124 549352 135136
rect 549404 135124 549410 135176
rect 561030 135124 561036 135176
rect 561088 135164 561094 135176
rect 564434 135164 564440 135176
rect 561088 135136 564440 135164
rect 561088 135124 561094 135136
rect 564434 135124 564440 135136
rect 564492 135124 564498 135176
rect 558454 135056 558460 135108
rect 558512 135096 558518 135108
rect 563054 135096 563060 135108
rect 558512 135068 563060 135096
rect 558512 135056 558518 135068
rect 563054 135056 563060 135068
rect 563112 135056 563118 135108
rect 549990 134580 549996 134632
rect 550048 134620 550054 134632
rect 560294 134620 560300 134632
rect 550048 134592 560300 134620
rect 550048 134580 550054 134592
rect 560294 134580 560300 134592
rect 560352 134580 560358 134632
rect 545022 134512 545028 134564
rect 545080 134552 545086 134564
rect 556154 134552 556160 134564
rect 545080 134524 556160 134552
rect 545080 134512 545086 134524
rect 556154 134512 556160 134524
rect 556212 134512 556218 134564
rect 58710 134376 58716 134428
rect 58768 134416 58774 134428
rect 59262 134416 59268 134428
rect 58768 134388 59268 134416
rect 58768 134376 58774 134388
rect 59262 134376 59268 134388
rect 59320 134376 59326 134428
rect 543642 134240 543648 134292
rect 543700 134280 543706 134292
rect 547874 134280 547880 134292
rect 543700 134252 547880 134280
rect 543700 134240 543706 134252
rect 547874 134240 547880 134252
rect 547932 134240 547938 134292
rect 540238 134036 540244 134088
rect 540296 134076 540302 134088
rect 541710 134076 541716 134088
rect 540296 134048 541716 134076
rect 540296 134036 540302 134048
rect 541710 134036 541716 134048
rect 541768 134036 541774 134088
rect 541618 133968 541624 134020
rect 541676 134008 541682 134020
rect 546586 134008 546592 134020
rect 541676 133980 546592 134008
rect 541676 133968 541682 133980
rect 546586 133968 546592 133980
rect 546644 133968 546650 134020
rect 558178 133968 558184 134020
rect 558236 134008 558242 134020
rect 563882 134008 563888 134020
rect 558236 133980 563888 134008
rect 558236 133968 558242 133980
rect 563882 133968 563888 133980
rect 563940 133968 563946 134020
rect 540606 133900 540612 133952
rect 540664 133940 540670 133952
rect 541434 133940 541440 133952
rect 540664 133912 541440 133940
rect 540664 133900 540670 133912
rect 541434 133900 541440 133912
rect 541492 133900 541498 133952
rect 43070 133832 43076 133884
rect 43128 133872 43134 133884
rect 57606 133872 57612 133884
rect 43128 133844 57612 133872
rect 43128 133832 43134 133844
rect 57606 133832 57612 133844
rect 57664 133832 57670 133884
rect 540422 133152 540428 133204
rect 540480 133192 540486 133204
rect 540974 133192 540980 133204
rect 540480 133164 540980 133192
rect 540480 133152 540486 133164
rect 540974 133152 540980 133164
rect 541032 133152 541038 133204
rect 542078 132744 542084 132796
rect 542136 132784 542142 132796
rect 546954 132784 546960 132796
rect 542136 132756 546960 132784
rect 542136 132744 542142 132756
rect 546954 132744 546960 132756
rect 547012 132744 547018 132796
rect 541986 132608 541992 132660
rect 542044 132648 542050 132660
rect 549254 132648 549260 132660
rect 542044 132620 549260 132648
rect 542044 132608 542050 132620
rect 549254 132608 549260 132620
rect 549312 132608 549318 132660
rect 541894 132472 541900 132524
rect 541952 132512 541958 132524
rect 542814 132512 542820 132524
rect 541952 132484 542820 132512
rect 541952 132472 541958 132484
rect 542814 132472 542820 132484
rect 542872 132472 542878 132524
rect 47394 132404 47400 132456
rect 47452 132444 47458 132456
rect 57606 132444 57612 132456
rect 47452 132416 57612 132444
rect 47452 132404 47458 132416
rect 57606 132404 57612 132416
rect 57664 132404 57670 132456
rect 542446 132404 542452 132456
rect 542504 132444 542510 132456
rect 578234 132444 578240 132456
rect 542504 132416 578240 132444
rect 542504 132404 542510 132416
rect 578234 132404 578240 132416
rect 578292 132404 578298 132456
rect 541342 131112 541348 131164
rect 541400 131152 541406 131164
rect 543734 131152 543740 131164
rect 541400 131124 543740 131152
rect 541400 131112 541406 131124
rect 543734 131112 543740 131124
rect 543792 131112 543798 131164
rect 36446 131044 36452 131096
rect 36504 131084 36510 131096
rect 57606 131084 57612 131096
rect 36504 131056 57612 131084
rect 36504 131044 36510 131056
rect 57606 131044 57612 131056
rect 57664 131044 57670 131096
rect 541066 131044 541072 131096
rect 541124 131084 541130 131096
rect 541526 131084 541532 131096
rect 541124 131056 541532 131084
rect 541124 131044 541130 131056
rect 541526 131044 541532 131056
rect 541584 131044 541590 131096
rect 542446 131044 542452 131096
rect 542504 131084 542510 131096
rect 568574 131084 568580 131096
rect 542504 131056 568580 131084
rect 542504 131044 542510 131056
rect 568574 131044 568580 131056
rect 568632 131044 568638 131096
rect 542170 130976 542176 131028
rect 542228 131016 542234 131028
rect 543458 131016 543464 131028
rect 542228 130988 543464 131016
rect 542228 130976 542234 130988
rect 543458 130976 543464 130988
rect 543516 130976 543522 131028
rect 541710 130840 541716 130892
rect 541768 130880 541774 130892
rect 542170 130880 542176 130892
rect 541768 130852 542176 130880
rect 541768 130840 541774 130852
rect 542170 130840 542176 130852
rect 542228 130840 542234 130892
rect 541710 130704 541716 130756
rect 541768 130744 541774 130756
rect 543642 130744 543648 130756
rect 541768 130716 543648 130744
rect 541768 130704 541774 130716
rect 543642 130704 543648 130716
rect 543700 130704 543706 130756
rect 541802 130364 541808 130416
rect 541860 130404 541866 130416
rect 541986 130404 541992 130416
rect 541860 130376 541992 130404
rect 541860 130364 541866 130376
rect 541986 130364 541992 130376
rect 542044 130364 542050 130416
rect 541342 130296 541348 130348
rect 541400 130336 541406 130348
rect 548518 130336 548524 130348
rect 541400 130308 548524 130336
rect 541400 130296 541406 130308
rect 548518 130296 548524 130308
rect 548576 130296 548582 130348
rect 540238 129820 540244 129872
rect 540296 129860 540302 129872
rect 545482 129860 545488 129872
rect 540296 129832 545488 129860
rect 540296 129820 540302 129832
rect 545482 129820 545488 129832
rect 545540 129820 545546 129872
rect 548058 129752 548064 129804
rect 548116 129792 548122 129804
rect 549346 129792 549352 129804
rect 548116 129764 549352 129792
rect 548116 129752 548122 129764
rect 549346 129752 549352 129764
rect 549404 129752 549410 129804
rect 549990 129752 549996 129804
rect 550048 129792 550054 129804
rect 550634 129792 550640 129804
rect 550048 129764 550640 129792
rect 550048 129752 550054 129764
rect 550634 129752 550640 129764
rect 550692 129752 550698 129804
rect 50062 129684 50068 129736
rect 50120 129724 50126 129736
rect 57606 129724 57612 129736
rect 50120 129696 57612 129724
rect 50120 129684 50126 129696
rect 57606 129684 57612 129696
rect 57664 129684 57670 129736
rect 540882 129684 540888 129736
rect 540940 129724 540946 129736
rect 541802 129724 541808 129736
rect 540940 129696 541808 129724
rect 540940 129684 540946 129696
rect 541802 129684 541808 129696
rect 541860 129684 541866 129736
rect 542446 129684 542452 129736
rect 542504 129724 542510 129736
rect 561674 129724 561680 129736
rect 542504 129696 561680 129724
rect 542504 129684 542510 129696
rect 561674 129684 561680 129696
rect 561732 129684 561738 129736
rect 546494 129616 546500 129668
rect 546552 129656 546558 129668
rect 548150 129656 548156 129668
rect 546552 129628 548156 129656
rect 546552 129616 546558 129628
rect 548150 129616 548156 129628
rect 548208 129616 548214 129668
rect 546402 129140 546408 129192
rect 546460 129180 546466 129192
rect 552014 129180 552020 129192
rect 546460 129152 552020 129180
rect 546460 129140 546466 129152
rect 552014 129140 552020 129152
rect 552072 129140 552078 129192
rect 542262 129072 542268 129124
rect 542320 129112 542326 129124
rect 549714 129112 549720 129124
rect 542320 129084 549720 129112
rect 542320 129072 542326 129084
rect 549714 129072 549720 129084
rect 549772 129072 549778 129124
rect 540330 129004 540336 129056
rect 540388 129044 540394 129056
rect 549346 129044 549352 129056
rect 540388 129016 549352 129044
rect 540388 129004 540394 129016
rect 549346 129004 549352 129016
rect 549404 129004 549410 129056
rect 56686 128800 56692 128852
rect 56744 128840 56750 128852
rect 58526 128840 58532 128852
rect 56744 128812 58532 128840
rect 56744 128800 56750 128812
rect 58526 128800 58532 128812
rect 58584 128800 58590 128852
rect 544286 128324 544292 128376
rect 544344 128364 544350 128376
rect 545114 128364 545120 128376
rect 544344 128336 545120 128364
rect 544344 128324 544350 128336
rect 545114 128324 545120 128336
rect 545172 128324 545178 128376
rect 548610 128324 548616 128376
rect 548668 128364 548674 128376
rect 549806 128364 549812 128376
rect 548668 128336 549812 128364
rect 548668 128324 548674 128336
rect 549806 128324 549812 128336
rect 549864 128324 549870 128376
rect 36814 128256 36820 128308
rect 36872 128296 36878 128308
rect 57606 128296 57612 128308
rect 36872 128268 57612 128296
rect 36872 128256 36878 128268
rect 57606 128256 57612 128268
rect 57664 128256 57670 128308
rect 543550 128256 543556 128308
rect 543608 128296 543614 128308
rect 543608 128268 557534 128296
rect 543608 128256 543614 128268
rect 547690 128188 547696 128240
rect 547748 128228 547754 128240
rect 547874 128228 547880 128240
rect 547748 128200 547880 128228
rect 547748 128188 547754 128200
rect 547874 128188 547880 128200
rect 547932 128188 547938 128240
rect 557506 128228 557534 128268
rect 567194 128228 567200 128240
rect 557506 128200 567200 128228
rect 567194 128188 567200 128200
rect 567252 128188 567258 128240
rect 543826 127644 543832 127696
rect 543884 127684 543890 127696
rect 544102 127684 544108 127696
rect 543884 127656 544108 127684
rect 543884 127644 543890 127656
rect 544102 127644 544108 127656
rect 544160 127644 544166 127696
rect 58342 127576 58348 127628
rect 58400 127616 58406 127628
rect 59354 127616 59360 127628
rect 58400 127588 59360 127616
rect 58400 127576 58406 127588
rect 59354 127576 59360 127588
rect 59412 127576 59418 127628
rect 541894 127576 541900 127628
rect 541952 127616 541958 127628
rect 541952 127588 542032 127616
rect 541952 127576 541958 127588
rect 542004 127424 542032 127588
rect 562410 127576 562416 127628
rect 562468 127616 562474 127628
rect 564526 127616 564532 127628
rect 562468 127588 564532 127616
rect 562468 127576 562474 127588
rect 564526 127576 564532 127588
rect 564584 127576 564590 127628
rect 541986 127372 541992 127424
rect 542044 127372 542050 127424
rect 545022 126964 545028 127016
rect 545080 127004 545086 127016
rect 546494 127004 546500 127016
rect 545080 126976 546500 127004
rect 545080 126964 545086 126976
rect 546494 126964 546500 126976
rect 546552 126964 546558 127016
rect 50982 126896 50988 126948
rect 51040 126936 51046 126948
rect 51718 126936 51724 126948
rect 51040 126908 51724 126936
rect 51040 126896 51046 126908
rect 51718 126896 51724 126908
rect 51776 126896 51782 126948
rect 54662 126896 54668 126948
rect 54720 126936 54726 126948
rect 57606 126936 57612 126948
rect 54720 126908 57612 126936
rect 54720 126896 54726 126908
rect 57606 126896 57612 126908
rect 57664 126896 57670 126948
rect 57790 126896 57796 126948
rect 57848 126936 57854 126948
rect 58710 126936 58716 126948
rect 57848 126908 58716 126936
rect 57848 126896 57854 126908
rect 58710 126896 58716 126908
rect 58768 126896 58774 126948
rect 543642 126896 543648 126948
rect 543700 126936 543706 126948
rect 546862 126936 546868 126948
rect 543700 126908 546868 126936
rect 543700 126896 543706 126908
rect 546862 126896 546868 126908
rect 546920 126896 546926 126948
rect 562502 126896 562508 126948
rect 562560 126936 562566 126948
rect 565814 126936 565820 126948
rect 562560 126908 565820 126936
rect 562560 126896 562566 126908
rect 565814 126896 565820 126908
rect 565872 126896 565878 126948
rect 544470 126828 544476 126880
rect 544528 126868 544534 126880
rect 548150 126868 548156 126880
rect 544528 126840 548156 126868
rect 544528 126828 544534 126840
rect 548150 126828 548156 126840
rect 548208 126828 548214 126880
rect 540790 126760 540796 126812
rect 540848 126800 540854 126812
rect 544930 126800 544936 126812
rect 540848 126772 544936 126800
rect 540848 126760 540854 126772
rect 544930 126760 544936 126772
rect 544988 126760 544994 126812
rect 55122 126352 55128 126404
rect 55180 126392 55186 126404
rect 56686 126392 56692 126404
rect 55180 126364 56692 126392
rect 55180 126352 55186 126364
rect 56686 126352 56692 126364
rect 56744 126352 56750 126404
rect 540790 126216 540796 126268
rect 540848 126256 540854 126268
rect 543090 126256 543096 126268
rect 540848 126228 543096 126256
rect 540848 126216 540854 126228
rect 543090 126216 543096 126228
rect 543148 126216 543154 126268
rect 540330 125808 540336 125860
rect 540388 125848 540394 125860
rect 541618 125848 541624 125860
rect 540388 125820 541624 125848
rect 540388 125808 540394 125820
rect 541618 125808 541624 125820
rect 541676 125808 541682 125860
rect 541342 125604 541348 125656
rect 541400 125644 541406 125656
rect 541710 125644 541716 125656
rect 541400 125616 541716 125644
rect 541400 125604 541406 125616
rect 541710 125604 541716 125616
rect 541768 125604 541774 125656
rect 542538 125536 542544 125588
rect 542596 125576 542602 125588
rect 544010 125576 544016 125588
rect 542596 125548 544016 125576
rect 542596 125536 542602 125548
rect 544010 125536 544016 125548
rect 544068 125536 544074 125588
rect 545206 125536 545212 125588
rect 545264 125576 545270 125588
rect 546862 125576 546868 125588
rect 545264 125548 546868 125576
rect 545264 125536 545270 125548
rect 546862 125536 546868 125548
rect 546920 125536 546926 125588
rect 543550 125468 543556 125520
rect 543608 125508 543614 125520
rect 570782 125508 570788 125520
rect 543608 125480 570788 125508
rect 543608 125468 543614 125480
rect 570782 125468 570788 125480
rect 570840 125468 570846 125520
rect 540882 125400 540888 125452
rect 540940 125440 540946 125452
rect 544470 125440 544476 125452
rect 540940 125412 544476 125440
rect 540940 125400 540946 125412
rect 544470 125400 544476 125412
rect 544528 125400 544534 125452
rect 542446 125332 542452 125384
rect 542504 125372 542510 125384
rect 544102 125372 544108 125384
rect 542504 125344 544108 125372
rect 542504 125332 542510 125344
rect 544102 125332 544108 125344
rect 544160 125332 544166 125384
rect 58710 125264 58716 125316
rect 58768 125304 58774 125316
rect 59446 125304 59452 125316
rect 58768 125276 59452 125304
rect 58768 125264 58774 125276
rect 59446 125264 59452 125276
rect 59504 125264 59510 125316
rect 540422 125264 540428 125316
rect 540480 125304 540486 125316
rect 543826 125304 543832 125316
rect 540480 125276 543832 125304
rect 540480 125264 540486 125276
rect 543826 125264 543832 125276
rect 543884 125264 543890 125316
rect 51718 125060 51724 125112
rect 51776 125100 51782 125112
rect 56594 125100 56600 125112
rect 51776 125072 56600 125100
rect 51776 125060 51782 125072
rect 56594 125060 56600 125072
rect 56652 125060 56658 125112
rect 50430 124924 50436 124976
rect 50488 124964 50494 124976
rect 56686 124964 56692 124976
rect 50488 124936 56692 124964
rect 50488 124924 50494 124936
rect 56686 124924 56692 124936
rect 56744 124924 56750 124976
rect 545942 124856 545948 124908
rect 546000 124896 546006 124908
rect 566458 124896 566464 124908
rect 546000 124868 566464 124896
rect 546000 124856 546006 124868
rect 566458 124856 566464 124868
rect 566516 124856 566522 124908
rect 57146 124584 57152 124636
rect 57204 124624 57210 124636
rect 58618 124624 58624 124636
rect 57204 124596 58624 124624
rect 57204 124584 57210 124596
rect 58618 124584 58624 124596
rect 58676 124584 58682 124636
rect 546034 124244 546040 124296
rect 546092 124284 546098 124296
rect 547966 124284 547972 124296
rect 546092 124256 547972 124284
rect 546092 124244 546098 124256
rect 547966 124244 547972 124256
rect 548024 124244 548030 124296
rect 544378 124216 544384 124228
rect 542004 124188 544384 124216
rect 23014 124108 23020 124160
rect 23072 124148 23078 124160
rect 57606 124148 57612 124160
rect 23072 124120 57612 124148
rect 23072 124108 23078 124120
rect 57606 124108 57612 124120
rect 57664 124108 57670 124160
rect 59078 124108 59084 124160
rect 59136 124148 59142 124160
rect 59354 124148 59360 124160
rect 59136 124120 59360 124148
rect 59136 124108 59142 124120
rect 59354 124108 59360 124120
rect 59412 124108 59418 124160
rect 542004 124024 542032 124188
rect 544378 124176 544384 124188
rect 544436 124176 544442 124228
rect 541986 123972 541992 124024
rect 542044 123972 542050 124024
rect 541342 123904 541348 123956
rect 541400 123944 541406 123956
rect 543734 123944 543740 123956
rect 541400 123916 543740 123944
rect 541400 123904 541406 123916
rect 543734 123904 543740 123916
rect 543792 123904 543798 123956
rect 53650 123564 53656 123616
rect 53708 123604 53714 123616
rect 57974 123604 57980 123616
rect 53708 123576 57980 123604
rect 53708 123564 53714 123576
rect 57974 123564 57980 123576
rect 58032 123564 58038 123616
rect 53282 123496 53288 123548
rect 53340 123536 53346 123548
rect 58618 123536 58624 123548
rect 53340 123508 58624 123536
rect 53340 123496 53346 123508
rect 58618 123496 58624 123508
rect 58676 123496 58682 123548
rect 52362 123428 52368 123480
rect 52420 123468 52426 123480
rect 57882 123468 57888 123480
rect 52420 123440 57888 123468
rect 52420 123428 52426 123440
rect 57882 123428 57888 123440
rect 57940 123428 57946 123480
rect 544378 123428 544384 123480
rect 544436 123468 544442 123480
rect 552750 123468 552756 123480
rect 544436 123440 552756 123468
rect 544436 123428 544442 123440
rect 552750 123428 552756 123440
rect 552808 123428 552814 123480
rect 53742 123224 53748 123276
rect 53800 123264 53806 123276
rect 54570 123264 54576 123276
rect 53800 123236 54576 123264
rect 53800 123224 53806 123236
rect 54570 123224 54576 123236
rect 54628 123224 54634 123276
rect 57606 123156 57612 123208
rect 57664 123196 57670 123208
rect 57790 123196 57796 123208
rect 57664 123168 57796 123196
rect 57664 123156 57670 123168
rect 57790 123156 57796 123168
rect 57848 123156 57854 123208
rect 547138 122816 547144 122868
rect 547196 122856 547202 122868
rect 547874 122856 547880 122868
rect 547196 122828 547880 122856
rect 547196 122816 547202 122828
rect 547874 122816 547880 122828
rect 547932 122816 547938 122868
rect 543642 122748 543648 122800
rect 543700 122788 543706 122800
rect 559466 122788 559472 122800
rect 543700 122760 559472 122788
rect 543700 122748 543706 122760
rect 559466 122748 559472 122760
rect 559524 122748 559530 122800
rect 57422 121524 57428 121576
rect 57480 121564 57486 121576
rect 57480 121536 57560 121564
rect 57480 121524 57486 121536
rect 38010 121388 38016 121440
rect 38068 121428 38074 121440
rect 57422 121428 57428 121440
rect 38068 121400 57428 121428
rect 38068 121388 38074 121400
rect 57422 121388 57428 121400
rect 57480 121388 57486 121440
rect 57532 121360 57560 121536
rect 540698 121456 540704 121508
rect 540756 121496 540762 121508
rect 541986 121496 541992 121508
rect 540756 121468 541992 121496
rect 540756 121456 540762 121468
rect 541986 121456 541992 121468
rect 542044 121456 542050 121508
rect 550082 121456 550088 121508
rect 550140 121496 550146 121508
rect 550634 121496 550640 121508
rect 550140 121468 550640 121496
rect 550140 121456 550146 121468
rect 550634 121456 550640 121468
rect 550692 121456 550698 121508
rect 57882 121388 57888 121440
rect 57940 121428 57946 121440
rect 58894 121428 58900 121440
rect 57940 121400 58900 121428
rect 57940 121388 57946 121400
rect 58894 121388 58900 121400
rect 58952 121388 58958 121440
rect 543550 121388 543556 121440
rect 543608 121428 543614 121440
rect 558086 121428 558092 121440
rect 543608 121400 558092 121428
rect 543608 121388 543614 121400
rect 558086 121388 558092 121400
rect 558144 121388 558150 121440
rect 59446 121360 59452 121372
rect 57532 121332 59452 121360
rect 59446 121320 59452 121332
rect 59504 121320 59510 121372
rect 542998 120708 543004 120760
rect 543056 120748 543062 120760
rect 546770 120748 546776 120760
rect 543056 120720 546776 120748
rect 543056 120708 543062 120720
rect 546770 120708 546776 120720
rect 546828 120708 546834 120760
rect 57330 120164 57336 120216
rect 57388 120204 57394 120216
rect 59630 120204 59636 120216
rect 57388 120176 59636 120204
rect 57388 120164 57394 120176
rect 59630 120164 59636 120176
rect 59688 120164 59694 120216
rect 57790 120096 57796 120148
rect 57848 120136 57854 120148
rect 59814 120136 59820 120148
rect 57848 120108 59820 120136
rect 57848 120096 57854 120108
rect 59814 120096 59820 120108
rect 59872 120096 59878 120148
rect 55122 120028 55128 120080
rect 55180 120068 55186 120080
rect 56686 120068 56692 120080
rect 55180 120040 56692 120068
rect 55180 120028 55186 120040
rect 56686 120028 56692 120040
rect 56744 120028 56750 120080
rect 54754 119960 54760 120012
rect 54812 120000 54818 120012
rect 57422 120000 57428 120012
rect 54812 119972 57428 120000
rect 54812 119960 54818 119972
rect 57422 119960 57428 119972
rect 57480 119960 57486 120012
rect 50982 119416 50988 119468
rect 51040 119456 51046 119468
rect 54570 119456 54576 119468
rect 51040 119428 54576 119456
rect 51040 119416 51046 119428
rect 54570 119416 54576 119428
rect 54628 119416 54634 119468
rect 51810 117988 51816 118040
rect 51868 118028 51874 118040
rect 53926 118028 53932 118040
rect 51868 118000 53932 118028
rect 51868 117988 51874 118000
rect 53926 117988 53932 118000
rect 53984 117988 53990 118040
rect 544286 117988 544292 118040
rect 544344 118028 544350 118040
rect 546586 118028 546592 118040
rect 544344 118000 546592 118028
rect 544344 117988 544350 118000
rect 546586 117988 546592 118000
rect 546644 117988 546650 118040
rect 53190 117648 53196 117700
rect 53248 117688 53254 117700
rect 54386 117688 54392 117700
rect 53248 117660 54392 117688
rect 53248 117648 53254 117660
rect 54386 117648 54392 117660
rect 54444 117648 54450 117700
rect 50430 117580 50436 117632
rect 50488 117620 50494 117632
rect 53834 117620 53840 117632
rect 50488 117592 53840 117620
rect 50488 117580 50494 117592
rect 53834 117580 53840 117592
rect 53892 117580 53898 117632
rect 543642 117308 543648 117360
rect 543700 117348 543706 117360
rect 547414 117348 547420 117360
rect 543700 117320 547420 117348
rect 543700 117308 543706 117320
rect 547414 117308 547420 117320
rect 547472 117308 547478 117360
rect 23106 117240 23112 117292
rect 23164 117280 23170 117292
rect 57054 117280 57060 117292
rect 23164 117252 57060 117280
rect 23164 117240 23170 117252
rect 57054 117240 57060 117252
rect 57112 117240 57118 117292
rect 59262 117240 59268 117292
rect 59320 117280 59326 117292
rect 59538 117280 59544 117292
rect 59320 117252 59544 117280
rect 59320 117240 59326 117252
rect 59538 117240 59544 117252
rect 59596 117240 59602 117292
rect 542446 117240 542452 117292
rect 542504 117280 542510 117292
rect 556890 117280 556896 117292
rect 542504 117252 556896 117280
rect 542504 117240 542510 117252
rect 556890 117240 556896 117252
rect 556948 117240 556954 117292
rect 544562 117172 544568 117224
rect 544620 117212 544626 117224
rect 545114 117212 545120 117224
rect 544620 117184 545120 117212
rect 544620 117172 544626 117184
rect 545114 117172 545120 117184
rect 545172 117172 545178 117224
rect 546126 117172 546132 117224
rect 546184 117212 546190 117224
rect 547690 117212 547696 117224
rect 546184 117184 547696 117212
rect 546184 117172 546190 117184
rect 547690 117172 547696 117184
rect 547748 117172 547754 117224
rect 547782 117172 547788 117224
rect 547840 117212 547846 117224
rect 549806 117212 549812 117224
rect 547840 117184 549812 117212
rect 547840 117172 547846 117184
rect 549806 117172 549812 117184
rect 549864 117172 549870 117224
rect 542722 117104 542728 117156
rect 542780 117144 542786 117156
rect 546770 117144 546776 117156
rect 542780 117116 546776 117144
rect 542780 117104 542786 117116
rect 546770 117104 546776 117116
rect 546828 117104 546834 117156
rect 57882 117036 57888 117088
rect 57940 117076 57946 117088
rect 59446 117076 59452 117088
rect 57940 117048 59452 117076
rect 57940 117036 57946 117048
rect 59446 117036 59452 117048
rect 59504 117036 59510 117088
rect 59262 116968 59268 117020
rect 59320 117008 59326 117020
rect 59630 117008 59636 117020
rect 59320 116980 59636 117008
rect 59320 116968 59326 116980
rect 59630 116968 59636 116980
rect 59688 116968 59694 117020
rect 53742 116560 53748 116612
rect 53800 116600 53806 116612
rect 57974 116600 57980 116612
rect 53800 116572 57980 116600
rect 53800 116560 53806 116572
rect 57974 116560 57980 116572
rect 58032 116560 58038 116612
rect 540514 115948 540520 116000
rect 540572 115988 540578 116000
rect 541066 115988 541072 116000
rect 540572 115960 541072 115988
rect 540572 115948 540578 115960
rect 541066 115948 541072 115960
rect 541124 115948 541130 116000
rect 44634 115880 44640 115932
rect 44692 115920 44698 115932
rect 57422 115920 57428 115932
rect 44692 115892 57428 115920
rect 44692 115880 44698 115892
rect 57422 115880 57428 115892
rect 57480 115880 57486 115932
rect 544470 115880 544476 115932
rect 544528 115920 544534 115932
rect 545574 115920 545580 115932
rect 544528 115892 545580 115920
rect 544528 115880 544534 115892
rect 545574 115880 545580 115892
rect 545632 115880 545638 115932
rect 555510 115880 555516 115932
rect 555568 115920 555574 115932
rect 556890 115920 556896 115932
rect 555568 115892 556896 115920
rect 555568 115880 555574 115892
rect 556890 115880 556896 115892
rect 556948 115880 556954 115932
rect 543274 115812 543280 115864
rect 543332 115852 543338 115864
rect 546034 115852 546040 115864
rect 543332 115824 546040 115852
rect 543332 115812 543338 115824
rect 546034 115812 546040 115824
rect 546092 115812 546098 115864
rect 542078 115744 542084 115796
rect 542136 115784 542142 115796
rect 545482 115784 545488 115796
rect 542136 115756 545488 115784
rect 542136 115744 542142 115756
rect 545482 115744 545488 115756
rect 545540 115744 545546 115796
rect 542722 114792 542728 114844
rect 542780 114832 542786 114844
rect 547322 114832 547328 114844
rect 542780 114804 547328 114832
rect 542780 114792 542786 114804
rect 547322 114792 547328 114804
rect 547380 114792 547386 114844
rect 547138 114520 547144 114572
rect 547196 114560 547202 114572
rect 549346 114560 549352 114572
rect 547196 114532 549352 114560
rect 547196 114520 547202 114532
rect 549346 114520 549352 114532
rect 549404 114520 549410 114572
rect 44726 114452 44732 114504
rect 44784 114492 44790 114504
rect 57422 114492 57428 114504
rect 44784 114464 57428 114492
rect 44784 114452 44790 114464
rect 57422 114452 57428 114464
rect 57480 114452 57486 114504
rect 552014 114452 552020 114504
rect 552072 114492 552078 114504
rect 555510 114492 555516 114504
rect 552072 114464 555516 114492
rect 552072 114452 552078 114464
rect 555510 114452 555516 114464
rect 555568 114452 555574 114504
rect 549346 114384 549352 114436
rect 549404 114424 549410 114436
rect 549714 114424 549720 114436
rect 549404 114396 549720 114424
rect 549404 114384 549410 114396
rect 549714 114384 549720 114396
rect 549772 114384 549778 114436
rect 543366 113840 543372 113892
rect 543424 113880 543430 113892
rect 553302 113880 553308 113892
rect 543424 113852 553308 113880
rect 543424 113840 543430 113852
rect 553302 113840 553308 113852
rect 553360 113840 553366 113892
rect 543090 113772 543096 113824
rect 543148 113812 543154 113824
rect 564434 113812 564440 113824
rect 543148 113784 564440 113812
rect 543148 113772 543154 113784
rect 564434 113772 564440 113784
rect 564492 113772 564498 113824
rect 542446 113568 542452 113620
rect 542504 113608 542510 113620
rect 548334 113608 548340 113620
rect 542504 113580 548340 113608
rect 542504 113568 542510 113580
rect 548334 113568 548340 113580
rect 548392 113568 548398 113620
rect 542262 113160 542268 113212
rect 542320 113200 542326 113212
rect 549254 113200 549260 113212
rect 542320 113172 549260 113200
rect 542320 113160 542326 113172
rect 549254 113160 549260 113172
rect 549312 113160 549318 113212
rect 543642 113092 543648 113144
rect 543700 113132 543706 113144
rect 545206 113132 545212 113144
rect 543700 113104 545212 113132
rect 543700 113092 543706 113104
rect 545206 113092 545212 113104
rect 545264 113092 545270 113144
rect 576210 113092 576216 113144
rect 576268 113132 576274 113144
rect 580534 113132 580540 113144
rect 576268 113104 580540 113132
rect 576268 113092 576274 113104
rect 580534 113092 580540 113104
rect 580592 113092 580598 113144
rect 548702 112480 548708 112532
rect 548760 112520 548766 112532
rect 560294 112520 560300 112532
rect 548760 112492 560300 112520
rect 548760 112480 548766 112492
rect 560294 112480 560300 112492
rect 560352 112480 560358 112532
rect 54570 112412 54576 112464
rect 54628 112452 54634 112464
rect 57238 112452 57244 112464
rect 54628 112424 57244 112452
rect 54628 112412 54634 112424
rect 57238 112412 57244 112424
rect 57296 112412 57302 112464
rect 550082 112412 550088 112464
rect 550140 112452 550146 112464
rect 563054 112452 563060 112464
rect 550140 112424 563060 112452
rect 550140 112412 550146 112424
rect 563054 112412 563060 112424
rect 563112 112412 563118 112464
rect 540422 112004 540428 112056
rect 540480 112044 540486 112056
rect 544102 112044 544108 112056
rect 540480 112016 544108 112044
rect 540480 112004 540486 112016
rect 544102 112004 544108 112016
rect 544160 112004 544166 112056
rect 547046 111868 547052 111920
rect 547104 111908 547110 111920
rect 549346 111908 549352 111920
rect 547104 111880 549352 111908
rect 547104 111868 547110 111880
rect 549346 111868 549352 111880
rect 549404 111868 549410 111920
rect 541802 111800 541808 111852
rect 541860 111840 541866 111852
rect 543734 111840 543740 111852
rect 541860 111812 543740 111840
rect 541860 111800 541866 111812
rect 543734 111800 543740 111812
rect 543792 111800 543798 111852
rect 547230 111800 547236 111852
rect 547288 111840 547294 111852
rect 547874 111840 547880 111852
rect 547288 111812 547880 111840
rect 547288 111800 547294 111812
rect 547874 111800 547880 111812
rect 547932 111800 547938 111852
rect 548886 111800 548892 111852
rect 548944 111840 548950 111852
rect 550634 111840 550640 111852
rect 548944 111812 550640 111840
rect 548944 111800 548950 111812
rect 550634 111800 550640 111812
rect 550692 111800 550698 111852
rect 565170 111800 565176 111852
rect 565228 111840 565234 111852
rect 565814 111840 565820 111852
rect 565228 111812 565820 111840
rect 565228 111800 565234 111812
rect 565814 111800 565820 111812
rect 565872 111800 565878 111852
rect 546126 111732 546132 111784
rect 546184 111772 546190 111784
rect 548794 111772 548800 111784
rect 546184 111744 548800 111772
rect 546184 111732 546190 111744
rect 548794 111732 548800 111744
rect 548852 111732 548858 111784
rect 549714 111732 549720 111784
rect 549772 111772 549778 111784
rect 551370 111772 551376 111784
rect 549772 111744 551376 111772
rect 549772 111732 549778 111744
rect 551370 111732 551376 111744
rect 551428 111732 551434 111784
rect 53742 111188 53748 111240
rect 53800 111228 53806 111240
rect 59354 111228 59360 111240
rect 53800 111200 59360 111228
rect 53800 111188 53806 111200
rect 59354 111188 59360 111200
rect 59412 111188 59418 111240
rect 53650 111120 53656 111172
rect 53708 111160 53714 111172
rect 59630 111160 59636 111172
rect 53708 111132 59636 111160
rect 53708 111120 53714 111132
rect 59630 111120 59636 111132
rect 59688 111120 59694 111172
rect 54754 111052 54760 111104
rect 54812 111092 54818 111104
rect 56686 111092 56692 111104
rect 54812 111064 56692 111092
rect 54812 111052 54818 111064
rect 56686 111052 56692 111064
rect 56744 111052 56750 111104
rect 543182 111052 543188 111104
rect 543240 111092 543246 111104
rect 548242 111092 548248 111104
rect 543240 111064 548248 111092
rect 543240 111052 543246 111064
rect 548242 111052 548248 111064
rect 548300 111052 548306 111104
rect 553302 110984 553308 111036
rect 553360 111024 553366 111036
rect 556154 111024 556160 111036
rect 553360 110996 556160 111024
rect 553360 110984 553366 110996
rect 556154 110984 556160 110996
rect 556212 110984 556218 111036
rect 541710 110508 541716 110560
rect 541768 110548 541774 110560
rect 546954 110548 546960 110560
rect 541768 110520 546960 110548
rect 541768 110508 541774 110520
rect 546954 110508 546960 110520
rect 547012 110508 547018 110560
rect 540422 110440 540428 110492
rect 540480 110480 540486 110492
rect 544930 110480 544936 110492
rect 540480 110452 544936 110480
rect 540480 110440 540486 110452
rect 544930 110440 544936 110452
rect 544988 110440 544994 110492
rect 51626 110372 51632 110424
rect 51684 110412 51690 110424
rect 57330 110412 57336 110424
rect 51684 110384 57336 110412
rect 51684 110372 51690 110384
rect 57330 110372 57336 110384
rect 57388 110372 57394 110424
rect 542446 110372 542452 110424
rect 542504 110412 542510 110424
rect 572162 110412 572168 110424
rect 542504 110384 572168 110412
rect 542504 110372 542510 110384
rect 572162 110372 572168 110384
rect 572220 110372 572226 110424
rect 542262 110304 542268 110356
rect 542320 110344 542326 110356
rect 542906 110344 542912 110356
rect 542320 110316 542912 110344
rect 542320 110304 542326 110316
rect 542906 110304 542912 110316
rect 542964 110304 542970 110356
rect 542998 110304 543004 110356
rect 543056 110344 543062 110356
rect 543642 110344 543648 110356
rect 543056 110316 543648 110344
rect 543056 110304 543062 110316
rect 543642 110304 543648 110316
rect 543700 110304 543706 110356
rect 545390 110304 545396 110356
rect 545448 110344 545454 110356
rect 546494 110344 546500 110356
rect 545448 110316 546500 110344
rect 545448 110304 545454 110316
rect 546494 110304 546500 110316
rect 546552 110304 546558 110356
rect 543734 110236 543740 110288
rect 543792 110276 543798 110288
rect 547874 110276 547880 110288
rect 543792 110248 547880 110276
rect 543792 110236 543798 110248
rect 547874 110236 547880 110248
rect 547932 110236 547938 110288
rect 540882 109896 540888 109948
rect 540940 109936 540946 109948
rect 541434 109936 541440 109948
rect 540940 109908 541440 109936
rect 540940 109896 540946 109908
rect 541434 109896 541440 109908
rect 541492 109896 541498 109948
rect 540790 109556 540796 109608
rect 540848 109596 540854 109608
rect 542446 109596 542452 109608
rect 540848 109568 542452 109596
rect 540848 109556 540854 109568
rect 542446 109556 542452 109568
rect 542504 109556 542510 109608
rect 542538 109420 542544 109472
rect 542596 109460 542602 109472
rect 548426 109460 548432 109472
rect 542596 109432 548432 109460
rect 542596 109420 542602 109432
rect 548426 109420 548432 109432
rect 548484 109420 548490 109472
rect 542630 109352 542636 109404
rect 542688 109352 542694 109404
rect 542648 109064 542676 109352
rect 542630 109012 542636 109064
rect 542688 109012 542694 109064
rect 543274 109012 543280 109064
rect 543332 109052 543338 109064
rect 546862 109052 546868 109064
rect 543332 109024 546868 109052
rect 543332 109012 543338 109024
rect 546862 109012 546868 109024
rect 546920 109012 546926 109064
rect 55766 108944 55772 108996
rect 55824 108984 55830 108996
rect 56594 108984 56600 108996
rect 55824 108956 56600 108984
rect 55824 108944 55830 108956
rect 56594 108944 56600 108956
rect 56652 108944 56658 108996
rect 48958 108876 48964 108928
rect 49016 108916 49022 108928
rect 57514 108916 57520 108928
rect 49016 108888 57520 108916
rect 49016 108876 49022 108888
rect 57514 108876 57520 108888
rect 57572 108876 57578 108928
rect 48866 108808 48872 108860
rect 48924 108848 48930 108860
rect 57422 108848 57428 108860
rect 48924 108820 57428 108848
rect 48924 108808 48930 108820
rect 57422 108808 57428 108820
rect 57480 108808 57486 108860
rect 540698 108808 540704 108860
rect 540756 108848 540762 108860
rect 543642 108848 543648 108860
rect 540756 108820 543648 108848
rect 540756 108808 540762 108820
rect 543642 108808 543648 108820
rect 543700 108808 543706 108860
rect 47854 107584 47860 107636
rect 47912 107624 47918 107636
rect 48958 107624 48964 107636
rect 47912 107596 48964 107624
rect 47912 107584 47918 107596
rect 48958 107584 48964 107596
rect 49016 107584 49022 107636
rect 543182 107584 543188 107636
rect 543240 107624 543246 107636
rect 562226 107624 562232 107636
rect 543240 107596 562232 107624
rect 543240 107584 543246 107596
rect 562226 107584 562232 107596
rect 562284 107584 562290 107636
rect 541894 106904 541900 106956
rect 541952 106944 541958 106956
rect 544562 106944 544568 106956
rect 541952 106916 544568 106944
rect 541952 106904 541958 106916
rect 544562 106904 544568 106916
rect 544620 106904 544626 106956
rect 545022 106224 545028 106276
rect 545080 106264 545086 106276
rect 546494 106264 546500 106276
rect 545080 106236 546500 106264
rect 545080 106224 545086 106236
rect 546494 106224 546500 106236
rect 546552 106224 546558 106276
rect 542262 106156 542268 106208
rect 542320 106196 542326 106208
rect 546954 106196 546960 106208
rect 542320 106168 546960 106196
rect 542320 106156 542326 106168
rect 546954 106156 546960 106168
rect 547012 106156 547018 106208
rect 543182 105544 543188 105596
rect 543240 105584 543246 105596
rect 546586 105584 546592 105596
rect 543240 105556 546592 105584
rect 543240 105544 543246 105556
rect 546586 105544 546592 105556
rect 546644 105544 546650 105596
rect 543366 104864 543372 104916
rect 543424 104904 543430 104916
rect 543424 104876 547874 104904
rect 543424 104864 543430 104876
rect 40586 104796 40592 104848
rect 40644 104836 40650 104848
rect 57514 104836 57520 104848
rect 40644 104808 57520 104836
rect 40644 104796 40650 104808
rect 57514 104796 57520 104808
rect 57572 104796 57578 104848
rect 547846 104836 547874 104876
rect 548242 104836 548248 104848
rect 547846 104808 548248 104836
rect 548242 104796 548248 104808
rect 548300 104796 548306 104848
rect 53374 104728 53380 104780
rect 53432 104768 53438 104780
rect 56870 104768 56876 104780
rect 53432 104740 56876 104768
rect 53432 104728 53438 104740
rect 56870 104728 56876 104740
rect 56928 104728 56934 104780
rect 543734 104592 543740 104644
rect 543792 104632 543798 104644
rect 549714 104632 549720 104644
rect 543792 104604 549720 104632
rect 543792 104592 543798 104604
rect 549714 104592 549720 104604
rect 549772 104592 549778 104644
rect 543274 103572 543280 103624
rect 543332 103612 543338 103624
rect 548886 103612 548892 103624
rect 543332 103584 548892 103612
rect 543332 103572 543338 103584
rect 548886 103572 548892 103584
rect 548944 103572 548950 103624
rect 547782 103504 547788 103556
rect 547840 103544 547846 103556
rect 549806 103544 549812 103556
rect 547840 103516 549812 103544
rect 547840 103504 547846 103516
rect 549806 103504 549812 103516
rect 549864 103504 549870 103556
rect 23198 103436 23204 103488
rect 23256 103476 23262 103488
rect 57514 103476 57520 103488
rect 23256 103448 57520 103476
rect 23256 103436 23262 103448
rect 57514 103436 57520 103448
rect 57572 103436 57578 103488
rect 27430 103368 27436 103420
rect 27488 103408 27494 103420
rect 57882 103408 57888 103420
rect 27488 103380 57888 103408
rect 27488 103368 27494 103380
rect 57882 103368 57888 103380
rect 57940 103368 57946 103420
rect 542170 102620 542176 102672
rect 542228 102660 542234 102672
rect 546862 102660 546868 102672
rect 542228 102632 546868 102660
rect 542228 102620 542234 102632
rect 546862 102620 546868 102632
rect 546920 102620 546926 102672
rect 50154 102212 50160 102264
rect 50212 102252 50218 102264
rect 52454 102252 52460 102264
rect 50212 102224 52460 102252
rect 50212 102212 50218 102224
rect 52454 102212 52460 102224
rect 52512 102212 52518 102264
rect 53282 102144 53288 102196
rect 53340 102184 53346 102196
rect 53926 102184 53932 102196
rect 53340 102156 53932 102184
rect 53340 102144 53346 102156
rect 53926 102144 53932 102156
rect 53984 102144 53990 102196
rect 543458 102144 543464 102196
rect 543516 102184 543522 102196
rect 544470 102184 544476 102196
rect 543516 102156 544476 102184
rect 543516 102144 543522 102156
rect 544470 102144 544476 102156
rect 544528 102144 544534 102196
rect 43254 102076 43260 102128
rect 43312 102116 43318 102128
rect 57514 102116 57520 102128
rect 43312 102088 57520 102116
rect 43312 102076 43318 102088
rect 57514 102076 57520 102088
rect 57572 102076 57578 102128
rect 552658 101396 552664 101448
rect 552716 101436 552722 101448
rect 565446 101436 565452 101448
rect 552716 101408 565452 101436
rect 552716 101396 552722 101408
rect 565446 101396 565452 101408
rect 565504 101396 565510 101448
rect 31662 100648 31668 100700
rect 31720 100688 31726 100700
rect 57514 100688 57520 100700
rect 31720 100660 57520 100688
rect 31720 100648 31726 100660
rect 57514 100648 57520 100660
rect 57572 100648 57578 100700
rect 58802 100104 58808 100156
rect 58860 100144 58866 100156
rect 59078 100144 59084 100156
rect 58860 100116 59084 100144
rect 58860 100104 58866 100116
rect 59078 100104 59084 100116
rect 59136 100104 59142 100156
rect 542078 99968 542084 100020
rect 542136 100008 542142 100020
rect 549254 100008 549260 100020
rect 542136 99980 549260 100008
rect 542136 99968 542142 99980
rect 549254 99968 549260 99980
rect 549312 99968 549318 100020
rect 59262 98676 59268 98728
rect 59320 98716 59326 98728
rect 59814 98716 59820 98728
rect 59320 98688 59820 98716
rect 59320 98676 59326 98688
rect 59814 98676 59820 98688
rect 59872 98676 59878 98728
rect 548794 98676 548800 98728
rect 548852 98716 548858 98728
rect 549254 98716 549260 98728
rect 548852 98688 549260 98716
rect 548852 98676 548858 98688
rect 549254 98676 549260 98688
rect 549312 98676 549318 98728
rect 58434 98608 58440 98660
rect 58492 98648 58498 98660
rect 59446 98648 59452 98660
rect 58492 98620 59452 98648
rect 58492 98608 58498 98620
rect 59446 98608 59452 98620
rect 59504 98608 59510 98660
rect 58710 98540 58716 98592
rect 58768 98580 58774 98592
rect 59538 98580 59544 98592
rect 58768 98552 59544 98580
rect 58768 98540 58774 98552
rect 59538 98540 59544 98552
rect 59596 98540 59602 98592
rect 543550 97928 543556 97980
rect 543608 97968 543614 97980
rect 575474 97968 575480 97980
rect 543608 97940 575480 97968
rect 543608 97928 543614 97940
rect 575474 97928 575480 97940
rect 575532 97928 575538 97980
rect 52454 97860 52460 97912
rect 52512 97900 52518 97912
rect 55858 97900 55864 97912
rect 52512 97872 55864 97900
rect 52512 97860 52518 97872
rect 55858 97860 55864 97872
rect 55916 97860 55922 97912
rect 2866 97724 2872 97776
rect 2924 97764 2930 97776
rect 4798 97764 4804 97776
rect 2924 97736 4804 97764
rect 2924 97724 2930 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 53374 96568 53380 96620
rect 53432 96608 53438 96620
rect 53834 96608 53840 96620
rect 53432 96580 53840 96608
rect 53432 96568 53438 96580
rect 53834 96568 53840 96580
rect 53892 96568 53898 96620
rect 540974 96568 540980 96620
rect 541032 96608 541038 96620
rect 543458 96608 543464 96620
rect 541032 96580 543464 96608
rect 541032 96568 541038 96580
rect 543458 96568 543464 96580
rect 543516 96568 543522 96620
rect 543642 96568 543648 96620
rect 543700 96608 543706 96620
rect 578786 96608 578792 96620
rect 543700 96580 578792 96608
rect 543700 96568 543706 96580
rect 578786 96568 578792 96580
rect 578844 96568 578850 96620
rect 543550 96500 543556 96552
rect 543608 96540 543614 96552
rect 577222 96540 577228 96552
rect 543608 96512 577228 96540
rect 543608 96500 543614 96512
rect 577222 96500 577228 96512
rect 577280 96500 577286 96552
rect 542170 95888 542176 95940
rect 542228 95928 542234 95940
rect 551186 95928 551192 95940
rect 542228 95900 551192 95928
rect 542228 95888 542234 95900
rect 551186 95888 551192 95900
rect 551244 95888 551250 95940
rect 30926 95140 30932 95192
rect 30984 95180 30990 95192
rect 57514 95180 57520 95192
rect 30984 95152 57520 95180
rect 30984 95140 30990 95152
rect 57514 95140 57520 95152
rect 57572 95140 57578 95192
rect 540606 95140 540612 95192
rect 540664 95180 540670 95192
rect 542262 95180 542268 95192
rect 540664 95152 542268 95180
rect 540664 95140 540670 95152
rect 542262 95140 542268 95152
rect 542320 95140 542326 95192
rect 543550 95140 543556 95192
rect 543608 95180 543614 95192
rect 581822 95180 581828 95192
rect 543608 95152 581828 95180
rect 543608 95140 543614 95152
rect 581822 95140 581828 95152
rect 581880 95140 581886 95192
rect 53190 95072 53196 95124
rect 53248 95112 53254 95124
rect 54570 95112 54576 95124
rect 53248 95084 54576 95112
rect 53248 95072 53254 95084
rect 54570 95072 54576 95084
rect 54628 95072 54634 95124
rect 50246 93780 50252 93832
rect 50304 93820 50310 93832
rect 57514 93820 57520 93832
rect 50304 93792 57520 93820
rect 50304 93780 50310 93792
rect 57514 93780 57520 93792
rect 57572 93780 57578 93832
rect 543550 93780 543556 93832
rect 543608 93820 543614 93832
rect 552566 93820 552572 93832
rect 543608 93792 552572 93820
rect 543608 93780 543614 93792
rect 552566 93780 552572 93792
rect 552624 93780 552630 93832
rect 541986 92624 541992 92676
rect 542044 92664 542050 92676
rect 542446 92664 542452 92676
rect 542044 92636 542452 92664
rect 542044 92624 542050 92636
rect 542446 92624 542452 92636
rect 542504 92624 542510 92676
rect 542262 92488 542268 92540
rect 542320 92528 542326 92540
rect 542446 92528 542452 92540
rect 542320 92500 542452 92528
rect 542320 92488 542326 92500
rect 542446 92488 542452 92500
rect 542504 92488 542510 92540
rect 551370 92488 551376 92540
rect 551428 92528 551434 92540
rect 552014 92528 552020 92540
rect 551428 92500 552020 92528
rect 551428 92488 551434 92500
rect 552014 92488 552020 92500
rect 552072 92488 552078 92540
rect 543550 92420 543556 92472
rect 543608 92460 543614 92472
rect 574922 92460 574928 92472
rect 543608 92432 574928 92460
rect 543608 92420 543614 92432
rect 574922 92420 574928 92432
rect 574980 92420 574986 92472
rect 542814 92216 542820 92268
rect 542872 92256 542878 92268
rect 547966 92256 547972 92268
rect 542872 92228 547972 92256
rect 542872 92216 542878 92228
rect 547966 92216 547972 92228
rect 548024 92216 548030 92268
rect 542630 92148 542636 92200
rect 542688 92188 542694 92200
rect 544286 92188 544292 92200
rect 542688 92160 544292 92188
rect 542688 92148 542694 92160
rect 544286 92148 544292 92160
rect 544344 92148 544350 92200
rect 546402 91740 546408 91792
rect 546460 91780 546466 91792
rect 551186 91780 551192 91792
rect 546460 91752 551192 91780
rect 546460 91740 546466 91752
rect 551186 91740 551192 91752
rect 551244 91740 551250 91792
rect 551370 91740 551376 91792
rect 551428 91780 551434 91792
rect 565170 91780 565176 91792
rect 551428 91752 565176 91780
rect 551428 91740 551434 91752
rect 565170 91740 565176 91752
rect 565228 91740 565234 91792
rect 542814 91128 542820 91180
rect 542872 91168 542878 91180
rect 547874 91168 547880 91180
rect 542872 91140 547880 91168
rect 542872 91128 542878 91140
rect 547874 91128 547880 91140
rect 547932 91128 547938 91180
rect 546034 90312 546040 90364
rect 546092 90352 546098 90364
rect 556154 90352 556160 90364
rect 546092 90324 556160 90352
rect 546092 90312 546098 90324
rect 556154 90312 556160 90324
rect 556212 90312 556218 90364
rect 543642 89700 543648 89752
rect 543700 89740 543706 89752
rect 545574 89740 545580 89752
rect 543700 89712 545580 89740
rect 543700 89700 543706 89712
rect 545574 89700 545580 89712
rect 545632 89700 545638 89752
rect 546126 89700 546132 89752
rect 546184 89740 546190 89752
rect 547046 89740 547052 89752
rect 546184 89712 547052 89740
rect 546184 89700 546190 89712
rect 547046 89700 547052 89712
rect 547104 89700 547110 89752
rect 34422 89632 34428 89684
rect 34480 89672 34486 89684
rect 57606 89672 57612 89684
rect 34480 89644 57612 89672
rect 34480 89632 34486 89644
rect 57606 89632 57612 89644
rect 57664 89632 57670 89684
rect 542722 89632 542728 89684
rect 542780 89672 542786 89684
rect 569310 89672 569316 89684
rect 542780 89644 569316 89672
rect 542780 89632 542786 89644
rect 569310 89632 569316 89644
rect 569368 89632 569374 89684
rect 545022 89428 545028 89480
rect 545080 89468 545086 89480
rect 547322 89468 547328 89480
rect 545080 89440 547328 89468
rect 545080 89428 545086 89440
rect 547322 89428 547328 89440
rect 547380 89428 547386 89480
rect 544470 89020 544476 89072
rect 544528 89060 544534 89072
rect 547414 89060 547420 89072
rect 544528 89032 547420 89060
rect 544528 89020 544534 89032
rect 547414 89020 547420 89032
rect 547472 89020 547478 89072
rect 547230 88380 547236 88392
rect 544396 88352 547236 88380
rect 541342 88272 541348 88324
rect 541400 88312 541406 88324
rect 544286 88312 544292 88324
rect 541400 88284 544292 88312
rect 541400 88272 541406 88284
rect 544286 88272 544292 88284
rect 544344 88272 544350 88324
rect 542262 88204 542268 88256
rect 542320 88244 542326 88256
rect 544396 88244 544424 88352
rect 547230 88340 547236 88352
rect 547288 88340 547294 88392
rect 542320 88216 544424 88244
rect 542320 88204 542326 88216
rect 38194 86912 38200 86964
rect 38252 86952 38258 86964
rect 57606 86952 57612 86964
rect 38252 86924 57612 86952
rect 38252 86912 38258 86924
rect 57606 86912 57612 86924
rect 57664 86912 57670 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 21358 85524 21364 85536
rect 3568 85496 21364 85524
rect 3568 85484 3574 85496
rect 21358 85484 21364 85496
rect 21416 85484 21422 85536
rect 58250 85484 58256 85536
rect 58308 85524 58314 85536
rect 58434 85524 58440 85536
rect 58308 85496 58440 85524
rect 58308 85484 58314 85496
rect 58434 85484 58440 85496
rect 58492 85484 58498 85536
rect 543642 85484 543648 85536
rect 543700 85524 543706 85536
rect 544930 85524 544936 85536
rect 543700 85496 544936 85524
rect 543700 85484 543706 85496
rect 544930 85484 544936 85496
rect 544988 85484 544994 85536
rect 57514 85416 57520 85468
rect 57572 85456 57578 85468
rect 58526 85456 58532 85468
rect 57572 85428 58532 85456
rect 57572 85416 57578 85428
rect 58526 85416 58532 85428
rect 58584 85416 58590 85468
rect 542630 85076 542636 85128
rect 542688 85116 542694 85128
rect 544194 85116 544200 85128
rect 542688 85088 544200 85116
rect 542688 85076 542694 85088
rect 544194 85076 544200 85088
rect 544252 85076 544258 85128
rect 542170 84940 542176 84992
rect 542228 84980 542234 84992
rect 549806 84980 549812 84992
rect 542228 84952 549812 84980
rect 542228 84940 542234 84952
rect 549806 84940 549812 84952
rect 549864 84940 549870 84992
rect 55122 84192 55128 84244
rect 55180 84232 55186 84244
rect 57054 84232 57060 84244
rect 55180 84204 57060 84232
rect 55180 84192 55186 84204
rect 57054 84192 57060 84204
rect 57112 84192 57118 84244
rect 547230 84192 547236 84244
rect 547288 84232 547294 84244
rect 550082 84232 550088 84244
rect 547288 84204 550088 84232
rect 547288 84192 547294 84204
rect 550082 84192 550088 84204
rect 550140 84192 550146 84244
rect 57146 84124 57152 84176
rect 57204 84164 57210 84176
rect 58250 84164 58256 84176
rect 57204 84136 58256 84164
rect 57204 84124 57210 84136
rect 58250 84124 58256 84136
rect 58308 84124 58314 84176
rect 57790 83920 57796 83972
rect 57848 83920 57854 83972
rect 57808 83768 57836 83920
rect 57790 83716 57796 83768
rect 57848 83716 57854 83768
rect 54662 83648 54668 83700
rect 54720 83688 54726 83700
rect 57698 83688 57704 83700
rect 54720 83660 57704 83688
rect 54720 83648 54726 83660
rect 57698 83648 57704 83660
rect 57756 83648 57762 83700
rect 548794 83444 548800 83496
rect 548852 83484 548858 83496
rect 561122 83484 561128 83496
rect 548852 83456 561128 83484
rect 548852 83444 548858 83456
rect 561122 83444 561128 83456
rect 561180 83444 561186 83496
rect 543458 82968 543464 83020
rect 543516 83008 543522 83020
rect 547966 83008 547972 83020
rect 543516 82980 547972 83008
rect 543516 82968 543522 82980
rect 547966 82968 547972 82980
rect 548024 82968 548030 83020
rect 543642 82900 543648 82952
rect 543700 82940 543706 82952
rect 546126 82940 546132 82952
rect 543700 82912 546132 82940
rect 543700 82900 543706 82912
rect 546126 82900 546132 82912
rect 546184 82900 546190 82952
rect 541434 82832 541440 82884
rect 541492 82872 541498 82884
rect 542446 82872 542452 82884
rect 541492 82844 542452 82872
rect 541492 82832 541498 82844
rect 542446 82832 542452 82844
rect 542504 82832 542510 82884
rect 542814 82832 542820 82884
rect 542872 82872 542878 82884
rect 544470 82872 544476 82884
rect 542872 82844 544476 82872
rect 542872 82832 542878 82844
rect 544470 82832 544476 82844
rect 544528 82832 544534 82884
rect 547414 82832 547420 82884
rect 547472 82872 547478 82884
rect 548886 82872 548892 82884
rect 547472 82844 548892 82872
rect 547472 82832 547478 82844
rect 548886 82832 548892 82844
rect 548944 82832 548950 82884
rect 17862 82764 17868 82816
rect 17920 82804 17926 82816
rect 57606 82804 57612 82816
rect 17920 82776 57612 82804
rect 17920 82764 17926 82776
rect 57606 82764 57612 82776
rect 57664 82764 57670 82816
rect 543550 82764 543556 82816
rect 543608 82804 543614 82816
rect 567746 82804 567752 82816
rect 543608 82776 567752 82804
rect 543608 82764 543614 82776
rect 567746 82764 567752 82776
rect 567804 82764 567810 82816
rect 47670 82696 47676 82748
rect 47728 82736 47734 82748
rect 57514 82736 57520 82748
rect 47728 82708 57520 82736
rect 47728 82696 47734 82708
rect 57514 82696 57520 82708
rect 57572 82696 57578 82748
rect 542078 82560 542084 82612
rect 542136 82600 542142 82612
rect 543826 82600 543832 82612
rect 542136 82572 543832 82600
rect 542136 82560 542142 82572
rect 543826 82560 543832 82572
rect 543884 82560 543890 82612
rect 544930 82152 544936 82204
rect 544988 82192 544994 82204
rect 547874 82192 547880 82204
rect 544988 82164 547880 82192
rect 544988 82152 544994 82164
rect 547874 82152 547880 82164
rect 547932 82152 547938 82204
rect 540606 82084 540612 82136
rect 540664 82124 540670 82136
rect 548242 82124 548248 82136
rect 540664 82096 548248 82124
rect 540664 82084 540670 82096
rect 548242 82084 548248 82096
rect 548300 82084 548306 82136
rect 552750 80044 552756 80096
rect 552808 80084 552814 80096
rect 555510 80084 555516 80096
rect 552808 80056 555516 80084
rect 552808 80044 552814 80056
rect 555510 80044 555516 80056
rect 555568 80044 555574 80096
rect 57882 79364 57888 79416
rect 57940 79404 57946 79416
rect 59630 79404 59636 79416
rect 57940 79376 59636 79404
rect 57940 79364 57946 79376
rect 59630 79364 59636 79376
rect 59688 79364 59694 79416
rect 57698 79296 57704 79348
rect 57756 79336 57762 79348
rect 57974 79336 57980 79348
rect 57756 79308 57980 79336
rect 57756 79296 57762 79308
rect 57974 79296 57980 79308
rect 58032 79296 58038 79348
rect 543550 78616 543556 78668
rect 543608 78656 543614 78668
rect 551278 78656 551284 78668
rect 543608 78628 551284 78656
rect 543608 78616 543614 78628
rect 551278 78616 551284 78628
rect 551336 78616 551342 78668
rect 543550 77188 543556 77240
rect 543608 77228 543614 77240
rect 580350 77228 580356 77240
rect 543608 77200 580356 77228
rect 543608 77188 543614 77200
rect 580350 77188 580356 77200
rect 580408 77188 580414 77240
rect 551278 76236 551284 76288
rect 551336 76276 551342 76288
rect 556890 76276 556896 76288
rect 551336 76248 556896 76276
rect 551336 76236 551342 76248
rect 556890 76236 556896 76248
rect 556948 76236 556954 76288
rect 51902 75828 51908 75880
rect 51960 75868 51966 75880
rect 57606 75868 57612 75880
rect 51960 75840 57612 75868
rect 51960 75828 51966 75840
rect 57606 75828 57612 75840
rect 57664 75828 57670 75880
rect 543550 75828 543556 75880
rect 543608 75868 543614 75880
rect 571886 75868 571892 75880
rect 543608 75840 571892 75868
rect 543608 75828 543614 75840
rect 571886 75828 571892 75840
rect 571944 75828 571950 75880
rect 55766 75760 55772 75812
rect 55824 75800 55830 75812
rect 57146 75800 57152 75812
rect 55824 75772 57152 75800
rect 55824 75760 55830 75772
rect 57146 75760 57152 75772
rect 57204 75760 57210 75812
rect 542630 75692 542636 75744
rect 542688 75732 542694 75744
rect 545850 75732 545856 75744
rect 542688 75704 545856 75732
rect 542688 75692 542694 75704
rect 545850 75692 545856 75704
rect 545908 75692 545914 75744
rect 57606 75556 57612 75608
rect 57664 75596 57670 75608
rect 57882 75596 57888 75608
rect 57664 75568 57888 75596
rect 57664 75556 57670 75568
rect 57882 75556 57888 75568
rect 57940 75556 57946 75608
rect 540514 75148 540520 75200
rect 540572 75188 540578 75200
rect 547874 75188 547880 75200
rect 540572 75160 547880 75188
rect 540572 75148 540578 75160
rect 547874 75148 547880 75160
rect 547932 75148 547938 75200
rect 574738 73108 574744 73160
rect 574796 73148 574802 73160
rect 580350 73148 580356 73160
rect 574796 73120 580356 73148
rect 574796 73108 574802 73120
rect 580350 73108 580356 73120
rect 580408 73108 580414 73160
rect 543550 71680 543556 71732
rect 543608 71720 543614 71732
rect 582650 71720 582656 71732
rect 543608 71692 582656 71720
rect 543608 71680 543614 71692
rect 582650 71680 582656 71692
rect 582708 71680 582714 71732
rect 547322 71612 547328 71664
rect 547380 71652 547386 71664
rect 550082 71652 550088 71664
rect 547380 71624 550088 71652
rect 547380 71612 547386 71624
rect 550082 71612 550088 71624
rect 550140 71612 550146 71664
rect 546494 71408 546500 71460
rect 546552 71448 546558 71460
rect 549254 71448 549260 71460
rect 546552 71420 549260 71448
rect 546552 71408 546558 71420
rect 549254 71408 549260 71420
rect 549312 71408 549318 71460
rect 543550 70320 543556 70372
rect 543608 70360 543614 70372
rect 566550 70360 566556 70372
rect 543608 70332 566556 70360
rect 543608 70320 543614 70332
rect 566550 70320 566556 70332
rect 566608 70320 566614 70372
rect 42610 69640 42616 69692
rect 42668 69680 42674 69692
rect 57054 69680 57060 69692
rect 42668 69652 57060 69680
rect 42668 69640 42674 69652
rect 57054 69640 57060 69652
rect 57112 69640 57118 69692
rect 542262 69232 542268 69284
rect 542320 69272 542326 69284
rect 543366 69272 543372 69284
rect 542320 69244 543372 69272
rect 542320 69232 542326 69244
rect 543366 69232 543372 69244
rect 543424 69232 543430 69284
rect 38286 68960 38292 69012
rect 38344 69000 38350 69012
rect 57882 69000 57888 69012
rect 38344 68972 57888 69000
rect 38344 68960 38350 68972
rect 57882 68960 57888 68972
rect 57940 68960 57946 69012
rect 39022 68892 39028 68944
rect 39080 68932 39086 68944
rect 57146 68932 57152 68944
rect 39080 68904 57152 68932
rect 39080 68892 39086 68904
rect 57146 68892 57152 68904
rect 57204 68892 57210 68944
rect 53282 68824 53288 68876
rect 53340 68864 53346 68876
rect 55950 68864 55956 68876
rect 53340 68836 55956 68864
rect 53340 68824 53346 68836
rect 55950 68824 55956 68836
rect 56008 68824 56014 68876
rect 40770 67532 40776 67584
rect 40828 67572 40834 67584
rect 57882 67572 57888 67584
rect 40828 67544 57888 67572
rect 40828 67532 40834 67544
rect 57882 67532 57888 67544
rect 57940 67532 57946 67584
rect 544562 67328 544568 67380
rect 544620 67368 544626 67380
rect 546494 67368 546500 67380
rect 544620 67340 546500 67368
rect 544620 67328 544626 67340
rect 546494 67328 546500 67340
rect 546552 67328 546558 67380
rect 542814 66172 542820 66224
rect 542872 66212 542878 66224
rect 582742 66212 582748 66224
rect 542872 66184 582748 66212
rect 542872 66172 542878 66184
rect 582742 66172 582748 66184
rect 582800 66172 582806 66224
rect 543550 66104 543556 66156
rect 543608 66144 543614 66156
rect 578326 66144 578332 66156
rect 543608 66116 578332 66144
rect 543608 66104 543614 66116
rect 578326 66104 578332 66116
rect 578384 66104 578390 66156
rect 543642 66036 543648 66088
rect 543700 66076 543706 66088
rect 547046 66076 547052 66088
rect 543700 66048 547052 66076
rect 543700 66036 543706 66048
rect 547046 66036 547052 66048
rect 547104 66036 547110 66088
rect 33778 64812 33784 64864
rect 33836 64852 33842 64864
rect 57882 64852 57888 64864
rect 33836 64824 57888 64852
rect 33836 64812 33842 64824
rect 57882 64812 57888 64824
rect 57940 64812 57946 64864
rect 543550 63928 543556 63980
rect 543608 63968 543614 63980
rect 549622 63968 549628 63980
rect 543608 63940 549628 63968
rect 543608 63928 543614 63940
rect 549622 63928 549628 63940
rect 549680 63928 549686 63980
rect 49050 63452 49056 63504
rect 49108 63492 49114 63504
rect 57882 63492 57888 63504
rect 49108 63464 57888 63492
rect 49108 63452 49114 63464
rect 57882 63452 57888 63464
rect 57940 63452 57946 63504
rect 548886 63316 548892 63368
rect 548944 63356 548950 63368
rect 549622 63356 549628 63368
rect 548944 63328 549628 63356
rect 548944 63316 548950 63328
rect 549622 63316 549628 63328
rect 549680 63316 549686 63368
rect 42702 62024 42708 62076
rect 42760 62064 42766 62076
rect 57882 62064 57888 62076
rect 42760 62036 57888 62064
rect 42760 62024 42766 62036
rect 57882 62024 57888 62036
rect 57940 62024 57946 62076
rect 543550 62024 543556 62076
rect 543608 62064 543614 62076
rect 560938 62064 560944 62076
rect 543608 62036 560944 62064
rect 543608 62024 543614 62036
rect 560938 62024 560944 62036
rect 560996 62024 561002 62076
rect 543642 61956 543648 62008
rect 543700 61996 543706 62008
rect 551094 61996 551100 62008
rect 543700 61968 551100 61996
rect 543700 61956 543706 61968
rect 551094 61956 551100 61968
rect 551152 61956 551158 62008
rect 571978 60664 571984 60716
rect 572036 60704 572042 60716
rect 580350 60704 580356 60716
rect 572036 60676 580356 60704
rect 572036 60664 572042 60676
rect 580350 60664 580356 60676
rect 580408 60664 580414 60716
rect 45002 59984 45008 60036
rect 45060 60024 45066 60036
rect 57054 60024 57060 60036
rect 45060 59996 57060 60024
rect 45060 59984 45066 59996
rect 57054 59984 57060 59996
rect 57112 59984 57118 60036
rect 24670 59304 24676 59356
rect 24728 59344 24734 59356
rect 57882 59344 57888 59356
rect 24728 59316 57888 59344
rect 24728 59304 24734 59316
rect 57882 59304 57888 59316
rect 57940 59304 57946 59356
rect 40402 57876 40408 57928
rect 40460 57916 40466 57928
rect 57882 57916 57888 57928
rect 40460 57888 57888 57916
rect 40460 57876 40466 57888
rect 57882 57876 57888 57888
rect 57940 57876 57946 57928
rect 543550 57876 543556 57928
rect 543608 57916 543614 57928
rect 572898 57916 572904 57928
rect 543608 57888 572904 57916
rect 543608 57876 543614 57888
rect 572898 57876 572904 57888
rect 572956 57876 572962 57928
rect 46014 56516 46020 56568
rect 46072 56556 46078 56568
rect 57882 56556 57888 56568
rect 46072 56528 57888 56556
rect 46072 56516 46078 56528
rect 57882 56516 57888 56528
rect 57940 56516 57946 56568
rect 543550 55836 543556 55888
rect 543608 55876 543614 55888
rect 562042 55876 562048 55888
rect 543608 55848 562048 55876
rect 543608 55836 543614 55848
rect 562042 55836 562048 55848
rect 562100 55836 562106 55888
rect 542722 53728 542728 53780
rect 542780 53768 542786 53780
rect 580258 53768 580264 53780
rect 542780 53740 580264 53768
rect 542780 53728 542786 53740
rect 580258 53728 580264 53740
rect 580316 53728 580322 53780
rect 542722 51008 542728 51060
rect 542780 51048 542786 51060
rect 551002 51048 551008 51060
rect 542780 51020 551008 51048
rect 542780 51008 542786 51020
rect 551002 51008 551008 51020
rect 551060 51008 551066 51060
rect 542722 49648 542728 49700
rect 542780 49688 542786 49700
rect 552474 49688 552480 49700
rect 542780 49660 552480 49688
rect 542780 49648 542786 49660
rect 552474 49648 552480 49660
rect 552532 49648 552538 49700
rect 47210 48968 47216 49020
rect 47268 49008 47274 49020
rect 57882 49008 57888 49020
rect 47268 48980 57888 49008
rect 47268 48968 47274 48980
rect 57882 48968 57888 48980
rect 57940 48968 57946 49020
rect 543642 48220 543648 48272
rect 543700 48260 543706 48272
rect 577130 48260 577136 48272
rect 543700 48232 577136 48260
rect 543700 48220 543706 48232
rect 577130 48220 577136 48232
rect 577188 48220 577194 48272
rect 543642 45500 543648 45552
rect 543700 45540 543706 45552
rect 582558 45540 582564 45552
rect 543700 45512 582564 45540
rect 543700 45500 543706 45512
rect 582558 45500 582564 45512
rect 582616 45500 582622 45552
rect 55582 45296 55588 45348
rect 55640 45336 55646 45348
rect 57146 45336 57152 45348
rect 55640 45308 57152 45336
rect 55640 45296 55646 45308
rect 57146 45296 57152 45308
rect 57204 45296 57210 45348
rect 543642 42780 543648 42832
rect 543700 42820 543706 42832
rect 547046 42820 547052 42832
rect 543700 42792 547052 42820
rect 543700 42780 543706 42792
rect 547046 42780 547052 42792
rect 547104 42780 547110 42832
rect 24762 41352 24768 41404
rect 24820 41392 24826 41404
rect 57882 41392 57888 41404
rect 24820 41364 57888 41392
rect 24820 41352 24826 41364
rect 57882 41352 57888 41364
rect 57940 41352 57946 41404
rect 543550 41352 543556 41404
rect 543608 41392 543614 41404
rect 557810 41392 557816 41404
rect 543608 41364 557816 41392
rect 543608 41352 543614 41364
rect 557810 41352 557816 41364
rect 557868 41352 557874 41404
rect 49326 41284 49332 41336
rect 49384 41324 49390 41336
rect 56686 41324 56692 41336
rect 49384 41296 56692 41324
rect 49384 41284 49390 41296
rect 56686 41284 56692 41296
rect 56744 41284 56750 41336
rect 543550 37204 543556 37256
rect 543608 37244 543614 37256
rect 560662 37244 560668 37256
rect 543608 37216 560668 37244
rect 543608 37204 543614 37216
rect 560662 37204 560668 37216
rect 560720 37204 560726 37256
rect 543642 35844 543648 35896
rect 543700 35884 543706 35896
rect 560570 35884 560576 35896
rect 543700 35856 560576 35884
rect 543700 35844 543706 35856
rect 560570 35844 560576 35856
rect 560628 35844 560634 35896
rect 25958 34416 25964 34468
rect 26016 34456 26022 34468
rect 57882 34456 57888 34468
rect 26016 34428 57888 34456
rect 26016 34416 26022 34428
rect 57882 34416 57888 34428
rect 57940 34416 57946 34468
rect 570690 33056 570696 33108
rect 570748 33096 570754 33108
rect 580258 33096 580264 33108
rect 570748 33068 580264 33096
rect 570748 33056 570754 33068
rect 580258 33056 580264 33068
rect 580316 33056 580322 33108
rect 36538 32988 36544 33040
rect 36596 33028 36602 33040
rect 57882 33028 57888 33040
rect 36596 33000 57888 33028
rect 36596 32988 36602 33000
rect 57882 32988 57888 33000
rect 57940 32988 57946 33040
rect 540698 31016 540704 31068
rect 540756 31056 540762 31068
rect 578602 31056 578608 31068
rect 540756 31028 578608 31056
rect 540756 31016 540762 31028
rect 578602 31016 578608 31028
rect 578660 31016 578666 31068
rect 156046 29860 156052 29912
rect 156104 29900 156110 29912
rect 157258 29900 157264 29912
rect 156104 29872 157264 29900
rect 156104 29860 156110 29872
rect 157258 29860 157264 29872
rect 157316 29860 157322 29912
rect 340874 29860 340880 29912
rect 340932 29900 340938 29912
rect 342086 29900 342092 29912
rect 340932 29872 342092 29900
rect 340932 29860 340938 29872
rect 342086 29860 342092 29872
rect 342144 29860 342150 29912
rect 361574 29860 361580 29912
rect 361632 29900 361638 29912
rect 362694 29900 362700 29912
rect 361632 29872 362700 29900
rect 361632 29860 361638 29872
rect 362694 29860 362700 29872
rect 362752 29860 362758 29912
rect 378134 29860 378140 29912
rect 378192 29900 378198 29912
rect 379438 29900 379444 29912
rect 378192 29872 379444 29900
rect 378192 29860 378198 29872
rect 379438 29860 379444 29872
rect 379496 29860 379502 29912
rect 458174 29860 458180 29912
rect 458232 29900 458238 29912
rect 459294 29900 459300 29912
rect 458232 29872 459300 29900
rect 458232 29860 458238 29872
rect 459294 29860 459300 29872
rect 459352 29860 459358 29912
rect 525794 29860 525800 29912
rect 525852 29900 525858 29912
rect 526914 29900 526920 29912
rect 525852 29872 526920 29900
rect 525852 29860 525858 29872
rect 526914 29860 526920 29872
rect 526972 29860 526978 29912
rect 521102 29724 521108 29776
rect 521160 29764 521166 29776
rect 521160 29736 528554 29764
rect 521160 29724 521166 29736
rect 54202 29656 54208 29708
rect 54260 29696 54266 29708
rect 63494 29696 63500 29708
rect 54260 29668 63500 29696
rect 54260 29656 54266 29668
rect 63494 29656 63500 29668
rect 63552 29656 63558 29708
rect 45186 29588 45192 29640
rect 45244 29628 45250 29640
rect 69014 29628 69020 29640
rect 45244 29600 69020 29628
rect 45244 29588 45250 29600
rect 69014 29588 69020 29600
rect 69072 29588 69078 29640
rect 528526 29628 528554 29736
rect 552198 29628 552204 29640
rect 528526 29600 552204 29628
rect 552198 29588 552204 29600
rect 552256 29588 552262 29640
rect 378042 29520 378048 29572
rect 378100 29560 378106 29572
rect 378226 29560 378232 29572
rect 378100 29532 378232 29560
rect 378100 29520 378106 29532
rect 378226 29520 378232 29532
rect 378284 29520 378290 29572
rect 523034 29520 523040 29572
rect 523092 29560 523098 29572
rect 566090 29560 566096 29572
rect 523092 29532 566096 29560
rect 523092 29520 523098 29532
rect 566090 29520 566096 29532
rect 566148 29520 566154 29572
rect 43162 29452 43168 29504
rect 43220 29492 43226 29504
rect 69658 29492 69664 29504
rect 43220 29464 69664 29492
rect 43220 29452 43226 29464
rect 69658 29452 69664 29464
rect 69716 29452 69722 29504
rect 476666 29452 476672 29504
rect 476724 29492 476730 29504
rect 525886 29492 525892 29504
rect 476724 29464 525892 29492
rect 476724 29452 476730 29464
rect 525886 29452 525892 29464
rect 525944 29452 525950 29504
rect 528186 29452 528192 29504
rect 528244 29492 528250 29504
rect 552382 29492 552388 29504
rect 528244 29464 552388 29492
rect 528244 29452 528250 29464
rect 552382 29452 552388 29464
rect 552440 29452 552446 29504
rect 43898 29384 43904 29436
rect 43956 29424 43962 29436
rect 123754 29424 123760 29436
rect 43956 29396 123760 29424
rect 43956 29384 43962 29396
rect 123754 29384 123760 29396
rect 123812 29384 123818 29436
rect 481818 29384 481824 29436
rect 481876 29424 481882 29436
rect 565262 29424 565268 29436
rect 481876 29396 565268 29424
rect 481876 29384 481882 29396
rect 565262 29384 565268 29396
rect 565320 29384 565326 29436
rect 47302 29316 47308 29368
rect 47360 29356 47366 29368
rect 199746 29356 199752 29368
rect 47360 29328 199752 29356
rect 47360 29316 47366 29328
rect 199746 29316 199752 29328
rect 199804 29316 199810 29368
rect 409690 29316 409696 29368
rect 409748 29356 409754 29368
rect 554130 29356 554136 29368
rect 409748 29328 554136 29356
rect 409748 29316 409754 29328
rect 554130 29316 554136 29328
rect 554188 29316 554194 29368
rect 42518 29248 42524 29300
rect 42576 29288 42582 29300
rect 195238 29288 195244 29300
rect 42576 29260 195244 29288
rect 42576 29248 42582 29260
rect 195238 29248 195244 29260
rect 195296 29248 195302 29300
rect 384574 29248 384580 29300
rect 384632 29288 384638 29300
rect 550266 29288 550272 29300
rect 384632 29260 550272 29288
rect 384632 29248 384638 29260
rect 550266 29248 550272 29260
rect 550324 29248 550330 29300
rect 39298 29180 39304 29232
rect 39356 29220 39362 29232
rect 193306 29220 193312 29232
rect 39356 29192 193312 29220
rect 39356 29180 39362 29192
rect 193306 29180 193312 29192
rect 193364 29180 193370 29232
rect 356882 29180 356888 29232
rect 356940 29220 356946 29232
rect 544746 29220 544752 29232
rect 356940 29192 544752 29220
rect 356940 29180 356946 29192
rect 544746 29180 544752 29192
rect 544804 29180 544810 29232
rect 43714 29112 43720 29164
rect 43772 29152 43778 29164
rect 205542 29152 205548 29164
rect 43772 29124 205548 29152
rect 43772 29112 43778 29124
rect 205542 29112 205548 29124
rect 205600 29112 205606 29164
rect 287330 29112 287336 29164
rect 287388 29152 287394 29164
rect 575474 29152 575480 29164
rect 287388 29124 575480 29152
rect 287388 29112 287394 29124
rect 575474 29112 575480 29124
rect 575532 29112 575538 29164
rect 39850 29044 39856 29096
rect 39908 29084 39914 29096
rect 217778 29084 217784 29096
rect 39908 29056 217784 29084
rect 39908 29044 39914 29056
rect 217778 29044 217784 29056
rect 217836 29044 217842 29096
rect 260926 29044 260932 29096
rect 260984 29084 260990 29096
rect 583018 29084 583024 29096
rect 260984 29056 583024 29084
rect 260984 29044 260990 29056
rect 583018 29044 583024 29056
rect 583076 29044 583082 29096
rect 28902 28976 28908 29028
rect 28960 29016 28966 29028
rect 159818 29016 159824 29028
rect 28960 28988 159824 29016
rect 28960 28976 28966 28988
rect 159818 28976 159824 28988
rect 159876 28976 159882 29028
rect 182358 28976 182364 29028
rect 182416 29016 182422 29028
rect 550358 29016 550364 29028
rect 182416 28988 550364 29016
rect 182416 28976 182422 28988
rect 550358 28976 550364 28988
rect 550416 28976 550422 29028
rect 47486 28908 47492 28960
rect 47544 28948 47550 28960
rect 325970 28948 325976 28960
rect 47544 28920 325976 28948
rect 47544 28908 47550 28920
rect 325970 28908 325976 28920
rect 326028 28908 326034 28960
rect 536558 28908 536564 28960
rect 536616 28948 536622 28960
rect 552106 28948 552112 28960
rect 536616 28920 552112 28948
rect 536616 28908 536622 28920
rect 552106 28908 552112 28920
rect 552164 28908 552170 28960
rect 52270 28840 52276 28892
rect 52328 28880 52334 28892
rect 67726 28880 67732 28892
rect 52328 28852 67732 28880
rect 52328 28840 52334 28852
rect 67726 28840 67732 28852
rect 67784 28840 67790 28892
rect 271230 28840 271236 28892
rect 271288 28880 271294 28892
rect 527818 28880 527824 28892
rect 271288 28852 527824 28880
rect 271288 28840 271294 28852
rect 527818 28840 527824 28852
rect 527876 28840 527882 28892
rect 537202 28840 537208 28892
rect 537260 28880 537266 28892
rect 550910 28880 550916 28892
rect 537260 28852 550916 28880
rect 537260 28840 537266 28852
rect 550910 28840 550916 28852
rect 550968 28840 550974 28892
rect 49510 28772 49516 28824
rect 49568 28812 49574 28824
rect 63218 28812 63224 28824
rect 49568 28784 63224 28812
rect 49568 28772 49574 28784
rect 63218 28772 63224 28784
rect 63276 28772 63282 28824
rect 295702 28772 295708 28824
rect 295760 28812 295766 28824
rect 473998 28812 474004 28824
rect 295760 28784 474004 28812
rect 295760 28772 295766 28784
rect 473998 28772 474004 28784
rect 474056 28772 474062 28824
rect 512086 28772 512092 28824
rect 512144 28812 512150 28824
rect 583478 28812 583484 28824
rect 512144 28784 583484 28812
rect 512144 28772 512150 28784
rect 583478 28772 583484 28784
rect 583536 28772 583542 28824
rect 50706 28704 50712 28756
rect 50764 28744 50770 28756
rect 62574 28744 62580 28756
rect 50764 28716 62580 28744
rect 50764 28704 50770 28716
rect 62574 28704 62580 28716
rect 62632 28704 62638 28756
rect 170858 28704 170864 28756
rect 170916 28744 170922 28756
rect 249978 28744 249984 28756
rect 170916 28716 249984 28744
rect 170916 28704 170922 28716
rect 249978 28704 249984 28716
rect 250036 28704 250042 28756
rect 338206 28704 338212 28756
rect 338264 28744 338270 28756
rect 524874 28744 524880 28756
rect 338264 28716 524880 28744
rect 338264 28704 338270 28716
rect 524874 28704 524880 28716
rect 524932 28704 524938 28756
rect 525886 28704 525892 28756
rect 525944 28744 525950 28756
rect 581086 28744 581092 28756
rect 525944 28716 581092 28744
rect 525944 28704 525950 28716
rect 581086 28704 581092 28716
rect 581144 28704 581150 28756
rect 19242 28636 19248 28688
rect 19300 28676 19306 28688
rect 82538 28676 82544 28688
rect 19300 28648 82544 28676
rect 19300 28636 19306 28648
rect 82538 28636 82544 28648
rect 82596 28636 82602 28688
rect 83458 28636 83464 28688
rect 83516 28676 83522 28688
rect 190730 28676 190736 28688
rect 83516 28648 190736 28676
rect 83516 28636 83522 28648
rect 190730 28636 190736 28648
rect 190788 28636 190794 28688
rect 443178 28636 443184 28688
rect 443236 28676 443242 28688
rect 563146 28676 563152 28688
rect 443236 28648 563152 28676
rect 443236 28636 443242 28648
rect 563146 28636 563152 28648
rect 563204 28636 563210 28688
rect 35342 28568 35348 28620
rect 35400 28608 35406 28620
rect 103790 28608 103796 28620
rect 35400 28580 103796 28608
rect 35400 28568 35406 28580
rect 103790 28568 103796 28580
rect 103848 28568 103854 28620
rect 143166 28568 143172 28620
rect 143224 28608 143230 28620
rect 251266 28608 251272 28620
rect 143224 28580 251272 28608
rect 143224 28568 143230 28580
rect 251266 28568 251272 28580
rect 251324 28568 251330 28620
rect 311158 28568 311164 28620
rect 311216 28608 311222 28620
rect 529934 28608 529940 28620
rect 311216 28580 529940 28608
rect 311216 28568 311222 28580
rect 529934 28568 529940 28580
rect 529992 28568 529998 28620
rect 532050 28568 532056 28620
rect 532108 28608 532114 28620
rect 581178 28608 581184 28620
rect 532108 28580 581184 28608
rect 532108 28568 532114 28580
rect 581178 28568 581184 28580
rect 581236 28568 581242 28620
rect 35802 28500 35808 28552
rect 35860 28540 35866 28552
rect 73522 28540 73528 28552
rect 35860 28512 73528 28540
rect 35860 28500 35866 28512
rect 73522 28500 73528 28512
rect 73580 28500 73586 28552
rect 78766 28500 78772 28552
rect 78824 28540 78830 28552
rect 188798 28540 188804 28552
rect 78824 28512 188804 28540
rect 78824 28500 78830 28512
rect 188798 28500 188804 28512
rect 188856 28500 188862 28552
rect 258994 28500 259000 28552
rect 259052 28540 259058 28552
rect 505738 28540 505744 28552
rect 259052 28512 505744 28540
rect 259052 28500 259058 28512
rect 505738 28500 505744 28512
rect 505796 28500 505802 28552
rect 506934 28500 506940 28552
rect 506992 28540 506998 28552
rect 565998 28540 566004 28552
rect 506992 28512 566004 28540
rect 506992 28500 506998 28512
rect 565998 28500 566004 28512
rect 566056 28500 566062 28552
rect 33594 28432 33600 28484
rect 33652 28472 33658 28484
rect 71590 28472 71596 28484
rect 33652 28444 71596 28472
rect 33652 28432 33658 28444
rect 71590 28432 71596 28444
rect 71648 28432 71654 28484
rect 72418 28432 72424 28484
rect 72476 28472 72482 28484
rect 141786 28472 141792 28484
rect 72476 28444 141792 28472
rect 72476 28432 72482 28444
rect 141786 28432 141792 28444
rect 141844 28432 141850 28484
rect 147674 28432 147680 28484
rect 147732 28472 147738 28484
rect 148870 28472 148876 28484
rect 147732 28444 148876 28472
rect 147732 28432 147738 28444
rect 148870 28432 148876 28444
rect 148928 28432 148934 28484
rect 157978 28432 157984 28484
rect 158036 28472 158042 28484
rect 272518 28472 272524 28484
rect 158036 28444 272524 28472
rect 158036 28432 158042 28444
rect 272518 28432 272524 28444
rect 272576 28432 272582 28484
rect 291838 28432 291844 28484
rect 291896 28472 291902 28484
rect 535454 28472 535460 28484
rect 291896 28444 535460 28472
rect 291896 28432 291902 28444
rect 535454 28432 535460 28444
rect 535512 28432 535518 28484
rect 29730 28364 29736 28416
rect 29788 28404 29794 28416
rect 92198 28404 92204 28416
rect 29788 28376 92204 28404
rect 29788 28364 29794 28376
rect 92198 28364 92204 28376
rect 92256 28364 92262 28416
rect 96798 28364 96804 28416
rect 96856 28404 96862 28416
rect 211338 28404 211344 28416
rect 96856 28376 211344 28404
rect 96856 28364 96862 28376
rect 211338 28364 211344 28376
rect 211396 28364 211402 28416
rect 505646 28364 505652 28416
rect 505704 28404 505710 28416
rect 574462 28404 574468 28416
rect 505704 28376 574468 28404
rect 505704 28364 505710 28376
rect 574462 28364 574468 28376
rect 574520 28364 574526 28416
rect 50890 28296 50896 28348
rect 50948 28336 50954 28348
rect 95418 28336 95424 28348
rect 50948 28308 95424 28336
rect 50948 28296 50954 28308
rect 95418 28296 95424 28308
rect 95476 28296 95482 28348
rect 130194 28296 130200 28348
rect 130252 28336 130258 28348
rect 252554 28336 252560 28348
rect 130252 28308 252560 28336
rect 130252 28296 130258 28308
rect 252554 28296 252560 28308
rect 252612 28296 252618 28348
rect 268010 28296 268016 28348
rect 268068 28336 268074 28348
rect 517514 28336 517520 28348
rect 268068 28308 517520 28336
rect 268068 28296 268074 28308
rect 517514 28296 517520 28308
rect 517572 28296 517578 28348
rect 529474 28296 529480 28348
rect 529532 28336 529538 28348
rect 575934 28336 575940 28348
rect 529532 28308 575940 28336
rect 529532 28296 529538 28308
rect 575934 28296 575940 28308
rect 575992 28296 575998 28348
rect 69934 28228 69940 28280
rect 69992 28268 69998 28280
rect 213270 28268 213276 28280
rect 69992 28240 213276 28268
rect 69992 28228 69998 28240
rect 213270 28228 213276 28240
rect 213328 28228 213334 28280
rect 266078 28228 266084 28280
rect 266136 28268 266142 28280
rect 451918 28268 451924 28280
rect 266136 28240 451924 28268
rect 266136 28228 266142 28240
rect 451918 28228 451924 28240
rect 451976 28228 451982 28280
rect 463694 28228 463700 28280
rect 463752 28268 463758 28280
rect 464430 28268 464436 28280
rect 463752 28240 464436 28268
rect 463752 28228 463758 28240
rect 464430 28228 464436 28240
rect 464488 28228 464494 28280
rect 476114 28228 476120 28280
rect 476172 28268 476178 28280
rect 477310 28268 477316 28280
rect 476172 28240 477316 28268
rect 476172 28228 476178 28240
rect 477310 28228 477316 28240
rect 477368 28228 477374 28280
rect 484486 28228 484492 28280
rect 484544 28268 484550 28280
rect 485682 28268 485688 28280
rect 484544 28240 485688 28268
rect 484544 28228 484550 28240
rect 485682 28228 485688 28240
rect 485740 28228 485746 28280
rect 505094 28228 505100 28280
rect 505152 28268 505158 28280
rect 506290 28268 506296 28280
rect 505152 28240 506296 28268
rect 505152 28228 505158 28240
rect 506290 28228 506296 28240
rect 506348 28228 506354 28280
rect 519170 28228 519176 28280
rect 519228 28268 519234 28280
rect 562594 28268 562600 28280
rect 519228 28240 562600 28268
rect 519228 28228 519234 28240
rect 562594 28228 562600 28240
rect 562652 28228 562658 28280
rect 40678 28160 40684 28212
rect 40736 28200 40742 28212
rect 72878 28200 72884 28212
rect 40736 28172 72884 28200
rect 40736 28160 40742 28172
rect 72878 28160 72884 28172
rect 72936 28160 72942 28212
rect 74534 28160 74540 28212
rect 74592 28200 74598 28212
rect 181070 28200 181076 28212
rect 74592 28172 181076 28200
rect 74592 28160 74598 28172
rect 181070 28160 181076 28172
rect 181128 28160 181134 28212
rect 186314 28160 186320 28212
rect 186372 28200 186378 28212
rect 187510 28200 187516 28212
rect 186372 28172 187516 28200
rect 186372 28160 186378 28172
rect 187510 28160 187516 28172
rect 187568 28160 187574 28212
rect 191834 28160 191840 28212
rect 191892 28200 191898 28212
rect 192662 28200 192668 28212
rect 191892 28172 192668 28200
rect 191892 28160 191898 28172
rect 192662 28160 192668 28172
rect 192720 28160 192726 28212
rect 215294 28160 215300 28212
rect 215352 28200 215358 28212
rect 216490 28200 216496 28212
rect 215352 28172 216496 28200
rect 215352 28160 215358 28172
rect 216490 28160 216496 28172
rect 216548 28160 216554 28212
rect 320174 28160 320180 28212
rect 320232 28200 320238 28212
rect 321462 28200 321468 28212
rect 320232 28172 321468 28200
rect 320232 28160 320238 28172
rect 321462 28160 321468 28172
rect 321520 28160 321526 28212
rect 321554 28160 321560 28212
rect 321612 28200 321618 28212
rect 322750 28200 322756 28212
rect 321612 28172 322756 28200
rect 321612 28160 321618 28172
rect 322750 28160 322756 28172
rect 322808 28160 322814 28212
rect 324314 28160 324320 28212
rect 324372 28200 324378 28212
rect 325326 28200 325332 28212
rect 324372 28172 325332 28200
rect 324372 28160 324378 28172
rect 325326 28160 325332 28172
rect 325384 28160 325390 28212
rect 329834 28160 329840 28212
rect 329892 28200 329898 28212
rect 331122 28200 331128 28212
rect 329892 28172 331128 28200
rect 329892 28160 329898 28172
rect 331122 28160 331128 28172
rect 331180 28160 331186 28212
rect 347774 28160 347780 28212
rect 347832 28200 347838 28212
rect 348510 28200 348516 28212
rect 347832 28172 348516 28200
rect 347832 28160 347838 28172
rect 348510 28160 348516 28172
rect 348568 28160 348574 28212
rect 354674 28160 354680 28212
rect 354732 28200 354738 28212
rect 355594 28200 355600 28212
rect 354732 28172 355600 28200
rect 354732 28160 354738 28172
rect 355594 28160 355600 28172
rect 355652 28160 355658 28212
rect 358814 28160 358820 28212
rect 358872 28200 358878 28212
rect 360102 28200 360108 28212
rect 358872 28172 360108 28200
rect 358872 28160 358878 28172
rect 360102 28160 360108 28172
rect 360160 28160 360166 28212
rect 367094 28160 367100 28212
rect 367152 28200 367158 28212
rect 367830 28200 367836 28212
rect 367152 28172 367836 28200
rect 367152 28160 367158 28172
rect 367830 28160 367836 28172
rect 367888 28160 367894 28212
rect 368474 28160 368480 28212
rect 368532 28200 368538 28212
rect 369762 28200 369768 28212
rect 368532 28172 369768 28200
rect 368532 28160 368538 28172
rect 369762 28160 369768 28172
rect 369820 28160 369826 28212
rect 389082 28160 389088 28212
rect 389140 28200 389146 28212
rect 536098 28200 536104 28212
rect 389140 28172 536104 28200
rect 389140 28160 389146 28172
rect 536098 28160 536104 28172
rect 536156 28160 536162 28212
rect 66346 28092 66352 28144
rect 66404 28132 66410 28144
rect 168190 28132 168196 28144
rect 66404 28104 168196 28132
rect 66404 28092 66410 28104
rect 168190 28092 168196 28104
rect 168248 28092 168254 28144
rect 300854 28092 300860 28144
rect 300912 28132 300918 28144
rect 302142 28132 302148 28144
rect 300912 28104 302148 28132
rect 300912 28092 300918 28104
rect 302142 28092 302148 28104
rect 302200 28092 302206 28144
rect 417418 28092 417424 28144
rect 417476 28132 417482 28144
rect 544838 28132 544844 28144
rect 417476 28104 544844 28132
rect 417476 28092 417482 28104
rect 544838 28092 544844 28104
rect 544896 28092 544902 28144
rect 63494 28024 63500 28076
rect 63552 28064 63558 28076
rect 63552 28036 84194 28064
rect 63552 28024 63558 28036
rect 84166 27996 84194 28036
rect 97994 28024 98000 28076
rect 98052 28064 98058 28076
rect 99282 28064 99288 28076
rect 98052 28036 99288 28064
rect 98052 28024 98058 28036
rect 99282 28024 99288 28036
rect 99340 28024 99346 28076
rect 99374 28024 99380 28076
rect 99432 28064 99438 28076
rect 100570 28064 100576 28076
rect 99432 28036 100576 28064
rect 99432 28024 99438 28036
rect 100570 28024 100576 28036
rect 100628 28024 100634 28076
rect 107746 28024 107752 28076
rect 107804 28064 107810 28076
rect 108942 28064 108948 28076
rect 107804 28036 108948 28064
rect 107804 28024 107810 28036
rect 108942 28024 108948 28036
rect 109000 28024 109006 28076
rect 109034 28024 109040 28076
rect 109092 28064 109098 28076
rect 201678 28064 201684 28076
rect 109092 28036 201684 28064
rect 109092 28024 109098 28036
rect 201678 28024 201684 28036
rect 201736 28024 201742 28076
rect 426434 28024 426440 28076
rect 426492 28064 426498 28076
rect 427722 28064 427728 28076
rect 426492 28036 427728 28064
rect 426492 28024 426498 28036
rect 427722 28024 427728 28036
rect 427780 28024 427786 28076
rect 427814 28024 427820 28076
rect 427872 28064 427878 28076
rect 429010 28064 429016 28076
rect 427872 28036 429016 28064
rect 427872 28024 427878 28036
rect 429010 28024 429016 28036
rect 429068 28024 429074 28076
rect 436094 28024 436100 28076
rect 436152 28064 436158 28076
rect 437382 28064 437388 28076
rect 436152 28036 437388 28064
rect 436152 28024 436158 28036
rect 437382 28024 437388 28036
rect 437440 28024 437446 28076
rect 445754 28024 445760 28076
rect 445812 28064 445818 28076
rect 447042 28064 447048 28076
rect 445812 28036 447048 28064
rect 445812 28024 445818 28036
rect 447042 28024 447048 28036
rect 447100 28024 447106 28076
rect 447134 28024 447140 28076
rect 447192 28064 447198 28076
rect 448330 28064 448336 28076
rect 447192 28036 448336 28064
rect 447192 28024 447198 28036
rect 448330 28024 448336 28036
rect 448388 28024 448394 28076
rect 448514 28024 448520 28076
rect 448572 28064 448578 28076
rect 449618 28064 449624 28076
rect 448572 28036 449624 28064
rect 448572 28024 448578 28036
rect 449618 28024 449624 28036
rect 449676 28024 449682 28076
rect 465074 28024 465080 28076
rect 465132 28064 465138 28076
rect 466362 28064 466368 28076
rect 465132 28036 466368 28064
rect 465132 28024 465138 28036
rect 466362 28024 466368 28036
rect 466420 28024 466426 28076
rect 484394 28024 484400 28076
rect 484452 28064 484458 28076
rect 485038 28064 485044 28076
rect 484452 28036 485044 28064
rect 484452 28024 484458 28036
rect 485038 28024 485044 28036
rect 485096 28024 485102 28076
rect 502426 28024 502432 28076
rect 502484 28064 502490 28076
rect 503070 28064 503076 28076
rect 502484 28036 503076 28064
rect 502484 28024 502490 28036
rect 503070 28024 503076 28036
rect 503128 28024 503134 28076
rect 503162 28024 503168 28076
rect 503220 28064 503226 28076
rect 569402 28064 569408 28076
rect 503220 28036 569408 28064
rect 503220 28024 503226 28036
rect 569402 28024 569408 28036
rect 569460 28024 569466 28076
rect 103146 27996 103152 28008
rect 84166 27968 103152 27996
rect 103146 27956 103152 27968
rect 103204 27956 103210 28008
rect 104158 27956 104164 28008
rect 104216 27996 104222 28008
rect 195882 27996 195888 28008
rect 104216 27968 195888 27996
rect 104216 27956 104222 27968
rect 195882 27956 195888 27968
rect 195940 27956 195946 28008
rect 327258 27956 327264 28008
rect 327316 27996 327322 28008
rect 562134 27996 562140 28008
rect 327316 27968 562140 27996
rect 327316 27956 327322 27968
rect 562134 27956 562140 27968
rect 562192 27956 562198 28008
rect 92566 27888 92572 27940
rect 92624 27928 92630 27940
rect 179782 27928 179788 27940
rect 92624 27900 179788 27928
rect 92624 27888 92630 27900
rect 179782 27888 179788 27900
rect 179840 27888 179846 27940
rect 344002 27888 344008 27940
rect 344060 27928 344066 27940
rect 563238 27928 563244 27940
rect 344060 27900 563244 27928
rect 344060 27888 344066 27900
rect 563238 27888 563244 27900
rect 563296 27888 563302 27940
rect 39574 27820 39580 27872
rect 39632 27860 39638 27872
rect 166902 27860 166908 27872
rect 39632 27832 166908 27860
rect 39632 27820 39638 27832
rect 166902 27820 166908 27832
rect 166960 27820 166966 27872
rect 275738 27820 275744 27872
rect 275796 27860 275802 27872
rect 510706 27860 510712 27872
rect 275796 27832 510712 27860
rect 275796 27820 275802 27832
rect 510706 27820 510712 27832
rect 510764 27820 510770 27872
rect 37642 27752 37648 27804
rect 37700 27792 37706 27804
rect 155954 27792 155960 27804
rect 37700 27764 155960 27792
rect 37700 27752 37706 27764
rect 155954 27752 155960 27764
rect 156012 27752 156018 27804
rect 18874 27684 18880 27736
rect 18932 27724 18938 27736
rect 128906 27724 128912 27736
rect 18932 27696 128912 27724
rect 18932 27684 18938 27696
rect 128906 27684 128912 27696
rect 128964 27684 128970 27736
rect 103514 27616 103520 27668
rect 103572 27656 103578 27668
rect 109034 27656 109040 27668
rect 103572 27628 109040 27656
rect 103572 27616 103578 27628
rect 109034 27616 109040 27628
rect 109092 27616 109098 27668
rect 170398 27616 170404 27668
rect 170456 27656 170462 27668
rect 170858 27656 170864 27668
rect 170456 27628 170864 27656
rect 170456 27616 170462 27628
rect 170858 27616 170864 27628
rect 170916 27616 170922 27668
rect 502334 27616 502340 27668
rect 502392 27656 502398 27668
rect 503162 27656 503168 27668
rect 502392 27628 503168 27656
rect 502392 27616 502398 27628
rect 503162 27616 503168 27628
rect 503220 27616 503226 27668
rect 35526 27548 35532 27600
rect 35584 27588 35590 27600
rect 70946 27588 70952 27600
rect 35584 27560 70952 27588
rect 35584 27548 35590 27560
rect 70946 27548 70952 27560
rect 71004 27548 71010 27600
rect 531406 27548 531412 27600
rect 531464 27588 531470 27600
rect 560478 27588 560484 27600
rect 531464 27560 560484 27588
rect 531464 27548 531470 27560
rect 560478 27548 560484 27560
rect 560536 27548 560542 27600
rect 50798 27480 50804 27532
rect 50856 27520 50862 27532
rect 70302 27520 70308 27532
rect 50856 27492 70308 27520
rect 50856 27480 50862 27492
rect 70302 27480 70308 27492
rect 70360 27480 70366 27532
rect 157334 27480 157340 27532
rect 157392 27520 157398 27532
rect 158530 27520 158536 27532
rect 157392 27492 158536 27520
rect 157392 27480 157398 27492
rect 158530 27480 158536 27492
rect 158588 27480 158594 27532
rect 493410 27480 493416 27532
rect 493468 27520 493474 27532
rect 570414 27520 570420 27532
rect 493468 27492 570420 27520
rect 493468 27480 493474 27492
rect 570414 27480 570420 27492
rect 570472 27480 570478 27532
rect 44266 27412 44272 27464
rect 44324 27452 44330 27464
rect 89622 27452 89628 27464
rect 44324 27424 89628 27452
rect 44324 27412 44330 27424
rect 89622 27412 89628 27424
rect 89680 27412 89686 27464
rect 535454 27412 535460 27464
rect 535512 27452 535518 27464
rect 563606 27452 563612 27464
rect 535512 27424 563612 27452
rect 535512 27412 535518 27424
rect 563606 27412 563612 27424
rect 563664 27412 563670 27464
rect 29914 27344 29920 27396
rect 29972 27384 29978 27396
rect 470870 27384 470876 27396
rect 29972 27356 470876 27384
rect 29972 27344 29978 27356
rect 470870 27344 470876 27356
rect 470928 27344 470934 27396
rect 510154 27344 510160 27396
rect 510212 27384 510218 27396
rect 573450 27384 573456 27396
rect 510212 27356 573456 27384
rect 510212 27344 510218 27356
rect 573450 27344 573456 27356
rect 573508 27344 573514 27396
rect 52546 27276 52552 27328
rect 52604 27316 52610 27328
rect 441246 27316 441252 27328
rect 52604 27288 441252 27316
rect 52604 27276 52610 27288
rect 441246 27276 441252 27288
rect 441304 27276 441310 27328
rect 491478 27276 491484 27328
rect 491536 27316 491542 27328
rect 553486 27316 553492 27328
rect 491536 27288 553492 27316
rect 491536 27276 491542 27288
rect 553486 27276 553492 27288
rect 553544 27276 553550 27328
rect 42426 27208 42432 27260
rect 42484 27248 42490 27260
rect 385218 27248 385224 27260
rect 42484 27220 385224 27248
rect 42484 27208 42490 27220
rect 385218 27208 385224 27220
rect 385276 27208 385282 27260
rect 398742 27208 398748 27260
rect 398800 27248 398806 27260
rect 583110 27248 583116 27260
rect 398800 27220 583116 27248
rect 398800 27208 398806 27220
rect 583110 27208 583116 27220
rect 583168 27208 583174 27260
rect 32766 27140 32772 27192
rect 32824 27180 32830 27192
rect 363966 27180 363972 27192
rect 32824 27152 363972 27180
rect 32824 27140 32830 27152
rect 363966 27140 363972 27152
rect 364024 27140 364030 27192
rect 381354 27140 381360 27192
rect 381412 27180 381418 27192
rect 561766 27180 561772 27192
rect 381412 27152 561772 27180
rect 381412 27140 381418 27152
rect 561766 27140 561772 27152
rect 561824 27140 561830 27192
rect 24394 27072 24400 27124
rect 24452 27112 24458 27124
rect 266722 27112 266728 27124
rect 24452 27084 266728 27112
rect 24452 27072 24458 27084
rect 266722 27072 266728 27084
rect 266780 27072 266786 27124
rect 268654 27072 268660 27124
rect 268712 27112 268718 27124
rect 577498 27112 577504 27124
rect 268712 27084 577504 27112
rect 268712 27072 268718 27084
rect 577498 27072 577504 27084
rect 577556 27072 577562 27124
rect 49142 27004 49148 27056
rect 49200 27044 49206 27056
rect 296990 27044 296996 27056
rect 49200 27016 296996 27044
rect 49200 27004 49206 27016
rect 296990 27004 296996 27016
rect 297048 27004 297054 27056
rect 410334 27004 410340 27056
rect 410392 27044 410398 27056
rect 576026 27044 576032 27056
rect 410392 27016 576032 27044
rect 410392 27004 410398 27016
rect 576026 27004 576032 27016
rect 576084 27004 576090 27056
rect 31110 26936 31116 26988
rect 31168 26976 31174 26988
rect 109586 26976 109592 26988
rect 31168 26948 109592 26976
rect 31168 26936 31174 26948
rect 109586 26936 109592 26948
rect 109644 26936 109650 26988
rect 390370 26936 390376 26988
rect 390428 26976 390434 26988
rect 540422 26976 540428 26988
rect 390428 26948 540428 26976
rect 390428 26936 390434 26948
rect 540422 26936 540428 26948
rect 540480 26936 540486 26988
rect 41046 26868 41052 26920
rect 41104 26908 41110 26920
rect 92474 26908 92480 26920
rect 41104 26880 92480 26908
rect 41104 26868 41110 26880
rect 92474 26868 92480 26880
rect 92532 26868 92538 26920
rect 515950 26868 515956 26920
rect 516008 26908 516014 26920
rect 549070 26908 549076 26920
rect 516008 26880 549076 26908
rect 516008 26868 516014 26880
rect 549070 26868 549076 26880
rect 549128 26868 549134 26920
rect 58618 26800 58624 26852
rect 58676 26840 58682 26852
rect 87690 26840 87696 26852
rect 58676 26812 87696 26840
rect 58676 26800 58682 26812
rect 87690 26800 87696 26812
rect 87748 26800 87754 26852
rect 514018 26800 514024 26852
rect 514076 26840 514082 26852
rect 549162 26840 549168 26852
rect 514076 26812 549168 26840
rect 514076 26800 514082 26812
rect 549162 26800 549168 26812
rect 549220 26800 549226 26852
rect 41874 26732 41880 26784
rect 41932 26772 41938 26784
rect 523678 26772 523684 26784
rect 41932 26744 523684 26772
rect 41932 26732 41938 26744
rect 523678 26732 523684 26744
rect 523736 26732 523742 26784
rect 69658 26664 69664 26716
rect 69716 26704 69722 26716
rect 520458 26704 520464 26716
rect 69716 26676 520464 26704
rect 69716 26664 69722 26676
rect 520458 26664 520464 26676
rect 520516 26664 520522 26716
rect 36998 26596 37004 26648
rect 37056 26636 37062 26648
rect 494054 26636 494060 26648
rect 37056 26608 494060 26636
rect 37056 26596 37062 26608
rect 494054 26596 494060 26608
rect 494112 26596 494118 26648
rect 516594 26596 516600 26648
rect 516652 26636 516658 26648
rect 549530 26636 549536 26648
rect 516652 26608 549536 26636
rect 516652 26596 516658 26608
rect 549530 26596 549536 26608
rect 549588 26596 549594 26648
rect 18966 26188 18972 26240
rect 19024 26228 19030 26240
rect 391934 26228 391940 26240
rect 19024 26200 391940 26228
rect 19024 26188 19030 26200
rect 391934 26188 391940 26200
rect 391992 26188 391998 26240
rect 536098 26188 536104 26240
rect 536156 26228 536162 26240
rect 547506 26228 547512 26240
rect 536156 26200 547512 26228
rect 536156 26188 536162 26200
rect 547506 26188 547512 26200
rect 547564 26188 547570 26240
rect 49234 26120 49240 26172
rect 49292 26160 49298 26172
rect 368474 26160 368480 26172
rect 49292 26132 368480 26160
rect 49292 26120 49298 26132
rect 368474 26120 368480 26132
rect 368532 26120 368538 26172
rect 492674 26120 492680 26172
rect 492732 26160 492738 26172
rect 560846 26160 560852 26172
rect 492732 26132 560852 26160
rect 492732 26120 492738 26132
rect 560846 26120 560852 26132
rect 560904 26120 560910 26172
rect 20622 26052 20628 26104
rect 20680 26092 20686 26104
rect 318794 26092 318800 26104
rect 20680 26064 318800 26092
rect 20680 26052 20686 26064
rect 318794 26052 318800 26064
rect 318852 26052 318858 26104
rect 322934 26052 322940 26104
rect 322992 26092 322998 26104
rect 578510 26092 578516 26104
rect 322992 26064 578516 26092
rect 322992 26052 322998 26064
rect 578510 26052 578516 26064
rect 578568 26052 578574 26104
rect 28718 25984 28724 26036
rect 28776 26024 28782 26036
rect 307754 26024 307760 26036
rect 28776 25996 307760 26024
rect 28776 25984 28782 25996
rect 307754 25984 307760 25996
rect 307812 25984 307818 26036
rect 325786 25984 325792 26036
rect 325844 26024 325850 26036
rect 578418 26024 578424 26036
rect 325844 25996 578424 26024
rect 325844 25984 325850 25996
rect 578418 25984 578424 25996
rect 578476 25984 578482 26036
rect 27338 25916 27344 25968
rect 27396 25956 27402 25968
rect 306374 25956 306380 25968
rect 27396 25928 306380 25956
rect 27396 25916 27402 25928
rect 306374 25916 306380 25928
rect 306432 25916 306438 25968
rect 520274 25916 520280 25968
rect 520332 25956 520338 25968
rect 571518 25956 571524 25968
rect 520332 25928 571524 25956
rect 520332 25916 520338 25928
rect 571518 25916 571524 25928
rect 571576 25916 571582 25968
rect 51994 25848 52000 25900
rect 52052 25888 52058 25900
rect 292574 25888 292580 25900
rect 52052 25860 292580 25888
rect 52052 25848 52058 25860
rect 292574 25848 292580 25860
rect 292632 25848 292638 25900
rect 513374 25848 513380 25900
rect 513432 25888 513438 25900
rect 567286 25888 567292 25900
rect 513432 25860 567292 25888
rect 513432 25848 513438 25860
rect 567286 25848 567292 25860
rect 567344 25848 567350 25900
rect 58710 25780 58716 25832
rect 58768 25820 58774 25832
rect 216674 25820 216680 25832
rect 58768 25792 216680 25820
rect 58768 25780 58774 25792
rect 216674 25780 216680 25792
rect 216732 25780 216738 25832
rect 516134 25780 516140 25832
rect 516192 25820 516198 25832
rect 571702 25820 571708 25832
rect 516192 25792 571708 25820
rect 516192 25780 516198 25792
rect 571702 25780 571708 25792
rect 571760 25780 571766 25832
rect 30742 25712 30748 25764
rect 30800 25752 30806 25764
rect 186314 25752 186320 25764
rect 30800 25724 186320 25752
rect 30800 25712 30806 25724
rect 186314 25712 186320 25724
rect 186372 25712 186378 25764
rect 396074 25712 396080 25764
rect 396132 25752 396138 25764
rect 545666 25752 545672 25764
rect 396132 25724 545672 25752
rect 396132 25712 396138 25724
rect 545666 25712 545672 25724
rect 545724 25712 545730 25764
rect 29822 25644 29828 25696
rect 29880 25684 29886 25696
rect 165706 25684 165712 25696
rect 29880 25656 165712 25684
rect 29880 25644 29886 25656
rect 165706 25644 165712 25656
rect 165764 25644 165770 25696
rect 416774 25644 416780 25696
rect 416832 25684 416838 25696
rect 575842 25684 575848 25696
rect 416832 25656 575848 25684
rect 416832 25644 416838 25656
rect 575842 25644 575848 25656
rect 575900 25644 575906 25696
rect 52822 25576 52828 25628
rect 52880 25616 52886 25628
rect 77294 25616 77300 25628
rect 52880 25588 77300 25616
rect 52880 25576 52886 25588
rect 77294 25576 77300 25588
rect 77352 25576 77358 25628
rect 342346 25576 342352 25628
rect 342404 25616 342410 25628
rect 573174 25616 573180 25628
rect 342404 25588 573180 25616
rect 342404 25576 342410 25588
rect 573174 25576 573180 25588
rect 573232 25576 573238 25628
rect 54846 25508 54852 25560
rect 54904 25548 54910 25560
rect 81434 25548 81440 25560
rect 54904 25520 81440 25548
rect 54904 25508 54910 25520
rect 81434 25508 81440 25520
rect 81492 25508 81498 25560
rect 321738 25508 321744 25560
rect 321796 25548 321802 25560
rect 563790 25548 563796 25560
rect 321796 25520 563796 25548
rect 321796 25508 321802 25520
rect 563790 25508 563796 25520
rect 563848 25508 563854 25560
rect 54938 25440 54944 25492
rect 54996 25480 55002 25492
rect 67634 25480 67640 25492
rect 54996 25452 67640 25480
rect 54996 25440 55002 25452
rect 67634 25440 67640 25452
rect 67692 25440 67698 25492
rect 502518 25440 502524 25492
rect 502576 25480 502582 25492
rect 546218 25480 546224 25492
rect 502576 25452 546224 25480
rect 502576 25440 502582 25452
rect 546218 25440 546224 25452
rect 546276 25440 546282 25492
rect 538214 25372 538220 25424
rect 538272 25412 538278 25424
rect 555694 25412 555700 25424
rect 538272 25384 555700 25412
rect 538272 25372 538278 25384
rect 555694 25372 555700 25384
rect 555752 25372 555758 25424
rect 461026 25304 461032 25356
rect 461084 25344 461090 25356
rect 540698 25344 540704 25356
rect 461084 25316 540704 25344
rect 461084 25304 461090 25316
rect 540698 25304 540704 25316
rect 540756 25304 540762 25356
rect 314654 24896 314660 24948
rect 314712 24936 314718 24948
rect 479058 24936 479064 24948
rect 314712 24908 479064 24936
rect 314712 24896 314718 24908
rect 479058 24896 479064 24908
rect 479116 24896 479122 24948
rect 53650 24828 53656 24880
rect 53708 24868 53714 24880
rect 85574 24868 85580 24880
rect 53708 24840 85580 24868
rect 53708 24828 53714 24840
rect 85574 24828 85580 24840
rect 85632 24828 85638 24880
rect 231854 24828 231860 24880
rect 231912 24868 231918 24880
rect 485038 24868 485044 24880
rect 231912 24840 485044 24868
rect 231912 24828 231918 24840
rect 485038 24828 485044 24840
rect 485096 24828 485102 24880
rect 32306 24760 32312 24812
rect 32364 24800 32370 24812
rect 444466 24800 444472 24812
rect 32364 24772 444472 24800
rect 32364 24760 32370 24772
rect 444466 24760 444472 24772
rect 444524 24760 444530 24812
rect 476114 24760 476120 24812
rect 476172 24800 476178 24812
rect 552290 24800 552296 24812
rect 476172 24772 552296 24800
rect 476172 24760 476178 24772
rect 552290 24760 552296 24772
rect 552348 24760 552354 24812
rect 50614 24692 50620 24744
rect 50672 24732 50678 24744
rect 397454 24732 397460 24744
rect 50672 24704 397460 24732
rect 50672 24692 50678 24704
rect 397454 24692 397460 24704
rect 397512 24692 397518 24744
rect 436094 24692 436100 24744
rect 436152 24732 436158 24744
rect 569218 24732 569224 24744
rect 436152 24704 569224 24732
rect 436152 24692 436158 24704
rect 569218 24692 569224 24704
rect 569276 24692 569282 24744
rect 26050 24624 26056 24676
rect 26108 24664 26114 24676
rect 354766 24664 354772 24676
rect 26108 24636 354772 24664
rect 26108 24624 26114 24636
rect 354766 24624 354772 24636
rect 354824 24624 354830 24676
rect 476022 24624 476028 24676
rect 476080 24664 476086 24676
rect 549990 24664 549996 24676
rect 476080 24636 549996 24664
rect 476080 24624 476086 24636
rect 549990 24624 549996 24636
rect 550048 24624 550054 24676
rect 21818 24556 21824 24608
rect 21876 24596 21882 24608
rect 333974 24596 333980 24608
rect 21876 24568 333980 24596
rect 21876 24556 21882 24568
rect 333974 24556 333980 24568
rect 334032 24556 334038 24608
rect 477494 24556 477500 24608
rect 477552 24596 477558 24608
rect 539962 24596 539968 24608
rect 477552 24568 539968 24596
rect 477552 24556 477558 24568
rect 539962 24556 539968 24568
rect 540020 24556 540026 24608
rect 31202 24488 31208 24540
rect 31260 24528 31266 24540
rect 256694 24528 256700 24540
rect 31260 24500 256700 24528
rect 31260 24488 31266 24500
rect 256694 24488 256700 24500
rect 256752 24488 256758 24540
rect 280154 24488 280160 24540
rect 280212 24528 280218 24540
rect 574370 24528 574376 24540
rect 280212 24500 574376 24528
rect 280212 24488 280218 24500
rect 574370 24488 574376 24500
rect 574428 24488 574434 24540
rect 21542 24420 21548 24472
rect 21600 24460 21606 24472
rect 311894 24460 311900 24472
rect 21600 24432 311900 24460
rect 21600 24420 21606 24432
rect 311894 24420 311900 24432
rect 311952 24420 311958 24472
rect 470594 24420 470600 24472
rect 470652 24460 470658 24472
rect 557626 24460 557632 24472
rect 470652 24432 557632 24460
rect 470652 24420 470658 24432
rect 557626 24420 557632 24432
rect 557684 24420 557690 24472
rect 38102 24352 38108 24404
rect 38160 24392 38166 24404
rect 204254 24392 204260 24404
rect 38160 24364 204260 24392
rect 38160 24352 38166 24364
rect 204254 24352 204260 24364
rect 204312 24352 204318 24404
rect 332594 24352 332600 24404
rect 332652 24392 332658 24404
rect 556338 24392 556344 24404
rect 332652 24364 556344 24392
rect 332652 24352 332658 24364
rect 556338 24352 556344 24364
rect 556396 24352 556402 24404
rect 50522 24284 50528 24336
rect 50580 24324 50586 24336
rect 191926 24324 191932 24336
rect 50580 24296 191932 24324
rect 50580 24284 50586 24296
rect 191926 24284 191932 24296
rect 191984 24284 191990 24336
rect 245654 24284 245660 24336
rect 245712 24324 245718 24336
rect 563698 24324 563704 24336
rect 245712 24296 563704 24324
rect 245712 24284 245718 24296
rect 563698 24284 563704 24296
rect 563756 24284 563762 24336
rect 41230 24216 41236 24268
rect 41288 24256 41294 24268
rect 182174 24256 182180 24268
rect 41288 24228 182180 24256
rect 41288 24216 41294 24228
rect 182174 24216 182180 24228
rect 182232 24216 182238 24268
rect 224954 24216 224960 24268
rect 225012 24256 225018 24268
rect 571426 24256 571432 24268
rect 225012 24228 571432 24256
rect 225012 24216 225018 24228
rect 571426 24216 571432 24228
rect 571484 24216 571490 24268
rect 25590 24148 25596 24200
rect 25648 24188 25654 24200
rect 131206 24188 131212 24200
rect 25648 24160 131212 24188
rect 25648 24148 25654 24160
rect 131206 24148 131212 24160
rect 131264 24148 131270 24200
rect 220814 24148 220820 24200
rect 220872 24188 220878 24200
rect 568666 24188 568672 24200
rect 220872 24160 568672 24188
rect 220872 24148 220878 24160
rect 568666 24148 568672 24160
rect 568724 24148 568730 24200
rect 21726 24080 21732 24132
rect 21784 24120 21790 24132
rect 124214 24120 124220 24132
rect 21784 24092 124220 24120
rect 21784 24080 21790 24092
rect 124214 24080 124220 24092
rect 124272 24080 124278 24132
rect 209866 24080 209872 24132
rect 209924 24120 209930 24132
rect 564710 24120 564716 24132
rect 209924 24092 564716 24120
rect 209924 24080 209930 24092
rect 564710 24080 564716 24092
rect 564768 24080 564774 24132
rect 52730 24012 52736 24064
rect 52788 24052 52794 24064
rect 142154 24052 142160 24064
rect 52788 24024 142160 24052
rect 52788 24012 52794 24024
rect 142154 24012 142160 24024
rect 142212 24012 142218 24064
rect 498194 24012 498200 24064
rect 498252 24052 498258 24064
rect 559834 24052 559840 24064
rect 498252 24024 559840 24052
rect 498252 24012 498258 24024
rect 559834 24012 559840 24024
rect 559892 24012 559898 24064
rect 42978 23944 42984 23996
rect 43036 23984 43042 23996
rect 99374 23984 99380 23996
rect 43036 23956 99380 23984
rect 43036 23944 43042 23956
rect 99374 23944 99380 23956
rect 99432 23944 99438 23996
rect 502426 23944 502432 23996
rect 502484 23984 502490 23996
rect 551462 23984 551468 23996
rect 502484 23956 551468 23984
rect 502484 23944 502490 23956
rect 551462 23944 551468 23956
rect 551520 23944 551526 23996
rect 51442 23876 51448 23928
rect 51500 23916 51506 23928
rect 98086 23916 98092 23928
rect 51500 23888 98092 23916
rect 51500 23876 51506 23888
rect 98086 23876 98092 23888
rect 98144 23876 98150 23928
rect 34146 23400 34152 23452
rect 34204 23440 34210 23452
rect 104894 23440 104900 23452
rect 34204 23412 104900 23440
rect 34204 23400 34210 23412
rect 104894 23400 104900 23412
rect 104952 23400 104958 23452
rect 517514 23400 517520 23452
rect 517572 23440 517578 23452
rect 540606 23440 540612 23452
rect 517572 23412 540612 23440
rect 517572 23400 517578 23412
rect 540606 23400 540612 23412
rect 540664 23400 540670 23452
rect 46658 23332 46664 23384
rect 46716 23372 46722 23384
rect 131114 23372 131120 23384
rect 46716 23344 131120 23372
rect 46716 23332 46722 23344
rect 131114 23332 131120 23344
rect 131172 23332 131178 23384
rect 184934 23332 184940 23384
rect 184992 23372 184998 23384
rect 581638 23372 581644 23384
rect 184992 23344 581644 23372
rect 184992 23332 184998 23344
rect 581638 23332 581644 23344
rect 581696 23332 581702 23384
rect 52914 23264 52920 23316
rect 52972 23304 52978 23316
rect 128446 23304 128452 23316
rect 52972 23276 128452 23304
rect 52972 23264 52978 23276
rect 128446 23264 128452 23276
rect 128504 23264 128510 23316
rect 529934 23264 529940 23316
rect 529992 23304 529998 23316
rect 562318 23304 562324 23316
rect 529992 23276 562324 23304
rect 529992 23264 529998 23276
rect 562318 23264 562324 23276
rect 562376 23264 562382 23316
rect 354674 23196 354680 23248
rect 354732 23236 354738 23248
rect 579614 23236 579620 23248
rect 354732 23208 579620 23236
rect 354732 23196 354738 23208
rect 579614 23196 579620 23208
rect 579672 23196 579678 23248
rect 21634 23128 21640 23180
rect 21692 23168 21698 23180
rect 342254 23168 342260 23180
rect 21692 23140 342260 23168
rect 21692 23128 21698 23140
rect 342254 23128 342260 23140
rect 342312 23128 342318 23180
rect 365714 23128 365720 23180
rect 365772 23168 365778 23180
rect 579798 23168 579804 23180
rect 365772 23140 579804 23168
rect 365772 23128 365778 23140
rect 579798 23128 579804 23140
rect 579856 23128 579862 23180
rect 36262 23060 36268 23112
rect 36320 23100 36326 23112
rect 321554 23100 321560 23112
rect 36320 23072 321560 23100
rect 36320 23060 36326 23072
rect 321554 23060 321560 23072
rect 321612 23060 321618 23112
rect 409966 23060 409972 23112
rect 410024 23100 410030 23112
rect 555326 23100 555332 23112
rect 410024 23072 555332 23100
rect 410024 23060 410030 23072
rect 555326 23060 555332 23072
rect 555384 23060 555390 23112
rect 24578 22992 24584 23044
rect 24636 23032 24642 23044
rect 285674 23032 285680 23044
rect 24636 23004 285680 23032
rect 24636 22992 24642 23004
rect 285674 22992 285680 23004
rect 285732 22992 285738 23044
rect 451274 22992 451280 23044
rect 451332 23032 451338 23044
rect 582926 23032 582932 23044
rect 451332 23004 582932 23032
rect 451332 22992 451338 23004
rect 582926 22992 582932 23004
rect 582984 22992 582990 23044
rect 45094 22924 45100 22976
rect 45152 22964 45158 22976
rect 303614 22964 303620 22976
rect 45152 22936 303620 22964
rect 45152 22924 45158 22936
rect 303614 22924 303620 22936
rect 303672 22924 303678 22976
rect 449894 22924 449900 22976
rect 449952 22964 449958 22976
rect 555418 22964 555424 22976
rect 449952 22936 555424 22964
rect 449952 22924 449958 22936
rect 555418 22924 555424 22936
rect 555476 22924 555482 22976
rect 23382 22856 23388 22908
rect 23440 22896 23446 22908
rect 270494 22896 270500 22908
rect 23440 22868 270500 22896
rect 23440 22856 23446 22868
rect 270494 22856 270500 22868
rect 270552 22856 270558 22908
rect 385034 22856 385040 22908
rect 385092 22896 385098 22908
rect 558546 22896 558552 22908
rect 385092 22868 558552 22896
rect 385092 22856 385098 22868
rect 558546 22856 558552 22868
rect 558604 22856 558610 22908
rect 22002 22788 22008 22840
rect 22060 22828 22066 22840
rect 72326 22828 72332 22840
rect 22060 22800 72332 22828
rect 22060 22788 22066 22800
rect 72326 22788 72332 22800
rect 72384 22788 72390 22840
rect 171134 22788 171140 22840
rect 171192 22828 171198 22840
rect 416682 22828 416688 22840
rect 171192 22800 416688 22828
rect 171192 22788 171198 22800
rect 416682 22788 416688 22800
rect 416740 22788 416746 22840
rect 456794 22788 456800 22840
rect 456852 22828 456858 22840
rect 556706 22828 556712 22840
rect 456852 22800 556712 22828
rect 456852 22788 456858 22800
rect 556706 22788 556712 22800
rect 556764 22788 556770 22840
rect 49418 22720 49424 22772
rect 49476 22760 49482 22772
rect 110414 22760 110420 22772
rect 49476 22732 110420 22760
rect 49476 22720 49482 22732
rect 110414 22720 110420 22732
rect 110472 22720 110478 22772
rect 168374 22720 168380 22772
rect 168432 22760 168438 22772
rect 553854 22760 553860 22772
rect 168432 22732 553860 22760
rect 168432 22720 168438 22732
rect 553854 22720 553860 22732
rect 553912 22720 553918 22772
rect 43990 22652 43996 22704
rect 44048 22692 44054 22704
rect 215294 22692 215300 22704
rect 44048 22664 215300 22692
rect 44048 22652 44054 22664
rect 215294 22652 215300 22664
rect 215352 22652 215358 22704
rect 465258 22652 465264 22704
rect 465316 22692 465322 22704
rect 554038 22692 554044 22704
rect 465316 22664 554044 22692
rect 465316 22652 465322 22664
rect 554038 22652 554044 22664
rect 554096 22652 554102 22704
rect 44082 22584 44088 22636
rect 44140 22624 44146 22636
rect 66346 22624 66352 22636
rect 44140 22596 66352 22624
rect 44140 22584 44146 22596
rect 66346 22584 66352 22596
rect 66404 22584 66410 22636
rect 107746 22584 107752 22636
rect 107804 22624 107810 22636
rect 554958 22624 554964 22636
rect 107804 22596 554964 22624
rect 107804 22584 107810 22596
rect 554958 22584 554964 22596
rect 555016 22584 555022 22636
rect 45370 22516 45376 22568
rect 45428 22556 45434 22568
rect 72418 22556 72424 22568
rect 45428 22528 72424 22556
rect 45428 22516 45434 22528
rect 72418 22516 72424 22528
rect 72476 22516 72482 22568
rect 160094 22516 160100 22568
rect 160152 22556 160158 22568
rect 548978 22556 548984 22568
rect 160152 22528 548984 22556
rect 160152 22516 160158 22528
rect 548978 22516 548984 22528
rect 549036 22516 549042 22568
rect 32674 22448 32680 22500
rect 32732 22488 32738 22500
rect 356054 22488 356060 22500
rect 32732 22460 356060 22488
rect 32732 22448 32738 22460
rect 356054 22448 356060 22460
rect 356112 22448 356118 22500
rect 58526 22040 58532 22092
rect 58584 22080 58590 22092
rect 78766 22080 78772 22092
rect 58584 22052 78772 22080
rect 58584 22040 58590 22052
rect 78766 22040 78772 22052
rect 78824 22040 78830 22092
rect 488534 22040 488540 22092
rect 488592 22080 488598 22092
rect 551554 22080 551560 22092
rect 488592 22052 551560 22080
rect 488592 22040 488598 22052
rect 551554 22040 551560 22052
rect 551612 22040 551618 22092
rect 47946 21972 47952 22024
rect 48004 22012 48010 22024
rect 411254 22012 411260 22024
rect 48004 21984 411260 22012
rect 48004 21972 48010 21984
rect 411254 21972 411260 21984
rect 411312 21972 411318 22024
rect 483014 21972 483020 22024
rect 483072 22012 483078 22024
rect 544378 22012 544384 22024
rect 483072 21984 544384 22012
rect 483072 21972 483078 21984
rect 544378 21972 544384 21984
rect 544436 21972 544442 22024
rect 54478 21904 54484 21956
rect 54536 21944 54542 21956
rect 400214 21944 400220 21956
rect 54536 21916 400220 21944
rect 54536 21904 54542 21916
rect 400214 21904 400220 21916
rect 400272 21904 400278 21956
rect 528554 21904 528560 21956
rect 528612 21944 528618 21956
rect 570598 21944 570604 21956
rect 528612 21916 570604 21944
rect 528612 21904 528618 21916
rect 570598 21904 570604 21916
rect 570656 21904 570662 21956
rect 52086 21836 52092 21888
rect 52144 21876 52150 21888
rect 209774 21876 209780 21888
rect 52144 21848 209780 21876
rect 52144 21836 52150 21848
rect 209774 21836 209780 21848
rect 209832 21836 209838 21888
rect 223574 21836 223580 21888
rect 223632 21876 223638 21888
rect 548610 21876 548616 21888
rect 223632 21848 548616 21876
rect 223632 21836 223638 21848
rect 548610 21836 548616 21848
rect 548668 21836 548674 21888
rect 51718 21768 51724 21820
rect 51776 21808 51782 21820
rect 364334 21808 364340 21820
rect 51776 21780 364340 21808
rect 51776 21768 51782 21780
rect 364334 21768 364340 21780
rect 364392 21768 364398 21820
rect 385126 21768 385132 21820
rect 385184 21808 385190 21820
rect 552658 21808 552664 21820
rect 385184 21780 552664 21808
rect 385184 21768 385190 21780
rect 552658 21768 552664 21780
rect 552716 21768 552722 21820
rect 46290 21700 46296 21752
rect 46348 21740 46354 21752
rect 255314 21740 255320 21752
rect 46348 21712 255320 21740
rect 46348 21700 46354 21712
rect 255314 21700 255320 21712
rect 255372 21700 255378 21752
rect 420914 21700 420920 21752
rect 420972 21740 420978 21752
rect 559098 21740 559104 21752
rect 420972 21712 559104 21740
rect 420972 21700 420978 21712
rect 559098 21700 559104 21712
rect 559156 21700 559162 21752
rect 56226 21632 56232 21684
rect 56284 21672 56290 21684
rect 197354 21672 197360 21684
rect 56284 21644 197360 21672
rect 56284 21632 56290 21644
rect 197354 21632 197360 21644
rect 197412 21632 197418 21684
rect 371234 21632 371240 21684
rect 371292 21672 371298 21684
rect 553670 21672 553676 21684
rect 371292 21644 553676 21672
rect 371292 21632 371298 21644
rect 553670 21632 553676 21644
rect 553728 21632 553734 21684
rect 51350 21564 51356 21616
rect 51408 21604 51414 21616
rect 169754 21604 169760 21616
rect 51408 21576 169760 21604
rect 51408 21564 51414 21576
rect 169754 21564 169760 21576
rect 169812 21564 169818 21616
rect 258074 21564 258080 21616
rect 258132 21604 258138 21616
rect 568850 21604 568856 21616
rect 258132 21576 568856 21604
rect 258132 21564 258138 21576
rect 568850 21564 568856 21576
rect 568908 21564 568914 21616
rect 54570 21496 54576 21548
rect 54628 21536 54634 21548
rect 156046 21536 156052 21548
rect 54628 21508 156052 21536
rect 54628 21496 54634 21508
rect 156046 21496 156052 21508
rect 156104 21496 156110 21548
rect 260834 21496 260840 21548
rect 260892 21536 260898 21548
rect 572990 21536 572996 21548
rect 260892 21508 572996 21536
rect 260892 21496 260898 21508
rect 572990 21496 572996 21508
rect 573048 21496 573054 21548
rect 46566 21428 46572 21480
rect 46624 21468 46630 21480
rect 147674 21468 147680 21480
rect 46624 21440 147680 21468
rect 46624 21428 46630 21440
rect 147674 21428 147680 21440
rect 147732 21428 147738 21480
rect 176654 21428 176660 21480
rect 176712 21468 176718 21480
rect 573082 21468 573088 21480
rect 176712 21440 573088 21468
rect 176712 21428 176718 21440
rect 573082 21428 573088 21440
rect 573140 21428 573146 21480
rect 43806 21360 43812 21412
rect 43864 21400 43870 21412
rect 103514 21400 103520 21412
rect 43864 21372 103520 21400
rect 43864 21360 43870 21372
rect 103514 21360 103520 21372
rect 103572 21360 103578 21412
rect 146386 21360 146392 21412
rect 146444 21400 146450 21412
rect 569586 21400 569592 21412
rect 146444 21372 569592 21400
rect 146444 21360 146450 21372
rect 569586 21360 569592 21372
rect 569644 21360 569650 21412
rect 49602 21292 49608 21344
rect 49660 21332 49666 21344
rect 92566 21332 92572 21344
rect 49660 21304 92572 21332
rect 49660 21292 49666 21304
rect 92566 21292 92572 21304
rect 92624 21292 92630 21344
rect 510706 21292 510712 21344
rect 510764 21332 510770 21344
rect 542170 21332 542176 21344
rect 510764 21304 542176 21332
rect 510764 21292 510770 21304
rect 542170 21292 542176 21304
rect 542228 21292 542234 21344
rect 57606 21224 57612 21276
rect 57664 21264 57670 21276
rect 96798 21264 96804 21276
rect 57664 21236 96804 21264
rect 57664 21224 57670 21236
rect 96798 21224 96804 21236
rect 96856 21224 96862 21276
rect 46382 21156 46388 21208
rect 46440 21196 46446 21208
rect 427814 21196 427820 21208
rect 46440 21168 427820 21196
rect 46440 21156 46446 21168
rect 427814 21156 427820 21168
rect 427872 21156 427878 21208
rect 58894 20612 58900 20664
rect 58952 20652 58958 20664
rect 69934 20652 69940 20664
rect 58952 20624 69940 20652
rect 58952 20612 58958 20624
rect 69934 20612 69940 20624
rect 69992 20612 69998 20664
rect 503714 20612 503720 20664
rect 503772 20652 503778 20664
rect 504358 20652 504364 20664
rect 503772 20624 504364 20652
rect 503772 20612 503778 20624
rect 504358 20612 504364 20624
rect 504416 20612 504422 20664
rect 524874 20612 524880 20664
rect 524932 20652 524938 20664
rect 551278 20652 551284 20664
rect 524932 20624 551284 20652
rect 524932 20612 524938 20624
rect 551278 20612 551284 20624
rect 551336 20612 551342 20664
rect 22646 20544 22652 20596
rect 22704 20584 22710 20596
rect 458174 20584 458180 20596
rect 22704 20556 458180 20584
rect 22704 20544 22710 20556
rect 458174 20544 458180 20556
rect 458232 20544 458238 20596
rect 480254 20544 480260 20596
rect 480312 20584 480318 20596
rect 556614 20584 556620 20596
rect 480312 20556 556620 20584
rect 480312 20544 480318 20556
rect 556614 20544 556620 20556
rect 556672 20544 556678 20596
rect 43622 20476 43628 20528
rect 43680 20516 43686 20528
rect 387794 20516 387800 20528
rect 43680 20488 387800 20516
rect 43680 20476 43686 20488
rect 387794 20476 387800 20488
rect 387852 20476 387858 20528
rect 423674 20476 423680 20528
rect 423732 20516 423738 20528
rect 580074 20516 580080 20528
rect 423732 20488 580080 20516
rect 423732 20476 423738 20488
rect 580074 20476 580080 20488
rect 580132 20476 580138 20528
rect 28534 20408 28540 20460
rect 28592 20448 28598 20460
rect 367094 20448 367100 20460
rect 28592 20420 367100 20448
rect 28592 20408 28598 20420
rect 367094 20408 367100 20420
rect 367152 20408 367158 20460
rect 421006 20408 421012 20460
rect 421064 20448 421070 20460
rect 546678 20448 546684 20460
rect 421064 20420 546684 20448
rect 421064 20408 421070 20420
rect 546678 20408 546684 20420
rect 546736 20408 546742 20460
rect 38378 20340 38384 20392
rect 38436 20380 38442 20392
rect 229094 20380 229100 20392
rect 38436 20352 229100 20380
rect 38436 20340 38442 20352
rect 229094 20340 229100 20352
rect 229152 20340 229158 20392
rect 231946 20340 231952 20392
rect 232004 20380 232010 20392
rect 564618 20380 564624 20392
rect 232004 20352 564624 20380
rect 232004 20340 232010 20352
rect 564618 20340 564624 20352
rect 564676 20340 564682 20392
rect 46198 20272 46204 20324
rect 46256 20312 46262 20324
rect 219526 20312 219532 20324
rect 46256 20284 219532 20312
rect 46256 20272 46262 20284
rect 219526 20272 219532 20284
rect 219584 20272 219590 20324
rect 251266 20272 251272 20324
rect 251324 20312 251330 20324
rect 583202 20312 583208 20324
rect 251324 20284 583208 20312
rect 251324 20272 251330 20284
rect 583202 20272 583208 20284
rect 583260 20272 583266 20324
rect 55122 20204 55128 20256
rect 55180 20244 55186 20256
rect 367186 20244 367192 20256
rect 55180 20216 367192 20244
rect 55180 20204 55186 20216
rect 367186 20204 367192 20216
rect 367244 20204 367250 20256
rect 434714 20204 434720 20256
rect 434772 20244 434778 20256
rect 559190 20244 559196 20256
rect 434772 20216 559196 20244
rect 434772 20204 434778 20216
rect 559190 20204 559196 20216
rect 559248 20204 559254 20256
rect 55766 20136 55772 20188
rect 55824 20176 55830 20188
rect 227714 20176 227720 20188
rect 55824 20148 227720 20176
rect 55824 20136 55830 20148
rect 227714 20136 227720 20148
rect 227772 20136 227778 20188
rect 292574 20136 292580 20188
rect 292632 20176 292638 20188
rect 554314 20176 554320 20188
rect 292632 20148 554320 20176
rect 292632 20136 292638 20148
rect 554314 20136 554320 20148
rect 554372 20136 554378 20188
rect 58342 20068 58348 20120
rect 58400 20108 58406 20120
rect 211246 20108 211252 20120
rect 58400 20080 211252 20108
rect 58400 20068 58406 20080
rect 211246 20068 211252 20080
rect 211304 20068 211310 20120
rect 253934 20068 253940 20120
rect 253992 20108 253998 20120
rect 548150 20108 548156 20120
rect 253992 20080 548156 20108
rect 253992 20068 253998 20080
rect 548150 20068 548156 20080
rect 548208 20068 548214 20120
rect 184934 20000 184940 20052
rect 184992 20040 184998 20052
rect 553578 20040 553584 20052
rect 184992 20012 553584 20040
rect 184992 20000 184998 20012
rect 553578 20000 553584 20012
rect 553636 20000 553642 20052
rect 39666 19932 39672 19984
rect 39724 19972 39730 19984
rect 139394 19972 139400 19984
rect 39724 19944 139400 19972
rect 39724 19932 39730 19944
rect 139394 19932 139400 19944
rect 139452 19932 139458 19984
rect 183646 19932 183652 19984
rect 183704 19972 183710 19984
rect 555234 19972 555240 19984
rect 183704 19944 555240 19972
rect 183704 19932 183710 19944
rect 555234 19932 555240 19944
rect 555292 19932 555298 19984
rect 55858 19864 55864 19916
rect 55916 19904 55922 19916
rect 153194 19904 153200 19916
rect 55916 19876 153200 19904
rect 55916 19864 55922 19876
rect 153194 19864 153200 19876
rect 153252 19864 153258 19916
rect 360194 19864 360200 19916
rect 360252 19904 360258 19916
rect 547598 19904 547604 19916
rect 360252 19876 547604 19904
rect 360252 19864 360258 19876
rect 547598 19864 547604 19876
rect 547656 19864 547662 19916
rect 57790 19796 57796 19848
rect 57848 19836 57854 19848
rect 130194 19836 130200 19848
rect 57848 19808 130200 19836
rect 57848 19796 57854 19808
rect 130194 19796 130200 19808
rect 130252 19796 130258 19848
rect 504358 19796 504364 19848
rect 504416 19836 504422 19848
rect 567654 19836 567660 19848
rect 504416 19808 567660 19836
rect 504416 19796 504422 19808
rect 567654 19796 567660 19808
rect 567712 19796 567718 19848
rect 22554 19728 22560 19780
rect 22612 19768 22618 19780
rect 462314 19768 462320 19780
rect 22612 19740 462320 19768
rect 22612 19728 22618 19740
rect 462314 19728 462320 19740
rect 462372 19728 462378 19780
rect 465074 19728 465080 19780
rect 465132 19768 465138 19780
rect 571794 19768 571800 19780
rect 465132 19740 571800 19768
rect 465132 19728 465138 19740
rect 571794 19728 571800 19740
rect 571852 19728 571858 19780
rect 44910 19660 44916 19712
rect 44968 19700 44974 19712
rect 189074 19700 189080 19712
rect 44968 19672 189080 19700
rect 44968 19660 44974 19672
rect 189074 19660 189080 19672
rect 189132 19660 189138 19712
rect 35710 19252 35716 19304
rect 35768 19292 35774 19304
rect 219434 19292 219440 19304
rect 35768 19264 219440 19292
rect 35768 19252 35774 19264
rect 219434 19252 219440 19264
rect 219492 19252 219498 19304
rect 247034 19252 247040 19304
rect 247092 19292 247098 19304
rect 573358 19292 573364 19304
rect 247092 19264 573364 19292
rect 247092 19252 247098 19264
rect 573358 19252 573364 19264
rect 573416 19252 573422 19304
rect 54754 19184 54760 19236
rect 54812 19224 54818 19236
rect 293954 19224 293960 19236
rect 54812 19196 293960 19224
rect 54812 19184 54818 19196
rect 293954 19184 293960 19196
rect 294012 19184 294018 19236
rect 358814 19184 358820 19236
rect 358872 19224 358878 19236
rect 551370 19224 551376 19236
rect 358872 19196 551376 19224
rect 358872 19184 358878 19196
rect 551370 19184 551376 19196
rect 551428 19184 551434 19236
rect 45278 19116 45284 19168
rect 45336 19156 45342 19168
rect 202874 19156 202880 19168
rect 45336 19128 202880 19156
rect 45336 19116 45342 19128
rect 202874 19116 202880 19128
rect 202932 19116 202938 19168
rect 419534 19116 419540 19168
rect 419592 19156 419598 19168
rect 565078 19156 565084 19168
rect 419592 19128 565084 19156
rect 419592 19116 419598 19128
rect 565078 19116 565084 19128
rect 565136 19116 565142 19168
rect 53374 19048 53380 19100
rect 53432 19088 53438 19100
rect 205634 19088 205640 19100
rect 53432 19060 205640 19088
rect 53432 19048 53438 19060
rect 205634 19048 205640 19060
rect 205692 19048 205698 19100
rect 463694 19048 463700 19100
rect 463752 19088 463758 19100
rect 574278 19088 574284 19100
rect 463752 19060 574284 19088
rect 463752 19048 463758 19060
rect 574278 19048 574284 19060
rect 574336 19048 574342 19100
rect 41322 18980 41328 19032
rect 41380 19020 41386 19032
rect 183554 19020 183560 19032
rect 41380 18992 183560 19020
rect 41380 18980 41386 18992
rect 183554 18980 183560 18992
rect 183612 18980 183618 19032
rect 459554 18980 459560 19032
rect 459612 19020 459618 19032
rect 563514 19020 563520 19032
rect 459612 18992 563520 19020
rect 459612 18980 459618 18992
rect 563514 18980 563520 18992
rect 563572 18980 563578 19032
rect 36630 18912 36636 18964
rect 36688 18952 36694 18964
rect 149054 18952 149060 18964
rect 36688 18924 149060 18952
rect 36688 18912 36694 18924
rect 149054 18912 149060 18924
rect 149112 18912 149118 18964
rect 317414 18912 317420 18964
rect 317472 18952 317478 18964
rect 557994 18952 558000 18964
rect 317472 18924 558000 18952
rect 317472 18912 317478 18924
rect 557994 18912 558000 18924
rect 558052 18912 558058 18964
rect 36906 18844 36912 18896
rect 36964 18884 36970 18896
rect 146294 18884 146300 18896
rect 36964 18856 146300 18884
rect 36964 18844 36970 18856
rect 146294 18844 146300 18856
rect 146352 18844 146358 18896
rect 271874 18844 271880 18896
rect 271932 18884 271938 18896
rect 567470 18884 567476 18896
rect 271932 18856 567476 18884
rect 271932 18844 271938 18856
rect 567470 18844 567476 18856
rect 567528 18844 567534 18896
rect 57422 18776 57428 18828
rect 57480 18816 57486 18828
rect 165614 18816 165620 18828
rect 57480 18788 165620 18816
rect 57480 18776 57486 18788
rect 165614 18776 165620 18788
rect 165672 18776 165678 18828
rect 251174 18776 251180 18828
rect 251232 18816 251238 18828
rect 561950 18816 561956 18828
rect 251232 18788 561956 18816
rect 251232 18776 251238 18788
rect 561950 18776 561956 18788
rect 562008 18776 562014 18828
rect 49970 18708 49976 18760
rect 50028 18748 50034 18760
rect 125594 18748 125600 18760
rect 50028 18720 125600 18748
rect 50028 18708 50034 18720
rect 125594 18708 125600 18720
rect 125652 18708 125658 18760
rect 136634 18708 136640 18760
rect 136692 18748 136698 18760
rect 570138 18748 570144 18760
rect 136692 18720 570144 18748
rect 136692 18708 136698 18720
rect 570138 18708 570144 18720
rect 570196 18708 570202 18760
rect 50338 18640 50344 18692
rect 50396 18680 50402 18692
rect 104158 18680 104164 18692
rect 50396 18652 104164 18680
rect 50396 18640 50402 18652
rect 104158 18640 104164 18652
rect 104216 18640 104222 18692
rect 113174 18640 113180 18692
rect 113232 18680 113238 18692
rect 549438 18680 549444 18692
rect 113232 18652 549444 18680
rect 113232 18640 113238 18652
rect 549438 18640 549444 18652
rect 549496 18640 549502 18692
rect 99374 18572 99380 18624
rect 99432 18612 99438 18624
rect 577406 18612 577412 18624
rect 99432 18584 577412 18612
rect 99432 18572 99438 18584
rect 577406 18572 577412 18584
rect 577464 18572 577470 18624
rect 46106 18504 46112 18556
rect 46164 18544 46170 18556
rect 147674 18544 147680 18556
rect 46164 18516 147680 18544
rect 46164 18504 46170 18516
rect 147674 18504 147680 18516
rect 147732 18504 147738 18556
rect 466454 18504 466460 18556
rect 466512 18544 466518 18556
rect 568758 18544 568764 18556
rect 466512 18516 568764 18544
rect 466512 18504 466518 18516
rect 568758 18504 568764 18516
rect 568816 18504 568822 18556
rect 55950 18436 55956 18488
rect 56008 18476 56014 18488
rect 154574 18476 154580 18488
rect 56008 18448 154580 18476
rect 56008 18436 56014 18448
rect 154574 18436 154580 18448
rect 154632 18436 154638 18488
rect 469214 18436 469220 18488
rect 469272 18476 469278 18488
rect 545298 18476 545304 18488
rect 469272 18448 545304 18476
rect 469272 18436 469278 18448
rect 545298 18436 545304 18448
rect 545356 18436 545362 18488
rect 45922 18368 45928 18420
rect 45980 18408 45986 18420
rect 83458 18408 83464 18420
rect 45980 18380 83464 18408
rect 45980 18368 45986 18380
rect 83458 18368 83464 18380
rect 83516 18368 83522 18420
rect 533338 18368 533344 18420
rect 533396 18408 533402 18420
rect 543274 18408 543280 18420
rect 533396 18380 543280 18408
rect 533396 18368 533402 18380
rect 543274 18368 543280 18380
rect 543332 18368 543338 18420
rect 46842 18300 46848 18352
rect 46900 18340 46906 18352
rect 120074 18340 120080 18352
rect 46900 18312 120080 18340
rect 46900 18300 46906 18312
rect 120074 18300 120080 18312
rect 120132 18300 120138 18352
rect 97994 17892 98000 17944
rect 98052 17932 98058 17944
rect 583386 17932 583392 17944
rect 98052 17904 583392 17932
rect 98052 17892 98058 17904
rect 583386 17892 583392 17904
rect 583444 17892 583450 17944
rect 106366 17824 106372 17876
rect 106424 17864 106430 17876
rect 581362 17864 581368 17876
rect 106424 17836 581368 17864
rect 106424 17824 106430 17836
rect 581362 17824 581368 17836
rect 581420 17824 581426 17876
rect 42058 17756 42064 17808
rect 42116 17796 42122 17808
rect 116026 17796 116032 17808
rect 42116 17768 116032 17796
rect 42116 17756 42122 17768
rect 116026 17756 116032 17768
rect 116084 17756 116090 17808
rect 157334 17756 157340 17808
rect 157392 17796 157398 17808
rect 583570 17796 583576 17808
rect 157392 17768 583576 17796
rect 157392 17756 157398 17768
rect 583570 17756 583576 17768
rect 583628 17756 583634 17808
rect 40954 17688 40960 17740
rect 41012 17728 41018 17740
rect 375374 17728 375380 17740
rect 41012 17700 375380 17728
rect 41012 17688 41018 17700
rect 375374 17688 375380 17700
rect 375432 17688 375438 17740
rect 378134 17688 378140 17740
rect 378192 17728 378198 17740
rect 546954 17728 546960 17740
rect 378192 17700 546960 17728
rect 378192 17688 378198 17700
rect 546954 17688 546960 17700
rect 547012 17688 547018 17740
rect 58066 17620 58072 17672
rect 58124 17660 58130 17672
rect 329834 17660 329840 17672
rect 58124 17632 329840 17660
rect 58124 17620 58130 17632
rect 329834 17620 329840 17632
rect 329892 17620 329898 17672
rect 340874 17620 340880 17672
rect 340932 17660 340938 17672
rect 577682 17660 577688 17672
rect 340932 17632 577688 17660
rect 340932 17620 340938 17632
rect 577682 17620 577688 17632
rect 577740 17620 577746 17672
rect 59906 17552 59912 17604
rect 59964 17592 59970 17604
rect 245746 17592 245752 17604
rect 59964 17564 245752 17592
rect 59964 17552 59970 17564
rect 245746 17552 245752 17564
rect 245804 17552 245810 17604
rect 460934 17552 460940 17604
rect 460992 17592 460998 17604
rect 573266 17592 573272 17604
rect 460992 17564 573272 17592
rect 460992 17552 460998 17564
rect 573266 17552 573272 17564
rect 573324 17552 573330 17604
rect 57698 17484 57704 17536
rect 57756 17524 57762 17536
rect 237374 17524 237380 17536
rect 57756 17496 237380 17524
rect 57756 17484 57762 17496
rect 237374 17484 237380 17496
rect 237432 17484 237438 17536
rect 527818 17484 527824 17536
rect 527876 17524 527882 17536
rect 544286 17524 544292 17536
rect 527876 17496 544292 17524
rect 527876 17484 527882 17496
rect 544286 17484 544292 17496
rect 544344 17484 544350 17536
rect 59814 17416 59820 17468
rect 59872 17456 59878 17468
rect 234614 17456 234620 17468
rect 59872 17428 234620 17456
rect 59872 17416 59878 17428
rect 234614 17416 234620 17428
rect 234672 17416 234678 17468
rect 427814 17416 427820 17468
rect 427872 17456 427878 17468
rect 571610 17456 571616 17468
rect 427872 17428 571616 17456
rect 427872 17416 427878 17428
rect 571610 17416 571616 17428
rect 571668 17416 571674 17468
rect 57330 17348 57336 17400
rect 57388 17388 57394 17400
rect 142798 17388 142804 17400
rect 57388 17360 142804 17388
rect 57388 17348 57394 17360
rect 142798 17348 142804 17360
rect 142856 17348 142862 17400
rect 414014 17348 414020 17400
rect 414072 17388 414078 17400
rect 571334 17388 571340 17400
rect 414072 17360 571340 17388
rect 414072 17348 414078 17360
rect 571334 17348 571340 17360
rect 571392 17348 571398 17400
rect 45462 17280 45468 17332
rect 45520 17320 45526 17332
rect 115934 17320 115940 17332
rect 45520 17292 115940 17320
rect 45520 17280 45526 17292
rect 115934 17280 115940 17292
rect 115992 17280 115998 17332
rect 259454 17280 259460 17332
rect 259512 17320 259518 17332
rect 541894 17320 541900 17332
rect 259512 17292 541900 17320
rect 259512 17280 259518 17292
rect 541894 17280 541900 17292
rect 541952 17280 541958 17332
rect 120074 17212 120080 17264
rect 120132 17252 120138 17264
rect 579982 17252 579988 17264
rect 120132 17224 579988 17252
rect 120132 17212 120138 17224
rect 579982 17212 579988 17224
rect 580040 17212 580046 17264
rect 52362 17144 52368 17196
rect 52420 17184 52426 17196
rect 170398 17184 170404 17196
rect 52420 17156 170404 17184
rect 52420 17144 52426 17156
rect 170398 17144 170404 17156
rect 170456 17144 170462 17196
rect 106274 16600 106280 16652
rect 106332 16640 106338 16652
rect 560294 16640 560300 16652
rect 106332 16612 560300 16640
rect 106332 16600 106338 16612
rect 560294 16600 560300 16612
rect 560352 16600 560358 16652
rect 48038 16532 48044 16584
rect 48096 16572 48102 16584
rect 164326 16572 164332 16584
rect 48096 16544 164332 16572
rect 48096 16532 48102 16544
rect 164326 16532 164332 16544
rect 164384 16532 164390 16584
rect 233234 16532 233240 16584
rect 233292 16572 233298 16584
rect 548794 16572 548800 16584
rect 233292 16544 548800 16572
rect 233292 16532 233298 16544
rect 548794 16532 548800 16544
rect 548852 16532 548858 16584
rect 48130 16464 48136 16516
rect 48188 16504 48194 16516
rect 161566 16504 161572 16516
rect 48188 16476 161572 16504
rect 48188 16464 48194 16476
rect 161566 16464 161572 16476
rect 161624 16464 161630 16516
rect 361574 16464 361580 16516
rect 361632 16504 361638 16516
rect 581730 16504 581736 16516
rect 361632 16476 581736 16504
rect 361632 16464 361638 16476
rect 581730 16464 581736 16476
rect 581788 16464 581794 16516
rect 58802 16396 58808 16448
rect 58860 16436 58866 16448
rect 157978 16436 157984 16448
rect 58860 16408 157984 16436
rect 58860 16396 58866 16408
rect 157978 16396 157984 16408
rect 158036 16396 158042 16448
rect 335446 16396 335452 16448
rect 335504 16436 335510 16448
rect 541434 16436 541440 16448
rect 335504 16408 541440 16436
rect 335504 16396 335510 16408
rect 541434 16396 541440 16408
rect 541492 16396 541498 16448
rect 347774 16328 347780 16380
rect 347832 16368 347838 16380
rect 544470 16368 544476 16380
rect 347832 16340 544476 16368
rect 347832 16328 347838 16340
rect 544470 16328 544476 16340
rect 544528 16328 544534 16380
rect 289814 16260 289820 16312
rect 289872 16300 289878 16312
rect 557074 16300 557080 16312
rect 289872 16272 557080 16300
rect 289872 16260 289878 16272
rect 557074 16260 557080 16272
rect 557132 16260 557138 16312
rect 264974 16192 264980 16244
rect 265032 16232 265038 16244
rect 564894 16232 564900 16244
rect 265032 16204 564900 16232
rect 265032 16192 265038 16204
rect 564894 16192 564900 16204
rect 564952 16192 564958 16244
rect 253474 16124 253480 16176
rect 253532 16164 253538 16176
rect 572806 16164 572812 16176
rect 253532 16136 572812 16164
rect 253532 16124 253538 16136
rect 572806 16124 572812 16136
rect 572864 16124 572870 16176
rect 228266 16056 228272 16108
rect 228324 16096 228330 16108
rect 558914 16096 558920 16108
rect 228324 16068 558920 16096
rect 228324 16056 228330 16068
rect 558914 16056 558920 16068
rect 558972 16056 558978 16108
rect 226334 15988 226340 16040
rect 226392 16028 226398 16040
rect 570046 16028 570052 16040
rect 226392 16000 570052 16028
rect 226392 15988 226398 16000
rect 570046 15988 570052 16000
rect 570104 15988 570110 16040
rect 33962 15920 33968 15972
rect 34020 15960 34026 15972
rect 130562 15960 130568 15972
rect 34020 15932 130568 15960
rect 34020 15920 34026 15932
rect 130562 15920 130568 15932
rect 130620 15920 130626 15972
rect 229370 15920 229376 15972
rect 229428 15960 229434 15972
rect 575750 15960 575756 15972
rect 229428 15932 575756 15960
rect 229428 15920 229434 15932
rect 575750 15920 575756 15932
rect 575808 15920 575814 15972
rect 35618 15852 35624 15904
rect 35676 15892 35682 15904
rect 158898 15892 158904 15904
rect 35676 15864 158904 15892
rect 35676 15852 35682 15864
rect 158898 15852 158904 15864
rect 158956 15852 158962 15904
rect 171962 15852 171968 15904
rect 172020 15892 172026 15904
rect 564802 15892 564808 15904
rect 172020 15864 564808 15892
rect 172020 15852 172026 15864
rect 564802 15852 564808 15864
rect 564860 15852 564866 15904
rect 398834 15784 398840 15836
rect 398892 15824 398898 15836
rect 544102 15824 544108 15836
rect 398892 15796 544108 15824
rect 398892 15784 398898 15796
rect 544102 15784 544108 15796
rect 544160 15784 544166 15836
rect 447134 15716 447140 15768
rect 447192 15756 447198 15768
rect 549806 15756 549812 15768
rect 447192 15728 549812 15756
rect 447192 15716 447198 15728
rect 549806 15716 549812 15728
rect 549864 15716 549870 15768
rect 522298 15648 522304 15700
rect 522356 15688 522362 15700
rect 567562 15688 567568 15700
rect 522356 15660 567568 15688
rect 522356 15648 522362 15660
rect 567562 15648 567568 15660
rect 567620 15648 567626 15700
rect 242894 15104 242900 15156
rect 242952 15144 242958 15156
rect 552750 15144 552756 15156
rect 242952 15116 552756 15144
rect 242952 15104 242958 15116
rect 552750 15104 552756 15116
rect 552808 15104 552814 15156
rect 380894 15036 380900 15088
rect 380952 15076 380958 15088
rect 540054 15076 540060 15088
rect 380952 15048 540060 15076
rect 380952 15036 380958 15048
rect 540054 15036 540060 15048
rect 540112 15036 540118 15088
rect 393314 14968 393320 15020
rect 393372 15008 393378 15020
rect 543734 15008 543740 15020
rect 393372 14980 543740 15008
rect 393372 14968 393378 14980
rect 543734 14968 543740 14980
rect 543792 14968 543798 15020
rect 404354 14900 404360 14952
rect 404412 14940 404418 14952
rect 546034 14940 546040 14952
rect 404412 14912 546040 14940
rect 404412 14900 404418 14912
rect 546034 14900 546040 14912
rect 546092 14900 546098 14952
rect 444374 14832 444380 14884
rect 444432 14872 444438 14884
rect 576118 14872 576124 14884
rect 444432 14844 576124 14872
rect 444432 14832 444438 14844
rect 576118 14832 576124 14844
rect 576176 14832 576182 14884
rect 426434 14764 426440 14816
rect 426492 14804 426498 14816
rect 544010 14804 544016 14816
rect 426492 14776 544016 14804
rect 426492 14764 426498 14776
rect 544010 14764 544016 14776
rect 544068 14764 544074 14816
rect 403618 14696 403624 14748
rect 403676 14736 403682 14748
rect 542262 14736 542268 14748
rect 403676 14708 542268 14736
rect 403676 14696 403682 14708
rect 542262 14696 542268 14708
rect 542320 14696 542326 14748
rect 398834 14628 398840 14680
rect 398892 14668 398898 14680
rect 541986 14668 541992 14680
rect 398892 14640 541992 14668
rect 398892 14628 398898 14640
rect 541986 14628 541992 14640
rect 542044 14628 542050 14680
rect 382366 14560 382372 14612
rect 382424 14600 382430 14612
rect 547230 14600 547236 14612
rect 382424 14572 547236 14600
rect 382424 14560 382430 14572
rect 547230 14560 547236 14572
rect 547288 14560 547294 14612
rect 378410 14492 378416 14544
rect 378468 14532 378474 14544
rect 548702 14532 548708 14544
rect 378468 14504 548708 14532
rect 378468 14492 378474 14504
rect 548702 14492 548708 14504
rect 548760 14492 548766 14544
rect 247586 14424 247592 14476
rect 247644 14464 247650 14476
rect 550082 14464 550088 14476
rect 247644 14436 550088 14464
rect 247644 14424 247650 14436
rect 550082 14424 550088 14436
rect 550140 14424 550146 14476
rect 430574 14356 430580 14408
rect 430632 14396 430638 14408
rect 543182 14396 543188 14408
rect 430632 14368 543188 14396
rect 430632 14356 430638 14368
rect 543182 14356 543188 14368
rect 543240 14356 543246 14408
rect 434806 14288 434812 14340
rect 434864 14328 434870 14340
rect 546770 14328 546776 14340
rect 434864 14300 546776 14328
rect 434864 14288 434870 14300
rect 546770 14288 546776 14300
rect 546828 14288 546834 14340
rect 433334 14220 433340 14272
rect 433392 14260 433398 14272
rect 541802 14260 541808 14272
rect 433392 14232 541808 14260
rect 433392 14220 433398 14232
rect 541802 14220 541808 14232
rect 541860 14220 541866 14272
rect 320174 13744 320180 13796
rect 320232 13784 320238 13796
rect 563422 13784 563428 13796
rect 320232 13756 563428 13784
rect 320232 13744 320238 13756
rect 563422 13744 563428 13756
rect 563480 13744 563486 13796
rect 372614 13676 372620 13728
rect 372672 13716 372678 13728
rect 583754 13716 583760 13728
rect 372672 13688 583760 13716
rect 372672 13676 372678 13688
rect 583754 13676 583760 13688
rect 583812 13676 583818 13728
rect 357526 13608 357532 13660
rect 357584 13648 357590 13660
rect 540330 13648 540336 13660
rect 357584 13620 540336 13648
rect 357584 13608 357590 13620
rect 540330 13608 540336 13620
rect 540388 13608 540394 13660
rect 349154 13540 349160 13592
rect 349212 13580 349218 13592
rect 542998 13580 543004 13592
rect 349212 13552 543004 13580
rect 349212 13540 349218 13552
rect 542998 13540 543004 13552
rect 543056 13540 543062 13592
rect 346946 13472 346952 13524
rect 347004 13512 347010 13524
rect 541618 13512 541624 13524
rect 347004 13484 541624 13512
rect 347004 13472 347010 13484
rect 541618 13472 541624 13484
rect 541676 13472 541682 13524
rect 367738 13404 367744 13456
rect 367796 13444 367802 13456
rect 579154 13444 579160 13456
rect 367796 13416 579160 13444
rect 367796 13404 367802 13416
rect 579154 13404 579160 13416
rect 579212 13404 579218 13456
rect 311434 13336 311440 13388
rect 311492 13376 311498 13388
rect 562410 13376 562416 13388
rect 311492 13348 562416 13376
rect 311492 13336 311498 13348
rect 562410 13336 562416 13348
rect 562468 13336 562474 13388
rect 297266 13268 297272 13320
rect 297324 13308 297330 13320
rect 558178 13308 558184 13320
rect 297324 13280 558184 13308
rect 297324 13268 297330 13280
rect 558178 13268 558184 13280
rect 558236 13268 558242 13320
rect 286594 13200 286600 13252
rect 286652 13240 286658 13252
rect 559558 13240 559564 13252
rect 286652 13212 559564 13240
rect 286652 13200 286658 13212
rect 559558 13200 559564 13212
rect 559616 13200 559622 13252
rect 234614 13132 234620 13184
rect 234672 13172 234678 13184
rect 553762 13172 553768 13184
rect 234672 13144 553768 13172
rect 234672 13132 234678 13144
rect 553762 13132 553768 13144
rect 553820 13132 553826 13184
rect 242894 13064 242900 13116
rect 242952 13104 242958 13116
rect 578694 13104 578700 13116
rect 242952 13076 578700 13104
rect 242952 13064 242958 13076
rect 578694 13064 578700 13076
rect 578752 13064 578758 13116
rect 364610 12996 364616 13048
rect 364668 13036 364674 13048
rect 545942 13036 545948 13048
rect 364668 13008 545948 13036
rect 364668 12996 364674 13008
rect 545942 12996 545948 13008
rect 546000 12996 546006 13048
rect 453298 12928 453304 12980
rect 453356 12968 453362 12980
rect 559006 12968 559012 12980
rect 453356 12940 559012 12968
rect 453356 12928 453362 12940
rect 559006 12928 559012 12940
rect 559064 12928 559070 12980
rect 473998 12860 474004 12912
rect 474056 12900 474062 12912
rect 549714 12900 549720 12912
rect 474056 12872 549720 12900
rect 474056 12860 474062 12872
rect 549714 12860 549720 12872
rect 549772 12860 549778 12912
rect 190546 12384 190552 12436
rect 190604 12424 190610 12436
rect 583662 12424 583668 12436
rect 190604 12396 583668 12424
rect 190604 12384 190610 12396
rect 583662 12384 583668 12396
rect 583720 12384 583726 12436
rect 313274 12316 313280 12368
rect 313332 12356 313338 12368
rect 543090 12356 543096 12368
rect 313332 12328 543096 12356
rect 313332 12316 313338 12328
rect 543090 12316 543096 12328
rect 543148 12316 543154 12368
rect 314746 12248 314752 12300
rect 314804 12288 314810 12300
rect 544562 12288 544568 12300
rect 314804 12260 544568 12288
rect 314804 12248 314810 12260
rect 544562 12248 544568 12260
rect 544620 12248 544626 12300
rect 321646 12180 321652 12232
rect 321704 12220 321710 12232
rect 540514 12220 540520 12232
rect 321704 12192 540520 12220
rect 321704 12180 321710 12192
rect 540514 12180 540520 12192
rect 540572 12180 540578 12232
rect 324314 12112 324320 12164
rect 324372 12152 324378 12164
rect 541710 12152 541716 12164
rect 324372 12124 541716 12152
rect 324372 12112 324378 12124
rect 541710 12112 541716 12124
rect 541768 12112 541774 12164
rect 328454 12044 328460 12096
rect 328512 12084 328518 12096
rect 543458 12084 543464 12096
rect 328512 12056 543464 12084
rect 328512 12044 328518 12056
rect 543458 12044 543464 12056
rect 543516 12044 543522 12096
rect 351914 11976 351920 12028
rect 351972 12016 351978 12028
rect 551186 12016 551192 12028
rect 351972 11988 551192 12016
rect 351972 11976 351978 11988
rect 551186 11976 551192 11988
rect 551244 11976 551250 12028
rect 346394 11908 346400 11960
rect 346452 11948 346458 11960
rect 543550 11948 543556 11960
rect 346452 11920 543556 11948
rect 346452 11908 346458 11920
rect 543550 11908 543556 11920
rect 543608 11908 543614 11960
rect 363046 11840 363052 11892
rect 363104 11880 363110 11892
rect 548058 11880 548064 11892
rect 363104 11852 548064 11880
rect 363104 11840 363110 11852
rect 548058 11840 548064 11852
rect 548116 11840 548122 11892
rect 256694 11772 256700 11824
rect 256752 11812 256758 11824
rect 577590 11812 577596 11824
rect 256752 11784 577596 11812
rect 256752 11772 256758 11784
rect 577590 11772 577596 11784
rect 577648 11772 577654 11824
rect 239306 11704 239312 11756
rect 239364 11744 239370 11756
rect 576302 11744 576308 11756
rect 239364 11716 576308 11744
rect 239364 11704 239370 11716
rect 576302 11704 576308 11716
rect 576360 11704 576366 11756
rect 357434 11636 357440 11688
rect 357492 11676 357498 11688
rect 542354 11676 542360 11688
rect 357492 11648 542360 11676
rect 357492 11636 357498 11648
rect 542354 11636 542360 11648
rect 542412 11636 542418 11688
rect 451918 11568 451924 11620
rect 451976 11608 451982 11620
rect 540238 11608 540244 11620
rect 451976 11580 540244 11608
rect 451976 11568 451982 11580
rect 540238 11568 540244 11580
rect 540296 11568 540302 11620
rect 505738 11500 505744 11552
rect 505796 11540 505802 11552
rect 543826 11540 543832 11552
rect 505796 11512 543832 11540
rect 505796 11500 505802 11512
rect 543826 11500 543832 11512
rect 543884 11500 543890 11552
rect 48958 10956 48964 11008
rect 49016 10996 49022 11008
rect 191834 10996 191840 11008
rect 49016 10968 191840 10996
rect 49016 10956 49022 10968
rect 191834 10956 191840 10968
rect 191892 10956 191898 11008
rect 303890 10344 303896 10396
rect 303948 10384 303954 10396
rect 557718 10384 557724 10396
rect 303948 10356 557724 10384
rect 303948 10344 303954 10356
rect 557718 10344 557724 10356
rect 557776 10344 557782 10396
rect 141234 10276 141240 10328
rect 141292 10316 141298 10328
rect 555142 10316 555148 10328
rect 141292 10288 555148 10316
rect 141292 10276 141298 10288
rect 555142 10276 555148 10288
rect 555200 10276 555206 10328
rect 307938 9052 307944 9104
rect 307996 9092 308002 9104
rect 550818 9092 550824 9104
rect 307996 9064 550824 9092
rect 307996 9052 308002 9064
rect 550818 9052 550824 9064
rect 550876 9052 550882 9104
rect 249978 8984 249984 9036
rect 250036 9024 250042 9036
rect 553394 9024 553400 9036
rect 250036 8996 553400 9024
rect 250036 8984 250042 8996
rect 553394 8984 553400 8996
rect 553452 8984 553458 9036
rect 208578 8916 208584 8968
rect 208636 8956 208642 8968
rect 556522 8956 556528 8968
rect 208636 8928 556528 8956
rect 208636 8916 208642 8928
rect 556522 8916 556528 8928
rect 556580 8916 556586 8968
rect 194410 7556 194416 7608
rect 194468 7596 194474 7608
rect 556246 7596 556252 7608
rect 194468 7568 556252 7596
rect 194468 7556 194474 7568
rect 556246 7556 556252 7568
rect 556304 7556 556310 7608
rect 567838 7556 567844 7608
rect 567896 7596 567902 7608
rect 579798 7596 579804 7608
rect 567896 7568 579804 7596
rect 567896 7556 567902 7568
rect 579798 7556 579804 7568
rect 579856 7556 579862 7608
rect 463970 6808 463976 6860
rect 464028 6848 464034 6860
rect 561214 6848 561220 6860
rect 464028 6820 561220 6848
rect 464028 6808 464034 6820
rect 561214 6808 561220 6820
rect 561272 6808 561278 6860
rect 446214 6740 446220 6792
rect 446272 6780 446278 6792
rect 545482 6780 545488 6792
rect 446272 6752 545488 6780
rect 446272 6740 446278 6752
rect 545482 6740 545488 6752
rect 545540 6740 545546 6792
rect 439130 6672 439136 6724
rect 439188 6712 439194 6724
rect 541066 6712 541072 6724
rect 439188 6684 541072 6712
rect 439188 6672 439194 6684
rect 541066 6672 541072 6684
rect 541124 6672 541130 6724
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 474550 6604 474556 6656
rect 474608 6644 474614 6656
rect 582374 6644 582380 6656
rect 474608 6616 582380 6644
rect 474608 6604 474614 6616
rect 582374 6604 582380 6616
rect 582432 6604 582438 6656
rect 460382 6536 460388 6588
rect 460440 6576 460446 6588
rect 569494 6576 569500 6588
rect 460440 6548 569500 6576
rect 460440 6536 460446 6548
rect 569494 6536 569500 6548
rect 569552 6536 569558 6588
rect 449802 6468 449808 6520
rect 449860 6508 449866 6520
rect 566366 6508 566372 6520
rect 449860 6480 566372 6508
rect 449860 6468 449866 6480
rect 566366 6468 566372 6480
rect 566424 6468 566430 6520
rect 442626 6400 442632 6452
rect 442684 6440 442690 6452
rect 575014 6440 575020 6452
rect 442684 6412 575020 6440
rect 442684 6400 442690 6412
rect 575014 6400 575020 6412
rect 575072 6400 575078 6452
rect 432046 6332 432052 6384
rect 432104 6372 432110 6384
rect 570506 6372 570512 6384
rect 432104 6344 570512 6372
rect 432104 6332 432110 6344
rect 570506 6332 570512 6344
rect 570564 6332 570570 6384
rect 424962 6264 424968 6316
rect 425020 6304 425026 6316
rect 564986 6304 564992 6316
rect 425020 6276 564992 6304
rect 425020 6264 425026 6276
rect 564986 6264 564992 6276
rect 565044 6264 565050 6316
rect 389450 6196 389456 6248
rect 389508 6236 389514 6248
rect 559282 6236 559288 6248
rect 389508 6208 559288 6236
rect 389508 6196 389514 6208
rect 559282 6196 559288 6208
rect 559340 6196 559346 6248
rect 300762 6128 300768 6180
rect 300820 6168 300826 6180
rect 545758 6168 545764 6180
rect 300820 6140 545764 6168
rect 300820 6128 300826 6140
rect 545758 6128 545764 6140
rect 545816 6128 545822 6180
rect 481726 6060 481732 6112
rect 481784 6100 481790 6112
rect 569954 6100 569960 6112
rect 481784 6072 569960 6100
rect 481784 6060 481790 6072
rect 569954 6060 569960 6072
rect 570012 6060 570018 6112
rect 488810 5992 488816 6044
rect 488868 6032 488874 6044
rect 561306 6032 561312 6044
rect 488868 6004 561312 6032
rect 488868 5992 488874 6004
rect 561306 5992 561312 6004
rect 561364 5992 561370 6044
rect 527818 5924 527824 5976
rect 527876 5964 527882 5976
rect 566182 5964 566188 5976
rect 527876 5936 566188 5964
rect 527876 5924 527882 5936
rect 566182 5924 566188 5936
rect 566240 5924 566246 5976
rect 288434 5448 288440 5500
rect 288492 5488 288498 5500
rect 546862 5488 546868 5500
rect 288492 5460 546868 5488
rect 288492 5448 288498 5460
rect 546862 5448 546868 5460
rect 546920 5448 546926 5500
rect 299474 5380 299480 5432
rect 299532 5420 299538 5432
rect 547138 5420 547144 5432
rect 299532 5392 547144 5420
rect 299532 5380 299538 5392
rect 547138 5380 547144 5392
rect 547196 5380 547202 5432
rect 478138 4768 478144 4820
rect 478196 4808 478202 4820
rect 557902 4808 557908 4820
rect 478196 4780 557908 4808
rect 478196 4768 478202 4780
rect 557902 4768 557908 4780
rect 557960 4768 557966 4820
rect 574830 4224 574836 4276
rect 574888 4264 574894 4276
rect 577406 4264 577412 4276
rect 574888 4236 577412 4264
rect 574888 4224 574894 4236
rect 577406 4224 577412 4236
rect 577464 4224 577470 4276
rect 48222 4088 48228 4140
rect 48280 4128 48286 4140
rect 117590 4128 117596 4140
rect 48280 4100 117596 4128
rect 48280 4088 48286 4100
rect 117590 4088 117596 4100
rect 117648 4088 117654 4140
rect 495894 4088 495900 4140
rect 495952 4128 495958 4140
rect 556430 4128 556436 4140
rect 495952 4100 556436 4128
rect 495952 4088 495958 4100
rect 556430 4088 556436 4100
rect 556488 4088 556494 4140
rect 42150 4020 42156 4072
rect 42208 4060 42214 4072
rect 182542 4060 182548 4072
rect 42208 4032 182548 4060
rect 42208 4020 42214 4032
rect 182542 4020 182548 4032
rect 182600 4020 182606 4072
rect 492306 4020 492312 4072
rect 492364 4060 492370 4072
rect 553946 4060 553952 4072
rect 492364 4032 553952 4060
rect 492364 4020 492370 4032
rect 553946 4020 553952 4032
rect 554004 4020 554010 4072
rect 556154 4020 556160 4072
rect 556212 4060 556218 4072
rect 563330 4060 563336 4072
rect 556212 4032 563336 4060
rect 556212 4020 556218 4032
rect 563330 4020 563336 4032
rect 563388 4020 563394 4072
rect 46750 3952 46756 4004
rect 46808 3992 46814 4004
rect 189718 3992 189724 4004
rect 46808 3964 189724 3992
rect 46808 3952 46814 3964
rect 189718 3952 189724 3964
rect 189776 3952 189782 4004
rect 222746 3952 222752 4004
rect 222804 3992 222810 4004
rect 526438 3992 526444 4004
rect 222804 3964 526444 3992
rect 222804 3952 222810 3964
rect 526438 3952 526444 3964
rect 526496 3952 526502 4004
rect 549070 3952 549076 4004
rect 549128 3992 549134 4004
rect 573634 3992 573640 4004
rect 549128 3964 573640 3992
rect 549128 3952 549134 3964
rect 573634 3952 573640 3964
rect 573692 3952 573698 4004
rect 50430 3884 50436 3936
rect 50488 3924 50494 3936
rect 193214 3924 193220 3936
rect 50488 3896 193220 3924
rect 50488 3884 50494 3896
rect 193214 3884 193220 3896
rect 193272 3884 193278 3936
rect 212166 3884 212172 3936
rect 212224 3924 212230 3936
rect 533338 3924 533344 3936
rect 212224 3896 533344 3924
rect 212224 3884 212230 3896
rect 533338 3884 533344 3896
rect 533396 3884 533402 3936
rect 534902 3884 534908 3936
rect 534960 3924 534966 3936
rect 565354 3924 565360 3936
rect 534960 3896 565360 3924
rect 534960 3884 534966 3896
rect 565354 3884 565360 3896
rect 565412 3884 565418 3936
rect 41138 3816 41144 3868
rect 41196 3856 41202 3868
rect 196802 3856 196808 3868
rect 41196 3828 196808 3856
rect 41196 3816 41202 3828
rect 196802 3816 196808 3828
rect 196860 3816 196866 3868
rect 240502 3816 240508 3868
rect 240560 3856 240566 3868
rect 574186 3856 574192 3868
rect 240560 3828 574192 3856
rect 240560 3816 240566 3828
rect 574186 3816 574192 3828
rect 574244 3816 574250 3868
rect 42242 3748 42248 3800
rect 42300 3788 42306 3800
rect 161290 3788 161296 3800
rect 42300 3760 161296 3788
rect 42300 3748 42306 3760
rect 161290 3748 161296 3760
rect 161348 3748 161354 3800
rect 175458 3748 175464 3800
rect 175516 3788 175522 3800
rect 522298 3788 522304 3800
rect 175516 3760 522304 3788
rect 175516 3748 175522 3760
rect 522298 3748 522304 3760
rect 522356 3748 522362 3800
rect 524230 3748 524236 3800
rect 524288 3788 524294 3800
rect 570230 3788 570236 3800
rect 524288 3760 570236 3788
rect 524288 3748 524294 3760
rect 570230 3748 570236 3760
rect 570288 3748 570294 3800
rect 34330 3680 34336 3732
rect 34388 3720 34394 3732
rect 197906 3720 197912 3732
rect 34388 3692 197912 3720
rect 34388 3680 34394 3692
rect 197906 3680 197912 3692
rect 197964 3680 197970 3732
rect 552658 3680 552664 3732
rect 552716 3720 552722 3732
rect 561858 3720 561864 3732
rect 552716 3692 561864 3720
rect 552716 3680 552722 3692
rect 561858 3680 561864 3692
rect 561916 3680 561922 3732
rect 565814 3680 565820 3732
rect 565872 3720 565878 3732
rect 566274 3720 566280 3732
rect 565872 3692 566280 3720
rect 565872 3680 565878 3692
rect 566274 3680 566280 3692
rect 566332 3680 566338 3732
rect 34238 3612 34244 3664
rect 34296 3652 34302 3664
rect 215662 3652 215668 3664
rect 34296 3624 215668 3652
rect 34296 3612 34302 3624
rect 215662 3612 215668 3624
rect 215720 3612 215726 3664
rect 218146 3612 218152 3664
rect 218204 3652 218210 3664
rect 574646 3652 574652 3664
rect 218204 3624 574652 3652
rect 218204 3612 218210 3624
rect 574646 3612 574652 3624
rect 574704 3612 574710 3664
rect 37090 3544 37096 3596
rect 37148 3584 37154 3596
rect 184842 3584 184848 3596
rect 37148 3556 184848 3584
rect 37148 3544 37154 3556
rect 184842 3544 184848 3556
rect 184900 3544 184906 3596
rect 184934 3544 184940 3596
rect 184992 3584 184998 3596
rect 186130 3584 186136 3596
rect 184992 3556 186136 3584
rect 184992 3544 184998 3556
rect 186130 3544 186136 3556
rect 186188 3544 186194 3596
rect 190822 3544 190828 3596
rect 190880 3584 190886 3596
rect 576854 3584 576860 3596
rect 190880 3556 576860 3584
rect 190880 3544 190886 3556
rect 576854 3544 576860 3556
rect 576912 3544 576918 3596
rect 39758 3476 39764 3528
rect 39816 3516 39822 3528
rect 134150 3516 134156 3528
rect 39816 3488 134156 3516
rect 39816 3476 39822 3488
rect 134150 3476 134156 3488
rect 134208 3476 134214 3528
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 136450 3516 136456 3528
rect 135312 3488 136456 3516
rect 135312 3476 135318 3488
rect 136450 3476 136456 3488
rect 136508 3476 136514 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144730 3516 144736 3528
rect 143592 3488 144736 3516
rect 143592 3476 143598 3488
rect 144730 3476 144736 3488
rect 144788 3476 144794 3528
rect 144822 3476 144828 3528
rect 144880 3516 144886 3528
rect 568022 3516 568028 3528
rect 144880 3488 568028 3516
rect 144880 3476 144886 3488
rect 568022 3476 568028 3488
rect 568080 3476 568086 3528
rect 36722 3408 36728 3460
rect 36780 3448 36786 3460
rect 57238 3448 57244 3460
rect 36780 3420 57244 3448
rect 36780 3408 36786 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 92750 3408 92756 3460
rect 92808 3448 92814 3460
rect 549898 3448 549904 3460
rect 92808 3420 549904 3448
rect 92808 3408 92814 3420
rect 549898 3408 549904 3420
rect 549956 3408 549962 3460
rect 559742 3408 559748 3460
rect 559800 3448 559806 3460
rect 575658 3448 575664 3460
rect 559800 3420 575664 3448
rect 559800 3408 559806 3420
rect 575658 3408 575664 3420
rect 575716 3408 575722 3460
rect 53006 3340 53012 3392
rect 53064 3380 53070 3392
rect 96246 3380 96252 3392
rect 53064 3352 96252 3380
rect 53064 3340 53070 3352
rect 96246 3340 96252 3352
rect 96304 3340 96310 3392
rect 184842 3340 184848 3392
rect 184900 3380 184906 3392
rect 187326 3380 187332 3392
rect 184900 3352 187332 3380
rect 184900 3340 184906 3352
rect 187326 3340 187332 3352
rect 187384 3340 187390 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219250 3380 219256 3392
rect 218112 3352 219256 3380
rect 218112 3340 218118 3352
rect 219250 3340 219256 3352
rect 219308 3340 219314 3392
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 235810 3380 235816 3392
rect 234672 3352 235816 3380
rect 234672 3340 234678 3352
rect 235810 3340 235816 3352
rect 235868 3340 235874 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260650 3380 260656 3392
rect 259512 3352 260656 3380
rect 259512 3340 259518 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 510062 3340 510068 3392
rect 510120 3380 510126 3392
rect 565814 3380 565820 3392
rect 510120 3352 565820 3380
rect 510120 3340 510126 3352
rect 565814 3340 565820 3352
rect 565872 3340 565878 3392
rect 499390 3272 499396 3324
rect 499448 3312 499454 3324
rect 555050 3312 555056 3324
rect 499448 3284 555056 3312
rect 499448 3272 499454 3284
rect 555050 3272 555056 3284
rect 555108 3272 555114 3324
rect 578970 3272 578976 3324
rect 579028 3312 579034 3324
rect 582190 3312 582196 3324
rect 579028 3284 582196 3312
rect 579028 3272 579034 3284
rect 582190 3272 582196 3284
rect 582248 3272 582254 3324
rect 545482 3204 545488 3256
rect 545540 3244 545546 3256
rect 567378 3244 567384 3256
rect 545540 3216 567384 3244
rect 545540 3204 545546 3216
rect 567378 3204 567384 3216
rect 567436 3204 567442 3256
rect 200298 3136 200304 3188
rect 200356 3176 200362 3188
rect 552842 3176 552848 3188
rect 200356 3148 552848 3176
rect 200356 3136 200362 3148
rect 552842 3136 552848 3148
rect 552900 3136 552906 3188
rect 572070 3000 572076 3052
rect 572128 3040 572134 3052
rect 573910 3040 573916 3052
rect 572128 3012 573916 3040
rect 572128 3000 572134 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 143534 2796 143540 2848
rect 143592 2836 143598 2848
rect 144822 2836 144828 2848
rect 143592 2808 144828 2836
rect 143592 2796 143598 2808
rect 144822 2796 144828 2808
rect 144880 2796 144886 2848
rect 276106 1300 276112 1352
rect 276164 1340 276170 1352
rect 549622 1340 549628 1352
rect 276164 1312 549628 1340
rect 276164 1300 276170 1312
rect 549622 1300 549628 1312
rect 549680 1300 549686 1352
rect 233786 8 233792 60
rect 233844 48 233850 60
rect 545206 48 545212 60
rect 233844 20 545212 48
rect 233844 8 233850 20
rect 545206 8 545212 20
rect 545264 8 545270 60
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 484400 700680 484452 700732
rect 543464 700680 543516 700732
rect 283840 700612 283892 700664
rect 381544 700612 381596 700664
rect 400128 700612 400180 700664
rect 527180 700612 527232 700664
rect 218980 700544 219032 700596
rect 347228 700544 347280 700596
rect 413652 700544 413704 700596
rect 551284 700544 551336 700596
rect 105452 700476 105504 700528
rect 347136 700476 347188 700528
rect 405004 700476 405056 700528
rect 559656 700476 559708 700528
rect 202788 700408 202840 700460
rect 498200 700408 498252 700460
rect 267648 700340 267700 700392
rect 564716 700340 564768 700392
rect 24308 700272 24360 700324
rect 567200 700272 567252 700324
rect 137836 698912 137888 698964
rect 374828 698912 374880 698964
rect 429844 698912 429896 698964
rect 550916 698912 550968 698964
rect 153200 694764 153252 694816
rect 552940 694764 552992 694816
rect 71780 690616 71832 690668
rect 399944 690616 399996 690668
rect 462320 690616 462372 690668
rect 550272 690616 550324 690668
rect 331220 689324 331272 689376
rect 400864 689324 400916 689376
rect 364340 689256 364392 689308
rect 550364 689256 550416 689308
rect 299480 687964 299532 688016
rect 551100 687964 551152 688016
rect 234620 687896 234672 687948
rect 538220 687896 538272 687948
rect 405096 687488 405148 687540
rect 554136 687488 554188 687540
rect 403992 687420 404044 687472
rect 553952 687420 554004 687472
rect 396908 687352 396960 687404
rect 554228 687352 554280 687404
rect 407028 687284 407080 687336
rect 569960 687284 570012 687336
rect 413468 687216 413520 687268
rect 582380 687216 582432 687268
rect 347780 686536 347832 686588
rect 568764 686536 568816 686588
rect 6920 686468 6972 686520
rect 549996 686468 550048 686520
rect 384948 686128 385000 686180
rect 446404 686128 446456 686180
rect 407672 686060 407724 686112
rect 553768 686060 553820 686112
rect 402796 685992 402848 686044
rect 554044 685992 554096 686044
rect 363604 685924 363656 685976
rect 528836 685924 528888 685976
rect 405188 685856 405240 685908
rect 580908 685856 580960 685908
rect 402336 685516 402388 685568
rect 468392 685516 468444 685568
rect 407580 685448 407632 685500
rect 456800 685448 456852 685500
rect 173164 685380 173216 685432
rect 514760 685380 514812 685432
rect 409696 685312 409748 685364
rect 450268 685312 450320 685364
rect 409052 685244 409104 685296
rect 454224 685244 454276 685296
rect 407764 685176 407816 685228
rect 470876 685176 470928 685228
rect 407856 685108 407908 685160
rect 509240 685108 509292 685160
rect 468300 685040 468352 685092
rect 571340 685040 571392 685092
rect 362224 684972 362276 685024
rect 473544 684972 473596 685024
rect 487620 684972 487672 685024
rect 582472 684972 582524 685024
rect 359464 684904 359516 684956
rect 470600 684904 470652 684956
rect 476488 684904 476540 684956
rect 581092 684904 581144 684956
rect 409144 684836 409196 684888
rect 523040 684836 523092 684888
rect 453856 684768 453908 684820
rect 576860 684768 576912 684820
rect 409328 684700 409380 684752
rect 535460 684700 535512 684752
rect 406660 684632 406712 684684
rect 552480 684632 552532 684684
rect 388720 684564 388772 684616
rect 539140 684564 539192 684616
rect 405280 684496 405332 684548
rect 437572 684496 437624 684548
rect 489552 684496 489604 684548
rect 581000 684496 581052 684548
rect 21364 684020 21416 684072
rect 502524 684020 502576 684072
rect 409236 683952 409288 684004
rect 497280 683952 497332 684004
rect 400036 683884 400088 683936
rect 521844 683884 521896 683936
rect 407948 683816 408000 683868
rect 436100 683816 436152 683868
rect 438676 683816 438728 683868
rect 567936 683816 567988 683868
rect 429016 683748 429068 683800
rect 563704 683748 563756 683800
rect 392584 683680 392636 683732
rect 429660 683680 429712 683732
rect 435456 683680 435508 683732
rect 572812 683680 572864 683732
rect 408132 683612 408184 683664
rect 550640 683612 550692 683664
rect 398104 683544 398156 683596
rect 545580 683544 545632 683596
rect 404268 683476 404320 683528
rect 555240 683476 555292 683528
rect 416688 683408 416740 683460
rect 573640 683408 573692 683460
rect 408316 683340 408368 683392
rect 581184 683340 581236 683392
rect 406844 683272 406896 683324
rect 580356 683272 580408 683324
rect 31024 683204 31076 683256
rect 509516 683204 509568 683256
rect 409420 683136 409472 683188
rect 424600 683136 424652 683188
rect 510528 683136 510580 683188
rect 579160 683136 579212 683188
rect 3424 682660 3476 682712
rect 550456 682660 550508 682712
rect 529664 682592 529716 682644
rect 551468 682592 551520 682644
rect 26148 682524 26200 682576
rect 532700 682524 532752 682576
rect 495164 682456 495216 682508
rect 551560 682456 551612 682508
rect 402244 682388 402296 682440
rect 440424 682388 440476 682440
rect 477500 682388 477552 682440
rect 567292 682388 567344 682440
rect 382924 682320 382976 682372
rect 422392 682320 422444 682372
rect 502248 682320 502300 682372
rect 561036 682320 561088 682372
rect 389824 682252 389876 682304
rect 480352 682252 480404 682304
rect 484860 682252 484912 682304
rect 575480 682252 575532 682304
rect 397368 682184 397420 682236
rect 442264 682184 442316 682236
rect 458180 682184 458232 682236
rect 554872 682184 554924 682236
rect 373908 682116 373960 682168
rect 416596 682116 416648 682168
rect 432880 682116 432932 682168
rect 570604 682116 570656 682168
rect 408040 682048 408092 682100
rect 547788 682048 547840 682100
rect 549904 682048 549956 682100
rect 574100 682048 574152 682100
rect 384396 681980 384448 682032
rect 530124 681980 530176 682032
rect 537852 681980 537904 682032
rect 565912 681980 565964 682032
rect 380164 681912 380216 681964
rect 545120 681912 545172 681964
rect 548800 681912 548852 681964
rect 576952 681912 577004 681964
rect 409512 681844 409564 681896
rect 580448 681844 580500 681896
rect 17776 681776 17828 681828
rect 411628 681776 411680 681828
rect 512736 681776 512788 681828
rect 577228 681776 577280 681828
rect 389088 681708 389140 681760
rect 412916 681708 412968 681760
rect 440056 681708 440108 681760
rect 458180 681708 458232 681760
rect 541716 681708 541768 681760
rect 577504 681708 577556 681760
rect 8944 681300 8996 681352
rect 552112 681300 552164 681352
rect 406568 681232 406620 681284
rect 457352 681232 457404 681284
rect 501788 681232 501840 681284
rect 574744 681232 574796 681284
rect 377404 681164 377456 681216
rect 420000 681164 420052 681216
rect 427820 681164 427872 681216
rect 504364 681164 504416 681216
rect 517244 681164 517296 681216
rect 572904 681164 572956 681216
rect 403716 681096 403768 681148
rect 463792 681096 463844 681148
rect 499212 681096 499264 681148
rect 580264 681096 580316 681148
rect 408224 681028 408276 681080
rect 400956 680960 401008 681012
rect 427912 680960 427964 681012
rect 439320 681028 439372 681080
rect 440056 680960 440108 681012
rect 440332 681028 440384 681080
rect 524420 681028 524472 681080
rect 547788 681028 547840 681080
rect 555332 681028 555384 681080
rect 551008 680960 551060 681012
rect 347044 680892 347096 680944
rect 432052 680892 432104 680944
rect 434628 680892 434680 680944
rect 550732 680892 550784 680944
rect 409604 680824 409656 680876
rect 552388 680824 552440 680876
rect 408960 680756 409012 680808
rect 552204 680756 552256 680808
rect 409880 680688 409932 680740
rect 553492 680688 553544 680740
rect 403808 680620 403860 680672
rect 553400 680620 553452 680672
rect 405464 680552 405516 680604
rect 580632 680552 580684 680604
rect 402520 680484 402572 680536
rect 580724 680484 580776 680536
rect 173256 680416 173308 680468
rect 461216 680416 461268 680468
rect 496636 680416 496688 680468
rect 577136 680416 577188 680468
rect 427084 680348 427136 680400
rect 440148 680348 440200 680400
rect 402428 679600 402480 679652
rect 427084 679600 427136 679652
rect 440148 679600 440200 679652
rect 580540 679600 580592 679652
rect 399484 679532 399536 679584
rect 553676 679532 553728 679584
rect 409788 679464 409840 679516
rect 449808 679464 449860 679516
rect 511448 679464 511500 679516
rect 577044 679464 577096 679516
rect 408408 679396 408460 679448
rect 553124 679396 553176 679448
rect 406476 679328 406528 679380
rect 551928 679328 551980 679380
rect 405556 679260 405608 679312
rect 551192 679260 551244 679312
rect 404912 679192 404964 679244
rect 552572 679192 552624 679244
rect 402612 679124 402664 679176
rect 553860 679124 553912 679176
rect 552020 679056 552072 679108
rect 582840 679056 582892 679108
rect 395436 678988 395488 679040
rect 580816 678988 580868 679040
rect 408040 678512 408092 678564
rect 408316 678512 408368 678564
rect 407856 678376 407908 678428
rect 408040 678376 408092 678428
rect 399852 678240 399904 678292
rect 409880 678240 409932 678292
rect 407580 678172 407632 678224
rect 407764 678172 407816 678224
rect 552020 678104 552072 678156
rect 552296 678104 552348 678156
rect 7564 677560 7616 677612
rect 407120 677560 407172 677612
rect 552020 677560 552072 677612
rect 579620 677560 579672 677612
rect 40040 676812 40092 676864
rect 397000 676812 397052 676864
rect 551560 676540 551612 676592
rect 552756 676540 552808 676592
rect 166908 676132 166960 676184
rect 169760 676132 169812 676184
rect 340880 676132 340932 676184
rect 340880 674976 340932 675028
rect 351184 674976 351236 675028
rect 328552 674908 328604 674960
rect 347780 674908 347832 674960
rect 154488 674840 154540 674892
rect 172704 674840 172756 674892
rect 329748 674840 329800 674892
rect 361580 674840 361632 674892
rect 552020 674840 552072 674892
rect 575664 674840 575716 674892
rect 552204 674160 552256 674212
rect 550180 674092 550232 674144
rect 550456 674092 550508 674144
rect 550824 674092 550876 674144
rect 551376 674092 551428 674144
rect 552204 673956 552256 674008
rect 552020 672052 552072 672104
rect 571616 672052 571668 672104
rect 347228 670624 347280 670676
rect 407120 670624 407172 670676
rect 383016 667904 383068 667956
rect 407120 667904 407172 667956
rect 553308 666544 553360 666596
rect 566740 666544 566792 666596
rect 385684 665184 385736 665236
rect 407120 665184 407172 665236
rect 397460 663688 397512 663740
rect 407212 663688 407264 663740
rect 393964 661172 394016 661224
rect 407304 661172 407356 661224
rect 387248 661104 387300 661156
rect 407212 661104 407264 661156
rect 348792 661036 348844 661088
rect 407396 661036 407448 661088
rect 404728 658248 404780 658300
rect 407304 658248 407356 658300
rect 3332 658180 3384 658232
rect 8944 658180 8996 658232
rect 553308 656888 553360 656940
rect 558920 656888 558972 656940
rect 347136 655460 347188 655512
rect 407212 655460 407264 655512
rect 404084 654168 404136 654220
rect 407212 654168 407264 654220
rect 552112 653216 552164 653268
rect 554964 653216 555016 653268
rect 376024 652740 376076 652792
rect 407212 652740 407264 652792
rect 351184 650632 351236 650684
rect 402704 650632 402756 650684
rect 407212 650632 407264 650684
rect 367836 648592 367888 648644
rect 407212 648592 407264 648644
rect 553308 648592 553360 648644
rect 564532 648592 564584 648644
rect 552572 645872 552624 645924
rect 556436 645872 556488 645924
rect 553216 644648 553268 644700
rect 556804 644648 556856 644700
rect 402888 644444 402940 644496
rect 407212 644444 407264 644496
rect 552112 644444 552164 644496
rect 565268 644444 565320 644496
rect 570696 643084 570748 643136
rect 579988 643084 580040 643136
rect 552020 642540 552072 642592
rect 554228 642540 554280 642592
rect 347136 641724 347188 641776
rect 407212 641724 407264 641776
rect 358084 640296 358136 640348
rect 407212 640296 407264 640348
rect 553308 640296 553360 640348
rect 574284 640296 574336 640348
rect 552112 637848 552164 637900
rect 557816 637848 557868 637900
rect 404176 637644 404228 637696
rect 407304 637644 407356 637696
rect 393228 637576 393280 637628
rect 407212 637576 407264 637628
rect 552020 637576 552072 637628
rect 562600 637576 562652 637628
rect 383568 636216 383620 636268
rect 407212 636216 407264 636268
rect 408316 635536 408368 635588
rect 408316 635332 408368 635384
rect 367744 633428 367796 633480
rect 407212 633428 407264 633480
rect 360844 632068 360896 632120
rect 407212 632068 407264 632120
rect 556804 632000 556856 632052
rect 580172 632000 580224 632052
rect 552020 631184 552072 631236
rect 554228 631184 554280 631236
rect 408224 628600 408276 628652
rect 408408 628600 408460 628652
rect 395344 627920 395396 627972
rect 407212 627920 407264 627972
rect 552020 625336 552072 625388
rect 557080 625336 557132 625388
rect 552020 623772 552072 623824
rect 582656 623772 582708 623824
rect 552572 619624 552624 619676
rect 576124 619624 576176 619676
rect 396724 618332 396776 618384
rect 407304 618332 407356 618384
rect 387432 618264 387484 618316
rect 407212 618264 407264 618316
rect 553308 616836 553360 616888
rect 576308 616836 576360 616888
rect 371884 615476 371936 615528
rect 407304 615476 407356 615528
rect 553308 612824 553360 612876
rect 558552 612824 558604 612876
rect 399760 612756 399812 612808
rect 407212 612756 407264 612808
rect 553216 612756 553268 612808
rect 578884 612756 578936 612808
rect 553308 611328 553360 611380
rect 569408 611328 569460 611380
rect 553308 609968 553360 610020
rect 571984 609968 572036 610020
rect 350448 608608 350500 608660
rect 368480 608608 368532 608660
rect 381636 608608 381688 608660
rect 407212 608608 407264 608660
rect 552480 608608 552532 608660
rect 555700 608608 555752 608660
rect 552204 607248 552256 607300
rect 555056 607248 555108 607300
rect 176568 607180 176620 607232
rect 209044 607180 209096 607232
rect 176568 605820 176620 605872
rect 203524 605820 203576 605872
rect 350448 605820 350500 605872
rect 371240 605820 371292 605872
rect 350448 604460 350500 604512
rect 364340 604460 364392 604512
rect 552020 603916 552072 603968
rect 554872 603916 554924 603968
rect 553308 603100 553360 603152
rect 582564 603100 582616 603152
rect 404268 603032 404320 603084
rect 407304 603032 407356 603084
rect 366364 601672 366416 601724
rect 407304 601672 407356 601724
rect 174544 598952 174596 599004
rect 207020 598952 207072 599004
rect 374644 598952 374696 599004
rect 407304 598952 407356 599004
rect 553308 598952 553360 599004
rect 560484 598952 560536 599004
rect 394608 596164 394660 596216
rect 407304 596164 407356 596216
rect 398748 594804 398800 594856
rect 407304 594804 407356 594856
rect 34152 593512 34204 593564
rect 34336 593512 34388 593564
rect 404268 592016 404320 592068
rect 407304 592016 407356 592068
rect 404820 590860 404872 590912
rect 405188 590860 405240 590912
rect 405188 590724 405240 590776
rect 407396 590724 407448 590776
rect 401508 590656 401560 590708
rect 407304 590656 407356 590708
rect 34152 589976 34204 590028
rect 209136 589976 209188 590028
rect 34060 589908 34112 589960
rect 36452 589908 36504 589960
rect 33968 589840 34020 589892
rect 36544 589840 36596 589892
rect 47584 589228 47636 589280
rect 207756 589228 207808 589280
rect 239312 589228 239364 589280
rect 402336 589228 402388 589280
rect 39856 589160 39908 589212
rect 207664 589160 207716 589212
rect 225144 589160 225196 589212
rect 404912 589160 404964 589212
rect 140780 589092 140832 589144
rect 349344 589092 349396 589144
rect 35624 589024 35676 589076
rect 78864 589024 78916 589076
rect 86040 589024 86092 589076
rect 402612 589024 402664 589076
rect 39396 588956 39448 589008
rect 402428 588956 402480 589008
rect 552112 588956 552164 589008
rect 554136 588956 554188 589008
rect 42064 588888 42116 588940
rect 405280 588888 405332 588940
rect 40776 588820 40828 588872
rect 405096 588820 405148 588872
rect 40868 588752 40920 588804
rect 405556 588752 405608 588804
rect 35348 588684 35400 588736
rect 405188 588684 405240 588736
rect 32772 588616 32824 588668
rect 406752 588616 406804 588668
rect 3516 588548 3568 588600
rect 399668 588548 399720 588600
rect 43720 588480 43772 588532
rect 172704 588480 172756 588532
rect 292764 588480 292816 588532
rect 399484 588480 399536 588532
rect 317420 588412 317472 588464
rect 347780 588412 347832 588464
rect 393136 587868 393188 587920
rect 407304 587868 407356 587920
rect 44732 587528 44784 587580
rect 264428 587528 264480 587580
rect 42524 587460 42576 587512
rect 407304 587460 407356 587512
rect 57888 587392 57940 587444
rect 82084 587392 82136 587444
rect 49056 587324 49108 587376
rect 78680 587324 78732 587376
rect 316040 587324 316092 587376
rect 350540 587324 350592 587376
rect 33048 587256 33100 587308
rect 71780 587256 71832 587308
rect 308496 587256 308548 587308
rect 354772 587256 354824 587308
rect 37188 587188 37240 587240
rect 81900 587188 81952 587240
rect 291016 587188 291068 587240
rect 352012 587188 352064 587240
rect 45376 587120 45428 587172
rect 95240 587120 95292 587172
rect 286324 587120 286376 587172
rect 348424 587120 348476 587172
rect 34244 587052 34296 587104
rect 101956 587052 102008 587104
rect 281080 587052 281132 587104
rect 350632 587052 350684 587104
rect 22836 586984 22888 587036
rect 106924 586984 106976 587036
rect 261024 586984 261076 587036
rect 356520 586984 356572 587036
rect 45008 586916 45060 586968
rect 131764 586916 131816 586968
rect 248144 586916 248196 586968
rect 348700 586916 348752 586968
rect 41328 586848 41380 586900
rect 139400 586848 139452 586900
rect 141976 586848 142028 586900
rect 163964 586848 164016 586900
rect 256608 586848 256660 586900
rect 359280 586848 359332 586900
rect 22928 586780 22980 586832
rect 124404 586780 124456 586832
rect 124864 586780 124916 586832
rect 133972 586780 134024 586832
rect 153844 586780 153896 586832
rect 227812 586780 227864 586832
rect 240784 586780 240836 586832
rect 348516 586780 348568 586832
rect 77208 586712 77260 586764
rect 180064 586712 180116 586764
rect 209780 586712 209832 586764
rect 238760 586712 238812 586764
rect 242440 586712 242492 586764
rect 357716 586712 357768 586764
rect 245568 586644 245620 586696
rect 361856 586644 361908 586696
rect 48964 586576 49016 586628
rect 245844 586576 245896 586628
rect 260656 586576 260708 586628
rect 361764 586576 361816 586628
rect 31576 586508 31628 586560
rect 81164 586508 81216 586560
rect 333888 586508 333940 586560
rect 348608 586508 348660 586560
rect 553308 586508 553360 586560
rect 578976 586508 579028 586560
rect 273536 586032 273588 586084
rect 306932 586032 306984 586084
rect 47216 585964 47268 586016
rect 240508 585964 240560 586016
rect 265072 585964 265124 586016
rect 298100 585964 298152 586016
rect 320456 585964 320508 586016
rect 348792 585964 348844 586016
rect 81808 585896 81860 585948
rect 349712 585896 349764 585948
rect 66352 585828 66404 585880
rect 356428 585828 356480 585880
rect 100852 585760 100904 585812
rect 405372 585760 405424 585812
rect 200672 585148 200724 585200
rect 376116 585148 376168 585200
rect 552572 585148 552624 585200
rect 571432 585148 571484 585200
rect 215484 584604 215536 584656
rect 282920 584604 282972 584656
rect 307760 584604 307812 584656
rect 349160 584604 349212 584656
rect 115204 584536 115256 584588
rect 211620 584536 211672 584588
rect 269764 584536 269816 584588
rect 346860 584536 346912 584588
rect 79784 584468 79836 584520
rect 350724 584468 350776 584520
rect 40960 584400 41012 584452
rect 349252 584400 349304 584452
rect 377496 583720 377548 583772
rect 407304 583720 407356 583772
rect 552940 583720 552992 583772
rect 560392 583720 560444 583772
rect 43904 583040 43956 583092
rect 87144 583040 87196 583092
rect 159088 583040 159140 583092
rect 270224 583040 270276 583092
rect 84384 582972 84436 583024
rect 349620 582972 349672 583024
rect 243544 581884 243596 581936
rect 349252 581884 349304 581936
rect 147220 581816 147272 581868
rect 274640 581816 274692 581868
rect 87328 581748 87380 581800
rect 248420 581748 248472 581800
rect 46756 581680 46808 581732
rect 253940 581680 253992 581732
rect 109040 581612 109092 581664
rect 330116 581612 330168 581664
rect 209136 580456 209188 580508
rect 250444 580456 250496 580508
rect 160100 580388 160152 580440
rect 258172 580388 258224 580440
rect 297916 580388 297968 580440
rect 367836 580388 367888 580440
rect 46204 580320 46256 580372
rect 209780 580320 209832 580372
rect 245752 580320 245804 580372
rect 347136 580320 347188 580372
rect 99472 580252 99524 580304
rect 355140 580252 355192 580304
rect 383384 579640 383436 579692
rect 407304 579640 407356 579692
rect 171692 579096 171744 579148
rect 238852 579096 238904 579148
rect 208032 579028 208084 579080
rect 347964 579028 348016 579080
rect 46480 578960 46532 579012
rect 302240 578960 302292 579012
rect 35440 578892 35492 578944
rect 306288 578892 306340 578944
rect 111800 577600 111852 577652
rect 219992 577600 220044 577652
rect 231676 577600 231728 577652
rect 355048 577600 355100 577652
rect 107660 577532 107712 577584
rect 234620 577532 234672 577584
rect 246948 577532 247000 577584
rect 281816 577532 281868 577584
rect 41236 577464 41288 577516
rect 53840 577464 53892 577516
rect 74448 577464 74500 577516
rect 351092 577464 351144 577516
rect 553308 577192 553360 577244
rect 557632 577192 557684 577244
rect 388444 576852 388496 576904
rect 407304 576852 407356 576904
rect 150532 576240 150584 576292
rect 172612 576240 172664 576292
rect 244188 576240 244240 576292
rect 350816 576240 350868 576292
rect 49148 576172 49200 576224
rect 224960 576172 225012 576224
rect 238668 576172 238720 576224
rect 348240 576172 348292 576224
rect 43812 576104 43864 576156
rect 63592 576104 63644 576156
rect 89628 576104 89680 576156
rect 350356 576104 350408 576156
rect 550180 575968 550232 576020
rect 550456 575968 550508 576020
rect 403900 575492 403952 575544
rect 407304 575492 407356 575544
rect 553308 575492 553360 575544
rect 560668 575492 560720 575544
rect 117320 574948 117372 575000
rect 237380 574948 237432 575000
rect 45284 574880 45336 574932
rect 136640 574880 136692 574932
rect 209044 574880 209096 574932
rect 349896 574880 349948 574932
rect 62028 574812 62080 574864
rect 350908 574812 350960 574864
rect 3608 574744 3660 574796
rect 365076 574744 365128 574796
rect 403992 573996 404044 574048
rect 407304 573996 407356 574048
rect 552112 573996 552164 574048
rect 554044 573996 554096 574048
rect 163412 573656 163464 573708
rect 236000 573656 236052 573708
rect 85488 573588 85540 573640
rect 147956 573588 148008 573640
rect 160008 573588 160060 573640
rect 349344 573588 349396 573640
rect 46664 573520 46716 573572
rect 264980 573520 265032 573572
rect 97908 573452 97960 573504
rect 331496 573452 331548 573504
rect 35532 573384 35584 573436
rect 349160 573384 349212 573436
rect 52644 573316 52696 573368
rect 405004 573316 405056 573368
rect 403992 572704 404044 572756
rect 407304 572704 407356 572756
rect 551376 572704 551428 572756
rect 552020 572704 552072 572756
rect 209688 572160 209740 572212
rect 278688 572160 278740 572212
rect 45100 572092 45152 572144
rect 91100 572092 91152 572144
rect 155224 572092 155276 572144
rect 255320 572092 255372 572144
rect 86868 572024 86920 572076
rect 237380 572024 237432 572076
rect 268936 572024 268988 572076
rect 354956 572024 355008 572076
rect 45744 571956 45796 572008
rect 300860 571956 300912 572008
rect 366456 571344 366508 571396
rect 407304 571344 407356 571396
rect 207940 570868 207992 570920
rect 351000 570868 351052 570920
rect 208124 570800 208176 570852
rect 356152 570800 356204 570852
rect 208308 570732 208360 570784
rect 363144 570732 363196 570784
rect 47768 570664 47820 570716
rect 258080 570664 258132 570716
rect 263508 570664 263560 570716
rect 353300 570664 353352 570716
rect 67548 570596 67600 570648
rect 353852 570596 353904 570648
rect 266268 569508 266320 569560
rect 347780 569508 347832 569560
rect 252468 569440 252520 569492
rect 353760 569440 353812 569492
rect 234528 569372 234580 569424
rect 352380 569372 352432 569424
rect 231768 569304 231820 569356
rect 354864 569304 354916 569356
rect 122748 569236 122800 569288
rect 352472 569236 352524 569288
rect 117228 569168 117280 569220
rect 353392 569168 353444 569220
rect 272892 568896 272944 568948
rect 370504 568896 370556 568948
rect 234896 568828 234948 568880
rect 357624 568828 357676 568880
rect 244556 568760 244608 568812
rect 374000 568760 374052 568812
rect 222016 568692 222068 568744
rect 361672 568692 361724 568744
rect 217508 568624 217560 568676
rect 357440 568624 357492 568676
rect 35072 568556 35124 568608
rect 407304 568556 407356 568608
rect 552572 568556 552624 568608
rect 574192 568556 574244 568608
rect 296628 568148 296680 568200
rect 348148 568148 348200 568200
rect 269028 568080 269080 568132
rect 351184 568080 351236 568132
rect 249708 568012 249760 568064
rect 351920 568012 351972 568064
rect 267648 567944 267700 567996
rect 369952 567944 370004 567996
rect 233148 567876 233200 567928
rect 352196 567876 352248 567928
rect 43536 567808 43588 567860
rect 128360 567808 128412 567860
rect 208216 567808 208268 567860
rect 360384 567808 360436 567860
rect 254860 567536 254912 567588
rect 365168 567536 365220 567588
rect 243268 567468 243320 567520
rect 385960 567468 386012 567520
rect 140228 567400 140280 567452
rect 359556 567400 359608 567452
rect 131212 567332 131264 567384
rect 353944 567332 353996 567384
rect 375104 567332 375156 567384
rect 407304 567332 407356 567384
rect 143448 567264 143500 567316
rect 384488 567264 384540 567316
rect 553308 567264 553360 567316
rect 560576 567264 560628 567316
rect 116400 567196 116452 567248
rect 401048 567196 401100 567248
rect 552480 567196 552532 567248
rect 563336 567196 563388 567248
rect 293868 566720 293920 566772
rect 350264 566720 350316 566772
rect 45928 566652 45980 566704
rect 174544 566652 174596 566704
rect 262036 566652 262088 566704
rect 348056 566652 348108 566704
rect 82084 566584 82136 566636
rect 226892 566584 226944 566636
rect 257988 566584 258040 566636
rect 349528 566584 349580 566636
rect 47032 566516 47084 566568
rect 118700 566516 118752 566568
rect 128268 566516 128320 566568
rect 359188 566516 359240 566568
rect 104808 566448 104860 566500
rect 349436 566448 349488 566500
rect 317788 566380 317840 566432
rect 367192 566380 367244 566432
rect 314936 566312 314988 566364
rect 373264 566312 373316 566364
rect 275008 566244 275060 566296
rect 392676 566244 392728 566296
rect 240968 566176 241020 566228
rect 358820 566176 358872 566228
rect 198464 566108 198516 566160
rect 357164 566108 357216 566160
rect 20628 566040 20680 566092
rect 121552 566040 121604 566092
rect 217048 566040 217100 566092
rect 381728 566040 381780 566092
rect 36820 565972 36872 566024
rect 376484 565972 376536 566024
rect 32588 565904 32640 565956
rect 405096 565904 405148 565956
rect 3240 565836 3292 565888
rect 17224 565836 17276 565888
rect 31300 565836 31352 565888
rect 405004 565836 405056 565888
rect 25964 565564 26016 565616
rect 311164 565564 311216 565616
rect 130752 565496 130804 565548
rect 353576 565496 353628 565548
rect 203524 565428 203576 565480
rect 243452 565428 243504 565480
rect 32956 565360 33008 565412
rect 93860 565360 93912 565412
rect 135904 565360 135956 565412
rect 252560 565360 252612 565412
rect 45192 565292 45244 565344
rect 175372 565292 175424 565344
rect 180064 565292 180116 565344
rect 225420 565292 225472 565344
rect 230388 565292 230440 565344
rect 310520 565292 310572 565344
rect 44640 565224 44692 565276
rect 78772 565224 78824 565276
rect 91008 565224 91060 565276
rect 253940 565224 253992 565276
rect 333796 565224 333848 565276
rect 347872 565224 347924 565276
rect 64788 565156 64840 565208
rect 249800 565156 249852 565208
rect 324688 565156 324740 565208
rect 354680 565156 354732 565208
rect 77116 565088 77168 565140
rect 295708 565088 295760 565140
rect 315948 565088 316000 565140
rect 374736 565088 374788 565140
rect 265992 565020 266044 565072
rect 358912 565020 358964 565072
rect 23388 564952 23440 565004
rect 82820 564952 82872 565004
rect 263416 564952 263468 565004
rect 360200 564952 360252 565004
rect 42432 564884 42484 564936
rect 104348 564884 104400 564936
rect 238668 564884 238720 564936
rect 360292 564884 360344 564936
rect 36912 564816 36964 564868
rect 111892 564816 111944 564868
rect 251824 564816 251876 564868
rect 379152 564816 379204 564868
rect 39304 564748 39356 564800
rect 168564 564748 168616 564800
rect 269856 564748 269908 564800
rect 399576 564748 399628 564800
rect 38108 564680 38160 564732
rect 191380 564680 191432 564732
rect 232504 564680 232556 564732
rect 368664 564680 368716 564732
rect 33968 564612 34020 564664
rect 244740 564612 244792 564664
rect 248328 564612 248380 564664
rect 396816 564612 396868 564664
rect 40592 564544 40644 564596
rect 124956 564544 125008 564596
rect 340144 564544 340196 564596
rect 383108 564544 383160 564596
rect 298928 564476 298980 564528
rect 402428 564476 402480 564528
rect 41052 564408 41104 564460
rect 382188 564408 382240 564460
rect 405556 564408 405608 564460
rect 407396 564408 407448 564460
rect 31392 564068 31444 564120
rect 339132 564068 339184 564120
rect 23204 564000 23256 564052
rect 255780 564000 255832 564052
rect 24308 563932 24360 563984
rect 56600 563932 56652 563984
rect 327816 563932 327868 563984
rect 352840 563932 352892 563984
rect 41880 563864 41932 563916
rect 74632 563864 74684 563916
rect 204168 563864 204220 563916
rect 247040 563864 247092 563916
rect 264888 563864 264940 563916
rect 343732 563864 343784 563916
rect 44824 563796 44876 563848
rect 88340 563796 88392 563848
rect 153936 563796 153988 563848
rect 175464 563796 175516 563848
rect 179696 563796 179748 563848
rect 262220 563796 262272 563848
rect 299388 563796 299440 563848
rect 389916 563796 389968 563848
rect 40684 563728 40736 563780
rect 87052 563728 87104 563780
rect 95148 563728 95200 563780
rect 222200 563728 222252 563780
rect 224776 563728 224828 563780
rect 355324 563728 355376 563780
rect 46388 563660 46440 563712
rect 175280 563660 175332 563712
rect 208032 563660 208084 563712
rect 353668 563660 353720 563712
rect 224224 563592 224276 563644
rect 398288 563592 398340 563644
rect 43444 563524 43496 563576
rect 162308 563524 162360 563576
rect 180708 563524 180760 563576
rect 378784 563524 378836 563576
rect 179144 563456 179196 563508
rect 385776 563456 385828 563508
rect 39212 563388 39264 563440
rect 181076 563388 181128 563440
rect 249708 563388 249760 563440
rect 389180 563388 389232 563440
rect 22008 563320 22060 563372
rect 301412 563320 301464 563372
rect 307668 563320 307720 563372
rect 402336 563320 402388 563372
rect 24768 563252 24820 563304
rect 325976 563252 326028 563304
rect 338764 563252 338816 563304
rect 365720 563252 365772 563304
rect 336648 563184 336700 563236
rect 364432 563184 364484 563236
rect 38476 563116 38528 563168
rect 401140 563116 401192 563168
rect 31116 563048 31168 563100
rect 395528 563048 395580 563100
rect 48228 562980 48280 563032
rect 49148 562980 49200 563032
rect 23020 562708 23072 562760
rect 113456 562708 113508 562760
rect 203616 562708 203668 562760
rect 340788 562708 340840 562760
rect 43352 562640 43404 562692
rect 405188 562640 405240 562692
rect 23112 562572 23164 562624
rect 65708 562572 65760 562624
rect 73068 562572 73120 562624
rect 91284 562572 91336 562624
rect 338028 562572 338080 562624
rect 347044 562572 347096 562624
rect 75828 562504 75880 562556
rect 124864 562504 124916 562556
rect 214472 562504 214524 562556
rect 249708 562504 249760 562556
rect 304080 562504 304132 562556
rect 369124 562504 369176 562556
rect 39764 562436 39816 562488
rect 81624 562436 81676 562488
rect 82820 562436 82872 562488
rect 148140 562436 148192 562488
rect 208768 562436 208820 562488
rect 338764 562436 338816 562488
rect 37004 562368 37056 562420
rect 83740 562368 83792 562420
rect 90824 562368 90876 562420
rect 173164 562368 173216 562420
rect 186872 562368 186924 562420
rect 335360 562368 335412 562420
rect 339132 562368 339184 562420
rect 382004 562368 382056 562420
rect 552020 562368 552072 562420
rect 556620 562368 556672 562420
rect 47400 562300 47452 562352
rect 74540 562300 74592 562352
rect 76656 562300 76708 562352
rect 173256 562300 173308 562352
rect 226800 562300 226852 562352
rect 406568 562300 406620 562352
rect 35532 562232 35584 562284
rect 94780 562232 94832 562284
rect 278320 562232 278372 562284
rect 346492 562232 346544 562284
rect 40500 562164 40552 562216
rect 99380 562164 99432 562216
rect 236368 562164 236420 562216
rect 336372 562164 336424 562216
rect 347688 562164 347740 562216
rect 378876 562164 378928 562216
rect 38384 562096 38436 562148
rect 105084 562096 105136 562148
rect 260288 562096 260340 562148
rect 367928 562096 367980 562148
rect 27436 562028 27488 562080
rect 51540 562028 51592 562080
rect 51632 562028 51684 562080
rect 138020 562028 138072 562080
rect 250444 562028 250496 562080
rect 372068 562028 372120 562080
rect 32864 561960 32916 562012
rect 138572 561960 138624 562012
rect 336280 561960 336332 562012
rect 381820 561960 381872 562012
rect 42340 561892 42392 561944
rect 193864 561892 193916 561944
rect 201408 561892 201460 561944
rect 366548 561892 366600 561944
rect 51080 561824 51132 561876
rect 181628 561824 181680 561876
rect 184848 561824 184900 561876
rect 368572 561824 368624 561876
rect 110144 561756 110196 561808
rect 391480 561756 391532 561808
rect 19156 561688 19208 561740
rect 50252 561688 50304 561740
rect 337568 561688 337620 561740
rect 346400 561688 346452 561740
rect 32680 561620 32732 561672
rect 407304 561620 407356 561672
rect 47124 561552 47176 561604
rect 67640 561552 67692 561604
rect 25688 561484 25740 561536
rect 52460 561484 52512 561536
rect 35440 561416 35492 561468
rect 63684 561416 63736 561468
rect 47308 561348 47360 561400
rect 77300 561348 77352 561400
rect 38200 561280 38252 561332
rect 69020 561280 69072 561332
rect 27160 561212 27212 561264
rect 59360 561212 59412 561264
rect 37096 561144 37148 561196
rect 70400 561144 70452 561196
rect 30012 561076 30064 561128
rect 63500 561076 63552 561128
rect 313096 561076 313148 561128
rect 352564 561076 352616 561128
rect 38292 561008 38344 561060
rect 83004 561008 83056 561060
rect 305920 561008 305972 561060
rect 364984 561008 365036 561060
rect 39488 560940 39540 560992
rect 86960 560940 87012 560992
rect 291200 560940 291252 560992
rect 352288 560940 352340 560992
rect 47492 560872 47544 560924
rect 62120 560872 62172 560924
rect 287888 560872 287940 560924
rect 382280 560872 382332 560924
rect 255688 560804 255740 560856
rect 359004 560804 359056 560856
rect 233792 560736 233844 560788
rect 351276 560736 351328 560788
rect 235816 560668 235868 560720
rect 399484 560668 399536 560720
rect 146208 560600 146260 560652
rect 352656 560600 352708 560652
rect 183008 560532 183060 560584
rect 403624 560532 403676 560584
rect 62488 560464 62540 560516
rect 392768 560464 392820 560516
rect 43628 560396 43680 560448
rect 405280 560396 405332 560448
rect 44088 560328 44140 560380
rect 407764 560328 407816 560380
rect 552940 560328 552992 560380
rect 569224 560328 569276 560380
rect 325608 560260 325660 560312
rect 357532 560260 357584 560312
rect 553308 560260 553360 560312
rect 582748 560260 582800 560312
rect 46848 560192 46900 560244
rect 49056 560192 49108 560244
rect 49608 560192 49660 560244
rect 59176 560192 59228 560244
rect 46572 560124 46624 560176
rect 48872 560124 48924 560176
rect 36636 559512 36688 559564
rect 39672 558900 39724 558952
rect 148876 559920 148928 559972
rect 277032 559920 277084 559972
rect 294788 560056 294840 560108
rect 294788 559920 294840 559972
rect 334992 559920 335044 559972
rect 339408 559920 339460 559972
rect 346492 559988 346544 560040
rect 348332 559988 348384 560040
rect 340696 559920 340748 559972
rect 340788 559920 340840 559972
rect 346400 559920 346452 559972
rect 347688 559852 347740 559904
rect 360568 559648 360620 559700
rect 347688 559580 347740 559632
rect 407948 559580 408000 559632
rect 348332 559512 348384 559564
rect 407580 559512 407632 559564
rect 347688 559444 347740 559496
rect 365812 559036 365864 559088
rect 347688 558968 347740 559020
rect 391296 558968 391348 559020
rect 352104 558900 352156 558952
rect 349436 558152 349488 558204
rect 349804 558152 349856 558204
rect 552940 557608 552992 557660
rect 561864 557608 561916 557660
rect 553308 557540 553360 557592
rect 568672 557540 568724 557592
rect 552020 556520 552072 556572
rect 554872 556520 554924 556572
rect 44548 556180 44600 556232
rect 46296 556180 46348 556232
rect 349436 554684 349488 554736
rect 351920 554684 351972 554736
rect 552020 553800 552072 553852
rect 553952 553800 554004 553852
rect 398564 552032 398616 552084
rect 407304 552032 407356 552084
rect 552388 552032 552440 552084
rect 579712 552032 579764 552084
rect 405280 551964 405332 552016
rect 407396 551964 407448 552016
rect 42708 551080 42760 551132
rect 46296 551080 46348 551132
rect 41144 550808 41196 550860
rect 46296 550808 46348 550860
rect 553308 550808 553360 550860
rect 559472 550808 559524 550860
rect 350448 550604 350500 550656
rect 388536 550604 388588 550656
rect 398656 550604 398708 550656
rect 407304 550604 407356 550656
rect 42616 549244 42668 549296
rect 46296 549244 46348 549296
rect 358268 549244 358320 549296
rect 407304 549244 407356 549296
rect 553308 549244 553360 549296
rect 575572 549244 575624 549296
rect 46112 549108 46164 549160
rect 46296 549108 46348 549160
rect 350172 546524 350224 546576
rect 366640 546524 366692 546576
rect 377588 546524 377640 546576
rect 407304 546524 407356 546576
rect 30196 546456 30248 546508
rect 46112 546456 46164 546508
rect 350448 546456 350500 546508
rect 388628 546456 388680 546508
rect 553308 546456 553360 546508
rect 560760 546456 560812 546508
rect 551468 545300 551520 545352
rect 552020 545300 552072 545352
rect 34060 545096 34112 545148
rect 46020 545096 46072 545148
rect 405372 543804 405424 543856
rect 407396 543804 407448 543856
rect 43168 543736 43220 543788
rect 46112 543736 46164 543788
rect 377680 543736 377732 543788
rect 407304 543736 407356 543788
rect 553308 543736 553360 543788
rect 561956 543736 562008 543788
rect 350448 542376 350500 542428
rect 363788 542376 363840 542428
rect 353944 542308 353996 542360
rect 407304 542308 407356 542360
rect 21916 540948 21968 541000
rect 46112 540948 46164 541000
rect 552572 539588 552624 539640
rect 567384 539588 567436 539640
rect 350448 538228 350500 538280
rect 367836 538228 367888 538280
rect 552572 538228 552624 538280
rect 559564 538228 559616 538280
rect 44088 538160 44140 538212
rect 46112 538160 46164 538212
rect 350448 536800 350500 536852
rect 372620 536800 372672 536852
rect 553308 535848 553360 535900
rect 559380 535848 559432 535900
rect 552388 534148 552440 534200
rect 570144 534148 570196 534200
rect 350448 534080 350500 534132
rect 380256 534080 380308 534132
rect 394148 534080 394200 534132
rect 407304 534080 407356 534132
rect 553308 534080 553360 534132
rect 581552 534080 581604 534132
rect 550180 533332 550232 533384
rect 550456 533332 550508 533384
rect 350172 532788 350224 532840
rect 359096 532788 359148 532840
rect 350448 532720 350500 532772
rect 381912 532720 381964 532772
rect 552020 532516 552072 532568
rect 553768 532516 553820 532568
rect 43076 531768 43128 531820
rect 46020 531768 46072 531820
rect 349436 531292 349488 531344
rect 351368 531292 351420 531344
rect 552020 530884 552072 530936
rect 553860 530884 553912 530936
rect 39028 529932 39080 529984
rect 46112 529932 46164 529984
rect 350448 529932 350500 529984
rect 380440 529932 380492 529984
rect 552664 529932 552716 529984
rect 563428 529932 563480 529984
rect 42248 528572 42300 528624
rect 45836 528572 45888 528624
rect 370596 528572 370648 528624
rect 407304 528572 407356 528624
rect 350448 527144 350500 527196
rect 376300 527144 376352 527196
rect 553308 527144 553360 527196
rect 564808 527144 564860 527196
rect 552020 526056 552072 526108
rect 553768 526056 553820 526108
rect 350448 525920 350500 525972
rect 356704 525920 356756 525972
rect 44732 525716 44784 525768
rect 46112 525716 46164 525768
rect 552020 525716 552072 525768
rect 553676 525716 553728 525768
rect 571984 525716 572036 525768
rect 579804 525716 579856 525768
rect 40776 525648 40828 525700
rect 45652 525648 45704 525700
rect 402612 525036 402664 525088
rect 407304 525036 407356 525088
rect 390376 524424 390428 524476
rect 407396 524424 407448 524476
rect 387340 523064 387392 523116
rect 407304 523064 407356 523116
rect 350448 522996 350500 523048
rect 378968 522996 379020 523048
rect 399944 522928 399996 522980
rect 407304 522928 407356 522980
rect 401232 521704 401284 521756
rect 407396 521704 407448 521756
rect 350080 521160 350132 521212
rect 352104 521160 352156 521212
rect 23296 520276 23348 520328
rect 46204 520276 46256 520328
rect 373540 520276 373592 520328
rect 407304 520276 407356 520328
rect 552020 520276 552072 520328
rect 571524 520276 571576 520328
rect 552020 519256 552072 519308
rect 553676 519256 553728 519308
rect 552020 518916 552072 518968
rect 564624 518916 564676 518968
rect 398472 517556 398524 517608
rect 407304 517556 407356 517608
rect 350448 517488 350500 517540
rect 383200 517488 383252 517540
rect 388996 517488 389048 517540
rect 407396 517488 407448 517540
rect 350448 516264 350500 516316
rect 367100 516264 367152 516316
rect 350080 516196 350132 516248
rect 384672 516196 384724 516248
rect 394516 516196 394568 516248
rect 407304 516196 407356 516248
rect 40408 516128 40460 516180
rect 46020 516128 46072 516180
rect 358176 516128 358228 516180
rect 407396 516128 407448 516180
rect 552020 516128 552072 516180
rect 570880 516128 570932 516180
rect 405188 516060 405240 516112
rect 407672 516060 407724 516112
rect 552020 514768 552072 514820
rect 567568 514768 567620 514820
rect 350080 513408 350132 513460
rect 354128 513408 354180 513460
rect 42156 513340 42208 513392
rect 45928 513340 45980 513392
rect 350448 513340 350500 513392
rect 368020 513340 368072 513392
rect 374828 513272 374880 513324
rect 407304 513272 407356 513324
rect 373448 511980 373500 512032
rect 407304 511980 407356 512032
rect 350448 511912 350500 511964
rect 353300 511912 353352 511964
rect 43996 510552 44048 510604
rect 46112 510552 46164 510604
rect 553308 509872 553360 509924
rect 559104 509872 559156 509924
rect 40500 509260 40552 509312
rect 46020 509260 46072 509312
rect 385868 509260 385920 509312
rect 407304 509260 407356 509312
rect 350448 509192 350500 509244
rect 399852 509192 399904 509244
rect 359556 509124 359608 509176
rect 407304 509124 407356 509176
rect 349988 506540 350040 506592
rect 352104 506540 352156 506592
rect 27528 506472 27580 506524
rect 46112 506472 46164 506524
rect 349896 506472 349948 506524
rect 351276 506472 351328 506524
rect 359556 506472 359608 506524
rect 407304 506472 407356 506524
rect 350448 506404 350500 506456
rect 403808 506404 403860 506456
rect 553124 506404 553176 506456
rect 570696 506404 570748 506456
rect 21824 505112 21876 505164
rect 46112 505112 46164 505164
rect 350080 505112 350132 505164
rect 380624 505112 380676 505164
rect 553308 505112 553360 505164
rect 572996 505112 573048 505164
rect 350448 503684 350500 503736
rect 360476 503684 360528 503736
rect 553308 503684 553360 503736
rect 566280 503684 566332 503736
rect 553308 502392 553360 502444
rect 559012 502392 559064 502444
rect 39396 501848 39448 501900
rect 46112 501848 46164 501900
rect 553124 501032 553176 501084
rect 566188 501032 566240 501084
rect 397276 500964 397328 501016
rect 407304 500964 407356 501016
rect 553308 500964 553360 501016
rect 572076 500964 572128 501016
rect 39856 500896 39908 500948
rect 45652 500896 45704 500948
rect 402152 500896 402204 500948
rect 407396 500896 407448 500948
rect 553308 499808 553360 499860
rect 557724 499808 557776 499860
rect 350448 499536 350500 499588
rect 380532 499536 380584 499588
rect 348700 498516 348752 498568
rect 349160 498516 349212 498568
rect 45928 498244 45980 498296
rect 46480 498244 46532 498296
rect 350448 498176 350500 498228
rect 355232 498176 355284 498228
rect 553308 498176 553360 498228
rect 577320 498176 577372 498228
rect 42064 498108 42116 498160
rect 46480 498108 46532 498160
rect 41052 496748 41104 496800
rect 46480 496748 46532 496800
rect 552204 496544 552256 496596
rect 555332 496544 555384 496596
rect 21732 495456 21784 495508
rect 46112 495456 46164 495508
rect 350448 495456 350500 495508
rect 387524 495456 387576 495508
rect 391848 495456 391900 495508
rect 407304 495456 407356 495508
rect 553308 495456 553360 495508
rect 563612 495456 563664 495508
rect 42524 495388 42576 495440
rect 46480 495388 46532 495440
rect 350448 494504 350500 494556
rect 355416 494504 355468 494556
rect 348608 493960 348660 494012
rect 349436 493960 349488 494012
rect 24216 492668 24268 492720
rect 46480 492668 46532 492720
rect 360936 492668 360988 492720
rect 407304 492668 407356 492720
rect 552572 492668 552624 492720
rect 581460 492668 581512 492720
rect 348976 491648 349028 491700
rect 349896 491648 349948 491700
rect 350356 491376 350408 491428
rect 353484 491376 353536 491428
rect 350448 491308 350500 491360
rect 372436 491308 372488 491360
rect 350356 491240 350408 491292
rect 352288 491240 352340 491292
rect 350448 489948 350500 490000
rect 374828 489948 374880 490000
rect 28632 489880 28684 489932
rect 46480 489880 46532 489932
rect 362316 489880 362368 489932
rect 407304 489880 407356 489932
rect 348516 488860 348568 488912
rect 349620 488860 349672 488912
rect 553308 488792 553360 488844
rect 559196 488792 559248 488844
rect 391756 488520 391808 488572
rect 407304 488520 407356 488572
rect 350448 488452 350500 488504
rect 387432 488452 387484 488504
rect 39212 487772 39264 487824
rect 45652 487772 45704 487824
rect 395988 487160 396040 487212
rect 407304 487160 407356 487212
rect 553308 487160 553360 487212
rect 573088 487160 573140 487212
rect 46480 486072 46532 486124
rect 46756 486072 46808 486124
rect 19248 485800 19300 485852
rect 46756 485800 46808 485852
rect 386328 485800 386380 485852
rect 407304 485800 407356 485852
rect 405464 485732 405516 485784
rect 407488 485732 407540 485784
rect 552848 484576 552900 484628
rect 556252 484576 556304 484628
rect 42064 484440 42116 484492
rect 46756 484440 46808 484492
rect 19064 484372 19116 484424
rect 45836 484372 45888 484424
rect 349988 484372 350040 484424
rect 352288 484372 352340 484424
rect 370688 484372 370740 484424
rect 407304 484372 407356 484424
rect 551284 484304 551336 484356
rect 552020 484304 552072 484356
rect 379060 483080 379112 483132
rect 407304 483080 407356 483132
rect 350448 483012 350500 483064
rect 386052 483012 386104 483064
rect 406016 483012 406068 483064
rect 407856 483012 407908 483064
rect 552572 483012 552624 483064
rect 575756 483012 575808 483064
rect 350448 481652 350500 481704
rect 367284 481652 367336 481704
rect 384856 481652 384908 481704
rect 407304 481652 407356 481704
rect 45008 481312 45060 481364
rect 46480 481312 46532 481364
rect 40960 480632 41012 480684
rect 46296 480632 46348 480684
rect 350080 480292 350132 480344
rect 362960 480292 363012 480344
rect 38568 480224 38620 480276
rect 46756 480224 46808 480276
rect 350448 480224 350500 480276
rect 368756 480224 368808 480276
rect 553308 478864 553360 478916
rect 577412 478864 577464 478916
rect 401416 477504 401468 477556
rect 407304 477504 407356 477556
rect 552572 477504 552624 477556
rect 563980 477504 564032 477556
rect 350080 476144 350132 476196
rect 364524 476144 364576 476196
rect 350448 476076 350500 476128
rect 377772 476076 377824 476128
rect 363880 474784 363932 474836
rect 407304 474784 407356 474836
rect 553308 474784 553360 474836
rect 563152 474784 563204 474836
rect 552940 474716 552992 474768
rect 582932 474716 582984 474768
rect 43352 474648 43404 474700
rect 46756 474648 46808 474700
rect 390468 473424 390520 473476
rect 407304 473424 407356 473476
rect 350448 473356 350500 473408
rect 356244 473356 356296 473408
rect 372252 473356 372304 473408
rect 407396 473356 407448 473408
rect 384764 471996 384816 472048
rect 407304 471996 407356 472048
rect 553308 470568 553360 470620
rect 567844 470568 567896 470620
rect 570788 470568 570840 470620
rect 580172 470568 580224 470620
rect 37648 469208 37700 469260
rect 46756 469208 46808 469260
rect 365260 469208 365312 469260
rect 407304 469208 407356 469260
rect 553308 469208 553360 469260
rect 578332 469208 578384 469260
rect 39396 467916 39448 467968
rect 46756 467916 46808 467968
rect 21640 467848 21692 467900
rect 46664 467848 46716 467900
rect 386236 467848 386288 467900
rect 407304 467848 407356 467900
rect 350448 466420 350500 466472
rect 391204 466420 391256 466472
rect 553308 466420 553360 466472
rect 567660 466420 567712 466472
rect 350080 466352 350132 466404
rect 396908 466352 396960 466404
rect 350448 465060 350500 465112
rect 371332 465060 371384 465112
rect 401324 465060 401376 465112
rect 407304 465060 407356 465112
rect 552020 465060 552072 465112
rect 574468 465060 574520 465112
rect 40960 464108 41012 464160
rect 46756 464108 46808 464160
rect 552020 463904 552072 463956
rect 556344 463904 556396 463956
rect 21548 463700 21600 463752
rect 46756 463700 46808 463752
rect 383292 463700 383344 463752
rect 407304 463700 407356 463752
rect 36820 463632 36872 463684
rect 46664 463632 46716 463684
rect 350080 462408 350132 462460
rect 369216 462408 369268 462460
rect 403808 462408 403860 462460
rect 407396 462408 407448 462460
rect 3516 462340 3568 462392
rect 19984 462340 20036 462392
rect 350448 462340 350500 462392
rect 386144 462340 386196 462392
rect 396908 462340 396960 462392
rect 407304 462340 407356 462392
rect 552020 462340 552072 462392
rect 574652 462340 574704 462392
rect 350448 460980 350500 461032
rect 363052 460980 363104 461032
rect 24584 460912 24636 460964
rect 46756 460912 46808 460964
rect 350080 460912 350132 460964
rect 371424 460912 371476 460964
rect 38476 460844 38528 460896
rect 46664 460844 46716 460896
rect 552204 459620 552256 459672
rect 573272 459620 573324 459672
rect 350448 459552 350500 459604
rect 373816 459552 373868 459604
rect 552020 459552 552072 459604
rect 581276 459552 581328 459604
rect 552020 459008 552072 459060
rect 553952 459008 554004 459060
rect 551284 458328 551336 458380
rect 553032 458328 553084 458380
rect 402704 458192 402756 458244
rect 407304 458192 407356 458244
rect 350448 457240 350500 457292
rect 356336 457240 356388 457292
rect 372344 456764 372396 456816
rect 407304 456764 407356 456816
rect 552020 456764 552072 456816
rect 576216 456764 576268 456816
rect 43628 456696 43680 456748
rect 46664 456696 46716 456748
rect 387524 456696 387576 456748
rect 407396 456696 407448 456748
rect 40868 456628 40920 456680
rect 46756 456628 46808 456680
rect 552020 456288 552072 456340
rect 553860 456288 553912 456340
rect 349068 456084 349120 456136
rect 352012 456084 352064 456136
rect 379152 455336 379204 455388
rect 407396 455336 407448 455388
rect 350448 454112 350500 454164
rect 380808 454112 380860 454164
rect 375288 454044 375340 454096
rect 407304 454044 407356 454096
rect 552480 454044 552532 454096
rect 566004 454044 566056 454096
rect 405464 452616 405516 452668
rect 407672 452616 407724 452668
rect 552572 452616 552624 452668
rect 559288 452616 559340 452668
rect 377864 451324 377916 451376
rect 407304 451324 407356 451376
rect 350448 451256 350500 451308
rect 380348 451256 380400 451308
rect 32588 451188 32640 451240
rect 46756 451188 46808 451240
rect 350448 451120 350500 451172
rect 353760 451120 353812 451172
rect 350448 449896 350500 449948
rect 374552 449896 374604 449948
rect 553308 448604 553360 448656
rect 561772 448604 561824 448656
rect 3148 448536 3200 448588
rect 20076 448536 20128 448588
rect 385592 448536 385644 448588
rect 407304 448536 407356 448588
rect 553032 448536 553084 448588
rect 570236 448536 570288 448588
rect 350448 447108 350500 447160
rect 365904 447108 365956 447160
rect 379428 447108 379480 447160
rect 407304 447108 407356 447160
rect 395528 447040 395580 447092
rect 407396 447040 407448 447092
rect 350448 445816 350500 445868
rect 366732 445816 366784 445868
rect 44732 445748 44784 445800
rect 46480 445748 46532 445800
rect 350080 445748 350132 445800
rect 375380 445748 375432 445800
rect 350448 445680 350500 445732
rect 400956 445680 401008 445732
rect 397000 445612 397052 445664
rect 407304 445612 407356 445664
rect 27068 444388 27120 444440
rect 45928 444388 45980 444440
rect 552572 444388 552624 444440
rect 583024 444388 583076 444440
rect 24492 442960 24544 443012
rect 46756 442960 46808 443012
rect 553308 442960 553360 443012
rect 573364 442960 573416 443012
rect 350448 441600 350500 441652
rect 368848 441600 368900 441652
rect 370780 441600 370832 441652
rect 407304 441600 407356 441652
rect 401140 441532 401192 441584
rect 407396 441532 407448 441584
rect 350448 440240 350500 440292
rect 382096 440240 382148 440292
rect 42524 438880 42576 438932
rect 45928 438880 45980 438932
rect 374920 438880 374972 438932
rect 407212 438880 407264 438932
rect 405004 438812 405056 438864
rect 407488 438812 407540 438864
rect 553308 438064 553360 438116
rect 558000 438064 558052 438116
rect 350080 437452 350132 437504
rect 387616 437452 387668 437504
rect 393044 437452 393096 437504
rect 407212 437452 407264 437504
rect 553308 437452 553360 437504
rect 562232 437452 562284 437504
rect 350448 437384 350500 437436
rect 403716 437384 403768 437436
rect 43628 436092 43680 436144
rect 46756 436092 46808 436144
rect 373632 436092 373684 436144
rect 407212 436092 407264 436144
rect 552664 436092 552716 436144
rect 563520 436092 563572 436144
rect 39856 434732 39908 434784
rect 46756 434732 46808 434784
rect 350448 434732 350500 434784
rect 372712 434732 372764 434784
rect 388812 434732 388864 434784
rect 407212 434732 407264 434784
rect 552664 434732 552716 434784
rect 581368 434732 581420 434784
rect 37924 433304 37976 433356
rect 46756 433304 46808 433356
rect 405280 432488 405332 432540
rect 407212 432488 407264 432540
rect 28908 431944 28960 431996
rect 46388 431944 46440 431996
rect 576308 431876 576360 431928
rect 580172 431876 580224 431928
rect 350448 430652 350500 430704
rect 361028 430652 361080 430704
rect 350080 430584 350132 430636
rect 363972 430584 364024 430636
rect 43904 430516 43956 430568
rect 46388 430516 46440 430568
rect 32588 429156 32640 429208
rect 46756 429156 46808 429208
rect 397184 427864 397236 427916
rect 407212 427864 407264 427916
rect 36728 427796 36780 427848
rect 46756 427796 46808 427848
rect 350448 427796 350500 427848
rect 405004 427796 405056 427848
rect 373724 426572 373776 426624
rect 407304 426572 407356 426624
rect 370872 426504 370924 426556
rect 407212 426504 407264 426556
rect 350448 426436 350500 426488
rect 403716 426436 403768 426488
rect 553032 426436 553084 426488
rect 574836 426436 574888 426488
rect 408408 426368 408460 426420
rect 409144 426368 409196 426420
rect 40868 425076 40920 425128
rect 46756 425076 46808 425128
rect 350448 425076 350500 425128
rect 360660 425076 360712 425128
rect 395896 425076 395948 425128
rect 407212 425076 407264 425128
rect 553032 425076 553084 425128
rect 568948 425076 569000 425128
rect 35256 425008 35308 425060
rect 46664 425008 46716 425060
rect 552940 423716 552992 423768
rect 569040 423716 569092 423768
rect 26976 423648 27028 423700
rect 46756 423648 46808 423700
rect 380716 423648 380768 423700
rect 407212 423648 407264 423700
rect 553032 423648 553084 423700
rect 570696 423648 570748 423700
rect 350448 422288 350500 422340
rect 365444 422288 365496 422340
rect 390284 422288 390336 422340
rect 407212 422288 407264 422340
rect 34980 421540 35032 421592
rect 40592 421540 40644 421592
rect 350080 420996 350132 421048
rect 353760 420996 353812 421048
rect 552296 420996 552348 421048
rect 555240 420996 555292 421048
rect 35256 420928 35308 420980
rect 46756 420928 46808 420980
rect 350448 420928 350500 420980
rect 369308 420928 369360 420980
rect 570880 420180 570932 420232
rect 580448 420180 580500 420232
rect 553032 419840 553084 419892
rect 558092 419840 558144 419892
rect 40592 419568 40644 419620
rect 46664 419568 46716 419620
rect 376392 419568 376444 419620
rect 407304 419568 407356 419620
rect 28448 419500 28500 419552
rect 46756 419500 46808 419552
rect 350448 419500 350500 419552
rect 361948 419500 362000 419552
rect 362408 419500 362460 419552
rect 407212 419500 407264 419552
rect 36820 418208 36872 418260
rect 46664 418208 46716 418260
rect 388904 418208 388956 418260
rect 407212 418208 407264 418260
rect 33692 418140 33744 418192
rect 46756 418140 46808 418192
rect 350448 418140 350500 418192
rect 400956 418140 401008 418192
rect 350448 416780 350500 416832
rect 377956 416780 378008 416832
rect 405096 416712 405148 416764
rect 407580 416712 407632 416764
rect 552020 416032 552072 416084
rect 559656 416032 559708 416084
rect 43904 415488 43956 415540
rect 46756 415488 46808 415540
rect 24400 415420 24452 415472
rect 46664 415420 46716 415472
rect 552020 415420 552072 415472
rect 566096 415420 566148 415472
rect 350448 414400 350500 414452
rect 356796 414400 356848 414452
rect 20444 413992 20496 414044
rect 46756 413992 46808 414044
rect 350448 413992 350500 414044
rect 383476 413992 383528 414044
rect 387708 413992 387760 414044
rect 407212 413992 407264 414044
rect 552020 412768 552072 412820
rect 555332 412768 555384 412820
rect 552204 412632 552256 412684
rect 578608 412632 578660 412684
rect 406200 411340 406252 411392
rect 407304 411340 407356 411392
rect 31484 411272 31536 411324
rect 46572 411272 46624 411324
rect 350448 411272 350500 411324
rect 390192 411272 390244 411324
rect 391664 411272 391716 411324
rect 407212 411272 407264 411324
rect 2964 411204 3016 411256
rect 31116 411204 31168 411256
rect 387524 409844 387576 409896
rect 407212 409844 407264 409896
rect 406292 408484 406344 408536
rect 408132 408484 408184 408536
rect 350448 407192 350500 407244
rect 375472 407192 375524 407244
rect 21456 407124 21508 407176
rect 46572 407124 46624 407176
rect 370964 407124 371016 407176
rect 407212 407124 407264 407176
rect 391388 405696 391440 405748
rect 407212 405696 407264 405748
rect 402520 405628 402572 405680
rect 407304 405628 407356 405680
rect 552940 405628 552992 405680
rect 579068 405628 579120 405680
rect 350448 404404 350500 404456
rect 358452 404404 358504 404456
rect 350080 404336 350132 404388
rect 367376 404336 367428 404388
rect 552940 403044 552992 403096
rect 562048 403044 562100 403096
rect 35164 402976 35216 403028
rect 45928 402976 45980 403028
rect 552848 402976 552900 403028
rect 575848 402976 575900 403028
rect 42432 401820 42484 401872
rect 43260 401820 43312 401872
rect 391572 401616 391624 401668
rect 407212 401616 407264 401668
rect 41972 400188 42024 400240
rect 46112 400188 46164 400240
rect 350448 400188 350500 400240
rect 365352 400188 365404 400240
rect 33784 398828 33836 398880
rect 46572 398828 46624 398880
rect 350448 398828 350500 398880
rect 359372 398828 359424 398880
rect 387432 397536 387484 397588
rect 407212 397536 407264 397588
rect 3516 397468 3568 397520
rect 17316 397468 17368 397520
rect 350448 397468 350500 397520
rect 397000 397468 397052 397520
rect 348516 397264 348568 397316
rect 351184 397264 351236 397316
rect 42432 396448 42484 396500
rect 46480 396448 46532 396500
rect 350448 396040 350500 396092
rect 382832 396040 382884 396092
rect 39580 394748 39632 394800
rect 45836 394748 45888 394800
rect 349804 394748 349856 394800
rect 352012 394748 352064 394800
rect 22744 394680 22796 394732
rect 46572 394680 46624 394732
rect 350080 394680 350132 394732
rect 351460 394680 351512 394732
rect 388352 394680 388404 394732
rect 407212 394680 407264 394732
rect 552940 394680 552992 394732
rect 581828 394680 581880 394732
rect 350448 394612 350500 394664
rect 399760 394612 399812 394664
rect 552020 393456 552072 393508
rect 554320 393456 554372 393508
rect 39580 393320 39632 393372
rect 46572 393320 46624 393372
rect 398380 393320 398432 393372
rect 407212 393320 407264 393372
rect 37832 392028 37884 392080
rect 46572 392028 46624 392080
rect 27344 391960 27396 392012
rect 46480 391960 46532 392012
rect 350448 391960 350500 392012
rect 356888 391960 356940 392012
rect 390100 390600 390152 390652
rect 407212 390600 407264 390652
rect 552848 390600 552900 390652
rect 560852 390600 560904 390652
rect 36268 390532 36320 390584
rect 46480 390532 46532 390584
rect 350080 390532 350132 390584
rect 352748 390532 352800 390584
rect 358360 390532 358412 390584
rect 407304 390532 407356 390584
rect 552940 390532 552992 390584
rect 568856 390532 568908 390584
rect 37188 390464 37240 390516
rect 46572 390464 46624 390516
rect 350448 390464 350500 390516
rect 395436 390464 395488 390516
rect 350080 390056 350132 390108
rect 350356 390056 350408 390108
rect 348884 389376 348936 389428
rect 349528 389376 349580 389428
rect 20536 389172 20588 389224
rect 46572 389172 46624 389224
rect 350356 389172 350408 389224
rect 401140 389172 401192 389224
rect 552296 389172 552348 389224
rect 578792 389172 578844 389224
rect 348884 388424 348936 388476
rect 357716 388424 357768 388476
rect 350448 387812 350500 387864
rect 397092 387812 397144 387864
rect 552940 387812 552992 387864
rect 579804 387812 579856 387864
rect 350356 387744 350408 387796
rect 377864 387744 377916 387796
rect 38016 387064 38068 387116
rect 45560 387064 45612 387116
rect 29920 386384 29972 386436
rect 46572 386384 46624 386436
rect 552940 386384 552992 386436
rect 560944 386384 560996 386436
rect 36452 386316 36504 386368
rect 46480 386316 46532 386368
rect 391480 386316 391532 386368
rect 407212 386316 407264 386368
rect 38016 385024 38068 385076
rect 46572 385024 46624 385076
rect 552940 385024 552992 385076
rect 563244 385024 563296 385076
rect 350080 384956 350132 385008
rect 351184 384956 351236 385008
rect 36452 384276 36504 384328
rect 45652 384276 45704 384328
rect 400680 383664 400732 383716
rect 407212 383664 407264 383716
rect 29644 382236 29696 382288
rect 46572 382236 46624 382288
rect 350448 382236 350500 382288
rect 394332 382236 394384 382288
rect 552940 381080 552992 381132
rect 559748 381080 559800 381132
rect 380072 381012 380124 381064
rect 407212 381012 407264 381064
rect 350356 380944 350408 380996
rect 387800 380944 387852 380996
rect 350448 380876 350500 380928
rect 392952 380876 393004 380928
rect 394424 380128 394476 380180
rect 407856 380128 407908 380180
rect 32496 379516 32548 379568
rect 46572 379516 46624 379568
rect 29552 378156 29604 378208
rect 46572 378156 46624 378208
rect 377864 378156 377916 378208
rect 407212 378156 407264 378208
rect 574928 378156 574980 378208
rect 580172 378156 580224 378208
rect 350448 376728 350500 376780
rect 375012 376728 375064 376780
rect 552940 376728 552992 376780
rect 583116 376728 583168 376780
rect 350356 375368 350408 375420
rect 395436 375368 395488 375420
rect 350448 375300 350500 375352
rect 375104 375300 375156 375352
rect 43444 374688 43496 374740
rect 47216 374688 47268 374740
rect 26884 374008 26936 374060
rect 46480 374008 46532 374060
rect 395712 374008 395764 374060
rect 407212 374008 407264 374060
rect 28356 372648 28408 372700
rect 46112 372648 46164 372700
rect 552940 372648 552992 372700
rect 556528 372648 556580 372700
rect 26792 372580 26844 372632
rect 46480 372580 46532 372632
rect 350448 372580 350500 372632
rect 379152 372580 379204 372632
rect 399944 372580 399996 372632
rect 407212 372580 407264 372632
rect 30748 371220 30800 371272
rect 46480 371220 46532 371272
rect 350448 371220 350500 371272
rect 375196 371220 375248 371272
rect 374552 371152 374604 371204
rect 407212 371152 407264 371204
rect 41880 369860 41932 369912
rect 43444 369860 43496 369912
rect 552940 369860 552992 369912
rect 562140 369860 562192 369912
rect 552940 368568 552992 368620
rect 557908 368568 557960 368620
rect 29736 368500 29788 368552
rect 46480 368500 46532 368552
rect 400772 368500 400824 368552
rect 407212 368500 407264 368552
rect 552848 368500 552900 368552
rect 571800 368500 571852 368552
rect 552020 368092 552072 368144
rect 553768 368092 553820 368144
rect 29828 367072 29880 367124
rect 46388 367072 46440 367124
rect 31392 367004 31444 367056
rect 46480 367004 46532 367056
rect 552940 365780 552992 365832
rect 566372 365780 566424 365832
rect 552848 365712 552900 365764
rect 578424 365712 578476 365764
rect 350448 365644 350500 365696
rect 353852 365644 353904 365696
rect 350448 364352 350500 364404
rect 383660 364352 383712 364404
rect 28724 362924 28776 362976
rect 46480 362924 46532 362976
rect 552848 362924 552900 362976
rect 555148 362924 555200 362976
rect 366732 361496 366784 361548
rect 407212 361496 407264 361548
rect 552204 360408 552256 360460
rect 555148 360408 555200 360460
rect 364064 360204 364116 360256
rect 407212 360204 407264 360256
rect 552940 360204 552992 360256
rect 571984 360204 572036 360256
rect 32680 358708 32732 358760
rect 46480 358708 46532 358760
rect 552940 358708 552992 358760
rect 574928 358708 574980 358760
rect 348792 358504 348844 358556
rect 352472 358504 352524 358556
rect 350448 357960 350500 358012
rect 355416 357960 355468 358012
rect 552664 357620 552716 357672
rect 556804 357620 556856 357672
rect 3148 357416 3200 357468
rect 24124 357416 24176 357468
rect 386972 357416 387024 357468
rect 407212 357416 407264 357468
rect 349988 356056 350040 356108
rect 352472 356056 352524 356108
rect 395528 356056 395580 356108
rect 407212 356056 407264 356108
rect 350448 355988 350500 356040
rect 388720 355988 388772 356040
rect 25504 354696 25556 354748
rect 46480 354696 46532 354748
rect 350448 354696 350500 354748
rect 375104 354696 375156 354748
rect 552940 354696 552992 354748
rect 571708 354696 571760 354748
rect 552940 354424 552992 354476
rect 553124 354424 553176 354476
rect 553124 353744 553176 353796
rect 558184 353744 558236 353796
rect 378048 353268 378100 353320
rect 407212 353268 407264 353320
rect 553124 353268 553176 353320
rect 574376 353268 574428 353320
rect 35072 353200 35124 353252
rect 46480 353200 46532 353252
rect 402520 351976 402572 352028
rect 407212 351976 407264 352028
rect 350356 351908 350408 351960
rect 352380 351908 352432 351960
rect 379336 351908 379388 351960
rect 407304 351908 407356 351960
rect 35072 351160 35124 351212
rect 39304 351160 39356 351212
rect 552020 350888 552072 350940
rect 554044 350888 554096 350940
rect 350172 350616 350224 350668
rect 352380 350616 352432 350668
rect 350448 350548 350500 350600
rect 362500 350548 362552 350600
rect 391480 350548 391532 350600
rect 407212 350548 407264 350600
rect 552296 350548 552348 350600
rect 583208 350548 583260 350600
rect 348976 349800 349028 349852
rect 349804 349800 349856 349852
rect 350448 349188 350500 349240
rect 368296 349188 368348 349240
rect 379244 349188 379296 349240
rect 407212 349188 407264 349240
rect 17684 349120 17736 349172
rect 46480 349120 46532 349172
rect 350356 349120 350408 349172
rect 388260 349120 388312 349172
rect 553124 349120 553176 349172
rect 583300 349120 583352 349172
rect 36360 348372 36412 348424
rect 47216 348372 47268 348424
rect 553124 346468 553176 346520
rect 573180 346468 573232 346520
rect 25412 346400 25464 346452
rect 46480 346400 46532 346452
rect 552664 346400 552716 346452
rect 578700 346400 578752 346452
rect 402796 346332 402848 346384
rect 407212 346332 407264 346384
rect 350356 345448 350408 345500
rect 353852 345448 353904 345500
rect 22652 345108 22704 345160
rect 45928 345108 45980 345160
rect 3332 345040 3384 345092
rect 29460 345040 29512 345092
rect 365444 344972 365496 345024
rect 407212 344972 407264 345024
rect 350356 343680 350408 343732
rect 381452 343680 381504 343732
rect 350172 343612 350224 343664
rect 385500 343612 385552 343664
rect 350356 343544 350408 343596
rect 363144 343544 363196 343596
rect 552020 342796 552072 342848
rect 553676 342796 553728 342848
rect 395252 342252 395304 342304
rect 407212 342252 407264 342304
rect 553124 342252 553176 342304
rect 567476 342252 567528 342304
rect 45192 342184 45244 342236
rect 46296 342184 46348 342236
rect 376668 339464 376720 339516
rect 407212 339464 407264 339516
rect 350356 338104 350408 338156
rect 366088 338104 366140 338156
rect 553124 338104 553176 338156
rect 573456 338104 573508 338156
rect 28264 336744 28316 336796
rect 46480 336744 46532 336796
rect 382188 336676 382240 336728
rect 407212 336676 407264 336728
rect 552940 335316 552992 335368
rect 566464 335316 566516 335368
rect 553124 335248 553176 335300
rect 564716 335248 564768 335300
rect 350356 333956 350408 334008
rect 382188 333956 382240 334008
rect 553124 333956 553176 334008
rect 580080 333956 580132 334008
rect 350356 332596 350408 332648
rect 366824 332596 366876 332648
rect 39304 332528 39356 332580
rect 45652 332528 45704 332580
rect 376576 331236 376628 331288
rect 407212 331236 407264 331288
rect 36636 331168 36688 331220
rect 46848 331168 46900 331220
rect 350356 329808 350408 329860
rect 363144 329808 363196 329860
rect 365536 329808 365588 329860
rect 407212 329808 407264 329860
rect 28172 328448 28224 328500
rect 45836 328448 45888 328500
rect 350356 328448 350408 328500
rect 369400 328448 369452 328500
rect 381360 328448 381412 328500
rect 407212 328448 407264 328500
rect 553124 327088 553176 327140
rect 577596 327088 577648 327140
rect 553124 325728 553176 325780
rect 569132 325728 569184 325780
rect 43720 325660 43772 325712
rect 45744 325660 45796 325712
rect 350356 325660 350408 325712
rect 363236 325660 363288 325712
rect 552940 325660 552992 325712
rect 581644 325660 581696 325712
rect 31300 325592 31352 325644
rect 46848 325592 46900 325644
rect 376484 325592 376536 325644
rect 407212 325592 407264 325644
rect 572076 325592 572128 325644
rect 580172 325592 580224 325644
rect 552940 323280 552992 323332
rect 556712 323280 556764 323332
rect 407120 323144 407172 323196
rect 407396 323144 407448 323196
rect 402152 323008 402204 323060
rect 407212 323008 407264 323060
rect 39212 322940 39264 322992
rect 46848 322940 46900 322992
rect 377312 322940 377364 322992
rect 407120 322940 407172 322992
rect 363236 322872 363288 322924
rect 407212 322872 407264 322924
rect 401048 322804 401100 322856
rect 407120 322804 407172 322856
rect 552020 321784 552072 321836
rect 553676 321784 553728 321836
rect 43352 321580 43404 321632
rect 46848 321580 46900 321632
rect 350356 321580 350408 321632
rect 378692 321580 378744 321632
rect 407856 320832 407908 320884
rect 408408 320832 408460 320884
rect 28080 320152 28132 320204
rect 46848 320152 46900 320204
rect 350356 320152 350408 320204
rect 371148 320152 371200 320204
rect 395804 320152 395856 320204
rect 407120 320152 407172 320204
rect 350172 320084 350224 320136
rect 383384 320084 383436 320136
rect 43720 318928 43772 318980
rect 46848 318928 46900 318980
rect 350356 318792 350408 318844
rect 382740 318792 382792 318844
rect 44640 318588 44692 318640
rect 46848 318588 46900 318640
rect 553124 317500 553176 317552
rect 564716 317500 564768 317552
rect 350356 317432 350408 317484
rect 393872 317432 393924 317484
rect 396632 317432 396684 317484
rect 407120 317432 407172 317484
rect 552940 317432 552992 317484
rect 579896 317432 579948 317484
rect 553124 316004 553176 316056
rect 576308 316004 576360 316056
rect 350356 315936 350408 315988
rect 398380 315936 398432 315988
rect 577504 315324 577556 315376
rect 580448 315324 580500 315376
rect 32680 314644 32732 314696
rect 46848 314644 46900 314696
rect 350172 314644 350224 314696
rect 392860 314644 392912 314696
rect 552940 313284 552992 313336
rect 583392 313284 583444 313336
rect 553124 313216 553176 313268
rect 567292 313216 567344 313268
rect 44364 313080 44416 313132
rect 46388 313080 46440 313132
rect 350356 311856 350408 311908
rect 388720 311856 388772 311908
rect 399852 311856 399904 311908
rect 407120 311856 407172 311908
rect 403532 310564 403584 310616
rect 407120 310564 407172 310616
rect 552940 310564 552992 310616
rect 574560 310564 574612 310616
rect 22560 310496 22612 310548
rect 46848 310496 46900 310548
rect 350356 310496 350408 310548
rect 368112 310496 368164 310548
rect 399760 310496 399812 310548
rect 407212 310496 407264 310548
rect 553124 310496 553176 310548
rect 577688 310496 577740 310548
rect 368020 310428 368072 310480
rect 407120 310428 407172 310480
rect 350172 309748 350224 309800
rect 357624 309748 357676 309800
rect 32404 309136 32456 309188
rect 46848 309136 46900 309188
rect 553124 309136 553176 309188
rect 575940 309136 575992 309188
rect 350356 307776 350408 307828
rect 353944 307776 353996 307828
rect 358544 307776 358596 307828
rect 407120 307776 407172 307828
rect 553124 307776 553176 307828
rect 572076 307776 572128 307828
rect 388260 307708 388312 307760
rect 407212 307708 407264 307760
rect 552020 307436 552072 307488
rect 553860 307436 553912 307488
rect 552296 305328 552348 305380
rect 555424 305328 555476 305380
rect 3516 304988 3568 305040
rect 26700 304988 26752 305040
rect 349896 304988 349948 305040
rect 350724 304988 350776 305040
rect 398012 304988 398064 305040
rect 407120 304988 407172 305040
rect 553124 304988 553176 305040
rect 583484 304988 583536 305040
rect 351184 304308 351236 304360
rect 352656 304308 352708 304360
rect 350356 303696 350408 303748
rect 374552 303696 374604 303748
rect 31300 303628 31352 303680
rect 46848 303628 46900 303680
rect 359648 303628 359700 303680
rect 407120 303628 407172 303680
rect 372804 302880 372856 302932
rect 379428 302880 379480 302932
rect 350356 302268 350408 302320
rect 354220 302268 354272 302320
rect 25596 302200 25648 302252
rect 46480 302200 46532 302252
rect 349804 302200 349856 302252
rect 350540 302200 350592 302252
rect 405188 302200 405240 302252
rect 407396 302200 407448 302252
rect 43536 302132 43588 302184
rect 46848 302132 46900 302184
rect 401048 300908 401100 300960
rect 407120 300908 407172 300960
rect 21272 300840 21324 300892
rect 46848 300840 46900 300892
rect 350356 300840 350408 300892
rect 365444 300840 365496 300892
rect 366732 300840 366784 300892
rect 407212 300840 407264 300892
rect 553124 300840 553176 300892
rect 570512 300840 570564 300892
rect 350080 300772 350132 300824
rect 353668 300772 353720 300824
rect 350356 299548 350408 299600
rect 379428 299548 379480 299600
rect 368020 299480 368072 299532
rect 407120 299480 407172 299532
rect 553124 299480 553176 299532
rect 571892 299480 571944 299532
rect 18972 298120 19024 298172
rect 46848 298120 46900 298172
rect 350356 298120 350408 298172
rect 354036 298120 354088 298172
rect 350080 297984 350132 298036
rect 350356 297984 350408 298036
rect 553124 297848 553176 297900
rect 556896 297848 556948 297900
rect 18880 296692 18932 296744
rect 46848 296692 46900 296744
rect 553124 296692 553176 296744
rect 572168 296692 572220 296744
rect 350080 295468 350132 295520
rect 350264 295468 350316 295520
rect 348424 295332 348476 295384
rect 349252 295332 349304 295384
rect 350264 295332 350316 295384
rect 379980 295332 380032 295384
rect 399392 295332 399444 295384
rect 407120 295332 407172 295384
rect 365168 294584 365220 294636
rect 384212 294584 384264 294636
rect 348976 294040 349028 294092
rect 350540 294040 350592 294092
rect 350264 293972 350316 294024
rect 368940 293972 368992 294024
rect 32772 293904 32824 293956
rect 46480 293904 46532 293956
rect 552020 293088 552072 293140
rect 553768 293088 553820 293140
rect 371056 292612 371108 292664
rect 407120 292612 407172 292664
rect 3516 292544 3568 292596
rect 20168 292544 20220 292596
rect 44640 292544 44692 292596
rect 46848 292544 46900 292596
rect 365168 292544 365220 292596
rect 407212 292544 407264 292596
rect 399668 292476 399720 292528
rect 407120 292476 407172 292528
rect 401232 292408 401284 292460
rect 407212 292408 407264 292460
rect 552204 291728 552256 291780
rect 555516 291728 555568 291780
rect 43536 291184 43588 291236
rect 46848 291184 46900 291236
rect 553124 291184 553176 291236
rect 562324 291184 562376 291236
rect 552020 290096 552072 290148
rect 553860 290096 553912 290148
rect 351184 288464 351236 288516
rect 356520 288464 356572 288516
rect 395620 288464 395672 288516
rect 407120 288464 407172 288516
rect 552940 288464 552992 288516
rect 563888 288464 563940 288516
rect 28540 288396 28592 288448
rect 46848 288396 46900 288448
rect 350264 288396 350316 288448
rect 386880 288396 386932 288448
rect 553124 288396 553176 288448
rect 578516 288396 578568 288448
rect 404912 287376 404964 287428
rect 407212 287376 407264 287428
rect 391112 287172 391164 287224
rect 407120 287172 407172 287224
rect 350264 287104 350316 287156
rect 357072 287104 357124 287156
rect 350264 286968 350316 287020
rect 356428 286968 356480 287020
rect 349344 286220 349396 286272
rect 350632 286220 350684 286272
rect 355508 285744 355560 285796
rect 399300 285744 399352 285796
rect 30932 285676 30984 285728
rect 46848 285676 46900 285728
rect 349804 285676 349856 285728
rect 407120 285676 407172 285728
rect 553124 285676 553176 285728
rect 569592 285676 569644 285728
rect 350264 285608 350316 285660
rect 365536 285608 365588 285660
rect 403900 285608 403952 285660
rect 407212 285608 407264 285660
rect 43444 284316 43496 284368
rect 44824 284316 44876 284368
rect 392492 284316 392544 284368
rect 407120 284316 407172 284368
rect 368296 284248 368348 284300
rect 407212 284248 407264 284300
rect 553124 283568 553176 283620
rect 564716 283568 564768 283620
rect 368204 282888 368256 282940
rect 407120 282888 407172 282940
rect 553124 282820 553176 282872
rect 568764 282820 568816 282872
rect 348424 282004 348476 282056
rect 349160 282004 349212 282056
rect 25320 281528 25372 281580
rect 46848 281528 46900 281580
rect 405096 281392 405148 281444
rect 409236 281392 409288 281444
rect 553124 280848 553176 280900
rect 558276 280848 558328 280900
rect 553124 280168 553176 280220
rect 564992 280168 565044 280220
rect 552940 280100 552992 280152
rect 564808 280100 564860 280152
rect 395160 278740 395212 278792
rect 407120 278740 407172 278792
rect 553124 278740 553176 278792
rect 570880 278740 570932 278792
rect 402060 277992 402112 278044
rect 408040 277992 408092 278044
rect 20352 277380 20404 277432
rect 46848 277380 46900 277432
rect 350264 277380 350316 277432
rect 403440 277380 403492 277432
rect 553124 277380 553176 277432
rect 563796 277380 563848 277432
rect 391296 277312 391348 277364
rect 407120 277312 407172 277364
rect 348884 276020 348936 276072
rect 350540 276020 350592 276072
rect 553124 276020 553176 276072
rect 576032 276020 576084 276072
rect 365076 275952 365128 276004
rect 407120 275952 407172 276004
rect 350264 275884 350316 275936
rect 387248 275884 387300 275936
rect 352564 275272 352616 275324
rect 357624 275272 357676 275324
rect 40776 274864 40828 274916
rect 46940 274864 46992 274916
rect 552296 274728 552348 274780
rect 555240 274728 555292 274780
rect 350264 273368 350316 273420
rect 355508 273368 355560 273420
rect 349988 273300 350040 273352
rect 353576 273300 353628 273352
rect 350172 273232 350224 273284
rect 391020 273232 391072 273284
rect 553124 273232 553176 273284
rect 579988 273232 580040 273284
rect 572076 273164 572128 273216
rect 580172 273164 580224 273216
rect 407488 272552 407540 272604
rect 407764 272552 407816 272604
rect 350264 271872 350316 271924
rect 353576 271872 353628 271924
rect 398380 271872 398432 271924
rect 407120 271872 407172 271924
rect 403992 271804 404044 271856
rect 407212 271804 407264 271856
rect 553124 270512 553176 270564
rect 577504 270512 577556 270564
rect 350264 270444 350316 270496
rect 395344 270444 395396 270496
rect 350080 270376 350132 270428
rect 350816 270376 350868 270428
rect 40500 270240 40552 270292
rect 43444 270240 43496 270292
rect 551928 270036 551980 270088
rect 552848 270036 552900 270088
rect 376484 269084 376536 269136
rect 407120 269084 407172 269136
rect 348884 269016 348936 269068
rect 350540 269016 350592 269068
rect 348976 268948 349028 269000
rect 349160 268948 349212 269000
rect 350264 268948 350316 269000
rect 355140 268948 355192 269000
rect 348976 268812 349028 268864
rect 349528 268812 349580 268864
rect 553124 268608 553176 268660
rect 556988 268608 557040 268660
rect 36636 268064 36688 268116
rect 39304 268064 39356 268116
rect 43444 267792 43496 267844
rect 46848 267792 46900 267844
rect 43260 267724 43312 267776
rect 44180 267724 44232 267776
rect 402796 267724 402848 267776
rect 407120 267724 407172 267776
rect 35072 266976 35124 267028
rect 39120 266976 39172 267028
rect 350264 266364 350316 266416
rect 389732 266364 389784 266416
rect 405648 266364 405700 266416
rect 407764 266364 407816 266416
rect 367928 265616 367980 265668
rect 396448 265616 396500 265668
rect 553124 264936 553176 264988
rect 570328 264936 570380 264988
rect 350264 263644 350316 263696
rect 367468 263644 367520 263696
rect 553124 263644 553176 263696
rect 567752 263644 567804 263696
rect 46296 263576 46348 263628
rect 46940 263576 46992 263628
rect 365628 263576 365680 263628
rect 407120 263576 407172 263628
rect 552940 263576 552992 263628
rect 568580 263576 568632 263628
rect 365536 262896 365588 262948
rect 367192 262896 367244 262948
rect 552020 262352 552072 262404
rect 554780 262352 554832 262404
rect 349436 262216 349488 262268
rect 351276 262216 351328 262268
rect 403900 262216 403952 262268
rect 407120 262216 407172 262268
rect 36360 262148 36412 262200
rect 43260 262148 43312 262200
rect 348976 262148 349028 262200
rect 349252 262148 349304 262200
rect 350264 262148 350316 262200
rect 365628 262148 365680 262200
rect 405004 262148 405056 262200
rect 406568 262148 406620 262200
rect 395068 261060 395120 261112
rect 396724 261060 396776 261112
rect 401232 260856 401284 260908
rect 407120 260856 407172 260908
rect 553124 260856 553176 260908
rect 564808 260856 564860 260908
rect 348976 260788 349028 260840
rect 349160 260788 349212 260840
rect 385500 260788 385552 260840
rect 387248 260788 387300 260840
rect 552940 259496 552992 259548
rect 567292 259496 567344 259548
rect 45468 259428 45520 259480
rect 46940 259428 46992 259480
rect 396540 259428 396592 259480
rect 407120 259428 407172 259480
rect 553124 259428 553176 259480
rect 583576 259428 583628 259480
rect 376300 259360 376352 259412
rect 377220 259360 377272 259412
rect 570604 259360 570656 259412
rect 580172 259360 580224 259412
rect 349528 258068 349580 258120
rect 385500 258068 385552 258120
rect 553124 258068 553176 258120
rect 560300 258068 560352 258120
rect 376300 256776 376352 256828
rect 407120 256776 407172 256828
rect 356980 256708 357032 256760
rect 407212 256708 407264 256760
rect 553124 256708 553176 256760
rect 564440 256708 564492 256760
rect 45284 255688 45336 255740
rect 45744 255688 45796 255740
rect 350172 255416 350224 255468
rect 350448 255416 350500 255468
rect 350448 255280 350500 255332
rect 393780 255280 393832 255332
rect 3148 255212 3200 255264
rect 31024 255212 31076 255264
rect 405372 255212 405424 255264
rect 407396 255212 407448 255264
rect 46388 254328 46440 254380
rect 46572 254328 46624 254380
rect 552940 253988 552992 254040
rect 564716 253988 564768 254040
rect 35072 253920 35124 253972
rect 46572 253920 46624 253972
rect 350448 253920 350500 253972
rect 355140 253920 355192 253972
rect 391296 253920 391348 253972
rect 407120 253920 407172 253972
rect 553124 253920 553176 253972
rect 570420 253920 570472 253972
rect 553124 252560 553176 252612
rect 569316 252560 569368 252612
rect 403992 251200 404044 251252
rect 407212 251200 407264 251252
rect 553124 251200 553176 251252
rect 573548 251200 573600 251252
rect 400128 251132 400180 251184
rect 407120 251132 407172 251184
rect 405372 251064 405424 251116
rect 408500 251064 408552 251116
rect 361120 249840 361172 249892
rect 407212 249840 407264 249892
rect 350448 249772 350500 249824
rect 397920 249772 397972 249824
rect 552940 249772 552992 249824
rect 568028 249772 568080 249824
rect 348792 249704 348844 249756
rect 349344 249704 349396 249756
rect 553124 249704 553176 249756
rect 567200 249704 567252 249756
rect 34980 249024 35032 249076
rect 46296 249024 46348 249076
rect 350448 248412 350500 248464
rect 400128 248412 400180 248464
rect 350080 248344 350132 248396
rect 355048 248344 355100 248396
rect 563704 247664 563756 247716
rect 575020 247664 575072 247716
rect 45376 247256 45428 247308
rect 46572 247256 46624 247308
rect 45100 247120 45152 247172
rect 45836 247120 45888 247172
rect 553124 247120 553176 247172
rect 562416 247120 562468 247172
rect 36360 247052 36412 247104
rect 46756 247052 46808 247104
rect 348608 247052 348660 247104
rect 352196 247052 352248 247104
rect 352564 247052 352616 247104
rect 353392 247052 353444 247104
rect 395896 246304 395948 246356
rect 406844 246304 406896 246356
rect 350448 245692 350500 245744
rect 357716 245760 357768 245812
rect 405004 245760 405056 245812
rect 406384 245760 406436 245812
rect 350356 245624 350408 245676
rect 363236 245692 363288 245744
rect 399668 245692 399720 245744
rect 407212 245692 407264 245744
rect 355876 245624 355928 245676
rect 359280 245624 359332 245676
rect 395344 245624 395396 245676
rect 407120 245624 407172 245676
rect 553124 245624 553176 245676
rect 563704 245624 563756 245676
rect 348884 244876 348936 244928
rect 359280 244876 359332 244928
rect 402612 244876 402664 244928
rect 407212 244876 407264 244928
rect 350172 244604 350224 244656
rect 352196 244604 352248 244656
rect 392400 244264 392452 244316
rect 407120 244264 407172 244316
rect 553124 244264 553176 244316
rect 583668 244264 583720 244316
rect 550180 243924 550232 243976
rect 550548 243924 550600 243976
rect 31024 242904 31076 242956
rect 45836 242904 45888 242956
rect 350448 242904 350500 242956
rect 396724 242904 396776 242956
rect 390192 242836 390244 242888
rect 407120 242836 407172 242888
rect 36636 242156 36688 242208
rect 47124 242156 47176 242208
rect 387248 241272 387300 241324
rect 581552 241272 581604 241324
rect 390008 241204 390060 241256
rect 563888 241204 563940 241256
rect 409512 241136 409564 241188
rect 571616 241136 571668 241188
rect 384948 240728 385000 240780
rect 409512 240592 409564 240644
rect 410156 240592 410208 240644
rect 410248 240592 410300 240644
rect 547328 240592 547380 240644
rect 562324 240796 562376 240848
rect 548708 240592 548760 240644
rect 574652 240728 574704 240780
rect 409236 240524 409288 240576
rect 412272 240524 412324 240576
rect 404084 240456 404136 240508
rect 410800 240456 410852 240508
rect 549996 240320 550048 240372
rect 552388 240320 552440 240372
rect 544292 240184 544344 240236
rect 544752 240184 544804 240236
rect 3056 240116 3108 240168
rect 30840 240116 30892 240168
rect 549536 240116 549588 240168
rect 550088 240116 550140 240168
rect 365628 240048 365680 240100
rect 577596 240048 577648 240100
rect 373816 239980 373868 240032
rect 567752 239980 567804 240032
rect 406752 239912 406804 239964
rect 580540 239912 580592 239964
rect 394516 239844 394568 239896
rect 564808 239844 564860 239896
rect 405648 239776 405700 239828
rect 573364 239776 573416 239828
rect 400128 239708 400180 239760
rect 567660 239708 567712 239760
rect 402612 239640 402664 239692
rect 564900 239640 564952 239692
rect 392952 239572 393004 239624
rect 548708 239572 548760 239624
rect 549904 239504 549956 239556
rect 564440 239504 564492 239556
rect 406200 239436 406252 239488
rect 551100 239436 551152 239488
rect 35808 239368 35860 239420
rect 45652 239368 45704 239420
rect 406844 239368 406896 239420
rect 549996 239368 550048 239420
rect 551468 239368 551520 239420
rect 560300 239368 560352 239420
rect 532056 239300 532108 239352
rect 554044 239300 554096 239352
rect 396632 239232 396684 239284
rect 550180 239232 550232 239284
rect 350356 238892 350408 238944
rect 499856 238892 499908 238944
rect 505652 238892 505704 238944
rect 570788 238892 570840 238944
rect 350448 238824 350500 238876
rect 392308 238824 392360 238876
rect 447048 238824 447100 238876
rect 551192 238824 551244 238876
rect 381544 238756 381596 238808
rect 509240 238756 509292 238808
rect 35348 238688 35400 238740
rect 46848 238688 46900 238740
rect 400864 238688 400916 238740
rect 427820 238688 427872 238740
rect 403716 238620 403768 238672
rect 440240 238620 440292 238672
rect 445116 238620 445168 238672
rect 570328 238620 570380 238672
rect 399300 238552 399352 238604
rect 428372 238552 428424 238604
rect 436744 238552 436796 238604
rect 559564 238552 559616 238604
rect 408960 238484 409012 238536
rect 504364 238484 504416 238536
rect 506664 238484 506716 238536
rect 555332 238484 555384 238536
rect 405556 238416 405608 238468
rect 514760 238416 514812 238468
rect 535276 238416 535328 238468
rect 550640 238416 550692 238468
rect 497924 238348 497976 238400
rect 558000 238348 558052 238400
rect 403440 238280 403492 238332
rect 463148 238280 463200 238332
rect 472624 238280 472676 238332
rect 551376 238280 551428 238332
rect 409144 238212 409196 238264
rect 442540 238212 442592 238264
rect 476396 238212 476448 238264
rect 554780 238212 554832 238264
rect 569224 238212 569276 238264
rect 570328 238212 570380 238264
rect 400036 238144 400088 238196
rect 432236 238144 432288 238196
rect 475384 238144 475436 238196
rect 571616 238144 571668 238196
rect 355324 238076 355376 238128
rect 416688 238076 416740 238128
rect 421288 238076 421340 238128
rect 547512 238076 547564 238128
rect 554044 238076 554096 238128
rect 561036 238076 561088 238128
rect 349896 238008 349948 238060
rect 540428 238008 540480 238060
rect 548064 238008 548116 238060
rect 558000 238008 558052 238060
rect 416688 237940 416740 237992
rect 490564 237940 490616 237992
rect 491116 237940 491168 237992
rect 501788 237940 501840 237992
rect 547604 237940 547656 237992
rect 372068 237872 372120 237924
rect 422852 237872 422904 237924
rect 482928 237872 482980 237924
rect 528192 237872 528244 237924
rect 544844 237872 544896 237924
rect 545856 237872 545908 237924
rect 552112 237872 552164 237924
rect 396816 237804 396868 237856
rect 515312 237804 515364 237856
rect 529848 237804 529900 237856
rect 545672 237804 545724 237856
rect 382832 237668 382884 237720
rect 567568 237668 567620 237720
rect 542084 237464 542136 237516
rect 549628 237464 549680 237516
rect 32772 237396 32824 237448
rect 46848 237396 46900 237448
rect 482928 237396 482980 237448
rect 483756 237396 483808 237448
rect 545764 237396 545816 237448
rect 548800 237396 548852 237448
rect 363788 237328 363840 237380
rect 552020 237328 552072 237380
rect 350448 237260 350500 237312
rect 376668 237260 376720 237312
rect 391756 237260 391808 237312
rect 578700 237260 578752 237312
rect 394332 237192 394384 237244
rect 574560 237192 574612 237244
rect 406568 237124 406620 237176
rect 580080 237124 580132 237176
rect 391572 237056 391624 237108
rect 563612 237056 563664 237108
rect 402060 236988 402112 237040
rect 573456 236988 573508 237040
rect 395712 236920 395764 236972
rect 566280 236920 566332 236972
rect 382004 236852 382056 236904
rect 550916 236852 550968 236904
rect 386880 236784 386932 236836
rect 545580 236784 545632 236836
rect 386144 236716 386196 236768
rect 532700 236716 532752 236768
rect 45376 236648 45428 236700
rect 46940 236648 46992 236700
rect 417424 236648 417476 236700
rect 553492 236648 553544 236700
rect 409328 236580 409380 236632
rect 419356 236580 419408 236632
rect 430304 236580 430356 236632
rect 556804 236580 556856 236632
rect 374828 236512 374880 236564
rect 454132 236512 454184 236564
rect 478604 236512 478656 236564
rect 556620 236512 556672 236564
rect 499212 236444 499264 236496
rect 571800 236444 571852 236496
rect 349896 235968 349948 236020
rect 350816 235968 350868 236020
rect 481548 235900 481600 235952
rect 564900 235900 564952 235952
rect 461216 235832 461268 235884
rect 550548 235832 550600 235884
rect 474648 235764 474700 235816
rect 568764 235764 568816 235816
rect 460940 235696 460992 235748
rect 564808 235696 564860 235748
rect 452568 235628 452620 235680
rect 563612 235628 563664 235680
rect 393872 235560 393924 235612
rect 511448 235560 511500 235612
rect 456708 235492 456760 235544
rect 573364 235492 573416 235544
rect 385592 235424 385644 235476
rect 551376 235424 551428 235476
rect 385040 235356 385092 235408
rect 554228 235356 554280 235408
rect 378140 235288 378192 235340
rect 558092 235288 558144 235340
rect 567660 235288 567712 235340
rect 569040 235288 569092 235340
rect 350172 235220 350224 235272
rect 541072 235220 541124 235272
rect 409420 235152 409472 235204
rect 491300 235152 491352 235204
rect 491116 235084 491168 235136
rect 562324 235084 562376 235136
rect 491208 235016 491260 235068
rect 552756 235016 552808 235068
rect 350448 234880 350500 234932
rect 356152 234880 356204 234932
rect 355508 234676 355560 234728
rect 363420 234676 363472 234728
rect 44456 234608 44508 234660
rect 45652 234608 45704 234660
rect 384764 234540 384816 234592
rect 580356 234540 580408 234592
rect 395160 234472 395212 234524
rect 545948 234472 546000 234524
rect 398472 234404 398524 234456
rect 555608 234404 555660 234456
rect 380624 234336 380676 234388
rect 540336 234336 540388 234388
rect 387708 234268 387760 234320
rect 548064 234268 548116 234320
rect 395252 234200 395304 234252
rect 566648 234200 566700 234252
rect 386236 234132 386288 234184
rect 561036 234132 561088 234184
rect 363972 234064 364024 234116
rect 544384 234064 544436 234116
rect 376760 233996 376812 234048
rect 559472 233996 559524 234048
rect 355600 233928 355652 233980
rect 555516 233928 555568 233980
rect 349068 233860 349120 233912
rect 349436 233860 349488 233912
rect 349988 233860 350040 233912
rect 580080 233860 580132 233912
rect 398012 233792 398064 233844
rect 547052 233792 547104 233844
rect 349068 233724 349120 233776
rect 352564 233724 352616 233776
rect 393136 233724 393188 233776
rect 541624 233724 541676 233776
rect 409972 233656 410024 233708
rect 410340 233656 410392 233708
rect 412640 233656 412692 233708
rect 412916 233656 412968 233708
rect 418804 233656 418856 233708
rect 420000 233656 420052 233708
rect 486976 233656 487028 233708
rect 496820 233656 496872 233708
rect 46664 233180 46716 233232
rect 47124 233180 47176 233232
rect 355876 233180 355928 233232
rect 356060 233180 356112 233232
rect 406936 233180 406988 233232
rect 580172 233180 580224 233232
rect 372436 233112 372488 233164
rect 540060 233112 540112 233164
rect 378692 233044 378744 233096
rect 547144 233044 547196 233096
rect 371148 232976 371200 233028
rect 541716 232976 541768 233028
rect 406292 232908 406344 232960
rect 578700 232908 578752 232960
rect 369216 232840 369268 232892
rect 542452 232840 542504 232892
rect 374552 232772 374604 232824
rect 547972 232772 548024 232824
rect 403808 232704 403860 232756
rect 577688 232704 577740 232756
rect 362500 232636 362552 232688
rect 540244 232636 540296 232688
rect 46848 232568 46900 232620
rect 47676 232568 47728 232620
rect 365444 232568 365496 232620
rect 548156 232568 548208 232620
rect 358452 232500 358504 232552
rect 541900 232500 541952 232552
rect 379428 232432 379480 232484
rect 471980 232432 472032 232484
rect 493416 232432 493468 232484
rect 563428 232432 563480 232484
rect 408868 232364 408920 232416
rect 470232 232364 470284 232416
rect 525616 232364 525668 232416
rect 554964 232364 555016 232416
rect 402888 232296 402940 232348
rect 416780 232296 416832 232348
rect 33600 231820 33652 231872
rect 46848 231820 46900 231872
rect 350448 231820 350500 231872
rect 353392 231820 353444 231872
rect 36452 231752 36504 231804
rect 45468 231752 45520 231804
rect 410800 231752 410852 231804
rect 538956 231752 539008 231804
rect 408224 231684 408276 231736
rect 544016 231684 544068 231736
rect 407764 231616 407816 231668
rect 546040 231616 546092 231668
rect 414020 231548 414072 231600
rect 558368 231548 558420 231600
rect 405004 231480 405056 231532
rect 549996 231480 550048 231532
rect 399392 231412 399444 231464
rect 548248 231412 548300 231464
rect 402152 231344 402204 231396
rect 562508 231344 562560 231396
rect 388352 231276 388404 231328
rect 552848 231276 552900 231328
rect 390376 231208 390428 231260
rect 563888 231208 563940 231260
rect 401324 231140 401376 231192
rect 583760 231140 583812 231192
rect 398564 231072 398616 231124
rect 581736 231072 581788 231124
rect 452660 231004 452712 231056
rect 574652 231004 574704 231056
rect 534724 230936 534776 230988
rect 536840 230936 536892 230988
rect 45284 230528 45336 230580
rect 45744 230528 45796 230580
rect 36636 230460 36688 230512
rect 46848 230460 46900 230512
rect 350448 230460 350500 230512
rect 543004 230460 543056 230512
rect 388720 229916 388772 229968
rect 448336 229916 448388 229968
rect 409052 229848 409104 229900
rect 503720 229848 503772 229900
rect 518164 229848 518216 229900
rect 543924 229848 543976 229900
rect 377772 229780 377824 229832
rect 497924 229780 497976 229832
rect 378968 229712 379020 229764
rect 401324 229712 401376 229764
rect 407948 229712 408000 229764
rect 543924 229712 543976 229764
rect 350448 229100 350500 229152
rect 366180 229100 366232 229152
rect 356796 228896 356848 228948
rect 411628 228896 411680 228948
rect 509332 228896 509384 228948
rect 572076 228896 572128 228948
rect 380532 228828 380584 228880
rect 543188 228828 543240 228880
rect 375196 228760 375248 228812
rect 541808 228760 541860 228812
rect 379980 228692 380032 228744
rect 549720 228692 549772 228744
rect 404912 228624 404964 228676
rect 576308 228624 576360 228676
rect 386972 228556 387024 228608
rect 559564 228556 559616 228608
rect 390284 228488 390336 228540
rect 563428 228488 563480 228540
rect 369400 228420 369452 228472
rect 546776 228420 546828 228472
rect 384856 228352 384908 228404
rect 577596 228352 577648 228404
rect 43260 227808 43312 227860
rect 47124 227808 47176 227860
rect 44088 227740 44140 227792
rect 46848 227740 46900 227792
rect 357072 227196 357124 227248
rect 418068 227196 418120 227248
rect 380808 227128 380860 227180
rect 512092 227128 512144 227180
rect 391020 227060 391072 227112
rect 527548 227060 527600 227112
rect 45376 226992 45428 227044
rect 46940 226992 46992 227044
rect 369308 226992 369360 227044
rect 525800 226992 525852 227044
rect 355324 226312 355376 226364
rect 360568 226312 360620 226364
rect 367836 225564 367888 225616
rect 481180 225564 481232 225616
rect 39304 225496 39356 225548
rect 46664 225496 46716 225548
rect 350448 224952 350500 225004
rect 360568 224952 360620 225004
rect 39120 224680 39172 224732
rect 44272 224680 44324 224732
rect 404176 224408 404228 224460
rect 444472 224408 444524 224460
rect 380256 224340 380308 224392
rect 459928 224340 459980 224392
rect 361028 224272 361080 224324
rect 429200 224272 429252 224324
rect 436744 224272 436796 224324
rect 563336 224272 563388 224324
rect 387616 224204 387668 224256
rect 521660 224204 521712 224256
rect 348792 223864 348844 223916
rect 349160 223864 349212 223916
rect 31116 223592 31168 223644
rect 46848 223592 46900 223644
rect 350448 223524 350500 223576
rect 388904 223524 388956 223576
rect 392308 222912 392360 222964
rect 413560 222912 413612 222964
rect 409880 222844 409932 222896
rect 472808 222844 472860 222896
rect 350172 222572 350224 222624
rect 352656 222572 352708 222624
rect 35348 222164 35400 222216
rect 46848 222164 46900 222216
rect 350264 222096 350316 222148
rect 351920 222096 351972 222148
rect 39948 221416 40000 221468
rect 40684 221416 40736 221468
rect 397920 221416 397972 221468
rect 477960 221416 478012 221468
rect 350448 221144 350500 221196
rect 356428 221144 356480 221196
rect 31208 220804 31260 220856
rect 46848 220804 46900 220856
rect 355968 220736 356020 220788
rect 356612 220736 356664 220788
rect 41052 220396 41104 220448
rect 46020 220396 46072 220448
rect 44272 220260 44324 220312
rect 46020 220260 46072 220312
rect 377956 220124 378008 220176
rect 435456 220124 435508 220176
rect 354036 220056 354088 220108
rect 494060 220056 494112 220108
rect 354588 219444 354640 219496
rect 356060 219444 356112 219496
rect 36912 218696 36964 218748
rect 46112 218696 46164 218748
rect 369124 218696 369176 218748
rect 476672 218696 476724 218748
rect 35808 218084 35860 218136
rect 46572 218084 46624 218136
rect 348976 218084 349028 218136
rect 349160 218084 349212 218136
rect 32312 218016 32364 218068
rect 46848 218016 46900 218068
rect 348700 218016 348752 218068
rect 349436 218016 349488 218068
rect 350448 218016 350500 218068
rect 355508 218016 355560 218068
rect 350264 217948 350316 218000
rect 354956 217948 355008 218000
rect 45928 217472 45980 217524
rect 45928 217268 45980 217320
rect 356704 217268 356756 217320
rect 445760 217268 445812 217320
rect 350448 217200 350500 217252
rect 355048 217200 355100 217252
rect 36912 216656 36964 216708
rect 46020 216656 46072 216708
rect 388628 215908 388680 215960
rect 535920 215908 535972 215960
rect 46388 215364 46440 215416
rect 47124 215364 47176 215416
rect 32220 215296 32272 215348
rect 46848 215296 46900 215348
rect 350448 215296 350500 215348
rect 353300 215296 353352 215348
rect 354588 215228 354640 215280
rect 356520 215228 356572 215280
rect 41788 214548 41840 214600
rect 44180 214548 44232 214600
rect 45100 214548 45152 214600
rect 45376 214548 45428 214600
rect 45836 214548 45888 214600
rect 47124 214548 47176 214600
rect 433340 214548 433392 214600
rect 581552 214548 581604 214600
rect 38108 213936 38160 213988
rect 46848 213936 46900 213988
rect 45376 213868 45428 213920
rect 45744 213868 45796 213920
rect 407028 213256 407080 213308
rect 485044 213256 485096 213308
rect 356888 213188 356940 213240
rect 542544 213188 542596 213240
rect 46572 213120 46624 213172
rect 47584 213120 47636 213172
rect 350448 212508 350500 212560
rect 508504 212508 508556 212560
rect 348976 212440 349028 212492
rect 349344 212440 349396 212492
rect 349068 212372 349120 212424
rect 349712 212372 349764 212424
rect 438676 211964 438728 212016
rect 477592 211964 477644 212016
rect 388536 211896 388588 211948
rect 441620 211896 441672 211948
rect 382740 211828 382792 211880
rect 524972 211828 525024 211880
rect 33876 211760 33928 211812
rect 47584 211760 47636 211812
rect 416964 211760 417016 211812
rect 583300 211760 583352 211812
rect 33876 211148 33928 211200
rect 46848 211148 46900 211200
rect 350448 208360 350500 208412
rect 539048 208360 539100 208412
rect 43812 208292 43864 208344
rect 46848 208292 46900 208344
rect 350448 207068 350500 207120
rect 541992 207068 542044 207120
rect 350264 207000 350316 207052
rect 566556 207000 566608 207052
rect 41236 206932 41288 206984
rect 46848 206932 46900 206984
rect 350448 206932 350500 206984
rect 376300 206932 376352 206984
rect 410064 206252 410116 206304
rect 507584 206252 507636 206304
rect 348976 206116 349028 206168
rect 352564 206116 352616 206168
rect 37188 205640 37240 205692
rect 46848 205640 46900 205692
rect 37004 205164 37056 205216
rect 37740 205164 37792 205216
rect 443000 204892 443052 204944
rect 508228 204892 508280 204944
rect 349988 204416 350040 204468
rect 351920 204416 351972 204468
rect 46848 204280 46900 204332
rect 47124 204280 47176 204332
rect 350264 204280 350316 204332
rect 389088 204280 389140 204332
rect 350448 204212 350500 204264
rect 418804 204212 418856 204264
rect 406476 203600 406528 203652
rect 519176 203600 519228 203652
rect 350080 203532 350132 203584
rect 545304 203532 545356 203584
rect 37004 202852 37056 202904
rect 45652 202852 45704 202904
rect 350448 202852 350500 202904
rect 414664 202852 414716 202904
rect 34888 202784 34940 202836
rect 45560 202784 45612 202836
rect 46388 202308 46440 202360
rect 47860 202308 47912 202360
rect 411352 202104 411404 202156
rect 476028 202104 476080 202156
rect 350448 201492 350500 201544
rect 383384 201492 383436 201544
rect 349068 200744 349120 200796
rect 359188 200744 359240 200796
rect 363328 200744 363380 200796
rect 507952 200744 508004 200796
rect 347688 200336 347740 200388
rect 42340 200064 42392 200116
rect 44272 200064 44324 200116
rect 46664 199928 46716 199980
rect 50344 199928 50396 199980
rect 347688 199860 347740 199912
rect 41052 199656 41104 199708
rect 75460 199656 75512 199708
rect 44548 199588 44600 199640
rect 90916 199588 90968 199640
rect 104072 199588 104124 199640
rect 104716 199588 104768 199640
rect 346308 199588 346360 199640
rect 348792 199588 348844 199640
rect 43444 199520 43496 199572
rect 92664 199520 92716 199572
rect 275836 199520 275888 199572
rect 340880 199520 340932 199572
rect 347504 199520 347556 199572
rect 350172 199520 350224 199572
rect 47032 199452 47084 199504
rect 108948 199452 109000 199504
rect 328184 199452 328236 199504
rect 348608 199452 348660 199504
rect 44824 199384 44876 199436
rect 158536 199384 158588 199436
rect 317236 199384 317288 199436
rect 348516 199384 348568 199436
rect 348976 199384 349028 199436
rect 354864 199384 354916 199436
rect 319812 199316 319864 199368
rect 360844 199316 360896 199368
rect 35440 199248 35492 199300
rect 106004 199248 106056 199300
rect 271512 199248 271564 199300
rect 358268 199248 358320 199300
rect 38200 199180 38252 199232
rect 118792 199180 118844 199232
rect 208400 199180 208452 199232
rect 366456 199180 366508 199232
rect 27160 199112 27212 199164
rect 127256 199112 127308 199164
rect 300492 199112 300544 199164
rect 560944 199112 560996 199164
rect 39488 199044 39540 199096
rect 104624 199044 104676 199096
rect 104716 199044 104768 199096
rect 370872 199044 370924 199096
rect 84108 198976 84160 199028
rect 371884 198976 371936 199028
rect 37096 198908 37148 198960
rect 167828 198908 167880 198960
rect 233516 198908 233568 198960
rect 542084 198908 542136 198960
rect 40500 198840 40552 198892
rect 221924 198840 221976 198892
rect 247040 198840 247092 198892
rect 559380 198840 559432 198892
rect 30012 198772 30064 198824
rect 160100 198772 160152 198824
rect 194232 198772 194284 198824
rect 559656 198772 559708 198824
rect 100852 198704 100904 198756
rect 467932 198704 467984 198756
rect 22928 198636 22980 198688
rect 48688 198636 48740 198688
rect 346216 198636 346268 198688
rect 360384 198636 360436 198688
rect 25688 198568 25740 198620
rect 101496 198568 101548 198620
rect 123392 198568 123444 198620
rect 570880 198568 570932 198620
rect 46572 198500 46624 198552
rect 168472 198500 168524 198552
rect 223856 198500 223908 198552
rect 553952 198500 554004 198552
rect 33048 198432 33100 198484
rect 67364 198432 67416 198484
rect 244464 198432 244516 198484
rect 558276 198432 558328 198484
rect 22836 198364 22888 198416
rect 55772 198364 55824 198416
rect 58624 198364 58676 198416
rect 77668 198364 77720 198416
rect 201960 198364 202012 198416
rect 491392 198364 491444 198416
rect 44732 198296 44784 198348
rect 88616 198296 88668 198348
rect 147864 198296 147916 198348
rect 254860 198296 254912 198348
rect 287612 198296 287664 198348
rect 551008 198296 551060 198348
rect 31576 198228 31628 198280
rect 64144 198228 64196 198280
rect 342996 198228 343048 198280
rect 365260 198228 365312 198280
rect 40408 198160 40460 198212
rect 145656 198160 145708 198212
rect 160744 198160 160796 198212
rect 166264 198160 166316 198212
rect 190368 198160 190420 198212
rect 383016 198160 383068 198212
rect 17776 198092 17828 198144
rect 49976 198092 50028 198144
rect 51908 198092 51960 198144
rect 165252 198092 165304 198144
rect 201316 198092 201368 198144
rect 268384 198092 268436 198144
rect 275376 198092 275428 198144
rect 364340 198092 364392 198144
rect 44088 198024 44140 198076
rect 208768 198024 208820 198076
rect 272156 198024 272208 198076
rect 307024 198024 307076 198076
rect 332048 198024 332100 198076
rect 401048 198024 401100 198076
rect 25780 197956 25832 198008
rect 48044 197956 48096 198008
rect 50068 197956 50120 198008
rect 50620 197956 50672 198008
rect 53012 197956 53064 198008
rect 395344 197956 395396 198008
rect 32864 197888 32916 197940
rect 63500 197888 63552 197940
rect 317880 197888 317932 197940
rect 385684 197888 385736 197940
rect 49516 197820 49568 197872
rect 72516 197820 72568 197872
rect 315304 197820 315356 197872
rect 349068 197820 349120 197872
rect 86684 197752 86736 197804
rect 346124 197752 346176 197804
rect 36912 197684 36964 197736
rect 487160 197684 487212 197736
rect 49332 197412 49384 197464
rect 54484 197412 54536 197464
rect 51264 197344 51316 197396
rect 53196 197344 53248 197396
rect 68284 197344 68336 197396
rect 71136 197344 71188 197396
rect 108580 197344 108632 197396
rect 109684 197344 109736 197396
rect 262496 197344 262548 197396
rect 264244 197344 264296 197396
rect 41328 197276 41380 197328
rect 73804 197276 73856 197328
rect 340420 197276 340472 197328
rect 369952 197276 370004 197328
rect 45376 197208 45428 197260
rect 89260 197208 89312 197260
rect 340880 197208 340932 197260
rect 349804 197208 349856 197260
rect 24124 197140 24176 197192
rect 422300 197140 422352 197192
rect 29460 197072 29512 197124
rect 412824 197072 412876 197124
rect 20076 197004 20128 197056
rect 392492 197004 392544 197056
rect 82176 196936 82228 196988
rect 379060 196936 379112 196988
rect 32956 196868 33008 196920
rect 295340 196868 295392 196920
rect 304356 196868 304408 196920
rect 371240 196868 371292 196920
rect 21456 196800 21508 196852
rect 275836 196800 275888 196852
rect 276664 196800 276716 196852
rect 352564 196800 352616 196852
rect 24308 196732 24360 196784
rect 246396 196732 246448 196784
rect 266084 196732 266136 196784
rect 351276 196732 351328 196784
rect 42248 196664 42300 196716
rect 220360 196664 220412 196716
rect 227720 196664 227772 196716
rect 361580 196664 361632 196716
rect 34244 196596 34296 196648
rect 75644 196596 75696 196648
rect 80152 196596 80204 196648
rect 556988 196596 557040 196648
rect 36728 196528 36780 196580
rect 135260 196528 135312 196580
rect 182640 196528 182692 196580
rect 354772 196528 354824 196580
rect 40592 196460 40644 196512
rect 125048 196460 125100 196512
rect 28448 196392 28500 196444
rect 551468 196392 551520 196444
rect 36636 196324 36688 196376
rect 463700 196324 463752 196376
rect 32404 195916 32456 195968
rect 519084 195916 519136 195968
rect 30840 195848 30892 195900
rect 465080 195848 465132 195900
rect 39948 195780 40000 195832
rect 121460 195780 121512 195832
rect 138204 195780 138256 195832
rect 569316 195780 569368 195832
rect 52276 195712 52328 195764
rect 128452 195712 128504 195764
rect 174268 195712 174320 195764
rect 549536 195712 549588 195764
rect 28080 195644 28132 195696
rect 395528 195644 395580 195696
rect 40776 195576 40828 195628
rect 228364 195576 228416 195628
rect 312728 195576 312780 195628
rect 573272 195576 573324 195628
rect 38384 195508 38436 195560
rect 86408 195508 86460 195560
rect 116952 195508 117004 195560
rect 363880 195508 363932 195560
rect 54760 195440 54812 195492
rect 247684 195440 247736 195492
rect 50896 195372 50948 195424
rect 266912 195440 266964 195492
rect 281172 195440 281224 195492
rect 348976 195440 349028 195492
rect 259460 195372 259512 195424
rect 260564 195372 260616 195424
rect 293960 195372 294012 195424
rect 294696 195372 294748 195424
rect 297916 195372 297968 195424
rect 356612 195372 356664 195424
rect 55588 195304 55640 195356
rect 350356 195304 350408 195356
rect 46756 195236 46808 195288
rect 452844 195236 452896 195288
rect 551928 195236 551980 195288
rect 556804 195236 556856 195288
rect 42156 195168 42208 195220
rect 175924 195168 175976 195220
rect 204536 195168 204588 195220
rect 361856 195168 361908 195220
rect 35532 195100 35584 195152
rect 69020 195100 69072 195152
rect 78680 195100 78732 195152
rect 79600 195100 79652 195152
rect 80060 195100 80112 195152
rect 80796 195100 80848 195152
rect 111800 195100 111852 195152
rect 113088 195100 113140 195152
rect 113180 195100 113232 195152
rect 114284 195100 114336 195152
rect 150532 195100 150584 195152
rect 151728 195100 151780 195152
rect 160100 195100 160152 195152
rect 161388 195100 161440 195152
rect 179512 195100 179564 195152
rect 180708 195100 180760 195152
rect 209780 195100 209832 195152
rect 210976 195100 211028 195152
rect 238760 195100 238812 195152
rect 239956 195100 240008 195152
rect 324320 195100 324372 195152
rect 324872 195100 324924 195152
rect 325700 195100 325752 195152
rect 326896 195100 326948 195152
rect 333980 195100 334032 195152
rect 335268 195100 335320 195152
rect 342720 195100 342772 195152
rect 355232 195100 355284 195152
rect 39764 195032 39816 195084
rect 73528 195032 73580 195084
rect 237380 194896 237432 194948
rect 238576 194896 238628 194948
rect 20444 194488 20496 194540
rect 572168 194488 572220 194540
rect 25320 194420 25372 194472
rect 566464 194420 566516 194472
rect 25412 194352 25464 194404
rect 566372 194352 566424 194404
rect 142068 194284 142120 194336
rect 529940 194284 529992 194336
rect 181352 194216 181404 194268
rect 449900 194216 449952 194268
rect 17224 194148 17276 194200
rect 281724 194148 281776 194200
rect 284760 194148 284812 194200
rect 364432 194148 364484 194200
rect 102140 194080 102192 194132
rect 364064 194080 364116 194132
rect 249616 194012 249668 194064
rect 390100 194012 390152 194064
rect 241244 193944 241296 193996
rect 370780 193944 370832 193996
rect 242992 193876 243044 193928
rect 365812 193876 365864 193928
rect 41144 193808 41196 193860
rect 141792 193808 141844 193860
rect 318892 193808 318944 193860
rect 562232 193808 562284 193860
rect 276020 193740 276072 193792
rect 352196 193740 352248 193792
rect 280528 193672 280580 193724
rect 351184 193672 351236 193724
rect 287980 193604 288032 193656
rect 358360 193604 358412 193656
rect 26700 193128 26752 193180
rect 478880 193128 478932 193180
rect 49608 193060 49660 193112
rect 189080 193060 189132 193112
rect 205180 193060 205232 193112
rect 575664 193060 575716 193112
rect 34152 192992 34204 193044
rect 337844 192992 337896 193044
rect 39672 192924 39724 192976
rect 87696 192924 87748 192976
rect 134340 192924 134392 192976
rect 346308 192924 346360 192976
rect 36912 192856 36964 192908
rect 154304 192856 154356 192908
rect 173624 192856 173676 192908
rect 361764 192856 361816 192908
rect 51448 192788 51500 192840
rect 194876 192788 194928 192840
rect 217784 192788 217836 192840
rect 349252 192788 349304 192840
rect 45468 192720 45520 192772
rect 243084 192720 243136 192772
rect 48964 192652 49016 192704
rect 263784 192652 263836 192704
rect 54208 192584 54260 192636
rect 355140 192584 355192 192636
rect 50804 192516 50856 192568
rect 356152 192516 356204 192568
rect 4804 192448 4856 192500
rect 506572 192448 506624 192500
rect 49976 192380 50028 192432
rect 172980 192380 173032 192432
rect 46848 192312 46900 192364
rect 151820 192312 151872 192364
rect 40592 192244 40644 192296
rect 85304 192244 85356 192296
rect 20168 191768 20220 191820
rect 574468 191768 574520 191820
rect 17316 191700 17368 191752
rect 391112 191700 391164 191752
rect 184572 191632 184624 191684
rect 359280 191632 359332 191684
rect 300860 191428 300912 191480
rect 348056 191428 348108 191480
rect 44640 191360 44692 191412
rect 202972 191360 203024 191412
rect 285404 191360 285456 191412
rect 353484 191360 353536 191412
rect 61568 191292 61620 191344
rect 307944 191292 307996 191344
rect 98644 191224 98696 191276
rect 366088 191224 366140 191276
rect 46848 191156 46900 191208
rect 333336 191156 333388 191208
rect 339500 191156 339552 191208
rect 351000 191156 351052 191208
rect 49424 191088 49476 191140
rect 472164 191088 472216 191140
rect 20352 190408 20404 190460
rect 578792 190408 578844 190460
rect 42064 190340 42116 190392
rect 275744 190340 275796 190392
rect 58808 190272 58860 190324
rect 341064 190272 341116 190324
rect 55956 190204 56008 190256
rect 349620 190204 349672 190256
rect 42248 190136 42300 190188
rect 380716 190136 380768 190188
rect 41328 190068 41380 190120
rect 392400 190068 392452 190120
rect 55036 190000 55088 190052
rect 409972 190000 410024 190052
rect 34152 189932 34204 189984
rect 169116 189932 169168 189984
rect 174636 189932 174688 189984
rect 560852 189932 560904 189984
rect 85764 189864 85816 189916
rect 556896 189864 556948 189916
rect 19340 189796 19392 189848
rect 556436 189796 556488 189848
rect 3516 189728 3568 189780
rect 567384 189728 567436 189780
rect 43812 189660 43864 189712
rect 216128 189660 216180 189712
rect 59452 189592 59504 189644
rect 226432 189592 226484 189644
rect 183928 188980 183980 189032
rect 582840 188980 582892 189032
rect 3424 188912 3476 188964
rect 396908 188912 396960 188964
rect 169760 188844 169812 188896
rect 356520 188844 356572 188896
rect 293132 188368 293184 188420
rect 352748 188368 352800 188420
rect 221280 188300 221332 188352
rect 252652 188300 252704 188352
rect 296352 188300 296404 188352
rect 379336 188300 379388 188352
rect 38200 187620 38252 187672
rect 179512 187620 179564 187672
rect 192024 187620 192076 187672
rect 360660 187620 360712 187672
rect 53472 187552 53524 187604
rect 236736 187552 236788 187604
rect 322112 187552 322164 187604
rect 559748 187552 559800 187604
rect 99932 187484 99984 187536
rect 370688 187484 370740 187536
rect 58716 187416 58768 187468
rect 357716 187416 357768 187468
rect 53564 187348 53616 187400
rect 354220 187348 354272 187400
rect 59728 187280 59780 187332
rect 363052 187280 363104 187332
rect 35532 187212 35584 187264
rect 349528 187212 349580 187264
rect 38292 187144 38344 187196
rect 370596 187144 370648 187196
rect 36544 187076 36596 187128
rect 371332 187076 371384 187128
rect 34336 187008 34388 187060
rect 377680 187008 377732 187060
rect 33692 186940 33744 186992
rect 490196 186940 490248 186992
rect 239036 186872 239088 186924
rect 353760 186872 353812 186924
rect 278964 186124 279016 186176
rect 366732 186124 366784 186176
rect 187516 186056 187568 186108
rect 354128 186056 354180 186108
rect 116676 185988 116728 186040
rect 351460 185988 351512 186040
rect 58256 185920 58308 185972
rect 303712 185920 303764 185972
rect 53380 185852 53432 185904
rect 356428 185852 356480 185904
rect 40776 185784 40828 185836
rect 359372 185784 359424 185836
rect 42156 185716 42208 185768
rect 381636 185716 381688 185768
rect 407120 185716 407172 185768
rect 438860 185716 438912 185768
rect 222292 185648 222344 185700
rect 561864 185648 561916 185700
rect 55864 185580 55916 185632
rect 408040 185580 408092 185632
rect 194968 184832 195020 184884
rect 201500 184832 201552 184884
rect 216496 184832 216548 184884
rect 347780 184832 347832 184884
rect 209872 184764 209924 184816
rect 352840 184764 352892 184816
rect 159180 184696 159232 184748
rect 352380 184696 352432 184748
rect 146944 184628 146996 184680
rect 351092 184628 351144 184680
rect 37832 184560 37884 184612
rect 245476 184560 245528 184612
rect 272524 184560 272576 184612
rect 383660 184560 383712 184612
rect 59820 184492 59872 184544
rect 355048 184492 355100 184544
rect 59636 184424 59688 184476
rect 357440 184424 357492 184476
rect 59084 184356 59136 184408
rect 363420 184356 363472 184408
rect 40960 184288 41012 184340
rect 183008 184288 183060 184340
rect 234528 184288 234580 184340
rect 560576 184288 560628 184340
rect 35716 184220 35768 184272
rect 367284 184220 367336 184272
rect 36636 184152 36688 184204
rect 371424 184152 371476 184204
rect 249984 184084 250036 184136
rect 352288 184084 352340 184136
rect 283472 184016 283524 184068
rect 347504 184016 347556 184068
rect 163044 183472 163096 183524
rect 348884 183472 348936 183524
rect 52184 183404 52236 183456
rect 359004 183404 359056 183456
rect 398840 183404 398892 183456
rect 402520 183404 402572 183456
rect 44088 183336 44140 183388
rect 353392 183336 353444 183388
rect 46020 183268 46072 183320
rect 360568 183268 360620 183320
rect 393780 183268 393832 183320
rect 407212 183268 407264 183320
rect 224224 183200 224276 183252
rect 552480 183200 552532 183252
rect 54668 183132 54720 183184
rect 399760 183132 399812 183184
rect 44732 183064 44784 183116
rect 407856 183064 407908 183116
rect 39672 182996 39724 183048
rect 459652 182996 459704 183048
rect 116032 182928 116084 182980
rect 558184 182928 558236 182980
rect 37924 182860 37976 182912
rect 529940 182860 529992 182912
rect 47860 182792 47912 182844
rect 573548 182792 573600 182844
rect 246120 182724 246172 182776
rect 351368 182724 351420 182776
rect 198096 182112 198148 182164
rect 302148 182112 302200 182164
rect 58900 182044 58952 182096
rect 364524 182044 364576 182096
rect 255780 181976 255832 182028
rect 561956 181976 562008 182028
rect 54944 181908 54996 181960
rect 376576 181908 376628 181960
rect 42064 181840 42116 181892
rect 368940 181840 368992 181892
rect 34244 181772 34296 181824
rect 373632 181772 373684 181824
rect 35624 181704 35676 181756
rect 381360 181704 381412 181756
rect 37096 181636 37148 181688
rect 387340 181636 387392 181688
rect 33968 181568 34020 181620
rect 391296 181568 391348 181620
rect 43536 181500 43588 181552
rect 412824 181500 412876 181552
rect 48872 181432 48924 181484
rect 426532 181432 426584 181484
rect 576124 181432 576176 181484
rect 580724 181432 580776 181484
rect 191840 180412 191892 180464
rect 274456 180412 274508 180464
rect 279608 180412 279660 180464
rect 357532 180412 357584 180464
rect 226800 180344 226852 180396
rect 358084 180344 358136 180396
rect 69664 180276 69716 180328
rect 197360 180276 197412 180328
rect 330484 180276 330536 180328
rect 552572 180276 552624 180328
rect 53104 180208 53156 180260
rect 65800 180208 65852 180260
rect 103796 180208 103848 180260
rect 347872 180208 347924 180260
rect 59912 180140 59964 180192
rect 372712 180140 372764 180192
rect 50252 180072 50304 180124
rect 400772 180072 400824 180124
rect 111984 179052 112036 179104
rect 130200 179052 130252 179104
rect 213920 179052 213972 179104
rect 346584 179052 346636 179104
rect 41972 178984 42024 179036
rect 345020 178984 345072 179036
rect 49332 178916 49384 178968
rect 367376 178916 367428 178968
rect 34060 178848 34112 178900
rect 401968 178848 402020 178900
rect 13820 178780 13872 178832
rect 432052 178780 432104 178832
rect 40500 178712 40552 178764
rect 460940 178712 460992 178764
rect 43260 178644 43312 178696
rect 488632 178644 488684 178696
rect 241612 177828 241664 177880
rect 375380 177828 375432 177880
rect 227720 177760 227772 177812
rect 469312 177760 469364 177812
rect 74816 177692 74868 177744
rect 378048 177692 378100 177744
rect 268660 177624 268712 177676
rect 578608 177624 578660 177676
rect 54576 177556 54628 177608
rect 368848 177556 368900 177608
rect 89812 177488 89864 177540
rect 99288 177488 99340 177540
rect 250628 177488 250680 177540
rect 571892 177488 571944 177540
rect 49056 177420 49108 177472
rect 391480 177420 391532 177472
rect 52644 177352 52696 177404
rect 398380 177352 398432 177404
rect 48228 177284 48280 177336
rect 399668 177284 399720 177336
rect 213276 176332 213328 176384
rect 273352 176332 273404 176384
rect 313096 176332 313148 176384
rect 380164 176332 380216 176384
rect 188160 176264 188212 176316
rect 362316 176264 362368 176316
rect 113364 176196 113416 176248
rect 379244 176196 379296 176248
rect 48136 176128 48188 176180
rect 353852 176128 353904 176180
rect 44456 176060 44508 176112
rect 360108 176060 360160 176112
rect 95240 175992 95292 176044
rect 443184 175992 443236 176044
rect 49792 175924 49844 175976
rect 526444 175924 526496 175976
rect 312452 175040 312504 175092
rect 352104 175040 352156 175092
rect 53288 174972 53340 175024
rect 349344 174972 349396 175024
rect 354312 174972 354364 175024
rect 467840 174972 467892 175024
rect 59544 174904 59596 174956
rect 380072 174904 380124 174956
rect 46756 174836 46808 174888
rect 385868 174836 385920 174888
rect 55680 174768 55732 174820
rect 401232 174768 401284 174820
rect 39764 174700 39816 174752
rect 391388 174700 391440 174752
rect 40408 174632 40460 174684
rect 483112 174632 483164 174684
rect 36728 174564 36780 174616
rect 552664 174564 552716 174616
rect 50068 174496 50120 174548
rect 574284 174496 574336 174548
rect 249340 173340 249392 173392
rect 352472 173340 352524 173392
rect 268384 173272 268436 173324
rect 506296 173272 506348 173324
rect 38660 173204 38712 173256
rect 368020 173204 368072 173256
rect 88432 173136 88484 173188
rect 480536 173136 480588 173188
rect 264152 172116 264204 172168
rect 353576 172116 353628 172168
rect 112168 172048 112220 172100
rect 129832 172048 129884 172100
rect 180800 172048 180852 172100
rect 327080 172048 327132 172100
rect 96712 171980 96764 172032
rect 242256 171980 242308 172032
rect 301044 171980 301096 172032
rect 468300 171980 468352 172032
rect 115940 171912 115992 171964
rect 343364 171912 343416 171964
rect 79324 171844 79376 171896
rect 355508 171844 355560 171896
rect 50712 171776 50764 171828
rect 375472 171776 375524 171828
rect 383384 171776 383436 171828
rect 386420 171776 386472 171828
rect 35256 170552 35308 170604
rect 193220 170552 193272 170604
rect 56416 170484 56468 170536
rect 230480 170484 230532 170536
rect 233884 170484 233936 170536
rect 389824 170484 389876 170536
rect 66444 170416 66496 170468
rect 347964 170416 348016 170468
rect 57888 170348 57940 170400
rect 387524 170348 387576 170400
rect 306472 169668 306524 169720
rect 367744 169668 367796 169720
rect 225512 169600 225564 169652
rect 365168 169600 365220 169652
rect 176660 169532 176712 169584
rect 294052 169532 294104 169584
rect 315304 169532 315356 169584
rect 484400 169532 484452 169584
rect 170772 169464 170824 169516
rect 355416 169464 355468 169516
rect 124404 169396 124456 169448
rect 363144 169396 363196 169448
rect 46572 169328 46624 169380
rect 325700 169328 325752 169380
rect 328736 169328 328788 169380
rect 394148 169328 394200 169380
rect 30104 169260 30156 169312
rect 335636 169260 335688 169312
rect 78036 169192 78088 169244
rect 388812 169192 388864 169244
rect 52828 169124 52880 169176
rect 371056 169124 371108 169176
rect 64512 169056 64564 169108
rect 563520 169056 563572 169108
rect 26792 168988 26844 169040
rect 552572 168988 552624 169040
rect 207480 167696 207532 167748
rect 402244 167696 402296 167748
rect 40868 167628 40920 167680
rect 314384 167628 314436 167680
rect 405280 167628 405332 167680
rect 565912 167628 565964 167680
rect 277400 166812 277452 166864
rect 356980 166812 357032 166864
rect 259000 166744 259052 166796
rect 350632 166744 350684 166796
rect 392860 166744 392912 166796
rect 549536 166744 549588 166796
rect 199752 166676 199804 166728
rect 372252 166676 372304 166728
rect 395068 166676 395120 166728
rect 561220 166676 561272 166728
rect 324412 166608 324464 166660
rect 563520 166608 563572 166660
rect 84200 166540 84252 166592
rect 367468 166540 367520 166592
rect 391204 166540 391256 166592
rect 560484 166540 560536 166592
rect 41144 166472 41196 166524
rect 377588 166472 377640 166524
rect 391848 166472 391900 166524
rect 566280 166472 566332 166524
rect 150532 166404 150584 166456
rect 539232 166404 539284 166456
rect 54852 166336 54904 166388
rect 470600 166336 470652 166388
rect 508504 166336 508556 166388
rect 514024 166336 514076 166388
rect 150440 166268 150492 166320
rect 567752 166268 567804 166320
rect 228732 165112 228784 165164
rect 374644 165112 374696 165164
rect 81900 165044 81952 165096
rect 231952 165044 232004 165096
rect 237380 165044 237432 165096
rect 506940 165044 506992 165096
rect 43352 164976 43404 165028
rect 350448 164976 350500 165028
rect 29552 164908 29604 164960
rect 376852 164908 376904 164960
rect 197176 164840 197228 164892
rect 560392 164840 560444 164892
rect 307024 164160 307076 164212
rect 309876 164160 309928 164212
rect 397276 164160 397328 164212
rect 548340 164160 548392 164212
rect 408132 164092 408184 164144
rect 560576 164092 560628 164144
rect 237748 164024 237800 164076
rect 384396 164024 384448 164076
rect 404728 164024 404780 164076
rect 570604 164024 570656 164076
rect 226156 163956 226208 164008
rect 324320 163956 324372 164008
rect 346400 163956 346452 164008
rect 560944 163956 560996 164008
rect 137284 163888 137336 163940
rect 360476 163888 360528 163940
rect 384488 163888 384540 163940
rect 552112 163888 552164 163940
rect 110880 163820 110932 163872
rect 278780 163820 278832 163872
rect 305092 163820 305144 163872
rect 550916 163820 550968 163872
rect 43628 163752 43680 163804
rect 260840 163752 260892 163804
rect 302240 163752 302292 163804
rect 551100 163752 551152 163804
rect 35164 163684 35216 163736
rect 214104 163684 214156 163736
rect 222200 163684 222252 163736
rect 546868 163684 546920 163736
rect 212540 163616 212592 163668
rect 541256 163616 541308 163668
rect 184940 163548 184992 163600
rect 540704 163548 540756 163600
rect 29644 163480 29696 163532
rect 460572 163480 460624 163532
rect 395620 163412 395672 163464
rect 510160 163412 510212 163464
rect 414664 162800 414716 162852
rect 420000 162800 420052 162852
rect 351092 162324 351144 162376
rect 377864 162324 377916 162376
rect 266360 162256 266412 162308
rect 356060 162256 356112 162308
rect 382188 162256 382240 162308
rect 400680 162256 400732 162308
rect 285680 162188 285732 162240
rect 403900 162188 403952 162240
rect 127072 162120 127124 162172
rect 383292 162120 383344 162172
rect 406660 162120 406712 162172
rect 551468 162120 551520 162172
rect 389732 161372 389784 161424
rect 549628 161372 549680 161424
rect 378876 161304 378928 161356
rect 545396 161304 545448 161356
rect 371976 161236 372028 161288
rect 552480 161236 552532 161288
rect 248420 161168 248472 161220
rect 376484 161168 376536 161220
rect 396724 161168 396776 161220
rect 580264 161168 580316 161220
rect 221648 161100 221700 161152
rect 356244 161100 356296 161152
rect 391664 161100 391716 161152
rect 578608 161100 578660 161152
rect 142436 161032 142488 161084
rect 361120 161032 361172 161084
rect 365352 161032 365404 161084
rect 560668 161032 560720 161084
rect 320180 160964 320232 161016
rect 578240 160964 578292 161016
rect 56784 160896 56836 160948
rect 358544 160896 358596 160948
rect 375104 160896 375156 160948
rect 578792 160896 578844 160948
rect 39396 160828 39448 160880
rect 240140 160828 240192 160880
rect 253940 160828 253992 160880
rect 581828 160828 581880 160880
rect 219716 160760 219768 160812
rect 566188 160760 566240 160812
rect 178132 160692 178184 160744
rect 553308 160692 553360 160744
rect 282828 160624 282880 160676
rect 426440 160624 426492 160676
rect 405096 160556 405148 160608
rect 548524 160556 548576 160608
rect 155316 159740 155368 159792
rect 388444 159740 388496 159792
rect 96712 159672 96764 159724
rect 366364 159672 366416 159724
rect 402796 159672 402848 159724
rect 549076 159672 549128 159724
rect 252560 159604 252612 159656
rect 546224 159604 546276 159656
rect 168380 159536 168432 159588
rect 480260 159536 480312 159588
rect 121460 159468 121512 159520
rect 454132 159468 454184 159520
rect 216772 159400 216824 159452
rect 553032 159400 553084 159452
rect 3424 159332 3476 159384
rect 359648 159332 359700 159384
rect 379152 159332 379204 159384
rect 539968 159332 540020 159384
rect 292580 158652 292632 158704
rect 439320 158652 439372 158704
rect 268016 158584 268068 158636
rect 349896 158584 349948 158636
rect 383108 158584 383160 158636
rect 540520 158584 540572 158636
rect 150164 158516 150216 158568
rect 359096 158516 359148 158568
rect 368112 158516 368164 158568
rect 539324 158516 539376 158568
rect 92572 158448 92624 158500
rect 320824 158448 320876 158500
rect 386052 158448 386104 158500
rect 559472 158448 559524 158500
rect 282920 158380 282972 158432
rect 540612 158380 540664 158432
rect 305000 158312 305052 158364
rect 571800 158312 571852 158364
rect 259552 158244 259604 158296
rect 552020 158244 552072 158296
rect 231860 158176 231912 158228
rect 539416 158176 539468 158228
rect 155960 158108 156012 158160
rect 481824 158108 481876 158160
rect 158720 158040 158772 158092
rect 551008 158040 551060 158092
rect 28172 157972 28224 158024
rect 559380 157972 559432 158024
rect 394608 157904 394660 157956
rect 537484 157904 537536 157956
rect 264244 157836 264296 157888
rect 406476 157836 406528 157888
rect 398656 157768 398708 157820
rect 537576 157768 537628 157820
rect 400956 157020 401008 157072
rect 551560 157020 551612 157072
rect 166264 156952 166316 157004
rect 188804 156952 188856 157004
rect 259644 156952 259696 157004
rect 309140 156952 309192 157004
rect 398748 156952 398800 157004
rect 556620 156952 556672 157004
rect 47584 156884 47636 156936
rect 204260 156884 204312 156936
rect 271880 156884 271932 156936
rect 368204 156884 368256 156936
rect 381452 156884 381504 156936
rect 571892 156884 571944 156936
rect 45928 156816 45980 156868
rect 361948 156816 362000 156868
rect 375012 156816 375064 156868
rect 574284 156816 574336 156868
rect 80244 156748 80296 156800
rect 281540 156748 281592 156800
rect 318248 156748 318300 156800
rect 328460 156748 328512 156800
rect 333980 156748 334032 156800
rect 541164 156748 541216 156800
rect 78772 156680 78824 156732
rect 323400 156680 323452 156732
rect 328552 156680 328604 156732
rect 558092 156680 558144 156732
rect 59360 156612 59412 156664
rect 59636 156612 59688 156664
rect 124312 156612 124364 156664
rect 574468 156612 574520 156664
rect 376760 156544 376812 156596
rect 377220 156544 377272 156596
rect 254584 155864 254636 155916
rect 369124 155864 369176 155916
rect 383476 155864 383528 155916
rect 537116 155864 537168 155916
rect 538956 155864 539008 155916
rect 539508 155864 539560 155916
rect 109684 155796 109736 155848
rect 161756 155796 161808 155848
rect 232596 155796 232648 155848
rect 348424 155796 348476 155848
rect 409788 155796 409840 155848
rect 565084 155796 565136 155848
rect 47952 155728 48004 155780
rect 136640 155728 136692 155780
rect 179420 155728 179472 155780
rect 229376 155728 229428 155780
rect 230020 155728 230072 155780
rect 355324 155728 355376 155780
rect 401416 155728 401468 155780
rect 557816 155728 557868 155780
rect 56048 155660 56100 155712
rect 154580 155660 154632 155712
rect 205640 155660 205692 155712
rect 360936 155660 360988 155712
rect 409604 155660 409656 155712
rect 567384 155660 567436 155712
rect 40960 155592 41012 155644
rect 238760 155592 238812 155644
rect 292488 155592 292540 155644
rect 349988 155592 350040 155644
rect 353944 155592 353996 155644
rect 554136 155592 554188 155644
rect 57612 155524 57664 155576
rect 361672 155524 361724 155576
rect 394424 155524 394476 155576
rect 555056 155524 555108 155576
rect 32220 155456 32272 155508
rect 284116 155456 284168 155508
rect 338120 155456 338172 155508
rect 562232 155456 562284 155508
rect 57704 155388 57756 155440
rect 372344 155388 372396 155440
rect 390468 155388 390520 155440
rect 565360 155388 565412 155440
rect 43628 155320 43680 155372
rect 368572 155320 368624 155372
rect 370504 155320 370556 155372
rect 576124 155320 576176 155372
rect 46388 155252 46440 155304
rect 162860 155252 162912 155304
rect 216680 155252 216732 155304
rect 547788 155252 547840 155304
rect 32588 155184 32640 155236
rect 396172 155184 396224 155236
rect 408316 155184 408368 155236
rect 570512 155184 570564 155236
rect 295708 155116 295760 155168
rect 350540 155116 350592 155168
rect 405372 155116 405424 155168
rect 556436 155116 556488 155168
rect 269120 155048 269172 155100
rect 322756 155048 322808 155100
rect 403992 155048 404044 155100
rect 553952 155048 554004 155100
rect 309232 154980 309284 155032
rect 357164 154980 357216 155032
rect 410156 154980 410208 155032
rect 538956 154980 539008 155032
rect 405188 154504 405240 154556
rect 542728 154504 542780 154556
rect 397000 154436 397052 154488
rect 542636 154436 542688 154488
rect 382096 154368 382148 154420
rect 539600 154368 539652 154420
rect 409696 154300 409748 154352
rect 569316 154300 569368 154352
rect 260288 154232 260340 154284
rect 299480 154232 299532 154284
rect 373264 154232 373316 154284
rect 542452 154232 542504 154284
rect 175280 154164 175332 154216
rect 289820 154164 289872 154216
rect 291200 154164 291252 154216
rect 340144 154164 340196 154216
rect 397092 154164 397144 154216
rect 573456 154164 573508 154216
rect 106280 154096 106332 154148
rect 308588 154096 308640 154148
rect 313740 154096 313792 154148
rect 377312 154096 377364 154148
rect 387064 154096 387116 154148
rect 572168 154096 572220 154148
rect 73252 154028 73304 154080
rect 223948 154028 224000 154080
rect 224868 154028 224920 154080
rect 581460 154028 581512 154080
rect 91100 153960 91152 154012
rect 166908 153960 166960 154012
rect 178040 153960 178092 154012
rect 544200 153960 544252 154012
rect 31024 153892 31076 153944
rect 519820 153892 519872 153944
rect 33876 153824 33928 153876
rect 548432 153824 548484 153876
rect 251916 153212 251968 153264
rect 259460 153212 259512 153264
rect 37740 153144 37792 153196
rect 129556 153144 129608 153196
rect 135996 153144 136048 153196
rect 224224 153144 224276 153196
rect 291200 153144 291252 153196
rect 348700 153144 348752 153196
rect 385776 153144 385828 153196
rect 391664 153144 391716 153196
rect 402704 153144 402756 153196
rect 580172 153144 580224 153196
rect 46112 153076 46164 153128
rect 141148 153076 141200 153128
rect 145012 153076 145064 153128
rect 178132 153076 178184 153128
rect 179788 153076 179840 153128
rect 216772 153076 216824 153128
rect 254492 153076 254544 153128
rect 373448 153076 373500 153128
rect 378784 153076 378836 153128
rect 414848 153076 414900 153128
rect 482928 153076 482980 153128
rect 555424 153076 555476 153128
rect 56600 153008 56652 153060
rect 208492 153008 208544 153060
rect 209412 153008 209464 153060
rect 354680 153008 354732 153060
rect 354772 153008 354824 153060
rect 363604 153008 363656 153060
rect 403624 153008 403676 153060
rect 448980 153008 449032 153060
rect 499672 153008 499724 153060
rect 580356 153008 580408 153060
rect 38384 152940 38436 152992
rect 209780 152940 209832 152992
rect 213920 152940 213972 152992
rect 384304 152940 384356 152992
rect 394056 152940 394108 152992
rect 447692 152940 447744 152992
rect 462412 152940 462464 152992
rect 563336 152940 563388 152992
rect 51356 152872 51408 152924
rect 126980 152872 127032 152924
rect 127624 152872 127676 152924
rect 315304 152872 315356 152924
rect 316592 152872 316644 152924
rect 360292 152872 360344 152924
rect 364984 152872 365036 152924
rect 421932 152872 421984 152924
rect 451280 152872 451332 152924
rect 561864 152872 561916 152924
rect 44916 152804 44968 152856
rect 160100 152804 160152 152856
rect 200396 152804 200448 152856
rect 392584 152804 392636 152856
rect 398196 152804 398248 152856
rect 529204 152804 529256 152856
rect 531412 152804 531464 152856
rect 534724 152804 534776 152856
rect 536104 152804 536156 152856
rect 539784 152804 539836 152856
rect 543096 152804 543148 152856
rect 561680 152804 561732 152856
rect 26976 152736 27028 152788
rect 107660 152736 107712 152788
rect 122748 152736 122800 152788
rect 330484 152736 330536 152788
rect 334992 152736 335044 152788
rect 354772 152736 354824 152788
rect 354864 152736 354916 152788
rect 358912 152736 358964 152788
rect 395436 152736 395488 152788
rect 543832 152736 543884 152788
rect 547236 152736 547288 152788
rect 566372 152736 566424 152788
rect 50344 152668 50396 152720
rect 82544 152668 82596 152720
rect 106372 152668 106424 152720
rect 358176 152668 358228 152720
rect 406016 152668 406068 152720
rect 555332 152668 555384 152720
rect 35072 152600 35124 152652
rect 297640 152600 297692 152652
rect 310520 152600 310572 152652
rect 354864 152600 354916 152652
rect 354956 152600 355008 152652
rect 362224 152600 362276 152652
rect 405464 152600 405516 152652
rect 560760 152600 560812 152652
rect 36360 152532 36412 152584
rect 326620 152532 326672 152584
rect 327264 152532 327316 152584
rect 357624 152532 357676 152584
rect 401508 152532 401560 152584
rect 561312 152532 561364 152584
rect 28356 152464 28408 152516
rect 67088 152464 67140 152516
rect 81256 152464 81308 152516
rect 377496 152464 377548 152516
rect 403532 152464 403584 152516
rect 580448 152464 580500 152516
rect 52000 152396 52052 152448
rect 57980 152396 58032 152448
rect 58164 152396 58216 152448
rect 111800 152396 111852 152448
rect 315028 152396 315080 152448
rect 359464 152396 359516 152448
rect 389916 152396 389968 152448
rect 425152 152396 425204 152448
rect 498200 152396 498252 152448
rect 557540 152396 557592 152448
rect 44364 152328 44416 152380
rect 76748 152328 76800 152380
rect 94780 152328 94832 152380
rect 121460 152328 121512 152380
rect 344008 152328 344060 152380
rect 360200 152328 360252 152380
rect 399484 152328 399536 152380
rect 434168 152328 434220 152380
rect 503076 152328 503128 152380
rect 538864 152328 538916 152380
rect 540428 152328 540480 152380
rect 543372 152328 543424 152380
rect 61292 152260 61344 152312
rect 68284 152260 68336 152312
rect 347872 152260 347924 152312
rect 358820 152260 358872 152312
rect 392768 152260 392820 152312
rect 410340 152260 410392 152312
rect 505652 152260 505704 152312
rect 518164 152260 518216 152312
rect 529204 152260 529256 152312
rect 534632 152260 534684 152312
rect 68744 152192 68796 152244
rect 69664 152192 69716 152244
rect 342076 152192 342128 152244
rect 350724 152192 350776 152244
rect 526444 151920 526496 151972
rect 528836 151920 528888 151972
rect 402336 151852 402388 151904
rect 403256 151852 403308 151904
rect 50620 151716 50672 151768
rect 96620 151716 96672 151768
rect 385500 151716 385552 151768
rect 549168 151716 549220 151768
rect 52736 151648 52788 151700
rect 113180 151648 113232 151700
rect 381912 151648 381964 151700
rect 540980 151648 541032 151700
rect 59452 151580 59504 151632
rect 198740 151580 198792 151632
rect 306380 151580 306432 151632
rect 543740 151580 543792 151632
rect 52092 151512 52144 151564
rect 113272 151512 113324 151564
rect 119896 151512 119948 151564
rect 366180 151512 366232 151564
rect 399852 151512 399904 151564
rect 564992 151512 565044 151564
rect 45284 151444 45336 151496
rect 356336 151444 356388 151496
rect 381820 151444 381872 151496
rect 549352 151444 549404 151496
rect 43996 151376 44048 151428
rect 368756 151376 368808 151428
rect 392676 151376 392728 151428
rect 569224 151376 569276 151428
rect 48044 151308 48096 151360
rect 387800 151308 387852 151360
rect 395804 151308 395856 151360
rect 573272 151308 573324 151360
rect 380348 151240 380400 151292
rect 559840 151240 559892 151292
rect 46112 151172 46164 151224
rect 412640 151172 412692 151224
rect 518900 151172 518952 151224
rect 556896 151172 556948 151224
rect 50528 151104 50580 151156
rect 75920 151104 75972 151156
rect 80060 151104 80112 151156
rect 552388 151104 552440 151156
rect 28264 151036 28316 151088
rect 572720 151036 572772 151088
rect 49148 150968 49200 151020
rect 70492 150968 70544 151020
rect 407304 150968 407356 151020
rect 567200 150968 567252 151020
rect 58992 150900 59044 150952
rect 78680 150900 78732 150952
rect 383200 150900 383252 150952
rect 537392 150900 537444 150952
rect 49240 150832 49292 150884
rect 60740 150832 60792 150884
rect 537116 150832 537168 150884
rect 540888 150832 540940 150884
rect 25504 150764 25556 150816
rect 380716 150764 380768 150816
rect 539048 150424 539100 150476
rect 540152 150424 540204 150476
rect 397184 150356 397236 150408
rect 538864 150356 538916 150408
rect 539508 150356 539560 150408
rect 539876 150356 539928 150408
rect 540704 150356 540756 150408
rect 542176 150356 542228 150408
rect 537484 150288 537536 150340
rect 540428 150288 540480 150340
rect 539416 150220 539468 150272
rect 545304 150356 545356 150408
rect 54392 150152 54444 150204
rect 59544 150152 59596 150204
rect 538956 150152 539008 150204
rect 545580 150152 545632 150204
rect 48780 150084 48832 150136
rect 59912 150084 59964 150136
rect 539600 150084 539652 150136
rect 551192 150084 551244 150136
rect 57336 150016 57388 150068
rect 255320 150016 255372 150068
rect 59268 149948 59320 150000
rect 293960 149948 294012 150000
rect 52920 149880 52972 149932
rect 313280 149880 313332 149932
rect 51264 149812 51316 149864
rect 366824 149880 366876 149932
rect 50160 149744 50212 149796
rect 387432 149880 387484 149932
rect 488540 149880 488592 149932
rect 523592 150016 523644 150068
rect 3332 149676 3384 149728
rect 523592 149880 523644 149932
rect 537392 149948 537444 150000
rect 543188 149948 543240 150000
rect 538772 149880 538824 149932
rect 539048 149880 539100 149932
rect 539416 149880 539468 149932
rect 550640 149880 550692 149932
rect 540704 149812 540756 149864
rect 546040 149812 546092 149864
rect 560392 149812 560444 149864
rect 549812 149744 549864 149796
rect 551376 149744 551428 149796
rect 565452 149744 565504 149796
rect 543556 149676 543608 149728
rect 565820 149676 565872 149728
rect 546132 148996 546184 149048
rect 548708 148996 548760 149048
rect 547788 148316 547840 148368
rect 568580 148316 568632 148368
rect 541900 148248 541952 148300
rect 545488 148248 545540 148300
rect 547144 147636 547196 147688
rect 547972 147636 548024 147688
rect 540704 147568 540756 147620
rect 542268 147568 542320 147620
rect 543464 147568 543516 147620
rect 564532 147568 564584 147620
rect 552848 147500 552900 147552
rect 559748 147500 559800 147552
rect 542176 146956 542228 147008
rect 542912 146956 542964 147008
rect 540888 146888 540940 146940
rect 545028 146888 545080 146940
rect 555608 146888 555660 146940
rect 564532 146888 564584 146940
rect 55128 146344 55180 146396
rect 59544 146344 59596 146396
rect 58532 146276 58584 146328
rect 59452 146276 59504 146328
rect 542820 146208 542872 146260
rect 543832 146208 543884 146260
rect 546500 146140 546552 146192
rect 548248 146140 548300 146192
rect 53472 146072 53524 146124
rect 58440 146072 58492 146124
rect 543280 146072 543332 146124
rect 547972 146072 548024 146124
rect 547236 146004 547288 146056
rect 548248 146004 548300 146056
rect 546960 145868 547012 145920
rect 547236 145868 547288 145920
rect 57428 144984 57480 145036
rect 59360 144984 59412 145036
rect 541348 144848 541400 144900
rect 542360 144848 542412 144900
rect 544384 144848 544436 144900
rect 546960 144848 547012 144900
rect 542268 144508 542320 144560
rect 546776 144508 546828 144560
rect 541716 144372 541768 144424
rect 546776 144372 546828 144424
rect 544568 144236 544620 144288
rect 560392 144236 560444 144288
rect 543004 144168 543056 144220
rect 560852 144168 560904 144220
rect 545028 144100 545080 144152
rect 547788 144100 547840 144152
rect 543096 144032 543148 144084
rect 546500 144032 546552 144084
rect 51632 143488 51684 143540
rect 55128 143556 55180 143608
rect 543280 143488 543332 143540
rect 558920 143488 558972 143540
rect 542544 143420 542596 143472
rect 543740 143420 543792 143472
rect 542912 143352 542964 143404
rect 545120 143352 545172 143404
rect 543372 142536 543424 142588
rect 548616 142536 548668 142588
rect 543464 142332 543516 142384
rect 548156 142332 548208 142384
rect 53840 142128 53892 142180
rect 55680 142128 55732 142180
rect 47860 142060 47912 142112
rect 56692 142060 56744 142112
rect 57796 142060 57848 142112
rect 59084 142060 59136 142112
rect 543556 142060 543608 142112
rect 569132 142060 569184 142112
rect 542912 141652 542964 141704
rect 545396 141652 545448 141704
rect 547420 141380 547472 141432
rect 550732 141380 550784 141432
rect 546592 140904 546644 140956
rect 547052 140904 547104 140956
rect 559564 140904 559616 140956
rect 561128 140904 561180 140956
rect 547236 140836 547288 140888
rect 547880 140836 547932 140888
rect 558276 140836 558328 140888
rect 560300 140836 560352 140888
rect 51264 140768 51316 140820
rect 55220 140768 55272 140820
rect 541808 140768 541860 140820
rect 547052 140768 547104 140820
rect 547788 140768 547840 140820
rect 548708 140768 548760 140820
rect 558368 140768 558420 140820
rect 558920 140768 558972 140820
rect 32496 140700 32548 140752
rect 56692 140700 56744 140752
rect 54576 140632 54628 140684
rect 57244 140632 57296 140684
rect 545948 140428 546000 140480
rect 548156 140428 548208 140480
rect 542820 140020 542872 140072
rect 544108 140020 544160 140072
rect 47860 139408 47912 139460
rect 48780 139408 48832 139460
rect 543372 139408 543424 139460
rect 544568 139408 544620 139460
rect 544936 139408 544988 139460
rect 545580 139408 545632 139460
rect 551928 139408 551980 139460
rect 555516 139408 555568 139460
rect 543556 139340 543608 139392
rect 559380 139340 559432 139392
rect 567936 139340 567988 139392
rect 580540 139340 580592 139392
rect 549720 139272 549772 139324
rect 555516 139272 555568 139324
rect 544660 139204 544712 139256
rect 547972 139204 548024 139256
rect 51724 138728 51776 138780
rect 52460 138728 52512 138780
rect 545028 137980 545080 138032
rect 545396 137980 545448 138032
rect 17684 137912 17736 137964
rect 57612 137912 57664 137964
rect 559748 137708 559800 137760
rect 566464 137708 566516 137760
rect 559564 137300 559616 137352
rect 566648 137300 566700 137352
rect 54576 137232 54628 137284
rect 55220 137232 55272 137284
rect 542452 136620 542504 136672
rect 542912 136620 542964 136672
rect 542820 136552 542872 136604
rect 564624 136552 564676 136604
rect 58716 136484 58768 136536
rect 58900 136484 58952 136536
rect 542452 136484 542504 136536
rect 557540 136484 557592 136536
rect 544384 136416 544436 136468
rect 547880 136416 547932 136468
rect 544936 136348 544988 136400
rect 549260 136348 549312 136400
rect 53564 135872 53616 135924
rect 57980 135872 58032 135924
rect 542268 135260 542320 135312
rect 544660 135260 544712 135312
rect 26148 135192 26200 135244
rect 57612 135192 57664 135244
rect 58440 135192 58492 135244
rect 59360 135192 59412 135244
rect 542452 135192 542504 135244
rect 572720 135192 572772 135244
rect 541992 135124 542044 135176
rect 546684 135124 546736 135176
rect 548616 135124 548668 135176
rect 549352 135124 549404 135176
rect 561036 135124 561088 135176
rect 564440 135124 564492 135176
rect 558460 135056 558512 135108
rect 563060 135056 563112 135108
rect 549996 134580 550048 134632
rect 560300 134580 560352 134632
rect 545028 134512 545080 134564
rect 556160 134512 556212 134564
rect 58716 134376 58768 134428
rect 59268 134376 59320 134428
rect 543648 134240 543700 134292
rect 547880 134240 547932 134292
rect 540244 134036 540296 134088
rect 541716 134036 541768 134088
rect 541624 133968 541676 134020
rect 546592 133968 546644 134020
rect 558184 133968 558236 134020
rect 563888 133968 563940 134020
rect 540612 133900 540664 133952
rect 541440 133900 541492 133952
rect 43076 133832 43128 133884
rect 57612 133832 57664 133884
rect 540428 133152 540480 133204
rect 540980 133152 541032 133204
rect 542084 132744 542136 132796
rect 546960 132744 547012 132796
rect 541992 132608 542044 132660
rect 549260 132608 549312 132660
rect 541900 132472 541952 132524
rect 542820 132472 542872 132524
rect 47400 132404 47452 132456
rect 57612 132404 57664 132456
rect 542452 132404 542504 132456
rect 578240 132404 578292 132456
rect 541348 131112 541400 131164
rect 543740 131112 543792 131164
rect 36452 131044 36504 131096
rect 57612 131044 57664 131096
rect 541072 131044 541124 131096
rect 541532 131044 541584 131096
rect 542452 131044 542504 131096
rect 568580 131044 568632 131096
rect 542176 130976 542228 131028
rect 543464 130976 543516 131028
rect 541716 130840 541768 130892
rect 542176 130840 542228 130892
rect 541716 130704 541768 130756
rect 543648 130704 543700 130756
rect 541808 130364 541860 130416
rect 541992 130364 542044 130416
rect 541348 130296 541400 130348
rect 548524 130296 548576 130348
rect 540244 129820 540296 129872
rect 545488 129820 545540 129872
rect 548064 129752 548116 129804
rect 549352 129752 549404 129804
rect 549996 129752 550048 129804
rect 550640 129752 550692 129804
rect 50068 129684 50120 129736
rect 57612 129684 57664 129736
rect 540888 129684 540940 129736
rect 541808 129684 541860 129736
rect 542452 129684 542504 129736
rect 561680 129684 561732 129736
rect 546500 129616 546552 129668
rect 548156 129616 548208 129668
rect 546408 129140 546460 129192
rect 552020 129140 552072 129192
rect 542268 129072 542320 129124
rect 549720 129072 549772 129124
rect 540336 129004 540388 129056
rect 549352 129004 549404 129056
rect 56692 128800 56744 128852
rect 58532 128800 58584 128852
rect 544292 128324 544344 128376
rect 545120 128324 545172 128376
rect 548616 128324 548668 128376
rect 549812 128324 549864 128376
rect 36820 128256 36872 128308
rect 57612 128256 57664 128308
rect 543556 128256 543608 128308
rect 547696 128188 547748 128240
rect 547880 128188 547932 128240
rect 567200 128188 567252 128240
rect 543832 127644 543884 127696
rect 544108 127644 544160 127696
rect 58348 127576 58400 127628
rect 59360 127576 59412 127628
rect 541900 127576 541952 127628
rect 562416 127576 562468 127628
rect 564532 127576 564584 127628
rect 541992 127372 542044 127424
rect 545028 126964 545080 127016
rect 546500 126964 546552 127016
rect 50988 126896 51040 126948
rect 51724 126896 51776 126948
rect 54668 126896 54720 126948
rect 57612 126896 57664 126948
rect 57796 126896 57848 126948
rect 58716 126896 58768 126948
rect 543648 126896 543700 126948
rect 546868 126896 546920 126948
rect 562508 126896 562560 126948
rect 565820 126896 565872 126948
rect 544476 126828 544528 126880
rect 548156 126828 548208 126880
rect 540796 126760 540848 126812
rect 544936 126760 544988 126812
rect 55128 126352 55180 126404
rect 56692 126352 56744 126404
rect 540796 126216 540848 126268
rect 543096 126216 543148 126268
rect 540336 125808 540388 125860
rect 541624 125808 541676 125860
rect 541348 125604 541400 125656
rect 541716 125604 541768 125656
rect 542544 125536 542596 125588
rect 544016 125536 544068 125588
rect 545212 125536 545264 125588
rect 546868 125536 546920 125588
rect 543556 125468 543608 125520
rect 570788 125468 570840 125520
rect 540888 125400 540940 125452
rect 544476 125400 544528 125452
rect 542452 125332 542504 125384
rect 544108 125332 544160 125384
rect 58716 125264 58768 125316
rect 59452 125264 59504 125316
rect 540428 125264 540480 125316
rect 543832 125264 543884 125316
rect 51724 125060 51776 125112
rect 56600 125060 56652 125112
rect 50436 124924 50488 124976
rect 56692 124924 56744 124976
rect 545948 124856 546000 124908
rect 566464 124856 566516 124908
rect 57152 124584 57204 124636
rect 58624 124584 58676 124636
rect 546040 124244 546092 124296
rect 547972 124244 548024 124296
rect 23020 124108 23072 124160
rect 57612 124108 57664 124160
rect 59084 124108 59136 124160
rect 59360 124108 59412 124160
rect 544384 124176 544436 124228
rect 541992 123972 542044 124024
rect 541348 123904 541400 123956
rect 543740 123904 543792 123956
rect 53656 123564 53708 123616
rect 57980 123564 58032 123616
rect 53288 123496 53340 123548
rect 58624 123496 58676 123548
rect 52368 123428 52420 123480
rect 57888 123428 57940 123480
rect 544384 123428 544436 123480
rect 552756 123428 552808 123480
rect 53748 123224 53800 123276
rect 54576 123224 54628 123276
rect 57612 123156 57664 123208
rect 57796 123156 57848 123208
rect 547144 122816 547196 122868
rect 547880 122816 547932 122868
rect 543648 122748 543700 122800
rect 559472 122748 559524 122800
rect 57428 121524 57480 121576
rect 38016 121388 38068 121440
rect 57428 121388 57480 121440
rect 540704 121456 540756 121508
rect 541992 121456 542044 121508
rect 550088 121456 550140 121508
rect 550640 121456 550692 121508
rect 57888 121388 57940 121440
rect 58900 121388 58952 121440
rect 543556 121388 543608 121440
rect 558092 121388 558144 121440
rect 59452 121320 59504 121372
rect 543004 120708 543056 120760
rect 546776 120708 546828 120760
rect 57336 120164 57388 120216
rect 59636 120164 59688 120216
rect 57796 120096 57848 120148
rect 59820 120096 59872 120148
rect 55128 120028 55180 120080
rect 56692 120028 56744 120080
rect 54760 119960 54812 120012
rect 57428 119960 57480 120012
rect 50988 119416 51040 119468
rect 54576 119416 54628 119468
rect 51816 117988 51868 118040
rect 53932 117988 53984 118040
rect 544292 117988 544344 118040
rect 546592 117988 546644 118040
rect 53196 117648 53248 117700
rect 54392 117648 54444 117700
rect 50436 117580 50488 117632
rect 53840 117580 53892 117632
rect 543648 117308 543700 117360
rect 547420 117308 547472 117360
rect 23112 117240 23164 117292
rect 57060 117240 57112 117292
rect 59268 117240 59320 117292
rect 59544 117240 59596 117292
rect 542452 117240 542504 117292
rect 556896 117240 556948 117292
rect 544568 117172 544620 117224
rect 545120 117172 545172 117224
rect 546132 117172 546184 117224
rect 547696 117172 547748 117224
rect 547788 117172 547840 117224
rect 549812 117172 549864 117224
rect 542728 117104 542780 117156
rect 546776 117104 546828 117156
rect 57888 117036 57940 117088
rect 59452 117036 59504 117088
rect 59268 116968 59320 117020
rect 59636 116968 59688 117020
rect 53748 116560 53800 116612
rect 57980 116560 58032 116612
rect 540520 115948 540572 116000
rect 541072 115948 541124 116000
rect 44640 115880 44692 115932
rect 57428 115880 57480 115932
rect 544476 115880 544528 115932
rect 545580 115880 545632 115932
rect 555516 115880 555568 115932
rect 556896 115880 556948 115932
rect 543280 115812 543332 115864
rect 546040 115812 546092 115864
rect 542084 115744 542136 115796
rect 545488 115744 545540 115796
rect 542728 114792 542780 114844
rect 547328 114792 547380 114844
rect 547144 114520 547196 114572
rect 549352 114520 549404 114572
rect 44732 114452 44784 114504
rect 57428 114452 57480 114504
rect 552020 114452 552072 114504
rect 555516 114452 555568 114504
rect 549352 114384 549404 114436
rect 549720 114384 549772 114436
rect 543372 113840 543424 113892
rect 553308 113840 553360 113892
rect 543096 113772 543148 113824
rect 564440 113772 564492 113824
rect 542452 113568 542504 113620
rect 548340 113568 548392 113620
rect 542268 113160 542320 113212
rect 549260 113160 549312 113212
rect 543648 113092 543700 113144
rect 545212 113092 545264 113144
rect 576216 113092 576268 113144
rect 580540 113092 580592 113144
rect 548708 112480 548760 112532
rect 560300 112480 560352 112532
rect 54576 112412 54628 112464
rect 57244 112412 57296 112464
rect 550088 112412 550140 112464
rect 563060 112412 563112 112464
rect 540428 112004 540480 112056
rect 544108 112004 544160 112056
rect 547052 111868 547104 111920
rect 549352 111868 549404 111920
rect 541808 111800 541860 111852
rect 543740 111800 543792 111852
rect 547236 111800 547288 111852
rect 547880 111800 547932 111852
rect 548892 111800 548944 111852
rect 550640 111800 550692 111852
rect 565176 111800 565228 111852
rect 565820 111800 565872 111852
rect 546132 111732 546184 111784
rect 548800 111732 548852 111784
rect 549720 111732 549772 111784
rect 551376 111732 551428 111784
rect 53748 111188 53800 111240
rect 59360 111188 59412 111240
rect 53656 111120 53708 111172
rect 59636 111120 59688 111172
rect 54760 111052 54812 111104
rect 56692 111052 56744 111104
rect 543188 111052 543240 111104
rect 548248 111052 548300 111104
rect 553308 110984 553360 111036
rect 556160 110984 556212 111036
rect 541716 110508 541768 110560
rect 546960 110508 547012 110560
rect 540428 110440 540480 110492
rect 544936 110440 544988 110492
rect 51632 110372 51684 110424
rect 57336 110372 57388 110424
rect 542452 110372 542504 110424
rect 572168 110372 572220 110424
rect 542268 110304 542320 110356
rect 542912 110304 542964 110356
rect 543004 110304 543056 110356
rect 543648 110304 543700 110356
rect 545396 110304 545448 110356
rect 546500 110304 546552 110356
rect 543740 110236 543792 110288
rect 547880 110236 547932 110288
rect 540888 109896 540940 109948
rect 541440 109896 541492 109948
rect 540796 109556 540848 109608
rect 542452 109556 542504 109608
rect 542544 109420 542596 109472
rect 548432 109420 548484 109472
rect 542636 109352 542688 109404
rect 542636 109012 542688 109064
rect 543280 109012 543332 109064
rect 546868 109012 546920 109064
rect 55772 108944 55824 108996
rect 56600 108944 56652 108996
rect 48964 108876 49016 108928
rect 57520 108876 57572 108928
rect 48872 108808 48924 108860
rect 57428 108808 57480 108860
rect 540704 108808 540756 108860
rect 543648 108808 543700 108860
rect 47860 107584 47912 107636
rect 48964 107584 49016 107636
rect 543188 107584 543240 107636
rect 562232 107584 562284 107636
rect 541900 106904 541952 106956
rect 544568 106904 544620 106956
rect 545028 106224 545080 106276
rect 546500 106224 546552 106276
rect 542268 106156 542320 106208
rect 546960 106156 547012 106208
rect 543188 105544 543240 105596
rect 546592 105544 546644 105596
rect 543372 104864 543424 104916
rect 40592 104796 40644 104848
rect 57520 104796 57572 104848
rect 548248 104796 548300 104848
rect 53380 104728 53432 104780
rect 56876 104728 56928 104780
rect 543740 104592 543792 104644
rect 549720 104592 549772 104644
rect 543280 103572 543332 103624
rect 548892 103572 548944 103624
rect 547788 103504 547840 103556
rect 549812 103504 549864 103556
rect 23204 103436 23256 103488
rect 57520 103436 57572 103488
rect 27436 103368 27488 103420
rect 57888 103368 57940 103420
rect 542176 102620 542228 102672
rect 546868 102620 546920 102672
rect 50160 102212 50212 102264
rect 52460 102212 52512 102264
rect 53288 102144 53340 102196
rect 53932 102144 53984 102196
rect 543464 102144 543516 102196
rect 544476 102144 544528 102196
rect 43260 102076 43312 102128
rect 57520 102076 57572 102128
rect 552664 101396 552716 101448
rect 565452 101396 565504 101448
rect 31668 100648 31720 100700
rect 57520 100648 57572 100700
rect 58808 100104 58860 100156
rect 59084 100104 59136 100156
rect 542084 99968 542136 100020
rect 549260 99968 549312 100020
rect 59268 98676 59320 98728
rect 59820 98676 59872 98728
rect 548800 98676 548852 98728
rect 549260 98676 549312 98728
rect 58440 98608 58492 98660
rect 59452 98608 59504 98660
rect 58716 98540 58768 98592
rect 59544 98540 59596 98592
rect 543556 97928 543608 97980
rect 575480 97928 575532 97980
rect 52460 97860 52512 97912
rect 55864 97860 55916 97912
rect 2872 97724 2924 97776
rect 4804 97724 4856 97776
rect 53380 96568 53432 96620
rect 53840 96568 53892 96620
rect 540980 96568 541032 96620
rect 543464 96568 543516 96620
rect 543648 96568 543700 96620
rect 578792 96568 578844 96620
rect 543556 96500 543608 96552
rect 577228 96500 577280 96552
rect 542176 95888 542228 95940
rect 551192 95888 551244 95940
rect 30932 95140 30984 95192
rect 57520 95140 57572 95192
rect 540612 95140 540664 95192
rect 542268 95140 542320 95192
rect 543556 95140 543608 95192
rect 581828 95140 581880 95192
rect 53196 95072 53248 95124
rect 54576 95072 54628 95124
rect 50252 93780 50304 93832
rect 57520 93780 57572 93832
rect 543556 93780 543608 93832
rect 552572 93780 552624 93832
rect 541992 92624 542044 92676
rect 542452 92624 542504 92676
rect 542268 92488 542320 92540
rect 542452 92488 542504 92540
rect 551376 92488 551428 92540
rect 552020 92488 552072 92540
rect 543556 92420 543608 92472
rect 574928 92420 574980 92472
rect 542820 92216 542872 92268
rect 547972 92216 548024 92268
rect 542636 92148 542688 92200
rect 544292 92148 544344 92200
rect 546408 91740 546460 91792
rect 551192 91740 551244 91792
rect 551376 91740 551428 91792
rect 565176 91740 565228 91792
rect 542820 91128 542872 91180
rect 547880 91128 547932 91180
rect 546040 90312 546092 90364
rect 556160 90312 556212 90364
rect 543648 89700 543700 89752
rect 545580 89700 545632 89752
rect 546132 89700 546184 89752
rect 547052 89700 547104 89752
rect 34428 89632 34480 89684
rect 57612 89632 57664 89684
rect 542728 89632 542780 89684
rect 569316 89632 569368 89684
rect 545028 89428 545080 89480
rect 547328 89428 547380 89480
rect 544476 89020 544528 89072
rect 547420 89020 547472 89072
rect 541348 88272 541400 88324
rect 544292 88272 544344 88324
rect 542268 88204 542320 88256
rect 547236 88340 547288 88392
rect 38200 86912 38252 86964
rect 57612 86912 57664 86964
rect 3516 85484 3568 85536
rect 21364 85484 21416 85536
rect 58256 85484 58308 85536
rect 58440 85484 58492 85536
rect 543648 85484 543700 85536
rect 544936 85484 544988 85536
rect 57520 85416 57572 85468
rect 58532 85416 58584 85468
rect 542636 85076 542688 85128
rect 544200 85076 544252 85128
rect 542176 84940 542228 84992
rect 549812 84940 549864 84992
rect 55128 84192 55180 84244
rect 57060 84192 57112 84244
rect 547236 84192 547288 84244
rect 550088 84192 550140 84244
rect 57152 84124 57204 84176
rect 58256 84124 58308 84176
rect 57796 83920 57848 83972
rect 57796 83716 57848 83768
rect 54668 83648 54720 83700
rect 57704 83648 57756 83700
rect 548800 83444 548852 83496
rect 561128 83444 561180 83496
rect 543464 82968 543516 83020
rect 547972 82968 548024 83020
rect 543648 82900 543700 82952
rect 546132 82900 546184 82952
rect 541440 82832 541492 82884
rect 542452 82832 542504 82884
rect 542820 82832 542872 82884
rect 544476 82832 544528 82884
rect 547420 82832 547472 82884
rect 548892 82832 548944 82884
rect 17868 82764 17920 82816
rect 57612 82764 57664 82816
rect 543556 82764 543608 82816
rect 567752 82764 567804 82816
rect 47676 82696 47728 82748
rect 57520 82696 57572 82748
rect 542084 82560 542136 82612
rect 543832 82560 543884 82612
rect 544936 82152 544988 82204
rect 547880 82152 547932 82204
rect 540612 82084 540664 82136
rect 548248 82084 548300 82136
rect 552756 80044 552808 80096
rect 555516 80044 555568 80096
rect 57888 79364 57940 79416
rect 59636 79364 59688 79416
rect 57704 79296 57756 79348
rect 57980 79296 58032 79348
rect 543556 78616 543608 78668
rect 551284 78616 551336 78668
rect 543556 77188 543608 77240
rect 580356 77188 580408 77240
rect 551284 76236 551336 76288
rect 556896 76236 556948 76288
rect 51908 75828 51960 75880
rect 57612 75828 57664 75880
rect 543556 75828 543608 75880
rect 571892 75828 571944 75880
rect 55772 75760 55824 75812
rect 57152 75760 57204 75812
rect 542636 75692 542688 75744
rect 545856 75692 545908 75744
rect 57612 75556 57664 75608
rect 57888 75556 57940 75608
rect 540520 75148 540572 75200
rect 547880 75148 547932 75200
rect 574744 73108 574796 73160
rect 580356 73108 580408 73160
rect 543556 71680 543608 71732
rect 582656 71680 582708 71732
rect 547328 71612 547380 71664
rect 550088 71612 550140 71664
rect 546500 71408 546552 71460
rect 549260 71408 549312 71460
rect 543556 70320 543608 70372
rect 566556 70320 566608 70372
rect 42616 69640 42668 69692
rect 57060 69640 57112 69692
rect 542268 69232 542320 69284
rect 543372 69232 543424 69284
rect 38292 68960 38344 69012
rect 57888 68960 57940 69012
rect 39028 68892 39080 68944
rect 57152 68892 57204 68944
rect 53288 68824 53340 68876
rect 55956 68824 56008 68876
rect 40776 67532 40828 67584
rect 57888 67532 57940 67584
rect 544568 67328 544620 67380
rect 546500 67328 546552 67380
rect 542820 66172 542872 66224
rect 582748 66172 582800 66224
rect 543556 66104 543608 66156
rect 578332 66104 578384 66156
rect 543648 66036 543700 66088
rect 547052 66036 547104 66088
rect 33784 64812 33836 64864
rect 57888 64812 57940 64864
rect 543556 63928 543608 63980
rect 549628 63928 549680 63980
rect 49056 63452 49108 63504
rect 57888 63452 57940 63504
rect 548892 63316 548944 63368
rect 549628 63316 549680 63368
rect 42708 62024 42760 62076
rect 57888 62024 57940 62076
rect 543556 62024 543608 62076
rect 560944 62024 560996 62076
rect 543648 61956 543700 62008
rect 551100 61956 551152 62008
rect 571984 60664 572036 60716
rect 580356 60664 580408 60716
rect 45008 59984 45060 60036
rect 57060 59984 57112 60036
rect 24676 59304 24728 59356
rect 57888 59304 57940 59356
rect 40408 57876 40460 57928
rect 57888 57876 57940 57928
rect 543556 57876 543608 57928
rect 572904 57876 572956 57928
rect 46020 56516 46072 56568
rect 57888 56516 57940 56568
rect 543556 55836 543608 55888
rect 562048 55836 562100 55888
rect 542728 53728 542780 53780
rect 580264 53728 580316 53780
rect 542728 51008 542780 51060
rect 551008 51008 551060 51060
rect 542728 49648 542780 49700
rect 552480 49648 552532 49700
rect 47216 48968 47268 49020
rect 57888 48968 57940 49020
rect 543648 48220 543700 48272
rect 577136 48220 577188 48272
rect 543648 45500 543700 45552
rect 582564 45500 582616 45552
rect 55588 45296 55640 45348
rect 57152 45296 57204 45348
rect 543648 42780 543700 42832
rect 547052 42780 547104 42832
rect 24768 41352 24820 41404
rect 57888 41352 57940 41404
rect 543556 41352 543608 41404
rect 557816 41352 557868 41404
rect 49332 41284 49384 41336
rect 56692 41284 56744 41336
rect 543556 37204 543608 37256
rect 560668 37204 560720 37256
rect 543648 35844 543700 35896
rect 560576 35844 560628 35896
rect 25964 34416 26016 34468
rect 57888 34416 57940 34468
rect 570696 33056 570748 33108
rect 580264 33056 580316 33108
rect 36544 32988 36596 33040
rect 57888 32988 57940 33040
rect 540704 31016 540756 31068
rect 578608 31016 578660 31068
rect 156052 29860 156104 29912
rect 157264 29860 157316 29912
rect 340880 29860 340932 29912
rect 342092 29860 342144 29912
rect 361580 29860 361632 29912
rect 362700 29860 362752 29912
rect 378140 29860 378192 29912
rect 379444 29860 379496 29912
rect 458180 29860 458232 29912
rect 459300 29860 459352 29912
rect 525800 29860 525852 29912
rect 526920 29860 526972 29912
rect 521108 29724 521160 29776
rect 54208 29656 54260 29708
rect 63500 29656 63552 29708
rect 45192 29588 45244 29640
rect 69020 29588 69072 29640
rect 552204 29588 552256 29640
rect 378048 29520 378100 29572
rect 378232 29520 378284 29572
rect 523040 29520 523092 29572
rect 566096 29520 566148 29572
rect 43168 29452 43220 29504
rect 69664 29452 69716 29504
rect 476672 29452 476724 29504
rect 525892 29452 525944 29504
rect 528192 29452 528244 29504
rect 552388 29452 552440 29504
rect 43904 29384 43956 29436
rect 123760 29384 123812 29436
rect 481824 29384 481876 29436
rect 565268 29384 565320 29436
rect 47308 29316 47360 29368
rect 199752 29316 199804 29368
rect 409696 29316 409748 29368
rect 554136 29316 554188 29368
rect 42524 29248 42576 29300
rect 195244 29248 195296 29300
rect 384580 29248 384632 29300
rect 550272 29248 550324 29300
rect 39304 29180 39356 29232
rect 193312 29180 193364 29232
rect 356888 29180 356940 29232
rect 544752 29180 544804 29232
rect 43720 29112 43772 29164
rect 205548 29112 205600 29164
rect 287336 29112 287388 29164
rect 575480 29112 575532 29164
rect 39856 29044 39908 29096
rect 217784 29044 217836 29096
rect 260932 29044 260984 29096
rect 583024 29044 583076 29096
rect 28908 28976 28960 29028
rect 159824 28976 159876 29028
rect 182364 28976 182416 29028
rect 550364 28976 550416 29028
rect 47492 28908 47544 28960
rect 325976 28908 326028 28960
rect 536564 28908 536616 28960
rect 552112 28908 552164 28960
rect 52276 28840 52328 28892
rect 67732 28840 67784 28892
rect 271236 28840 271288 28892
rect 527824 28840 527876 28892
rect 537208 28840 537260 28892
rect 550916 28840 550968 28892
rect 49516 28772 49568 28824
rect 63224 28772 63276 28824
rect 295708 28772 295760 28824
rect 474004 28772 474056 28824
rect 512092 28772 512144 28824
rect 583484 28772 583536 28824
rect 50712 28704 50764 28756
rect 62580 28704 62632 28756
rect 170864 28704 170916 28756
rect 249984 28704 250036 28756
rect 338212 28704 338264 28756
rect 524880 28704 524932 28756
rect 525892 28704 525944 28756
rect 581092 28704 581144 28756
rect 19248 28636 19300 28688
rect 82544 28636 82596 28688
rect 83464 28636 83516 28688
rect 190736 28636 190788 28688
rect 443184 28636 443236 28688
rect 563152 28636 563204 28688
rect 35348 28568 35400 28620
rect 103796 28568 103848 28620
rect 143172 28568 143224 28620
rect 251272 28568 251324 28620
rect 311164 28568 311216 28620
rect 529940 28568 529992 28620
rect 532056 28568 532108 28620
rect 581184 28568 581236 28620
rect 35808 28500 35860 28552
rect 73528 28500 73580 28552
rect 78772 28500 78824 28552
rect 188804 28500 188856 28552
rect 259000 28500 259052 28552
rect 505744 28500 505796 28552
rect 506940 28500 506992 28552
rect 566004 28500 566056 28552
rect 33600 28432 33652 28484
rect 71596 28432 71648 28484
rect 72424 28432 72476 28484
rect 141792 28432 141844 28484
rect 147680 28432 147732 28484
rect 148876 28432 148928 28484
rect 157984 28432 158036 28484
rect 272524 28432 272576 28484
rect 291844 28432 291896 28484
rect 535460 28432 535512 28484
rect 29736 28364 29788 28416
rect 92204 28364 92256 28416
rect 96804 28364 96856 28416
rect 211344 28364 211396 28416
rect 505652 28364 505704 28416
rect 574468 28364 574520 28416
rect 50896 28296 50948 28348
rect 95424 28296 95476 28348
rect 130200 28296 130252 28348
rect 252560 28296 252612 28348
rect 268016 28296 268068 28348
rect 517520 28296 517572 28348
rect 529480 28296 529532 28348
rect 575940 28296 575992 28348
rect 69940 28228 69992 28280
rect 213276 28228 213328 28280
rect 266084 28228 266136 28280
rect 451924 28228 451976 28280
rect 463700 28228 463752 28280
rect 464436 28228 464488 28280
rect 476120 28228 476172 28280
rect 477316 28228 477368 28280
rect 484492 28228 484544 28280
rect 485688 28228 485740 28280
rect 505100 28228 505152 28280
rect 506296 28228 506348 28280
rect 519176 28228 519228 28280
rect 562600 28228 562652 28280
rect 40684 28160 40736 28212
rect 72884 28160 72936 28212
rect 74540 28160 74592 28212
rect 181076 28160 181128 28212
rect 186320 28160 186372 28212
rect 187516 28160 187568 28212
rect 191840 28160 191892 28212
rect 192668 28160 192720 28212
rect 215300 28160 215352 28212
rect 216496 28160 216548 28212
rect 320180 28160 320232 28212
rect 321468 28160 321520 28212
rect 321560 28160 321612 28212
rect 322756 28160 322808 28212
rect 324320 28160 324372 28212
rect 325332 28160 325384 28212
rect 329840 28160 329892 28212
rect 331128 28160 331180 28212
rect 347780 28160 347832 28212
rect 348516 28160 348568 28212
rect 354680 28160 354732 28212
rect 355600 28160 355652 28212
rect 358820 28160 358872 28212
rect 360108 28160 360160 28212
rect 367100 28160 367152 28212
rect 367836 28160 367888 28212
rect 368480 28160 368532 28212
rect 369768 28160 369820 28212
rect 389088 28160 389140 28212
rect 536104 28160 536156 28212
rect 66352 28092 66404 28144
rect 168196 28092 168248 28144
rect 300860 28092 300912 28144
rect 302148 28092 302200 28144
rect 417424 28092 417476 28144
rect 544844 28092 544896 28144
rect 63500 28024 63552 28076
rect 98000 28024 98052 28076
rect 99288 28024 99340 28076
rect 99380 28024 99432 28076
rect 100576 28024 100628 28076
rect 107752 28024 107804 28076
rect 108948 28024 109000 28076
rect 109040 28024 109092 28076
rect 201684 28024 201736 28076
rect 426440 28024 426492 28076
rect 427728 28024 427780 28076
rect 427820 28024 427872 28076
rect 429016 28024 429068 28076
rect 436100 28024 436152 28076
rect 437388 28024 437440 28076
rect 445760 28024 445812 28076
rect 447048 28024 447100 28076
rect 447140 28024 447192 28076
rect 448336 28024 448388 28076
rect 448520 28024 448572 28076
rect 449624 28024 449676 28076
rect 465080 28024 465132 28076
rect 466368 28024 466420 28076
rect 484400 28024 484452 28076
rect 485044 28024 485096 28076
rect 502432 28024 502484 28076
rect 503076 28024 503128 28076
rect 503168 28024 503220 28076
rect 569408 28024 569460 28076
rect 103152 27956 103204 28008
rect 104164 27956 104216 28008
rect 195888 27956 195940 28008
rect 327264 27956 327316 28008
rect 562140 27956 562192 28008
rect 92572 27888 92624 27940
rect 179788 27888 179840 27940
rect 344008 27888 344060 27940
rect 563244 27888 563296 27940
rect 39580 27820 39632 27872
rect 166908 27820 166960 27872
rect 275744 27820 275796 27872
rect 510712 27820 510764 27872
rect 37648 27752 37700 27804
rect 155960 27752 156012 27804
rect 18880 27684 18932 27736
rect 128912 27684 128964 27736
rect 103520 27616 103572 27668
rect 109040 27616 109092 27668
rect 170404 27616 170456 27668
rect 170864 27616 170916 27668
rect 502340 27616 502392 27668
rect 503168 27616 503220 27668
rect 35532 27548 35584 27600
rect 70952 27548 71004 27600
rect 531412 27548 531464 27600
rect 560484 27548 560536 27600
rect 50804 27480 50856 27532
rect 70308 27480 70360 27532
rect 157340 27480 157392 27532
rect 158536 27480 158588 27532
rect 493416 27480 493468 27532
rect 570420 27480 570472 27532
rect 44272 27412 44324 27464
rect 89628 27412 89680 27464
rect 535460 27412 535512 27464
rect 563612 27412 563664 27464
rect 29920 27344 29972 27396
rect 470876 27344 470928 27396
rect 510160 27344 510212 27396
rect 573456 27344 573508 27396
rect 52552 27276 52604 27328
rect 441252 27276 441304 27328
rect 491484 27276 491536 27328
rect 553492 27276 553544 27328
rect 42432 27208 42484 27260
rect 385224 27208 385276 27260
rect 398748 27208 398800 27260
rect 583116 27208 583168 27260
rect 32772 27140 32824 27192
rect 363972 27140 364024 27192
rect 381360 27140 381412 27192
rect 561772 27140 561824 27192
rect 24400 27072 24452 27124
rect 266728 27072 266780 27124
rect 268660 27072 268712 27124
rect 577504 27072 577556 27124
rect 49148 27004 49200 27056
rect 296996 27004 297048 27056
rect 410340 27004 410392 27056
rect 576032 27004 576084 27056
rect 31116 26936 31168 26988
rect 109592 26936 109644 26988
rect 390376 26936 390428 26988
rect 540428 26936 540480 26988
rect 41052 26868 41104 26920
rect 92480 26868 92532 26920
rect 515956 26868 516008 26920
rect 549076 26868 549128 26920
rect 58624 26800 58676 26852
rect 87696 26800 87748 26852
rect 514024 26800 514076 26852
rect 549168 26800 549220 26852
rect 41880 26732 41932 26784
rect 523684 26732 523736 26784
rect 69664 26664 69716 26716
rect 520464 26664 520516 26716
rect 37004 26596 37056 26648
rect 494060 26596 494112 26648
rect 516600 26596 516652 26648
rect 549536 26596 549588 26648
rect 18972 26188 19024 26240
rect 391940 26188 391992 26240
rect 536104 26188 536156 26240
rect 547512 26188 547564 26240
rect 49240 26120 49292 26172
rect 368480 26120 368532 26172
rect 492680 26120 492732 26172
rect 560852 26120 560904 26172
rect 20628 26052 20680 26104
rect 318800 26052 318852 26104
rect 322940 26052 322992 26104
rect 578516 26052 578568 26104
rect 28724 25984 28776 26036
rect 307760 25984 307812 26036
rect 325792 25984 325844 26036
rect 578424 25984 578476 26036
rect 27344 25916 27396 25968
rect 306380 25916 306432 25968
rect 520280 25916 520332 25968
rect 571524 25916 571576 25968
rect 52000 25848 52052 25900
rect 292580 25848 292632 25900
rect 513380 25848 513432 25900
rect 567292 25848 567344 25900
rect 58716 25780 58768 25832
rect 216680 25780 216732 25832
rect 516140 25780 516192 25832
rect 571708 25780 571760 25832
rect 30748 25712 30800 25764
rect 186320 25712 186372 25764
rect 396080 25712 396132 25764
rect 545672 25712 545724 25764
rect 29828 25644 29880 25696
rect 165712 25644 165764 25696
rect 416780 25644 416832 25696
rect 575848 25644 575900 25696
rect 52828 25576 52880 25628
rect 77300 25576 77352 25628
rect 342352 25576 342404 25628
rect 573180 25576 573232 25628
rect 54852 25508 54904 25560
rect 81440 25508 81492 25560
rect 321744 25508 321796 25560
rect 563796 25508 563848 25560
rect 54944 25440 54996 25492
rect 67640 25440 67692 25492
rect 502524 25440 502576 25492
rect 546224 25440 546276 25492
rect 538220 25372 538272 25424
rect 555700 25372 555752 25424
rect 461032 25304 461084 25356
rect 540704 25304 540756 25356
rect 314660 24896 314712 24948
rect 479064 24896 479116 24948
rect 53656 24828 53708 24880
rect 85580 24828 85632 24880
rect 231860 24828 231912 24880
rect 485044 24828 485096 24880
rect 32312 24760 32364 24812
rect 444472 24760 444524 24812
rect 476120 24760 476172 24812
rect 552296 24760 552348 24812
rect 50620 24692 50672 24744
rect 397460 24692 397512 24744
rect 436100 24692 436152 24744
rect 569224 24692 569276 24744
rect 26056 24624 26108 24676
rect 354772 24624 354824 24676
rect 476028 24624 476080 24676
rect 549996 24624 550048 24676
rect 21824 24556 21876 24608
rect 333980 24556 334032 24608
rect 477500 24556 477552 24608
rect 539968 24556 540020 24608
rect 31208 24488 31260 24540
rect 256700 24488 256752 24540
rect 280160 24488 280212 24540
rect 574376 24488 574428 24540
rect 21548 24420 21600 24472
rect 311900 24420 311952 24472
rect 470600 24420 470652 24472
rect 557632 24420 557684 24472
rect 38108 24352 38160 24404
rect 204260 24352 204312 24404
rect 332600 24352 332652 24404
rect 556344 24352 556396 24404
rect 50528 24284 50580 24336
rect 191932 24284 191984 24336
rect 245660 24284 245712 24336
rect 563704 24284 563756 24336
rect 41236 24216 41288 24268
rect 182180 24216 182232 24268
rect 224960 24216 225012 24268
rect 571432 24216 571484 24268
rect 25596 24148 25648 24200
rect 131212 24148 131264 24200
rect 220820 24148 220872 24200
rect 568672 24148 568724 24200
rect 21732 24080 21784 24132
rect 124220 24080 124272 24132
rect 209872 24080 209924 24132
rect 564716 24080 564768 24132
rect 52736 24012 52788 24064
rect 142160 24012 142212 24064
rect 498200 24012 498252 24064
rect 559840 24012 559892 24064
rect 42984 23944 43036 23996
rect 99380 23944 99432 23996
rect 502432 23944 502484 23996
rect 551468 23944 551520 23996
rect 51448 23876 51500 23928
rect 98092 23876 98144 23928
rect 34152 23400 34204 23452
rect 104900 23400 104952 23452
rect 517520 23400 517572 23452
rect 540612 23400 540664 23452
rect 46664 23332 46716 23384
rect 131120 23332 131172 23384
rect 184940 23332 184992 23384
rect 581644 23332 581696 23384
rect 52920 23264 52972 23316
rect 128452 23264 128504 23316
rect 529940 23264 529992 23316
rect 562324 23264 562376 23316
rect 354680 23196 354732 23248
rect 579620 23196 579672 23248
rect 21640 23128 21692 23180
rect 342260 23128 342312 23180
rect 365720 23128 365772 23180
rect 579804 23128 579856 23180
rect 36268 23060 36320 23112
rect 321560 23060 321612 23112
rect 409972 23060 410024 23112
rect 555332 23060 555384 23112
rect 24584 22992 24636 23044
rect 285680 22992 285732 23044
rect 451280 22992 451332 23044
rect 582932 22992 582984 23044
rect 45100 22924 45152 22976
rect 303620 22924 303672 22976
rect 449900 22924 449952 22976
rect 555424 22924 555476 22976
rect 23388 22856 23440 22908
rect 270500 22856 270552 22908
rect 385040 22856 385092 22908
rect 558552 22856 558604 22908
rect 22008 22788 22060 22840
rect 72332 22788 72384 22840
rect 171140 22788 171192 22840
rect 416688 22788 416740 22840
rect 456800 22788 456852 22840
rect 556712 22788 556764 22840
rect 49424 22720 49476 22772
rect 110420 22720 110472 22772
rect 168380 22720 168432 22772
rect 553860 22720 553912 22772
rect 43996 22652 44048 22704
rect 215300 22652 215352 22704
rect 465264 22652 465316 22704
rect 554044 22652 554096 22704
rect 44088 22584 44140 22636
rect 66352 22584 66404 22636
rect 107752 22584 107804 22636
rect 554964 22584 555016 22636
rect 45376 22516 45428 22568
rect 72424 22516 72476 22568
rect 160100 22516 160152 22568
rect 548984 22516 549036 22568
rect 32680 22448 32732 22500
rect 356060 22448 356112 22500
rect 58532 22040 58584 22092
rect 78772 22040 78824 22092
rect 488540 22040 488592 22092
rect 551560 22040 551612 22092
rect 47952 21972 48004 22024
rect 411260 21972 411312 22024
rect 483020 21972 483072 22024
rect 544384 21972 544436 22024
rect 54484 21904 54536 21956
rect 400220 21904 400272 21956
rect 528560 21904 528612 21956
rect 570604 21904 570656 21956
rect 52092 21836 52144 21888
rect 209780 21836 209832 21888
rect 223580 21836 223632 21888
rect 548616 21836 548668 21888
rect 51724 21768 51776 21820
rect 364340 21768 364392 21820
rect 385132 21768 385184 21820
rect 552664 21768 552716 21820
rect 46296 21700 46348 21752
rect 255320 21700 255372 21752
rect 420920 21700 420972 21752
rect 559104 21700 559156 21752
rect 56232 21632 56284 21684
rect 197360 21632 197412 21684
rect 371240 21632 371292 21684
rect 553676 21632 553728 21684
rect 51356 21564 51408 21616
rect 169760 21564 169812 21616
rect 258080 21564 258132 21616
rect 568856 21564 568908 21616
rect 54576 21496 54628 21548
rect 156052 21496 156104 21548
rect 260840 21496 260892 21548
rect 572996 21496 573048 21548
rect 46572 21428 46624 21480
rect 147680 21428 147732 21480
rect 176660 21428 176712 21480
rect 573088 21428 573140 21480
rect 43812 21360 43864 21412
rect 103520 21360 103572 21412
rect 146392 21360 146444 21412
rect 569592 21360 569644 21412
rect 49608 21292 49660 21344
rect 92572 21292 92624 21344
rect 510712 21292 510764 21344
rect 542176 21292 542228 21344
rect 57612 21224 57664 21276
rect 96804 21224 96856 21276
rect 46388 21156 46440 21208
rect 427820 21156 427872 21208
rect 58900 20612 58952 20664
rect 69940 20612 69992 20664
rect 503720 20612 503772 20664
rect 504364 20612 504416 20664
rect 524880 20612 524932 20664
rect 551284 20612 551336 20664
rect 22652 20544 22704 20596
rect 458180 20544 458232 20596
rect 480260 20544 480312 20596
rect 556620 20544 556672 20596
rect 43628 20476 43680 20528
rect 387800 20476 387852 20528
rect 423680 20476 423732 20528
rect 580080 20476 580132 20528
rect 28540 20408 28592 20460
rect 367100 20408 367152 20460
rect 421012 20408 421064 20460
rect 546684 20408 546736 20460
rect 38384 20340 38436 20392
rect 229100 20340 229152 20392
rect 231952 20340 232004 20392
rect 564624 20340 564676 20392
rect 46204 20272 46256 20324
rect 219532 20272 219584 20324
rect 251272 20272 251324 20324
rect 583208 20272 583260 20324
rect 55128 20204 55180 20256
rect 367192 20204 367244 20256
rect 434720 20204 434772 20256
rect 559196 20204 559248 20256
rect 55772 20136 55824 20188
rect 227720 20136 227772 20188
rect 292580 20136 292632 20188
rect 554320 20136 554372 20188
rect 58348 20068 58400 20120
rect 211252 20068 211304 20120
rect 253940 20068 253992 20120
rect 548156 20068 548208 20120
rect 184940 20000 184992 20052
rect 553584 20000 553636 20052
rect 39672 19932 39724 19984
rect 139400 19932 139452 19984
rect 183652 19932 183704 19984
rect 555240 19932 555292 19984
rect 55864 19864 55916 19916
rect 153200 19864 153252 19916
rect 360200 19864 360252 19916
rect 547604 19864 547656 19916
rect 57796 19796 57848 19848
rect 130200 19796 130252 19848
rect 504364 19796 504416 19848
rect 567660 19796 567712 19848
rect 22560 19728 22612 19780
rect 462320 19728 462372 19780
rect 465080 19728 465132 19780
rect 571800 19728 571852 19780
rect 44916 19660 44968 19712
rect 189080 19660 189132 19712
rect 35716 19252 35768 19304
rect 219440 19252 219492 19304
rect 247040 19252 247092 19304
rect 573364 19252 573416 19304
rect 54760 19184 54812 19236
rect 293960 19184 294012 19236
rect 358820 19184 358872 19236
rect 551376 19184 551428 19236
rect 45284 19116 45336 19168
rect 202880 19116 202932 19168
rect 419540 19116 419592 19168
rect 565084 19116 565136 19168
rect 53380 19048 53432 19100
rect 205640 19048 205692 19100
rect 463700 19048 463752 19100
rect 574284 19048 574336 19100
rect 41328 18980 41380 19032
rect 183560 18980 183612 19032
rect 459560 18980 459612 19032
rect 563520 18980 563572 19032
rect 36636 18912 36688 18964
rect 149060 18912 149112 18964
rect 317420 18912 317472 18964
rect 558000 18912 558052 18964
rect 36912 18844 36964 18896
rect 146300 18844 146352 18896
rect 271880 18844 271932 18896
rect 567476 18844 567528 18896
rect 57428 18776 57480 18828
rect 165620 18776 165672 18828
rect 251180 18776 251232 18828
rect 561956 18776 562008 18828
rect 49976 18708 50028 18760
rect 125600 18708 125652 18760
rect 136640 18708 136692 18760
rect 570144 18708 570196 18760
rect 50344 18640 50396 18692
rect 104164 18640 104216 18692
rect 113180 18640 113232 18692
rect 549444 18640 549496 18692
rect 99380 18572 99432 18624
rect 577412 18572 577464 18624
rect 46112 18504 46164 18556
rect 147680 18504 147732 18556
rect 466460 18504 466512 18556
rect 568764 18504 568816 18556
rect 55956 18436 56008 18488
rect 154580 18436 154632 18488
rect 469220 18436 469272 18488
rect 545304 18436 545356 18488
rect 45928 18368 45980 18420
rect 83464 18368 83516 18420
rect 533344 18368 533396 18420
rect 543280 18368 543332 18420
rect 46848 18300 46900 18352
rect 120080 18300 120132 18352
rect 98000 17892 98052 17944
rect 583392 17892 583444 17944
rect 106372 17824 106424 17876
rect 581368 17824 581420 17876
rect 42064 17756 42116 17808
rect 116032 17756 116084 17808
rect 157340 17756 157392 17808
rect 583576 17756 583628 17808
rect 40960 17688 41012 17740
rect 375380 17688 375432 17740
rect 378140 17688 378192 17740
rect 546960 17688 547012 17740
rect 58072 17620 58124 17672
rect 329840 17620 329892 17672
rect 340880 17620 340932 17672
rect 577688 17620 577740 17672
rect 59912 17552 59964 17604
rect 245752 17552 245804 17604
rect 460940 17552 460992 17604
rect 573272 17552 573324 17604
rect 57704 17484 57756 17536
rect 237380 17484 237432 17536
rect 527824 17484 527876 17536
rect 544292 17484 544344 17536
rect 59820 17416 59872 17468
rect 234620 17416 234672 17468
rect 427820 17416 427872 17468
rect 571616 17416 571668 17468
rect 57336 17348 57388 17400
rect 142804 17348 142856 17400
rect 414020 17348 414072 17400
rect 571340 17348 571392 17400
rect 45468 17280 45520 17332
rect 115940 17280 115992 17332
rect 259460 17280 259512 17332
rect 541900 17280 541952 17332
rect 120080 17212 120132 17264
rect 579988 17212 580040 17264
rect 52368 17144 52420 17196
rect 170404 17144 170456 17196
rect 106280 16600 106332 16652
rect 560300 16600 560352 16652
rect 48044 16532 48096 16584
rect 164332 16532 164384 16584
rect 233240 16532 233292 16584
rect 548800 16532 548852 16584
rect 48136 16464 48188 16516
rect 161572 16464 161624 16516
rect 361580 16464 361632 16516
rect 581736 16464 581788 16516
rect 58808 16396 58860 16448
rect 157984 16396 158036 16448
rect 335452 16396 335504 16448
rect 541440 16396 541492 16448
rect 347780 16328 347832 16380
rect 544476 16328 544528 16380
rect 289820 16260 289872 16312
rect 557080 16260 557132 16312
rect 264980 16192 265032 16244
rect 564900 16192 564952 16244
rect 253480 16124 253532 16176
rect 572812 16124 572864 16176
rect 228272 16056 228324 16108
rect 558920 16056 558972 16108
rect 226340 15988 226392 16040
rect 570052 15988 570104 16040
rect 33968 15920 34020 15972
rect 130568 15920 130620 15972
rect 229376 15920 229428 15972
rect 575756 15920 575808 15972
rect 35624 15852 35676 15904
rect 158904 15852 158956 15904
rect 171968 15852 172020 15904
rect 564808 15852 564860 15904
rect 398840 15784 398892 15836
rect 544108 15784 544160 15836
rect 447140 15716 447192 15768
rect 549812 15716 549864 15768
rect 522304 15648 522356 15700
rect 567568 15648 567620 15700
rect 242900 15104 242952 15156
rect 552756 15104 552808 15156
rect 380900 15036 380952 15088
rect 540060 15036 540112 15088
rect 393320 14968 393372 15020
rect 543740 14968 543792 15020
rect 404360 14900 404412 14952
rect 546040 14900 546092 14952
rect 444380 14832 444432 14884
rect 576124 14832 576176 14884
rect 426440 14764 426492 14816
rect 544016 14764 544068 14816
rect 403624 14696 403676 14748
rect 542268 14696 542320 14748
rect 398840 14628 398892 14680
rect 541992 14628 542044 14680
rect 382372 14560 382424 14612
rect 547236 14560 547288 14612
rect 378416 14492 378468 14544
rect 548708 14492 548760 14544
rect 247592 14424 247644 14476
rect 550088 14424 550140 14476
rect 430580 14356 430632 14408
rect 543188 14356 543240 14408
rect 434812 14288 434864 14340
rect 546776 14288 546828 14340
rect 433340 14220 433392 14272
rect 541808 14220 541860 14272
rect 320180 13744 320232 13796
rect 563428 13744 563480 13796
rect 372620 13676 372672 13728
rect 583760 13676 583812 13728
rect 357532 13608 357584 13660
rect 540336 13608 540388 13660
rect 349160 13540 349212 13592
rect 543004 13540 543056 13592
rect 346952 13472 347004 13524
rect 541624 13472 541676 13524
rect 367744 13404 367796 13456
rect 579160 13404 579212 13456
rect 311440 13336 311492 13388
rect 562416 13336 562468 13388
rect 297272 13268 297324 13320
rect 558184 13268 558236 13320
rect 286600 13200 286652 13252
rect 559564 13200 559616 13252
rect 234620 13132 234672 13184
rect 553768 13132 553820 13184
rect 242900 13064 242952 13116
rect 578700 13064 578752 13116
rect 364616 12996 364668 13048
rect 545948 12996 546000 13048
rect 453304 12928 453356 12980
rect 559012 12928 559064 12980
rect 474004 12860 474056 12912
rect 549720 12860 549772 12912
rect 190552 12384 190604 12436
rect 583668 12384 583720 12436
rect 313280 12316 313332 12368
rect 543096 12316 543148 12368
rect 314752 12248 314804 12300
rect 544568 12248 544620 12300
rect 321652 12180 321704 12232
rect 540520 12180 540572 12232
rect 324320 12112 324372 12164
rect 541716 12112 541768 12164
rect 328460 12044 328512 12096
rect 543464 12044 543516 12096
rect 351920 11976 351972 12028
rect 551192 11976 551244 12028
rect 346400 11908 346452 11960
rect 543556 11908 543608 11960
rect 363052 11840 363104 11892
rect 548064 11840 548116 11892
rect 256700 11772 256752 11824
rect 577596 11772 577648 11824
rect 239312 11704 239364 11756
rect 576308 11704 576360 11756
rect 357440 11636 357492 11688
rect 542360 11636 542412 11688
rect 451924 11568 451976 11620
rect 540244 11568 540296 11620
rect 505744 11500 505796 11552
rect 543832 11500 543884 11552
rect 48964 10956 49016 11008
rect 191840 10956 191892 11008
rect 303896 10344 303948 10396
rect 557724 10344 557776 10396
rect 141240 10276 141292 10328
rect 555148 10276 555200 10328
rect 307944 9052 307996 9104
rect 550824 9052 550876 9104
rect 249984 8984 250036 9036
rect 553400 8984 553452 9036
rect 208584 8916 208636 8968
rect 556528 8916 556580 8968
rect 194416 7556 194468 7608
rect 556252 7556 556304 7608
rect 567844 7556 567896 7608
rect 579804 7556 579856 7608
rect 463976 6808 464028 6860
rect 561220 6808 561272 6860
rect 446220 6740 446272 6792
rect 545488 6740 545540 6792
rect 439136 6672 439188 6724
rect 541072 6672 541124 6724
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 474556 6604 474608 6656
rect 582380 6604 582432 6656
rect 460388 6536 460440 6588
rect 569500 6536 569552 6588
rect 449808 6468 449860 6520
rect 566372 6468 566424 6520
rect 442632 6400 442684 6452
rect 575020 6400 575072 6452
rect 432052 6332 432104 6384
rect 570512 6332 570564 6384
rect 424968 6264 425020 6316
rect 564992 6264 565044 6316
rect 389456 6196 389508 6248
rect 559288 6196 559340 6248
rect 300768 6128 300820 6180
rect 545764 6128 545816 6180
rect 481732 6060 481784 6112
rect 569960 6060 570012 6112
rect 488816 5992 488868 6044
rect 561312 5992 561364 6044
rect 527824 5924 527876 5976
rect 566188 5924 566240 5976
rect 288440 5448 288492 5500
rect 546868 5448 546920 5500
rect 299480 5380 299532 5432
rect 547144 5380 547196 5432
rect 478144 4768 478196 4820
rect 557908 4768 557960 4820
rect 574836 4224 574888 4276
rect 577412 4224 577464 4276
rect 48228 4088 48280 4140
rect 117596 4088 117648 4140
rect 495900 4088 495952 4140
rect 556436 4088 556488 4140
rect 42156 4020 42208 4072
rect 182548 4020 182600 4072
rect 492312 4020 492364 4072
rect 553952 4020 554004 4072
rect 556160 4020 556212 4072
rect 563336 4020 563388 4072
rect 46756 3952 46808 4004
rect 189724 3952 189776 4004
rect 222752 3952 222804 4004
rect 526444 3952 526496 4004
rect 549076 3952 549128 4004
rect 573640 3952 573692 4004
rect 50436 3884 50488 3936
rect 193220 3884 193272 3936
rect 212172 3884 212224 3936
rect 533344 3884 533396 3936
rect 534908 3884 534960 3936
rect 565360 3884 565412 3936
rect 41144 3816 41196 3868
rect 196808 3816 196860 3868
rect 240508 3816 240560 3868
rect 574192 3816 574244 3868
rect 42248 3748 42300 3800
rect 161296 3748 161348 3800
rect 175464 3748 175516 3800
rect 522304 3748 522356 3800
rect 524236 3748 524288 3800
rect 570236 3748 570288 3800
rect 34336 3680 34388 3732
rect 197912 3680 197964 3732
rect 552664 3680 552716 3732
rect 561864 3680 561916 3732
rect 565820 3680 565872 3732
rect 566280 3680 566332 3732
rect 34244 3612 34296 3664
rect 215668 3612 215720 3664
rect 218152 3612 218204 3664
rect 574652 3612 574704 3664
rect 37096 3544 37148 3596
rect 184848 3544 184900 3596
rect 184940 3544 184992 3596
rect 186136 3544 186188 3596
rect 190828 3544 190880 3596
rect 576860 3544 576912 3596
rect 39764 3476 39816 3528
rect 134156 3476 134208 3528
rect 135260 3476 135312 3528
rect 136456 3476 136508 3528
rect 143540 3476 143592 3528
rect 144736 3476 144788 3528
rect 144828 3476 144880 3528
rect 568028 3476 568080 3528
rect 36728 3408 36780 3460
rect 57244 3408 57296 3460
rect 92756 3408 92808 3460
rect 549904 3408 549956 3460
rect 559748 3408 559800 3460
rect 575664 3408 575716 3460
rect 53012 3340 53064 3392
rect 96252 3340 96304 3392
rect 184848 3340 184900 3392
rect 187332 3340 187384 3392
rect 218060 3340 218112 3392
rect 219256 3340 219308 3392
rect 234620 3340 234672 3392
rect 235816 3340 235868 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 259460 3340 259512 3392
rect 260656 3340 260708 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 510068 3340 510120 3392
rect 565820 3340 565872 3392
rect 499396 3272 499448 3324
rect 555056 3272 555108 3324
rect 578976 3272 579028 3324
rect 582196 3272 582248 3324
rect 545488 3204 545540 3256
rect 567384 3204 567436 3256
rect 200304 3136 200356 3188
rect 552848 3136 552900 3188
rect 572076 3000 572128 3052
rect 573916 3000 573968 3052
rect 143540 2796 143592 2848
rect 144828 2796 144880 2848
rect 276112 1300 276164 1352
rect 549628 1300 549680 1352
rect 233792 8 233844 60
rect 545212 8 545264 60
<< metal2 >>
rect 6932 703582 7972 703610
rect 6932 686526 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 6920 686520 6972 686526
rect 6920 686462 6972 686468
rect 21364 684072 21416 684078
rect 21364 684014 21416 684020
rect 3424 682712 3476 682718
rect 3424 682654 3476 682660
rect 3332 658232 3384 658238
rect 3330 658200 3332 658209
rect 3384 658200 3386 658209
rect 3330 658135 3386 658144
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3436 553897 3464 682654
rect 17776 681828 17828 681834
rect 17776 681770 17828 681776
rect 8944 681352 8996 681358
rect 8944 681294 8996 681300
rect 7564 677612 7616 677618
rect 7564 677554 7616 677560
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 588606 3556 671191
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3516 588600 3568 588606
rect 3516 588542 3568 588548
rect 3620 574802 3648 619103
rect 3698 606112 3754 606121
rect 3698 606047 3754 606056
rect 3712 588577 3740 606047
rect 3698 588568 3754 588577
rect 3698 588503 3754 588512
rect 3608 574796 3660 574802
rect 3608 574738 3660 574744
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3436 197305 3464 501735
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4066 201920 4122 201929
rect 4066 201855 4122 201864
rect 3422 197296 3478 197305
rect 3422 197231 3478 197240
rect 4080 194449 4108 201855
rect 4066 194440 4122 194449
rect 4066 194375 4122 194384
rect 1398 192536 1454 192545
rect 1398 192471 1454 192480
rect 4804 192500 4856 192506
rect 542 -960 654 480
rect 1412 354 1440 192471
rect 4804 192442 4856 192448
rect 2778 191040 2834 191049
rect 2778 190975 2834 190984
rect 2792 16574 2820 190975
rect 3516 189780 3568 189786
rect 3516 189722 3568 189728
rect 3424 188964 3476 188970
rect 3424 188906 3476 188912
rect 3436 188873 3464 188906
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3424 159384 3476 159390
rect 3424 159326 3476 159332
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 149734 3372 149767
rect 3332 149728 3384 149734
rect 3332 149670 3384 149676
rect 2872 97776 2924 97782
rect 2872 97718 2924 97724
rect 2884 97617 2912 97718
rect 2870 97608 2926 97617
rect 2870 97543 2926 97552
rect 3436 58585 3464 159326
rect 3528 136785 3556 189722
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 4816 97782 4844 192442
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 7576 6662 7604 677554
rect 8956 658238 8984 681294
rect 9678 680096 9734 680105
rect 9678 680031 9734 680040
rect 8944 658232 8996 658238
rect 8944 658174 8996 658180
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 680031
rect 17224 565888 17276 565894
rect 17224 565830 17276 565836
rect 17236 194206 17264 565830
rect 17316 397520 17368 397526
rect 17316 397462 17368 397468
rect 17224 194200 17276 194206
rect 17224 194142 17276 194148
rect 17328 191758 17356 397462
rect 17684 349172 17736 349178
rect 17684 349114 17736 349120
rect 17316 191752 17368 191758
rect 17316 191694 17368 191700
rect 13820 178832 13872 178838
rect 13820 178774 13872 178780
rect 13832 16574 13860 178774
rect 17696 137970 17724 349114
rect 17788 198150 17816 681770
rect 17866 584352 17922 584361
rect 17866 584287 17922 584296
rect 17776 198144 17828 198150
rect 17776 198086 17828 198092
rect 17684 137964 17736 137970
rect 17684 137906 17736 137912
rect 17880 82822 17908 584287
rect 20628 566092 20680 566098
rect 20628 566034 20680 566040
rect 19156 561740 19208 561746
rect 19156 561682 19208 561688
rect 19064 484424 19116 484430
rect 19064 484366 19116 484372
rect 18972 298172 19024 298178
rect 18972 298114 19024 298120
rect 18880 296744 18932 296750
rect 18880 296686 18932 296692
rect 17868 82816 17920 82822
rect 17868 82758 17920 82764
rect 18892 27742 18920 296686
rect 18880 27736 18932 27742
rect 18880 27678 18932 27684
rect 18984 26246 19012 298114
rect 19076 156641 19104 484366
rect 19062 156632 19118 156641
rect 19062 156567 19118 156576
rect 19168 152697 19196 561682
rect 19248 485852 19300 485858
rect 19248 485794 19300 485800
rect 19154 152688 19210 152697
rect 19154 152623 19210 152632
rect 19260 28694 19288 485794
rect 19984 462392 20036 462398
rect 19984 462334 20036 462340
rect 19996 198665 20024 462334
rect 20076 448588 20128 448594
rect 20076 448530 20128 448536
rect 19982 198656 20038 198665
rect 19982 198591 20038 198600
rect 20088 197062 20116 448530
rect 20444 414044 20496 414050
rect 20444 413986 20496 413992
rect 20168 292596 20220 292602
rect 20168 292538 20220 292544
rect 20076 197056 20128 197062
rect 20076 196998 20128 197004
rect 20180 191826 20208 292538
rect 20352 277432 20404 277438
rect 20352 277374 20404 277380
rect 20168 191820 20220 191826
rect 20168 191762 20220 191768
rect 20364 190466 20392 277374
rect 20456 194546 20484 413986
rect 20536 389224 20588 389230
rect 20536 389166 20588 389172
rect 20444 194540 20496 194546
rect 20444 194482 20496 194488
rect 20352 190460 20404 190466
rect 20352 190402 20404 190408
rect 19340 189848 19392 189854
rect 19340 189790 19392 189796
rect 19248 28688 19300 28694
rect 19248 28630 19300 28636
rect 18972 26240 19024 26246
rect 18972 26182 19024 26188
rect 19352 16574 19380 189790
rect 20548 20369 20576 389166
rect 20640 26110 20668 566034
rect 21272 300892 21324 300898
rect 21272 300834 21324 300840
rect 21284 198529 21312 300834
rect 21270 198520 21326 198529
rect 21270 198455 21326 198464
rect 21376 85542 21404 684014
rect 31024 683256 31076 683262
rect 31024 683198 31076 683204
rect 26148 682576 26200 682582
rect 26148 682518 26200 682524
rect 25778 587480 25834 587489
rect 25778 587415 25834 587424
rect 22836 587036 22888 587042
rect 22836 586978 22888 586984
rect 22008 563372 22060 563378
rect 22008 563314 22060 563320
rect 21916 541000 21968 541006
rect 21916 540942 21968 540948
rect 21824 505164 21876 505170
rect 21824 505106 21876 505112
rect 21732 495508 21784 495514
rect 21732 495450 21784 495456
rect 21640 467900 21692 467906
rect 21640 467842 21692 467848
rect 21548 463752 21600 463758
rect 21548 463694 21600 463700
rect 21456 407176 21508 407182
rect 21456 407118 21508 407124
rect 21468 196858 21496 407118
rect 21456 196852 21508 196858
rect 21456 196794 21508 196800
rect 21364 85536 21416 85542
rect 21364 85478 21416 85484
rect 20628 26104 20680 26110
rect 20628 26046 20680 26052
rect 21560 24478 21588 463694
rect 21548 24472 21600 24478
rect 21548 24414 21600 24420
rect 21652 23186 21680 467842
rect 21744 24138 21772 495450
rect 21836 24614 21864 505106
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21732 24132 21784 24138
rect 21732 24074 21784 24080
rect 21928 23225 21956 540942
rect 21914 23216 21970 23225
rect 21640 23180 21692 23186
rect 21914 23151 21970 23160
rect 21640 23122 21692 23128
rect 22020 22846 22048 563314
rect 22744 394732 22796 394738
rect 22744 394674 22796 394680
rect 22652 345160 22704 345166
rect 22652 345102 22704 345108
rect 22560 310548 22612 310554
rect 22560 310490 22612 310496
rect 22008 22840 22060 22846
rect 22008 22782 22060 22788
rect 20534 20360 20590 20369
rect 20534 20295 20590 20304
rect 22572 19786 22600 310490
rect 22664 20602 22692 345102
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22756 20505 22784 394674
rect 22848 198422 22876 586978
rect 22928 586832 22980 586838
rect 22928 586774 22980 586780
rect 22940 198694 22968 586774
rect 24674 565856 24730 565865
rect 24674 565791 24730 565800
rect 23388 565004 23440 565010
rect 23388 564946 23440 564952
rect 23204 564052 23256 564058
rect 23204 563994 23256 564000
rect 23020 562760 23072 562766
rect 23020 562702 23072 562708
rect 22928 198688 22980 198694
rect 22928 198630 22980 198636
rect 22836 198416 22888 198422
rect 22836 198358 22888 198364
rect 23032 124166 23060 562702
rect 23112 562624 23164 562630
rect 23112 562566 23164 562572
rect 23020 124160 23072 124166
rect 23020 124102 23072 124108
rect 23124 117298 23152 562566
rect 23112 117292 23164 117298
rect 23112 117234 23164 117240
rect 23216 103494 23244 563994
rect 23296 520328 23348 520334
rect 23296 520270 23348 520276
rect 23204 103488 23256 103494
rect 23204 103430 23256 103436
rect 23308 22817 23336 520270
rect 23400 22914 23428 564946
rect 24308 563984 24360 563990
rect 24308 563926 24360 563932
rect 24216 492720 24268 492726
rect 24216 492662 24268 492668
rect 24124 357468 24176 357474
rect 24124 357410 24176 357416
rect 24136 197198 24164 357410
rect 24124 197192 24176 197198
rect 24124 197134 24176 197140
rect 24228 153785 24256 492662
rect 24320 196790 24348 563926
rect 24584 460964 24636 460970
rect 24584 460906 24636 460912
rect 24492 443012 24544 443018
rect 24492 442954 24544 442960
rect 24400 415472 24452 415478
rect 24400 415414 24452 415420
rect 24308 196784 24360 196790
rect 24308 196726 24360 196732
rect 24214 153776 24270 153785
rect 24214 153711 24270 153720
rect 24412 27130 24440 415414
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24504 22953 24532 442954
rect 24596 23050 24624 460906
rect 24688 59362 24716 565791
rect 24768 563304 24820 563310
rect 24768 563246 24820 563252
rect 24676 59356 24728 59362
rect 24676 59298 24728 59304
rect 24780 41410 24808 563246
rect 25688 561536 25740 561542
rect 25688 561478 25740 561484
rect 25504 354748 25556 354754
rect 25504 354690 25556 354696
rect 25412 346452 25464 346458
rect 25412 346394 25464 346400
rect 25320 281580 25372 281586
rect 25320 281522 25372 281528
rect 25332 194478 25360 281522
rect 25320 194472 25372 194478
rect 25320 194414 25372 194420
rect 25424 194410 25452 346394
rect 25412 194404 25464 194410
rect 25412 194346 25464 194352
rect 25516 150822 25544 354690
rect 25596 302252 25648 302258
rect 25596 302194 25648 302200
rect 25504 150816 25556 150822
rect 25504 150758 25556 150764
rect 24768 41404 24820 41410
rect 24768 41346 24820 41352
rect 25608 24206 25636 302194
rect 25700 198626 25728 561478
rect 25688 198620 25740 198626
rect 25688 198562 25740 198568
rect 25792 198014 25820 587415
rect 25870 587344 25926 587353
rect 25870 587279 25926 587288
rect 25884 198257 25912 587279
rect 25964 565616 26016 565622
rect 25964 565558 26016 565564
rect 25870 198248 25926 198257
rect 25870 198183 25926 198192
rect 25780 198008 25832 198014
rect 25780 197950 25832 197956
rect 25976 34474 26004 565558
rect 26054 562048 26110 562057
rect 26054 561983 26110 561992
rect 25964 34468 26016 34474
rect 25964 34410 26016 34416
rect 26068 24682 26096 561983
rect 26160 135250 26188 682518
rect 30102 562184 30158 562193
rect 30102 562119 30158 562128
rect 27436 562080 27488 562086
rect 27436 562022 27488 562028
rect 27160 561264 27212 561270
rect 27160 561206 27212 561212
rect 27068 444440 27120 444446
rect 27068 444382 27120 444388
rect 26976 423700 27028 423706
rect 26976 423642 27028 423648
rect 26884 374060 26936 374066
rect 26884 374002 26936 374008
rect 26792 372632 26844 372638
rect 26792 372574 26844 372580
rect 26700 305040 26752 305046
rect 26700 304982 26752 304988
rect 26712 193186 26740 304982
rect 26700 193180 26752 193186
rect 26700 193122 26752 193128
rect 26804 169046 26832 372574
rect 26792 169040 26844 169046
rect 26792 168982 26844 168988
rect 26896 158137 26924 374002
rect 26882 158128 26938 158137
rect 26882 158063 26938 158072
rect 26988 152794 27016 423642
rect 27080 158001 27108 444382
rect 27172 199170 27200 561206
rect 27250 560960 27306 560969
rect 27250 560895 27306 560904
rect 27160 199164 27212 199170
rect 27160 199106 27212 199112
rect 27264 194313 27292 560895
rect 27344 392012 27396 392018
rect 27344 391954 27396 391960
rect 27250 194304 27306 194313
rect 27250 194239 27306 194248
rect 27066 157992 27122 158001
rect 27066 157927 27122 157936
rect 26976 152788 27028 152794
rect 26976 152730 27028 152736
rect 26148 135244 26200 135250
rect 26148 135186 26200 135192
rect 27356 25974 27384 391954
rect 27448 103426 27476 562022
rect 28814 561776 28870 561785
rect 28814 561711 28870 561720
rect 27528 506524 27580 506530
rect 27528 506466 27580 506472
rect 27436 103420 27488 103426
rect 27436 103362 27488 103368
rect 27540 29209 27568 506466
rect 28632 489932 28684 489938
rect 28632 489874 28684 489880
rect 28448 419552 28500 419558
rect 28448 419494 28500 419500
rect 28356 372700 28408 372706
rect 28356 372642 28408 372648
rect 28264 336796 28316 336802
rect 28264 336738 28316 336744
rect 28172 328500 28224 328506
rect 28172 328442 28224 328448
rect 28080 320204 28132 320210
rect 28080 320146 28132 320152
rect 28092 195702 28120 320146
rect 28080 195696 28132 195702
rect 28080 195638 28132 195644
rect 27618 192808 27674 192817
rect 27618 192743 27674 192752
rect 27526 29200 27582 29209
rect 27526 29135 27582 29144
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 24584 23044 24636 23050
rect 24584 22986 24636 22992
rect 24490 22944 24546 22953
rect 23388 22908 23440 22914
rect 24490 22879 24546 22888
rect 23388 22850 23440 22856
rect 23294 22808 23350 22817
rect 23294 22743 23350 22752
rect 22742 20496 22798 20505
rect 22742 20431 22798 20440
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 27632 16574 27660 192743
rect 28184 158030 28212 328442
rect 28172 158024 28224 158030
rect 28172 157966 28224 157972
rect 28276 151094 28304 336738
rect 28368 152522 28396 372642
rect 28460 196450 28488 419494
rect 28540 288448 28592 288454
rect 28540 288390 28592 288396
rect 28448 196444 28500 196450
rect 28448 196386 28500 196392
rect 28356 152516 28408 152522
rect 28356 152458 28408 152464
rect 28264 151088 28316 151094
rect 28264 151030 28316 151036
rect 28552 20466 28580 288390
rect 28644 152561 28672 489874
rect 28724 362976 28776 362982
rect 28724 362918 28776 362924
rect 28630 152552 28686 152561
rect 28630 152487 28686 152496
rect 28736 26042 28764 362918
rect 28828 160721 28856 561711
rect 30012 561128 30064 561134
rect 30012 561070 30064 561076
rect 28908 431996 28960 432002
rect 28908 431938 28960 431944
rect 28814 160712 28870 160721
rect 28814 160647 28870 160656
rect 28920 29034 28948 431938
rect 29920 386436 29972 386442
rect 29920 386378 29972 386384
rect 29644 382288 29696 382294
rect 29644 382230 29696 382236
rect 29552 378208 29604 378214
rect 29552 378150 29604 378156
rect 29460 345092 29512 345098
rect 29460 345034 29512 345040
rect 29472 197130 29500 345034
rect 29460 197124 29512 197130
rect 29460 197066 29512 197072
rect 29564 164966 29592 378150
rect 29552 164960 29604 164966
rect 29552 164902 29604 164908
rect 29656 163538 29684 382230
rect 29736 368552 29788 368558
rect 29736 368494 29788 368500
rect 29644 163532 29696 163538
rect 29644 163474 29696 163480
rect 28908 29028 28960 29034
rect 28908 28970 28960 28976
rect 29748 28422 29776 368494
rect 29828 367124 29880 367130
rect 29828 367066 29880 367072
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 28724 26036 28776 26042
rect 28724 25978 28776 25984
rect 29840 25702 29868 367066
rect 29932 27402 29960 386378
rect 30024 198830 30052 561070
rect 30012 198824 30064 198830
rect 30012 198766 30064 198772
rect 30116 169318 30144 562119
rect 30286 560280 30342 560289
rect 30286 560215 30342 560224
rect 30196 546508 30248 546514
rect 30196 546450 30248 546456
rect 30104 169312 30156 169318
rect 30104 169254 30156 169260
rect 30208 27441 30236 546450
rect 30194 27432 30250 27441
rect 29920 27396 29972 27402
rect 30194 27367 30250 27376
rect 29920 27338 29972 27344
rect 29828 25696 29880 25702
rect 29828 25638 29880 25644
rect 30300 24721 30328 560215
rect 30748 371272 30800 371278
rect 30748 371214 30800 371220
rect 30760 25770 30788 371214
rect 30932 285728 30984 285734
rect 30932 285670 30984 285676
rect 30840 240168 30892 240174
rect 30840 240110 30892 240116
rect 30852 195906 30880 240110
rect 30840 195900 30892 195906
rect 30840 195842 30892 195848
rect 30944 95198 30972 285670
rect 31036 255270 31064 683198
rect 35254 679552 35310 679561
rect 35254 679487 35310 679496
rect 34242 625968 34298 625977
rect 34242 625903 34298 625912
rect 34150 622840 34206 622849
rect 34150 622775 34206 622784
rect 34164 605834 34192 622775
rect 34072 605806 34192 605834
rect 34072 596174 34100 605806
rect 34256 601066 34284 625903
rect 34426 623792 34482 623801
rect 34426 623727 34482 623736
rect 33980 596146 34100 596174
rect 34164 601038 34284 601066
rect 33980 589898 34008 596146
rect 34164 593722 34192 601038
rect 34334 598360 34390 598369
rect 34334 598295 34390 598304
rect 34242 598088 34298 598097
rect 34242 598023 34298 598032
rect 34072 593694 34192 593722
rect 34072 589966 34100 593694
rect 34152 593564 34204 593570
rect 34152 593506 34204 593512
rect 34164 590034 34192 593506
rect 34256 593450 34284 598023
rect 34348 593570 34376 598295
rect 34336 593564 34388 593570
rect 34336 593506 34388 593512
rect 34256 593422 34376 593450
rect 34152 590028 34204 590034
rect 34152 589970 34204 589976
rect 34060 589960 34112 589966
rect 34060 589902 34112 589908
rect 33968 589892 34020 589898
rect 33968 589834 34020 589840
rect 32772 588668 32824 588674
rect 32772 588610 32824 588616
rect 31576 586560 31628 586566
rect 31576 586502 31628 586508
rect 31300 565888 31352 565894
rect 31300 565830 31352 565836
rect 31116 563100 31168 563106
rect 31116 563042 31168 563048
rect 31128 411262 31156 563042
rect 31116 411256 31168 411262
rect 31116 411198 31168 411204
rect 31312 325650 31340 565830
rect 31392 564120 31444 564126
rect 31392 564062 31444 564068
rect 31404 367062 31432 564062
rect 31484 411324 31536 411330
rect 31484 411266 31536 411272
rect 31392 367056 31444 367062
rect 31392 366998 31444 367004
rect 31300 325644 31352 325650
rect 31300 325586 31352 325592
rect 31300 303680 31352 303686
rect 31300 303622 31352 303628
rect 31024 255264 31076 255270
rect 31024 255206 31076 255212
rect 31024 242956 31076 242962
rect 31024 242898 31076 242904
rect 31036 153950 31064 242898
rect 31116 223644 31168 223650
rect 31116 223586 31168 223592
rect 31024 153944 31076 153950
rect 31024 153886 31076 153892
rect 30932 95192 30984 95198
rect 30932 95134 30984 95140
rect 31128 26994 31156 223586
rect 31208 220856 31260 220862
rect 31208 220798 31260 220804
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 30748 25764 30800 25770
rect 30748 25706 30800 25712
rect 30286 24712 30342 24721
rect 30286 24647 30342 24656
rect 31220 24546 31248 220798
rect 31312 29073 31340 303622
rect 31496 29345 31524 411266
rect 31588 198286 31616 586502
rect 32588 565956 32640 565962
rect 32588 565898 32640 565904
rect 31666 560688 31722 560697
rect 31666 560623 31722 560632
rect 31576 198280 31628 198286
rect 31576 198222 31628 198228
rect 31680 100706 31708 560623
rect 32600 451246 32628 565898
rect 32680 561672 32732 561678
rect 32680 561614 32732 561620
rect 32588 451240 32640 451246
rect 32588 451182 32640 451188
rect 32588 429208 32640 429214
rect 32588 429150 32640 429156
rect 32496 379568 32548 379574
rect 32496 379510 32548 379516
rect 32404 309188 32456 309194
rect 32404 309130 32456 309136
rect 32312 218068 32364 218074
rect 32312 218010 32364 218016
rect 32220 215348 32272 215354
rect 32220 215290 32272 215296
rect 31758 171864 31814 171873
rect 31758 171799 31814 171808
rect 31668 100700 31720 100706
rect 31668 100642 31720 100648
rect 31482 29336 31538 29345
rect 31482 29271 31538 29280
rect 31298 29064 31354 29073
rect 31298 28999 31354 29008
rect 31208 24540 31260 24546
rect 31208 24482 31260 24488
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 31772 16574 31800 171799
rect 32232 155514 32260 215290
rect 32220 155508 32272 155514
rect 32220 155450 32272 155456
rect 32324 24818 32352 218010
rect 32416 195974 32444 309130
rect 32404 195968 32456 195974
rect 32404 195910 32456 195916
rect 32508 140758 32536 379510
rect 32600 155242 32628 429150
rect 32692 358766 32720 561614
rect 32680 358760 32732 358766
rect 32680 358702 32732 358708
rect 32680 314696 32732 314702
rect 32680 314638 32732 314644
rect 32588 155236 32640 155242
rect 32588 155178 32640 155184
rect 32496 140752 32548 140758
rect 32496 140694 32548 140700
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32692 22506 32720 314638
rect 32784 293962 32812 588610
rect 33048 587308 33100 587314
rect 33048 587250 33100 587256
rect 32956 565412 33008 565418
rect 32956 565354 33008 565360
rect 32864 562012 32916 562018
rect 32864 561954 32916 561960
rect 32772 293956 32824 293962
rect 32772 293898 32824 293904
rect 32772 237448 32824 237454
rect 32772 237390 32824 237396
rect 32784 27198 32812 237390
rect 32876 197946 32904 561954
rect 32864 197940 32916 197946
rect 32864 197882 32916 197888
rect 32968 196926 32996 565354
rect 33060 198490 33088 587250
rect 34244 587104 34296 587110
rect 34244 587046 34296 587052
rect 33968 564664 34020 564670
rect 33968 564606 34020 564612
rect 33874 558784 33930 558793
rect 33874 558719 33930 558728
rect 33692 418192 33744 418198
rect 33692 418134 33744 418140
rect 33600 231872 33652 231878
rect 33600 231814 33652 231820
rect 33048 198484 33100 198490
rect 33048 198426 33100 198432
rect 32956 196920 33008 196926
rect 32956 196862 33008 196868
rect 33612 28490 33640 231814
rect 33704 186998 33732 418134
rect 33784 398880 33836 398886
rect 33784 398822 33836 398828
rect 33692 186992 33744 186998
rect 33692 186934 33744 186940
rect 33796 64870 33824 398822
rect 33888 211818 33916 558719
rect 33876 211812 33928 211818
rect 33876 211754 33928 211760
rect 33876 211200 33928 211206
rect 33876 211142 33928 211148
rect 33888 153882 33916 211142
rect 33980 203561 34008 564606
rect 34150 561096 34206 561105
rect 34150 561031 34206 561040
rect 34060 545148 34112 545154
rect 34060 545090 34112 545096
rect 33966 203552 34022 203561
rect 33966 203487 34022 203496
rect 33968 181620 34020 181626
rect 33968 181562 34020 181568
rect 33876 153876 33928 153882
rect 33876 153818 33928 153824
rect 33784 64864 33836 64870
rect 33784 64806 33836 64812
rect 33600 28484 33652 28490
rect 33600 28426 33652 28432
rect 32772 27192 32824 27198
rect 32772 27134 32824 27140
rect 32680 22500 32732 22506
rect 32680 22442 32732 22448
rect 13832 16546 14320 16574
rect 19352 16546 19472 16574
rect 27632 16546 28488 16574
rect 31772 16546 31984 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 19444 480 19472 16546
rect 24214 3496 24270 3505
rect 24214 3431 24270 3440
rect 24228 480 24256 3431
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 33980 15978 34008 181562
rect 34072 178906 34100 545090
rect 34164 193050 34192 561031
rect 34256 196654 34284 587046
rect 34348 196897 34376 593422
rect 34440 570625 34468 623727
rect 34886 619984 34942 619993
rect 34886 619919 34942 619928
rect 34426 570616 34482 570625
rect 34426 570551 34482 570560
rect 34426 560824 34482 560833
rect 34426 560759 34482 560768
rect 34334 196888 34390 196897
rect 34334 196823 34390 196832
rect 34244 196648 34296 196654
rect 34244 196590 34296 196596
rect 34152 193044 34204 193050
rect 34152 192986 34204 192992
rect 34152 189984 34204 189990
rect 34152 189926 34204 189932
rect 34060 178900 34112 178906
rect 34060 178842 34112 178848
rect 34164 23458 34192 189926
rect 34336 187060 34388 187066
rect 34336 187002 34388 187008
rect 34244 181824 34296 181830
rect 34244 181766 34296 181772
rect 34152 23452 34204 23458
rect 34152 23394 34204 23400
rect 33968 15972 34020 15978
rect 33968 15914 34020 15920
rect 34256 3670 34284 181766
rect 34348 3738 34376 187002
rect 34440 89690 34468 560759
rect 34900 202842 34928 619919
rect 35072 568608 35124 568614
rect 35072 568550 35124 568556
rect 34980 421592 35032 421598
rect 34980 421534 35032 421540
rect 34992 249082 35020 421534
rect 35084 353258 35112 568550
rect 35268 425066 35296 679487
rect 40052 676870 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 690674 71820 702986
rect 89180 700369 89208 703520
rect 105464 700534 105492 703520
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 89166 700360 89222 700369
rect 89166 700295 89222 700304
rect 137848 698970 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 698964 137888 698970
rect 137836 698906 137888 698912
rect 153212 694822 153240 702406
rect 153200 694816 153252 694822
rect 153200 694758 153252 694764
rect 71780 690668 71832 690674
rect 71780 690610 71832 690616
rect 40040 676864 40092 676870
rect 40040 676806 40092 676812
rect 169772 676190 169800 702406
rect 202800 700466 202828 703520
rect 218992 700602 219020 703520
rect 218980 700596 219032 700602
rect 218980 700538 219032 700544
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 234632 687954 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700398 267688 703520
rect 283852 700670 283880 703520
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 267648 700392 267700 700398
rect 267648 700334 267700 700340
rect 299492 688022 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 689382 331260 702986
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 347228 700596 347280 700602
rect 347228 700538 347280 700544
rect 347136 700528 347188 700534
rect 347136 700470 347188 700476
rect 331220 689376 331272 689382
rect 331220 689318 331272 689324
rect 299480 688016 299532 688022
rect 299480 687958 299532 687964
rect 234620 687948 234672 687954
rect 234620 687890 234672 687896
rect 173164 685432 173216 685438
rect 173164 685374 173216 685380
rect 166908 676184 166960 676190
rect 166906 676152 166908 676161
rect 169760 676184 169812 676190
rect 166960 676152 166962 676161
rect 169760 676126 169812 676132
rect 166906 676087 166962 676096
rect 154486 674928 154542 674937
rect 154486 674863 154488 674872
rect 154540 674863 154542 674872
rect 172704 674892 172756 674898
rect 154488 674834 154540 674840
rect 172704 674834 172756 674840
rect 172610 668672 172666 668681
rect 172610 668607 172666 668616
rect 35622 626920 35678 626929
rect 35622 626855 35678 626864
rect 35438 621072 35494 621081
rect 35438 621007 35494 621016
rect 35348 588736 35400 588742
rect 35348 588678 35400 588684
rect 35256 425060 35308 425066
rect 35256 425002 35308 425008
rect 35256 420980 35308 420986
rect 35256 420922 35308 420928
rect 35164 403028 35216 403034
rect 35164 402970 35216 402976
rect 35072 353252 35124 353258
rect 35072 353194 35124 353200
rect 35072 351212 35124 351218
rect 35072 351154 35124 351160
rect 35084 267034 35112 351154
rect 35072 267028 35124 267034
rect 35072 266970 35124 266976
rect 35072 253972 35124 253978
rect 35072 253914 35124 253920
rect 34980 249076 35032 249082
rect 34980 249018 35032 249024
rect 34888 202836 34940 202842
rect 34888 202778 34940 202784
rect 35084 152658 35112 253914
rect 35176 163742 35204 402970
rect 35268 170610 35296 420922
rect 35360 238746 35388 588678
rect 35452 578950 35480 621007
rect 35530 618216 35586 618225
rect 35530 618151 35586 618160
rect 35440 578944 35492 578950
rect 35440 578886 35492 578892
rect 35544 573442 35572 618151
rect 35636 589082 35664 626855
rect 35714 599992 35770 600001
rect 35714 599927 35770 599936
rect 35624 589076 35676 589082
rect 35624 589018 35676 589024
rect 35622 587208 35678 587217
rect 35622 587143 35678 587152
rect 35532 573436 35584 573442
rect 35532 573378 35584 573384
rect 35532 562284 35584 562290
rect 35532 562226 35584 562232
rect 35440 561468 35492 561474
rect 35440 561410 35492 561416
rect 35348 238740 35400 238746
rect 35348 238682 35400 238688
rect 35348 222216 35400 222222
rect 35348 222158 35400 222164
rect 35256 170604 35308 170610
rect 35256 170546 35308 170552
rect 35164 163736 35216 163742
rect 35164 163678 35216 163684
rect 35072 152652 35124 152658
rect 35072 152594 35124 152600
rect 34428 89684 34480 89690
rect 34428 89626 34480 89632
rect 35360 28626 35388 222158
rect 35452 199306 35480 561410
rect 35440 199300 35492 199306
rect 35440 199242 35492 199248
rect 35544 195158 35572 562226
rect 35636 198393 35664 587143
rect 35728 199073 35756 599927
rect 36452 589960 36504 589966
rect 36452 589902 36504 589908
rect 36268 390584 36320 390590
rect 36268 390526 36320 390532
rect 35808 239420 35860 239426
rect 35808 239362 35860 239368
rect 35820 220153 35848 239362
rect 35806 220144 35862 220153
rect 35806 220079 35862 220088
rect 35808 218136 35860 218142
rect 35808 218078 35860 218084
rect 35714 199064 35770 199073
rect 35714 198999 35770 199008
rect 35622 198384 35678 198393
rect 35622 198319 35678 198328
rect 35532 195152 35584 195158
rect 35532 195094 35584 195100
rect 35532 187264 35584 187270
rect 35532 187206 35584 187212
rect 35348 28620 35400 28626
rect 35348 28562 35400 28568
rect 35544 27606 35572 187206
rect 35716 184272 35768 184278
rect 35716 184214 35768 184220
rect 35624 181756 35676 181762
rect 35624 181698 35676 181704
rect 35532 27600 35584 27606
rect 35532 27542 35584 27548
rect 35636 15910 35664 181698
rect 35728 19310 35756 184214
rect 35820 28558 35848 218078
rect 35808 28552 35860 28558
rect 35808 28494 35860 28500
rect 36280 23118 36308 390526
rect 36464 386374 36492 589902
rect 36544 589892 36596 589898
rect 36544 589834 36596 589840
rect 36452 386368 36504 386374
rect 36452 386310 36504 386316
rect 36452 384328 36504 384334
rect 36452 384270 36504 384276
rect 36360 348424 36412 348430
rect 36360 348366 36412 348372
rect 36372 262206 36400 348366
rect 36360 262200 36412 262206
rect 36360 262142 36412 262148
rect 36360 247104 36412 247110
rect 36360 247046 36412 247052
rect 36372 152590 36400 247046
rect 36464 231810 36492 384270
rect 36452 231804 36504 231810
rect 36452 231746 36504 231752
rect 36556 198121 36584 589834
rect 84382 589520 84438 589529
rect 84382 589455 84438 589464
rect 47584 589280 47636 589286
rect 47584 589222 47636 589228
rect 39856 589212 39908 589218
rect 39856 589154 39908 589160
rect 39396 589008 39448 589014
rect 39396 588950 39448 588956
rect 37188 587240 37240 587246
rect 37188 587182 37240 587188
rect 36820 566024 36872 566030
rect 36820 565966 36872 565972
rect 36636 559564 36688 559570
rect 36636 559506 36688 559512
rect 36648 331226 36676 559506
rect 36832 463690 36860 565966
rect 36912 564868 36964 564874
rect 36912 564810 36964 564816
rect 36820 463684 36872 463690
rect 36820 463626 36872 463632
rect 36728 427848 36780 427854
rect 36728 427790 36780 427796
rect 36636 331220 36688 331226
rect 36636 331162 36688 331168
rect 36636 268116 36688 268122
rect 36636 268058 36688 268064
rect 36648 242214 36676 268058
rect 36636 242208 36688 242214
rect 36636 242150 36688 242156
rect 36636 230512 36688 230518
rect 36636 230454 36688 230460
rect 36542 198112 36598 198121
rect 36542 198047 36598 198056
rect 36648 196382 36676 230454
rect 36740 196586 36768 427790
rect 36820 418260 36872 418266
rect 36820 418202 36872 418208
rect 36728 196580 36780 196586
rect 36728 196522 36780 196528
rect 36636 196376 36688 196382
rect 36636 196318 36688 196324
rect 36544 187128 36596 187134
rect 36544 187070 36596 187076
rect 36450 184512 36506 184521
rect 36450 184447 36506 184456
rect 36360 152584 36412 152590
rect 36360 152526 36412 152532
rect 36464 131102 36492 184447
rect 36452 131096 36504 131102
rect 36452 131038 36504 131044
rect 36556 33046 36584 187070
rect 36636 184204 36688 184210
rect 36636 184146 36688 184152
rect 36544 33040 36596 33046
rect 36544 32982 36596 32988
rect 36268 23112 36320 23118
rect 36268 23054 36320 23060
rect 35716 19304 35768 19310
rect 35716 19246 35768 19252
rect 36648 18970 36676 184146
rect 36728 174616 36780 174622
rect 36728 174558 36780 174564
rect 36636 18964 36688 18970
rect 36636 18906 36688 18912
rect 35624 15904 35676 15910
rect 35624 15846 35676 15852
rect 34336 3732 34388 3738
rect 34336 3674 34388 3680
rect 34244 3664 34296 3670
rect 34244 3606 34296 3612
rect 35990 3496 36046 3505
rect 36740 3466 36768 174558
rect 36832 128314 36860 418202
rect 36924 218754 36952 564810
rect 37004 562420 37056 562426
rect 37004 562362 37056 562368
rect 36912 218748 36964 218754
rect 36912 218690 36964 218696
rect 36912 216708 36964 216714
rect 36912 216650 36964 216656
rect 36924 197742 36952 216650
rect 37016 205222 37044 562362
rect 37096 561196 37148 561202
rect 37096 561138 37148 561144
rect 37004 205216 37056 205222
rect 37004 205158 37056 205164
rect 37004 202904 37056 202910
rect 37004 202846 37056 202852
rect 36912 197736 36964 197742
rect 36912 197678 36964 197684
rect 36912 192908 36964 192914
rect 36912 192850 36964 192856
rect 36820 128308 36872 128314
rect 36820 128250 36872 128256
rect 36924 18902 36952 192850
rect 37016 26654 37044 202846
rect 37108 198966 37136 561138
rect 37200 390522 37228 587182
rect 39304 564800 39356 564806
rect 39304 564742 39356 564748
rect 38108 564732 38160 564738
rect 38108 564674 38160 564680
rect 38014 560008 38070 560017
rect 38014 559943 38070 559952
rect 37648 469260 37700 469266
rect 37648 469202 37700 469208
rect 37188 390516 37240 390522
rect 37188 390458 37240 390464
rect 37188 205692 37240 205698
rect 37188 205634 37240 205640
rect 37200 199753 37228 205634
rect 37186 199744 37242 199753
rect 37186 199679 37242 199688
rect 37096 198960 37148 198966
rect 37096 198902 37148 198908
rect 37096 181688 37148 181694
rect 37096 181630 37148 181636
rect 37004 26648 37056 26654
rect 37004 26590 37056 26596
rect 36912 18896 36964 18902
rect 36912 18838 36964 18844
rect 37108 3602 37136 181630
rect 37660 27810 37688 469202
rect 37924 433356 37976 433362
rect 37924 433298 37976 433304
rect 37832 392080 37884 392086
rect 37832 392022 37884 392028
rect 37738 220824 37794 220833
rect 37738 220759 37794 220768
rect 37752 205737 37780 220759
rect 37738 205728 37794 205737
rect 37738 205663 37794 205672
rect 37740 205216 37792 205222
rect 37740 205158 37792 205164
rect 37752 153202 37780 205158
rect 37844 184618 37872 392022
rect 37832 184612 37884 184618
rect 37832 184554 37884 184560
rect 37936 182918 37964 433298
rect 38028 387122 38056 559943
rect 38016 387116 38068 387122
rect 38016 387058 38068 387064
rect 38016 385076 38068 385082
rect 38016 385018 38068 385024
rect 37924 182912 37976 182918
rect 37924 182854 37976 182860
rect 37740 153196 37792 153202
rect 37740 153138 37792 153144
rect 38028 121446 38056 385018
rect 38120 218113 38148 564674
rect 39212 563440 39264 563446
rect 39212 563382 39264 563388
rect 38476 563168 38528 563174
rect 38476 563110 38528 563116
rect 38384 562148 38436 562154
rect 38384 562090 38436 562096
rect 38200 561332 38252 561338
rect 38200 561274 38252 561280
rect 38106 218104 38162 218113
rect 38106 218039 38162 218048
rect 38108 213988 38160 213994
rect 38108 213930 38160 213936
rect 38016 121440 38068 121446
rect 38016 121382 38068 121388
rect 37648 27804 37700 27810
rect 37648 27746 37700 27752
rect 38120 24410 38148 213930
rect 38212 199238 38240 561274
rect 38292 561060 38344 561066
rect 38292 561002 38344 561008
rect 38200 199232 38252 199238
rect 38200 199174 38252 199180
rect 38304 198937 38332 561002
rect 38290 198928 38346 198937
rect 38290 198863 38346 198872
rect 38396 195566 38424 562090
rect 38488 460902 38516 563110
rect 39028 529984 39080 529990
rect 39028 529926 39080 529932
rect 38568 480276 38620 480282
rect 38568 480218 38620 480224
rect 38476 460896 38528 460902
rect 38476 460838 38528 460844
rect 38384 195560 38436 195566
rect 38384 195502 38436 195508
rect 38200 187672 38252 187678
rect 38200 187614 38252 187620
rect 38212 86970 38240 187614
rect 38292 187196 38344 187202
rect 38292 187138 38344 187144
rect 38200 86964 38252 86970
rect 38200 86906 38252 86912
rect 38304 69018 38332 187138
rect 38384 152992 38436 152998
rect 38384 152934 38436 152940
rect 38292 69012 38344 69018
rect 38292 68954 38344 68960
rect 38108 24404 38160 24410
rect 38108 24346 38160 24352
rect 38396 20398 38424 152934
rect 38580 28665 38608 480218
rect 38660 173256 38712 173262
rect 38660 173198 38712 173204
rect 38566 28656 38622 28665
rect 38566 28591 38622 28600
rect 38384 20392 38436 20398
rect 38384 20334 38436 20340
rect 38672 16574 38700 173198
rect 39040 68950 39068 529926
rect 39224 487830 39252 563382
rect 39212 487824 39264 487830
rect 39212 487766 39264 487772
rect 39316 351218 39344 564742
rect 39408 501906 39436 588950
rect 39764 562488 39816 562494
rect 39764 562430 39816 562436
rect 39488 560992 39540 560998
rect 39488 560934 39540 560940
rect 39396 501900 39448 501906
rect 39396 501842 39448 501848
rect 39396 467968 39448 467974
rect 39396 467910 39448 467916
rect 39304 351212 39356 351218
rect 39304 351154 39356 351160
rect 39304 332580 39356 332586
rect 39304 332522 39356 332528
rect 39212 322992 39264 322998
rect 39212 322934 39264 322940
rect 39120 267028 39172 267034
rect 39120 266970 39172 266976
rect 39132 224738 39160 266970
rect 39120 224732 39172 224738
rect 39120 224674 39172 224680
rect 39224 199889 39252 322934
rect 39316 268122 39344 332522
rect 39304 268116 39356 268122
rect 39304 268058 39356 268064
rect 39304 225548 39356 225554
rect 39304 225490 39356 225496
rect 39210 199880 39266 199889
rect 39210 199815 39266 199824
rect 39028 68944 39080 68950
rect 39028 68886 39080 68892
rect 39316 29238 39344 225490
rect 39408 160886 39436 467910
rect 39500 199102 39528 560934
rect 39578 560144 39634 560153
rect 39578 560079 39634 560088
rect 39592 394806 39620 560079
rect 39672 558952 39724 558958
rect 39672 558894 39724 558900
rect 39580 394800 39632 394806
rect 39580 394742 39632 394748
rect 39580 393372 39632 393378
rect 39580 393314 39632 393320
rect 39488 199096 39540 199102
rect 39488 199038 39540 199044
rect 39396 160880 39448 160886
rect 39396 160822 39448 160828
rect 39304 29232 39356 29238
rect 39304 29174 39356 29180
rect 39592 27878 39620 393314
rect 39684 192982 39712 558894
rect 39776 195090 39804 562430
rect 39868 500954 39896 589154
rect 42064 588940 42116 588946
rect 42064 588882 42116 588888
rect 40776 588872 40828 588878
rect 40776 588814 40828 588820
rect 40592 564596 40644 564602
rect 40592 564538 40644 564544
rect 40500 562216 40552 562222
rect 40500 562158 40552 562164
rect 40408 516180 40460 516186
rect 40408 516122 40460 516128
rect 39856 500948 39908 500954
rect 39856 500890 39908 500896
rect 39856 434784 39908 434790
rect 39856 434726 39908 434732
rect 39764 195084 39816 195090
rect 39764 195026 39816 195032
rect 39672 192976 39724 192982
rect 39672 192918 39724 192924
rect 39672 183048 39724 183054
rect 39672 182990 39724 182996
rect 39580 27872 39632 27878
rect 39580 27814 39632 27820
rect 39684 19990 39712 182990
rect 39764 174752 39816 174758
rect 39764 174694 39816 174700
rect 39672 19984 39724 19990
rect 39672 19926 39724 19932
rect 38672 16546 39160 16574
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 35990 3431 36046 3440
rect 36728 3460 36780 3466
rect 36004 480 36032 3431
rect 36728 3402 36780 3408
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39776 3534 39804 174694
rect 39868 29102 39896 434726
rect 39948 221468 40000 221474
rect 39948 221410 40000 221416
rect 39960 195838 39988 221410
rect 40420 198218 40448 516122
rect 40512 509318 40540 562158
rect 40500 509312 40552 509318
rect 40500 509254 40552 509260
rect 40604 421598 40632 564538
rect 40684 563780 40736 563786
rect 40684 563722 40736 563728
rect 40592 421592 40644 421598
rect 40592 421534 40644 421540
rect 40592 419620 40644 419626
rect 40592 419562 40644 419568
rect 40500 270292 40552 270298
rect 40500 270234 40552 270240
rect 40512 198898 40540 270234
rect 40500 198892 40552 198898
rect 40500 198834 40552 198840
rect 40408 198212 40460 198218
rect 40408 198154 40460 198160
rect 40604 196518 40632 419562
rect 40696 221474 40724 563722
rect 40788 525706 40816 588814
rect 40868 588804 40920 588810
rect 40868 588746 40920 588752
rect 40776 525700 40828 525706
rect 40776 525642 40828 525648
rect 40774 510504 40830 510513
rect 40774 510439 40830 510448
rect 40788 276049 40816 510439
rect 40880 456686 40908 588746
rect 41328 586900 41380 586906
rect 41328 586842 41380 586848
rect 40960 584452 41012 584458
rect 40960 584394 41012 584400
rect 40972 480690 41000 584394
rect 41236 577516 41288 577522
rect 41236 577458 41288 577464
rect 41052 564460 41104 564466
rect 41052 564402 41104 564408
rect 41064 496806 41092 564402
rect 41144 550860 41196 550866
rect 41144 550802 41196 550808
rect 41052 496800 41104 496806
rect 41052 496742 41104 496748
rect 40960 480684 41012 480690
rect 40960 480626 41012 480632
rect 40960 464160 41012 464166
rect 40960 464102 41012 464108
rect 40868 456680 40920 456686
rect 40868 456622 40920 456628
rect 40868 425128 40920 425134
rect 40868 425070 40920 425076
rect 40774 276040 40830 276049
rect 40774 275975 40830 275984
rect 40776 274916 40828 274922
rect 40776 274858 40828 274864
rect 40684 221468 40736 221474
rect 40684 221410 40736 221416
rect 40682 204912 40738 204921
rect 40682 204847 40738 204856
rect 40592 196512 40644 196518
rect 40592 196454 40644 196460
rect 39948 195832 40000 195838
rect 39948 195774 40000 195780
rect 40592 192296 40644 192302
rect 40592 192238 40644 192244
rect 40500 178764 40552 178770
rect 40500 178706 40552 178712
rect 40408 174684 40460 174690
rect 40408 174626 40460 174632
rect 40420 57934 40448 174626
rect 40512 100065 40540 178706
rect 40604 104854 40632 192238
rect 40592 104848 40644 104854
rect 40592 104790 40644 104796
rect 40498 100056 40554 100065
rect 40498 99991 40554 100000
rect 40408 57928 40460 57934
rect 40408 57870 40460 57876
rect 39856 29096 39908 29102
rect 39856 29038 39908 29044
rect 40696 28218 40724 204847
rect 40788 195634 40816 274858
rect 40776 195628 40828 195634
rect 40776 195570 40828 195576
rect 40776 185836 40828 185842
rect 40776 185778 40828 185784
rect 40788 67590 40816 185778
rect 40880 167686 40908 425070
rect 40972 184346 41000 464102
rect 41052 220448 41104 220454
rect 41052 220390 41104 220396
rect 41064 199714 41092 220390
rect 41052 199708 41104 199714
rect 41052 199650 41104 199656
rect 41156 193866 41184 550802
rect 41248 206990 41276 577458
rect 41236 206984 41288 206990
rect 41236 206926 41288 206932
rect 41340 197334 41368 586842
rect 41880 563916 41932 563922
rect 41880 563858 41932 563864
rect 41892 369918 41920 563858
rect 42076 498166 42104 588882
rect 43720 588532 43772 588538
rect 43720 588474 43772 588480
rect 42524 587512 42576 587518
rect 42524 587454 42576 587460
rect 42432 564936 42484 564942
rect 42432 564878 42484 564884
rect 42340 561944 42392 561950
rect 42340 561886 42392 561892
rect 42248 528624 42300 528630
rect 42248 528566 42300 528572
rect 42156 513392 42208 513398
rect 42156 513334 42208 513340
rect 42064 498160 42116 498166
rect 42064 498102 42116 498108
rect 42064 484492 42116 484498
rect 42064 484434 42116 484440
rect 41972 400240 42024 400246
rect 41972 400182 42024 400188
rect 41880 369912 41932 369918
rect 41880 369854 41932 369860
rect 41788 214600 41840 214606
rect 41788 214542 41840 214548
rect 41328 197328 41380 197334
rect 41328 197270 41380 197276
rect 41144 193860 41196 193866
rect 41144 193802 41196 193808
rect 41328 190120 41380 190126
rect 41328 190062 41380 190068
rect 41234 189952 41290 189961
rect 41234 189887 41290 189896
rect 40960 184340 41012 184346
rect 40960 184282 41012 184288
rect 41050 180296 41106 180305
rect 41050 180231 41106 180240
rect 40868 167680 40920 167686
rect 40868 167622 40920 167628
rect 40960 155644 41012 155650
rect 40960 155586 41012 155592
rect 40776 67584 40828 67590
rect 40776 67526 40828 67532
rect 40684 28212 40736 28218
rect 40684 28154 40736 28160
rect 40972 17746 41000 155586
rect 41064 26926 41092 180231
rect 41144 166524 41196 166530
rect 41144 166466 41196 166472
rect 41052 26920 41104 26926
rect 41052 26862 41104 26868
rect 40960 17740 41012 17746
rect 40960 17682 41012 17688
rect 41156 3874 41184 166466
rect 41248 24274 41276 189887
rect 41236 24268 41288 24274
rect 41236 24210 41288 24216
rect 41340 19038 41368 190062
rect 41800 24857 41828 214542
rect 41878 200016 41934 200025
rect 41878 199951 41934 199960
rect 41892 26790 41920 199951
rect 41984 179042 42012 400182
rect 42076 190398 42104 484434
rect 42168 195226 42196 513334
rect 42260 196722 42288 528566
rect 42352 200122 42380 561886
rect 42444 401878 42472 564878
rect 42536 495446 42564 587454
rect 43536 567860 43588 567866
rect 43536 567802 43588 567808
rect 43444 563576 43496 563582
rect 43444 563518 43496 563524
rect 43352 562692 43404 562698
rect 43352 562634 43404 562640
rect 42708 551132 42760 551138
rect 42708 551074 42760 551080
rect 42616 549296 42668 549302
rect 42616 549238 42668 549244
rect 42524 495440 42576 495446
rect 42524 495382 42576 495388
rect 42524 438932 42576 438938
rect 42524 438874 42576 438880
rect 42432 401872 42484 401878
rect 42432 401814 42484 401820
rect 42432 396500 42484 396506
rect 42432 396442 42484 396448
rect 42340 200116 42392 200122
rect 42340 200058 42392 200064
rect 42248 196716 42300 196722
rect 42248 196658 42300 196664
rect 42156 195220 42208 195226
rect 42156 195162 42208 195168
rect 42064 190392 42116 190398
rect 42064 190334 42116 190340
rect 42248 190188 42300 190194
rect 42248 190130 42300 190136
rect 42156 185768 42208 185774
rect 42156 185710 42208 185716
rect 42064 181892 42116 181898
rect 42064 181834 42116 181840
rect 41972 179036 42024 179042
rect 41972 178978 42024 178984
rect 41880 26784 41932 26790
rect 41880 26726 41932 26732
rect 41786 24848 41842 24857
rect 41786 24783 41842 24792
rect 41328 19032 41380 19038
rect 41328 18974 41380 18980
rect 42076 17814 42104 181834
rect 42064 17808 42116 17814
rect 42064 17750 42116 17756
rect 42168 4078 42196 185710
rect 42156 4072 42208 4078
rect 42156 4014 42208 4020
rect 41144 3868 41196 3874
rect 41144 3810 41196 3816
rect 42260 3806 42288 190130
rect 42444 27266 42472 396442
rect 42536 29306 42564 438874
rect 42628 69698 42656 549238
rect 42616 69692 42668 69698
rect 42616 69634 42668 69640
rect 42720 62082 42748 551074
rect 43168 543788 43220 543794
rect 43168 543730 43220 543736
rect 43076 531820 43128 531826
rect 43076 531762 43128 531768
rect 42982 205728 43038 205737
rect 42982 205663 43038 205672
rect 42708 62076 42760 62082
rect 42708 62018 42760 62024
rect 42524 29300 42576 29306
rect 42524 29242 42576 29248
rect 42432 27260 42484 27266
rect 42432 27202 42484 27208
rect 42996 24002 43024 205663
rect 43088 133890 43116 531762
rect 43076 133884 43128 133890
rect 43076 133826 43128 133832
rect 43180 29510 43208 543730
rect 43364 474706 43392 562634
rect 43352 474700 43404 474706
rect 43352 474642 43404 474648
rect 43260 401872 43312 401878
rect 43260 401814 43312 401820
rect 43272 267782 43300 401814
rect 43456 374746 43484 563518
rect 43444 374740 43496 374746
rect 43444 374682 43496 374688
rect 43444 369912 43496 369918
rect 43444 369854 43496 369860
rect 43352 321632 43404 321638
rect 43352 321574 43404 321580
rect 43260 267776 43312 267782
rect 43260 267718 43312 267724
rect 43260 262200 43312 262206
rect 43260 262142 43312 262148
rect 43272 227866 43300 262142
rect 43260 227860 43312 227866
rect 43260 227802 43312 227808
rect 43260 178696 43312 178702
rect 43260 178638 43312 178644
rect 43272 102134 43300 178638
rect 43364 165034 43392 321574
rect 43456 317393 43484 369854
rect 43442 317384 43498 317393
rect 43442 317319 43498 317328
rect 43548 302190 43576 567802
rect 43628 560448 43680 560454
rect 43628 560390 43680 560396
rect 43640 456754 43668 560390
rect 43628 456748 43680 456754
rect 43628 456690 43680 456696
rect 43628 436144 43680 436150
rect 43628 436086 43680 436092
rect 43536 302184 43588 302190
rect 43536 302126 43588 302132
rect 43536 291236 43588 291242
rect 43536 291178 43588 291184
rect 43444 284368 43496 284374
rect 43444 284310 43496 284316
rect 43456 270298 43484 284310
rect 43444 270292 43496 270298
rect 43444 270234 43496 270240
rect 43444 267844 43496 267850
rect 43444 267786 43496 267792
rect 43456 199578 43484 267786
rect 43444 199572 43496 199578
rect 43444 199514 43496 199520
rect 43548 181558 43576 291178
rect 43536 181552 43588 181558
rect 43536 181494 43588 181500
rect 43352 165028 43404 165034
rect 43352 164970 43404 164976
rect 43640 163810 43668 436086
rect 43732 325718 43760 588474
rect 44732 587580 44784 587586
rect 44732 587522 44784 587528
rect 43904 583092 43956 583098
rect 43904 583034 43956 583040
rect 43812 576156 43864 576162
rect 43812 576098 43864 576104
rect 43720 325712 43772 325718
rect 43720 325654 43772 325660
rect 43720 318980 43772 318986
rect 43720 318922 43772 318928
rect 43628 163804 43680 163810
rect 43628 163746 43680 163752
rect 43628 155372 43680 155378
rect 43628 155314 43680 155320
rect 43260 102128 43312 102134
rect 43260 102070 43312 102076
rect 43168 29504 43220 29510
rect 43168 29446 43220 29452
rect 42984 23996 43036 24002
rect 42984 23938 43036 23944
rect 43640 20534 43668 155314
rect 43732 29170 43760 318922
rect 43824 208350 43852 576098
rect 43916 430574 43944 583034
rect 44640 565276 44692 565282
rect 44640 565218 44692 565224
rect 43994 563136 44050 563145
rect 43994 563071 44050 563080
rect 44008 510610 44036 563071
rect 44088 560380 44140 560386
rect 44088 560322 44140 560328
rect 44100 538218 44128 560322
rect 44548 556232 44600 556238
rect 44548 556174 44600 556180
rect 44088 538212 44140 538218
rect 44088 538154 44140 538160
rect 43996 510604 44048 510610
rect 43996 510546 44048 510552
rect 43904 430568 43956 430574
rect 43904 430510 43956 430516
rect 43904 415540 43956 415546
rect 43904 415482 43956 415488
rect 43812 208344 43864 208350
rect 43812 208286 43864 208292
rect 43812 189712 43864 189718
rect 43812 189654 43864 189660
rect 43720 29164 43772 29170
rect 43720 29106 43772 29112
rect 43824 21418 43852 189654
rect 43916 29442 43944 415482
rect 44364 313132 44416 313138
rect 44364 313074 44416 313080
rect 44180 267776 44232 267782
rect 44180 267718 44232 267724
rect 44192 264897 44220 267718
rect 44178 264888 44234 264897
rect 44178 264823 44234 264832
rect 44088 227792 44140 227798
rect 44088 227734 44140 227740
rect 44100 198082 44128 227734
rect 44272 224732 44324 224738
rect 44272 224674 44324 224680
rect 44178 220824 44234 220833
rect 44178 220759 44234 220768
rect 44192 214606 44220 220759
rect 44284 220318 44312 224674
rect 44272 220312 44324 220318
rect 44272 220254 44324 220260
rect 44180 214600 44232 214606
rect 44180 214542 44232 214548
rect 44272 200116 44324 200122
rect 44272 200058 44324 200064
rect 44088 198076 44140 198082
rect 44088 198018 44140 198024
rect 44088 183388 44140 183394
rect 44088 183330 44140 183336
rect 43996 151428 44048 151434
rect 43996 151370 44048 151376
rect 43904 29436 43956 29442
rect 43904 29378 43956 29384
rect 44008 22710 44036 151370
rect 43996 22704 44048 22710
rect 43996 22646 44048 22652
rect 44100 22642 44128 183330
rect 44284 27470 44312 200058
rect 44376 152386 44404 313074
rect 44456 234660 44508 234666
rect 44456 234602 44508 234608
rect 44468 176118 44496 234602
rect 44560 199646 44588 556174
rect 44652 318646 44680 565218
rect 44744 525774 44772 587522
rect 45376 587172 45428 587178
rect 45376 587114 45428 587120
rect 45008 586968 45060 586974
rect 45008 586910 45060 586916
rect 44824 563848 44876 563854
rect 44824 563790 44876 563796
rect 44732 525768 44784 525774
rect 44732 525710 44784 525716
rect 44732 445800 44784 445806
rect 44732 445742 44784 445748
rect 44640 318640 44692 318646
rect 44640 318582 44692 318588
rect 44640 292596 44692 292602
rect 44640 292538 44692 292544
rect 44548 199640 44600 199646
rect 44548 199582 44600 199588
rect 44652 191418 44680 292538
rect 44744 198354 44772 445742
rect 44836 284374 44864 563790
rect 44914 561368 44970 561377
rect 44914 561303 44970 561312
rect 44928 310321 44956 561303
rect 45020 481370 45048 586910
rect 45284 574932 45336 574938
rect 45284 574874 45336 574880
rect 45100 572144 45152 572150
rect 45100 572086 45152 572092
rect 45008 481364 45060 481370
rect 45008 481306 45060 481312
rect 45006 359408 45062 359417
rect 45006 359343 45062 359352
rect 44914 310312 44970 310321
rect 44914 310247 44970 310256
rect 44824 284368 44876 284374
rect 44824 284310 44876 284316
rect 44822 283248 44878 283257
rect 44822 283183 44878 283192
rect 44836 199442 44864 283183
rect 44824 199436 44876 199442
rect 44824 199378 44876 199384
rect 44732 198348 44784 198354
rect 44732 198290 44784 198296
rect 44640 191412 44692 191418
rect 44640 191354 44692 191360
rect 44732 183116 44784 183122
rect 44732 183058 44784 183064
rect 44638 177712 44694 177721
rect 44638 177647 44694 177656
rect 44456 176112 44508 176118
rect 44456 176054 44508 176060
rect 44364 152380 44416 152386
rect 44364 152322 44416 152328
rect 44652 115938 44680 177647
rect 44640 115932 44692 115938
rect 44640 115874 44692 115880
rect 44744 114510 44772 183058
rect 44916 152856 44968 152862
rect 44916 152798 44968 152804
rect 44732 114504 44784 114510
rect 44732 114446 44784 114452
rect 44272 27464 44324 27470
rect 44272 27406 44324 27412
rect 44088 22636 44140 22642
rect 44088 22578 44140 22584
rect 43812 21412 43864 21418
rect 43812 21354 43864 21360
rect 43628 20528 43680 20534
rect 43628 20470 43680 20476
rect 44928 19718 44956 152798
rect 45020 60042 45048 359343
rect 45112 264761 45140 572086
rect 45192 565344 45244 565350
rect 45192 565286 45244 565292
rect 45204 342242 45232 565286
rect 45192 342236 45244 342242
rect 45192 342178 45244 342184
rect 45190 339552 45246 339561
rect 45190 339487 45246 339496
rect 45098 264752 45154 264761
rect 45098 264687 45154 264696
rect 45100 247172 45152 247178
rect 45100 247114 45152 247120
rect 45112 244361 45140 247114
rect 45098 244352 45154 244361
rect 45098 244287 45154 244296
rect 45100 214600 45152 214606
rect 45100 214542 45152 214548
rect 45112 200569 45140 214542
rect 45098 200560 45154 200569
rect 45098 200495 45154 200504
rect 45098 155408 45154 155417
rect 45098 155343 45154 155352
rect 45008 60036 45060 60042
rect 45008 59978 45060 59984
rect 45112 22982 45140 155343
rect 45204 29646 45232 339487
rect 45296 257961 45324 574874
rect 45282 257952 45338 257961
rect 45282 257887 45338 257896
rect 45284 255740 45336 255746
rect 45284 255682 45336 255688
rect 45296 230586 45324 255682
rect 45388 247314 45416 587114
rect 47216 586016 47268 586022
rect 47216 585958 47268 585964
rect 46756 581732 46808 581738
rect 46756 581674 46808 581680
rect 46204 580372 46256 580378
rect 46204 580314 46256 580320
rect 45744 572008 45796 572014
rect 45744 571950 45796 571956
rect 45652 525700 45704 525706
rect 45652 525642 45704 525648
rect 45664 525201 45692 525642
rect 45650 525192 45706 525201
rect 45650 525127 45706 525136
rect 45756 510921 45784 571950
rect 45928 566704 45980 566710
rect 45928 566646 45980 566652
rect 45940 544241 45968 566646
rect 46110 556200 46166 556209
rect 46110 556135 46166 556144
rect 46124 549166 46152 556135
rect 46112 549160 46164 549166
rect 46112 549102 46164 549108
rect 46110 546544 46166 546553
rect 46110 546479 46112 546488
rect 46164 546479 46166 546488
rect 46112 546450 46164 546456
rect 46018 545728 46074 545737
rect 46018 545663 46074 545672
rect 46032 545154 46060 545663
rect 46020 545148 46072 545154
rect 46020 545090 46072 545096
rect 46110 544368 46166 544377
rect 46110 544303 46166 544312
rect 45926 544232 45982 544241
rect 45926 544167 45982 544176
rect 46124 543794 46152 544303
rect 46112 543788 46164 543794
rect 46112 543730 46164 543736
rect 46110 541104 46166 541113
rect 46110 541039 46166 541048
rect 46124 541006 46152 541039
rect 46112 541000 46164 541006
rect 46112 540942 46164 540948
rect 46112 538212 46164 538218
rect 46112 538154 46164 538160
rect 46124 538121 46152 538154
rect 46110 538112 46166 538121
rect 46110 538047 46166 538056
rect 46018 532264 46074 532273
rect 46018 532199 46074 532208
rect 46032 531826 46060 532199
rect 46020 531820 46072 531826
rect 46020 531762 46072 531768
rect 46112 529984 46164 529990
rect 46110 529952 46112 529961
rect 46164 529952 46166 529961
rect 46110 529887 46166 529896
rect 45834 529000 45890 529009
rect 45834 528935 45890 528944
rect 45848 528630 45876 528935
rect 45836 528624 45888 528630
rect 45836 528566 45888 528572
rect 46216 526561 46244 580314
rect 46480 579012 46532 579018
rect 46480 578954 46532 578960
rect 46388 563712 46440 563718
rect 46388 563654 46440 563660
rect 46294 556608 46350 556617
rect 46294 556543 46350 556552
rect 46308 556238 46336 556543
rect 46296 556232 46348 556238
rect 46296 556174 46348 556180
rect 46294 551440 46350 551449
rect 46294 551375 46350 551384
rect 46308 551138 46336 551375
rect 46296 551132 46348 551138
rect 46296 551074 46348 551080
rect 46294 550896 46350 550905
rect 46294 550831 46296 550840
rect 46348 550831 46350 550840
rect 46296 550802 46348 550808
rect 46294 549808 46350 549817
rect 46294 549743 46350 549752
rect 46308 549302 46336 549743
rect 46296 549296 46348 549302
rect 46296 549238 46348 549244
rect 46296 549160 46348 549166
rect 46296 549102 46348 549108
rect 46202 526552 46258 526561
rect 46202 526487 46258 526496
rect 46112 525768 46164 525774
rect 46112 525710 46164 525716
rect 46124 518894 46152 525710
rect 46202 520432 46258 520441
rect 46202 520367 46258 520376
rect 46216 520334 46244 520367
rect 46204 520328 46256 520334
rect 46204 520270 46256 520276
rect 46124 518866 46244 518894
rect 46018 516624 46074 516633
rect 46018 516559 46074 516568
rect 46032 516186 46060 516559
rect 46020 516180 46072 516186
rect 46020 516122 46072 516128
rect 45926 513904 45982 513913
rect 45926 513839 45982 513848
rect 45940 513398 45968 513839
rect 45928 513392 45980 513398
rect 45928 513334 45980 513340
rect 45742 510912 45798 510921
rect 45742 510847 45798 510856
rect 46112 510604 46164 510610
rect 46112 510546 46164 510552
rect 46124 509561 46152 510546
rect 46110 509552 46166 509561
rect 46110 509487 46166 509496
rect 46020 509312 46072 509318
rect 46020 509254 46072 509260
rect 45652 500948 45704 500954
rect 45652 500890 45704 500896
rect 45664 500721 45692 500890
rect 45650 500712 45706 500721
rect 45650 500647 45706 500656
rect 45928 498296 45980 498302
rect 45928 498238 45980 498244
rect 45940 494601 45968 498238
rect 45926 494592 45982 494601
rect 45926 494527 45982 494536
rect 45652 487824 45704 487830
rect 45652 487766 45704 487772
rect 45560 387116 45612 387122
rect 45560 387058 45612 387064
rect 45572 345014 45600 387058
rect 45664 384334 45692 487766
rect 45834 484528 45890 484537
rect 45834 484463 45890 484472
rect 45848 484430 45876 484463
rect 45836 484424 45888 484430
rect 45836 484366 45888 484372
rect 45926 445088 45982 445097
rect 45926 445023 45982 445032
rect 45940 444446 45968 445023
rect 45928 444440 45980 444446
rect 45928 444382 45980 444388
rect 45926 439648 45982 439657
rect 45926 439583 45982 439592
rect 45940 438938 45968 439583
rect 45928 438932 45980 438938
rect 45928 438874 45980 438880
rect 45926 403608 45982 403617
rect 45926 403543 45982 403552
rect 45940 403034 45968 403543
rect 45928 403028 45980 403034
rect 45928 402970 45980 402976
rect 45836 394800 45888 394806
rect 45836 394742 45888 394748
rect 45652 384328 45704 384334
rect 45652 384270 45704 384276
rect 45848 373994 45876 394742
rect 45756 373966 45876 373994
rect 45572 344986 45692 345014
rect 45664 332586 45692 344986
rect 45652 332580 45704 332586
rect 45652 332522 45704 332528
rect 45756 330562 45784 373966
rect 45926 345400 45982 345409
rect 45926 345335 45982 345344
rect 45940 345166 45968 345335
rect 45928 345160 45980 345166
rect 45928 345102 45980 345108
rect 45664 330534 45784 330562
rect 45468 259480 45520 259486
rect 45468 259422 45520 259428
rect 45480 253858 45508 259422
rect 45480 253830 45600 253858
rect 45572 247466 45600 253830
rect 45480 247438 45600 247466
rect 45376 247308 45428 247314
rect 45376 247250 45428 247256
rect 45480 238754 45508 247438
rect 45664 239426 45692 330534
rect 45834 328808 45890 328817
rect 45834 328743 45890 328752
rect 45848 328506 45876 328743
rect 45836 328500 45888 328506
rect 45836 328442 45888 328448
rect 45744 325712 45796 325718
rect 45744 325654 45796 325660
rect 45756 255746 45784 325654
rect 45834 264616 45890 264625
rect 45834 264551 45890 264560
rect 45744 255740 45796 255746
rect 45744 255682 45796 255688
rect 45848 247178 45876 264551
rect 45926 256728 45982 256737
rect 45926 256663 45982 256672
rect 45836 247172 45888 247178
rect 45836 247114 45888 247120
rect 45834 242992 45890 243001
rect 45834 242927 45836 242936
rect 45888 242927 45890 242936
rect 45836 242898 45888 242904
rect 45652 239420 45704 239426
rect 45652 239362 45704 239368
rect 45388 238726 45508 238754
rect 45388 236706 45416 238726
rect 45376 236700 45428 236706
rect 45376 236642 45428 236648
rect 45650 234696 45706 234705
rect 45650 234631 45652 234640
rect 45704 234631 45706 234640
rect 45652 234602 45704 234608
rect 45468 231804 45520 231810
rect 45468 231746 45520 231752
rect 45284 230580 45336 230586
rect 45284 230522 45336 230528
rect 45376 227044 45428 227050
rect 45376 226986 45428 226992
rect 45388 214606 45416 226986
rect 45480 226250 45508 231746
rect 45744 230580 45796 230586
rect 45744 230522 45796 230528
rect 45480 226222 45692 226250
rect 45376 214600 45428 214606
rect 45376 214542 45428 214548
rect 45376 213920 45428 213926
rect 45376 213862 45428 213868
rect 45388 197266 45416 213862
rect 45664 205634 45692 226222
rect 45756 213926 45784 230522
rect 45940 217530 45968 256663
rect 46032 220454 46060 509254
rect 46110 506968 46166 506977
rect 46110 506903 46166 506912
rect 46124 506530 46152 506903
rect 46112 506524 46164 506530
rect 46112 506466 46164 506472
rect 46110 505200 46166 505209
rect 46110 505135 46112 505144
rect 46164 505135 46166 505144
rect 46112 505106 46164 505112
rect 46112 501900 46164 501906
rect 46112 501842 46164 501848
rect 46124 501401 46152 501842
rect 46110 501392 46166 501401
rect 46110 501327 46166 501336
rect 46110 496088 46166 496097
rect 46110 496023 46166 496032
rect 46124 495514 46152 496023
rect 46112 495508 46164 495514
rect 46112 495450 46164 495456
rect 46110 400344 46166 400353
rect 46110 400279 46166 400288
rect 46124 400246 46152 400279
rect 46112 400240 46164 400246
rect 46112 400182 46164 400188
rect 46110 373144 46166 373153
rect 46110 373079 46166 373088
rect 46124 372706 46152 373079
rect 46112 372700 46164 372706
rect 46112 372642 46164 372648
rect 46020 220448 46072 220454
rect 46020 220390 46072 220396
rect 46020 220312 46072 220318
rect 46020 220254 46072 220260
rect 45928 217524 45980 217530
rect 45928 217466 45980 217472
rect 46032 217410 46060 220254
rect 46112 218748 46164 218754
rect 46112 218690 46164 218696
rect 45848 217382 46060 217410
rect 45848 214606 45876 217382
rect 45928 217320 45980 217326
rect 45928 217262 45980 217268
rect 46018 217288 46074 217297
rect 45836 214600 45888 214606
rect 45836 214542 45888 214548
rect 45744 213920 45796 213926
rect 45744 213862 45796 213868
rect 45664 205606 45784 205634
rect 45650 203688 45706 203697
rect 45650 203623 45706 203632
rect 45664 202910 45692 203623
rect 45652 202904 45704 202910
rect 45558 202872 45614 202881
rect 45652 202846 45704 202852
rect 45558 202807 45560 202816
rect 45612 202807 45614 202816
rect 45560 202778 45612 202784
rect 45756 201521 45784 205606
rect 45742 201512 45798 201521
rect 45742 201447 45798 201456
rect 45376 197260 45428 197266
rect 45376 197202 45428 197208
rect 45940 195401 45968 217262
rect 46018 217223 46074 217232
rect 46032 216714 46060 217223
rect 46020 216708 46072 216714
rect 46020 216650 46072 216656
rect 45926 195392 45982 195401
rect 45926 195327 45982 195336
rect 45468 192772 45520 192778
rect 45468 192714 45520 192720
rect 45374 181520 45430 181529
rect 45374 181455 45430 181464
rect 45284 151496 45336 151502
rect 45284 151438 45336 151444
rect 45192 29640 45244 29646
rect 45192 29582 45244 29588
rect 45100 22976 45152 22982
rect 45100 22918 45152 22924
rect 44916 19712 44968 19718
rect 44916 19654 44968 19660
rect 45296 19174 45324 151438
rect 45388 22574 45416 181455
rect 45376 22568 45428 22574
rect 45376 22510 45428 22516
rect 45284 19168 45336 19174
rect 45284 19110 45336 19116
rect 45480 17338 45508 192714
rect 46020 183320 46072 183326
rect 46020 183262 46072 183268
rect 45928 156868 45980 156874
rect 45928 156810 45980 156816
rect 45940 18426 45968 156810
rect 46032 56574 46060 183262
rect 46124 153134 46152 218690
rect 46216 204377 46244 518866
rect 46308 489841 46336 549102
rect 46294 489832 46350 489841
rect 46294 489767 46350 489776
rect 46296 480684 46348 480690
rect 46296 480626 46348 480632
rect 46308 438841 46336 480626
rect 46400 480321 46428 563654
rect 46492 498302 46520 578954
rect 46664 573572 46716 573578
rect 46664 573514 46716 573520
rect 46572 560176 46624 560182
rect 46572 560118 46624 560124
rect 46480 498296 46532 498302
rect 46480 498238 46532 498244
rect 46480 498160 46532 498166
rect 46480 498102 46532 498108
rect 46492 497321 46520 498102
rect 46478 497312 46534 497321
rect 46478 497247 46534 497256
rect 46480 496800 46532 496806
rect 46480 496742 46532 496748
rect 46492 495961 46520 496742
rect 46478 495952 46534 495961
rect 46478 495887 46534 495896
rect 46480 495440 46532 495446
rect 46480 495382 46532 495388
rect 46492 495281 46520 495382
rect 46478 495272 46534 495281
rect 46478 495207 46534 495216
rect 46478 493232 46534 493241
rect 46478 493167 46534 493176
rect 46492 492726 46520 493167
rect 46480 492720 46532 492726
rect 46480 492662 46532 492668
rect 46478 489968 46534 489977
rect 46478 489903 46480 489912
rect 46532 489903 46534 489912
rect 46480 489874 46532 489880
rect 46480 486124 46532 486130
rect 46480 486066 46532 486072
rect 46492 482361 46520 486066
rect 46478 482352 46534 482361
rect 46478 482287 46534 482296
rect 46480 481364 46532 481370
rect 46480 481306 46532 481312
rect 46386 480312 46442 480321
rect 46386 480247 46442 480256
rect 46492 460934 46520 481306
rect 46584 474201 46612 560118
rect 46676 475561 46704 573514
rect 46768 486130 46796 581674
rect 47032 566568 47084 566574
rect 47032 566510 47084 566516
rect 46848 560244 46900 560250
rect 46848 560186 46900 560192
rect 46756 486124 46808 486130
rect 46756 486066 46808 486072
rect 46754 485888 46810 485897
rect 46754 485823 46756 485832
rect 46808 485823 46810 485832
rect 46756 485794 46808 485800
rect 46754 485208 46810 485217
rect 46754 485143 46810 485152
rect 46768 484498 46796 485143
rect 46756 484492 46808 484498
rect 46756 484434 46808 484440
rect 46754 480584 46810 480593
rect 46754 480519 46810 480528
rect 46768 480282 46796 480519
rect 46756 480276 46808 480282
rect 46756 480218 46808 480224
rect 46662 475552 46718 475561
rect 46662 475487 46718 475496
rect 46756 474700 46808 474706
rect 46756 474642 46808 474648
rect 46570 474192 46626 474201
rect 46570 474127 46626 474136
rect 46768 473521 46796 474642
rect 46754 473512 46810 473521
rect 46754 473447 46810 473456
rect 46754 469704 46810 469713
rect 46754 469639 46810 469648
rect 46768 469266 46796 469639
rect 46756 469260 46808 469266
rect 46756 469202 46808 469208
rect 46662 468344 46718 468353
rect 46662 468279 46718 468288
rect 46676 467906 46704 468279
rect 46754 468072 46810 468081
rect 46754 468007 46810 468016
rect 46768 467974 46796 468007
rect 46756 467968 46808 467974
rect 46756 467910 46808 467916
rect 46664 467900 46716 467906
rect 46664 467842 46716 467848
rect 46754 464264 46810 464273
rect 46754 464199 46810 464208
rect 46768 464166 46796 464199
rect 46756 464160 46808 464166
rect 46756 464102 46808 464108
rect 46754 463856 46810 463865
rect 46754 463791 46810 463800
rect 46768 463758 46796 463791
rect 46756 463752 46808 463758
rect 46756 463694 46808 463700
rect 46664 463684 46716 463690
rect 46664 463626 46716 463632
rect 46676 463321 46704 463626
rect 46662 463312 46718 463321
rect 46662 463247 46718 463256
rect 46754 461000 46810 461009
rect 46754 460935 46756 460944
rect 46492 460906 46612 460934
rect 46808 460935 46810 460944
rect 46756 460906 46808 460912
rect 46478 446040 46534 446049
rect 46478 445975 46534 445984
rect 46492 445806 46520 445975
rect 46480 445800 46532 445806
rect 46480 445742 46532 445748
rect 46584 442921 46612 460906
rect 46664 460896 46716 460902
rect 46664 460838 46716 460844
rect 46676 459921 46704 460838
rect 46662 459912 46718 459921
rect 46662 459847 46718 459856
rect 46664 456748 46716 456754
rect 46664 456690 46716 456696
rect 46676 455841 46704 456690
rect 46756 456680 46808 456686
rect 46756 456622 46808 456628
rect 46768 456521 46796 456622
rect 46754 456512 46810 456521
rect 46754 456447 46810 456456
rect 46662 455832 46718 455841
rect 46662 455767 46718 455776
rect 46756 451240 46808 451246
rect 46756 451182 46808 451188
rect 46768 450401 46796 451182
rect 46754 450392 46810 450401
rect 46754 450327 46810 450336
rect 46754 443320 46810 443329
rect 46754 443255 46810 443264
rect 46768 443018 46796 443255
rect 46756 443012 46808 443018
rect 46756 442954 46808 442960
rect 46570 442912 46626 442921
rect 46570 442847 46626 442856
rect 46294 438832 46350 438841
rect 46294 438767 46350 438776
rect 46754 436520 46810 436529
rect 46754 436455 46810 436464
rect 46768 436150 46796 436455
rect 46756 436144 46808 436150
rect 46756 436086 46808 436092
rect 46756 434784 46808 434790
rect 46754 434752 46756 434761
rect 46808 434752 46810 434761
rect 46754 434687 46810 434696
rect 46754 433664 46810 433673
rect 46754 433599 46810 433608
rect 46768 433362 46796 433599
rect 46756 433356 46808 433362
rect 46756 433298 46808 433304
rect 46386 432032 46442 432041
rect 46386 431967 46388 431976
rect 46440 431967 46442 431976
rect 46388 431938 46440 431944
rect 46388 430568 46440 430574
rect 46388 430510 46440 430516
rect 46400 430001 46428 430510
rect 46386 429992 46442 430001
rect 46386 429927 46442 429936
rect 46754 429312 46810 429321
rect 46754 429247 46810 429256
rect 46768 429214 46796 429247
rect 46756 429208 46808 429214
rect 46756 429150 46808 429156
rect 46754 427952 46810 427961
rect 46754 427887 46810 427896
rect 46768 427854 46796 427887
rect 46756 427848 46808 427854
rect 46756 427790 46808 427796
rect 46570 425368 46626 425377
rect 46570 425303 46626 425312
rect 46478 421288 46534 421297
rect 46478 421223 46534 421232
rect 46492 412634 46520 421223
rect 46584 413930 46612 425303
rect 46754 425232 46810 425241
rect 46754 425167 46810 425176
rect 46768 425134 46796 425167
rect 46756 425128 46808 425134
rect 46756 425070 46808 425076
rect 46664 425060 46716 425066
rect 46664 425002 46716 425008
rect 46676 424561 46704 425002
rect 46662 424552 46718 424561
rect 46662 424487 46718 424496
rect 46754 423736 46810 423745
rect 46754 423671 46756 423680
rect 46808 423671 46810 423680
rect 46756 423642 46808 423648
rect 46754 421016 46810 421025
rect 46754 420951 46756 420960
rect 46808 420951 46810 420960
rect 46756 420922 46808 420928
rect 46662 420064 46718 420073
rect 46662 419999 46718 420008
rect 46676 419626 46704 419999
rect 46754 419656 46810 419665
rect 46664 419620 46716 419626
rect 46754 419591 46810 419600
rect 46664 419562 46716 419568
rect 46768 419558 46796 419591
rect 46756 419552 46808 419558
rect 46756 419494 46808 419500
rect 46662 418704 46718 418713
rect 46662 418639 46718 418648
rect 46676 418266 46704 418639
rect 46754 418296 46810 418305
rect 46664 418260 46716 418266
rect 46754 418231 46810 418240
rect 46664 418202 46716 418208
rect 46768 418198 46796 418231
rect 46756 418192 46808 418198
rect 46756 418134 46808 418140
rect 46662 415984 46718 415993
rect 46662 415919 46718 415928
rect 46676 415478 46704 415919
rect 46754 415576 46810 415585
rect 46754 415511 46756 415520
rect 46808 415511 46810 415520
rect 46756 415482 46808 415488
rect 46664 415472 46716 415478
rect 46664 415414 46716 415420
rect 46754 414080 46810 414089
rect 46754 414015 46756 414024
rect 46808 414015 46810 414024
rect 46756 413986 46808 413992
rect 46584 413902 46796 413930
rect 46492 412606 46704 412634
rect 46570 411360 46626 411369
rect 46570 411295 46572 411304
rect 46624 411295 46626 411304
rect 46572 411266 46624 411272
rect 46570 407688 46626 407697
rect 46570 407623 46626 407632
rect 46584 407182 46612 407623
rect 46572 407176 46624 407182
rect 46572 407118 46624 407124
rect 46570 399528 46626 399537
rect 46570 399463 46626 399472
rect 46584 398886 46612 399463
rect 46572 398880 46624 398886
rect 46572 398822 46624 398828
rect 46478 396672 46534 396681
rect 46478 396607 46534 396616
rect 46492 396506 46520 396607
rect 46480 396500 46532 396506
rect 46480 396442 46532 396448
rect 46570 395040 46626 395049
rect 46570 394975 46626 394984
rect 46584 394738 46612 394975
rect 46572 394732 46624 394738
rect 46572 394674 46624 394680
rect 46570 393680 46626 393689
rect 46570 393615 46626 393624
rect 46584 393378 46612 393615
rect 46572 393372 46624 393378
rect 46572 393314 46624 393320
rect 46478 392728 46534 392737
rect 46478 392663 46534 392672
rect 46492 392018 46520 392663
rect 46570 392184 46626 392193
rect 46570 392119 46626 392128
rect 46584 392086 46612 392119
rect 46572 392080 46624 392086
rect 46572 392022 46624 392028
rect 46480 392012 46532 392018
rect 46480 391954 46532 391960
rect 46478 390960 46534 390969
rect 46478 390895 46534 390904
rect 46492 390590 46520 390895
rect 46480 390584 46532 390590
rect 46480 390526 46532 390532
rect 46570 390552 46626 390561
rect 46570 390487 46572 390496
rect 46624 390487 46626 390496
rect 46572 390458 46624 390464
rect 46570 389600 46626 389609
rect 46570 389535 46626 389544
rect 46584 389230 46612 389535
rect 46572 389224 46624 389230
rect 46572 389166 46624 389172
rect 46570 386472 46626 386481
rect 46570 386407 46572 386416
rect 46624 386407 46626 386416
rect 46572 386378 46624 386384
rect 46480 386368 46532 386374
rect 46480 386310 46532 386316
rect 46492 385801 46520 386310
rect 46478 385792 46534 385801
rect 46478 385727 46534 385736
rect 46570 385112 46626 385121
rect 46570 385047 46572 385056
rect 46624 385047 46626 385056
rect 46572 385018 46624 385024
rect 46570 382392 46626 382401
rect 46570 382327 46626 382336
rect 46584 382294 46612 382327
rect 46572 382288 46624 382294
rect 46572 382230 46624 382236
rect 46478 381032 46534 381041
rect 46478 380967 46534 380976
rect 46492 377482 46520 380967
rect 46570 379944 46626 379953
rect 46570 379879 46626 379888
rect 46584 379574 46612 379879
rect 46572 379568 46624 379574
rect 46572 379510 46624 379516
rect 46570 378312 46626 378321
rect 46570 378247 46626 378256
rect 46584 378214 46612 378247
rect 46572 378208 46624 378214
rect 46572 378150 46624 378156
rect 46492 377454 46612 377482
rect 46478 374096 46534 374105
rect 46478 374031 46480 374040
rect 46532 374031 46534 374040
rect 46480 374002 46532 374008
rect 46478 372736 46534 372745
rect 46478 372671 46534 372680
rect 46492 372638 46520 372671
rect 46480 372632 46532 372638
rect 46480 372574 46532 372580
rect 46478 371512 46534 371521
rect 46478 371447 46534 371456
rect 46492 371278 46520 371447
rect 46480 371272 46532 371278
rect 46480 371214 46532 371220
rect 46478 369064 46534 369073
rect 46478 368999 46534 369008
rect 46492 368558 46520 368999
rect 46480 368552 46532 368558
rect 46480 368494 46532 368500
rect 46386 367704 46442 367713
rect 46386 367639 46442 367648
rect 46400 367130 46428 367639
rect 46388 367124 46440 367130
rect 46388 367066 46440 367072
rect 46480 367056 46532 367062
rect 46480 366998 46532 367004
rect 46492 366081 46520 366998
rect 46478 366072 46534 366081
rect 46478 366007 46534 366016
rect 46478 363488 46534 363497
rect 46478 363423 46534 363432
rect 46492 362982 46520 363423
rect 46480 362976 46532 362982
rect 46480 362918 46532 362924
rect 46480 358760 46532 358766
rect 46480 358702 46532 358708
rect 46492 357921 46520 358702
rect 46478 357912 46534 357921
rect 46478 357847 46534 357856
rect 46478 354784 46534 354793
rect 46478 354719 46480 354728
rect 46532 354719 46534 354728
rect 46480 354690 46532 354696
rect 46480 353252 46532 353258
rect 46480 353194 46532 353200
rect 46492 353161 46520 353194
rect 46478 353152 46534 353161
rect 46478 353087 46534 353096
rect 46478 349480 46534 349489
rect 46478 349415 46534 349424
rect 46492 349178 46520 349415
rect 46480 349172 46532 349178
rect 46480 349114 46532 349120
rect 46478 347168 46534 347177
rect 46478 347103 46534 347112
rect 46492 346458 46520 347103
rect 46480 346452 46532 346458
rect 46480 346394 46532 346400
rect 46296 342236 46348 342242
rect 46296 342178 46348 342184
rect 46308 263634 46336 342178
rect 46478 336832 46534 336841
rect 46478 336767 46480 336776
rect 46532 336767 46534 336776
rect 46480 336738 46532 336744
rect 46386 329896 46442 329905
rect 46386 329831 46442 329840
rect 46400 313138 46428 329831
rect 46388 313132 46440 313138
rect 46388 313074 46440 313080
rect 46478 302968 46534 302977
rect 46478 302903 46534 302912
rect 46492 302258 46520 302903
rect 46480 302252 46532 302258
rect 46480 302194 46532 302200
rect 46480 293956 46532 293962
rect 46480 293898 46532 293904
rect 46492 292641 46520 293898
rect 46478 292632 46534 292641
rect 46478 292567 46534 292576
rect 46478 284336 46534 284345
rect 46478 284271 46534 284280
rect 46296 263628 46348 263634
rect 46296 263570 46348 263576
rect 46388 254380 46440 254386
rect 46388 254322 46440 254328
rect 46400 252521 46428 254322
rect 46386 252512 46442 252521
rect 46386 252447 46442 252456
rect 46296 249076 46348 249082
rect 46296 249018 46348 249024
rect 46202 204368 46258 204377
rect 46202 204303 46258 204312
rect 46202 201648 46258 201657
rect 46202 201583 46258 201592
rect 46112 153128 46164 153134
rect 46112 153070 46164 153076
rect 46112 151224 46164 151230
rect 46112 151166 46164 151172
rect 46020 56568 46072 56574
rect 46020 56510 46072 56516
rect 46124 18562 46152 151166
rect 46216 20330 46244 201583
rect 46308 21758 46336 249018
rect 46386 245440 46442 245449
rect 46386 245375 46442 245384
rect 46400 222193 46428 245375
rect 46386 222184 46442 222193
rect 46386 222119 46442 222128
rect 46388 215416 46440 215422
rect 46388 215358 46440 215364
rect 46400 202366 46428 215358
rect 46388 202360 46440 202366
rect 46388 202302 46440 202308
rect 46386 188864 46442 188873
rect 46386 188799 46442 188808
rect 46400 155961 46428 188799
rect 46492 156777 46520 284271
rect 46584 254386 46612 377454
rect 46572 254380 46624 254386
rect 46572 254322 46624 254328
rect 46570 254280 46626 254289
rect 46570 254215 46626 254224
rect 46584 253978 46612 254215
rect 46572 253972 46624 253978
rect 46572 253914 46624 253920
rect 46572 247308 46624 247314
rect 46572 247250 46624 247256
rect 46584 226681 46612 247250
rect 46676 244361 46704 412606
rect 46768 247625 46796 413902
rect 46860 331378 46888 560186
rect 46860 331350 46980 331378
rect 46848 331220 46900 331226
rect 46848 331162 46900 331168
rect 46860 330721 46888 331162
rect 46846 330712 46902 330721
rect 46846 330647 46902 330656
rect 46952 330562 46980 331350
rect 46860 330534 46980 330562
rect 46860 328001 46888 330534
rect 46846 327992 46902 328001
rect 46846 327927 46902 327936
rect 46848 325644 46900 325650
rect 46848 325586 46900 325592
rect 46860 325281 46888 325586
rect 46846 325272 46902 325281
rect 46846 325207 46902 325216
rect 46846 323096 46902 323105
rect 46846 323031 46902 323040
rect 46860 322998 46888 323031
rect 46848 322992 46900 322998
rect 46848 322934 46900 322940
rect 46846 321736 46902 321745
rect 46846 321671 46902 321680
rect 46860 321638 46888 321671
rect 46848 321632 46900 321638
rect 46848 321574 46900 321580
rect 46846 320240 46902 320249
rect 46846 320175 46848 320184
rect 46900 320175 46902 320184
rect 46848 320146 46900 320152
rect 46846 319016 46902 319025
rect 46846 318951 46848 318960
rect 46900 318951 46902 318960
rect 46848 318922 46900 318928
rect 46848 318640 46900 318646
rect 46848 318582 46900 318588
rect 46860 318481 46888 318582
rect 46846 318472 46902 318481
rect 46846 318407 46902 318416
rect 46846 314800 46902 314809
rect 46846 314735 46902 314744
rect 46860 314702 46888 314735
rect 46848 314696 46900 314702
rect 46848 314638 46900 314644
rect 46846 310992 46902 311001
rect 46846 310927 46902 310936
rect 46860 310554 46888 310927
rect 46848 310548 46900 310554
rect 46848 310490 46900 310496
rect 46846 309224 46902 309233
rect 46846 309159 46848 309168
rect 46900 309159 46902 309168
rect 46848 309130 46900 309136
rect 46846 303784 46902 303793
rect 46846 303719 46902 303728
rect 46860 303686 46888 303719
rect 46848 303680 46900 303686
rect 46848 303622 46900 303628
rect 46848 302184 46900 302190
rect 46846 302152 46848 302161
rect 46900 302152 46902 302161
rect 46846 302087 46902 302096
rect 46846 300928 46902 300937
rect 46846 300863 46848 300872
rect 46900 300863 46902 300872
rect 46848 300834 46900 300840
rect 46846 298208 46902 298217
rect 46846 298143 46848 298152
rect 46900 298143 46902 298152
rect 46848 298114 46900 298120
rect 46846 296848 46902 296857
rect 46846 296783 46902 296792
rect 46860 296750 46888 296783
rect 46848 296744 46900 296750
rect 46848 296686 46900 296692
rect 46846 292904 46902 292913
rect 46846 292839 46902 292848
rect 46860 292602 46888 292839
rect 46848 292596 46900 292602
rect 46848 292538 46900 292544
rect 46846 291544 46902 291553
rect 46846 291479 46902 291488
rect 46860 291242 46888 291479
rect 46848 291236 46900 291242
rect 46848 291178 46900 291184
rect 46846 288552 46902 288561
rect 46846 288487 46902 288496
rect 46860 288454 46888 288487
rect 46848 288448 46900 288454
rect 46848 288390 46900 288396
rect 46846 285832 46902 285841
rect 46846 285767 46902 285776
rect 46860 285734 46888 285767
rect 46848 285728 46900 285734
rect 46848 285670 46900 285676
rect 46938 285288 46994 285297
rect 46938 285223 46994 285232
rect 46846 281616 46902 281625
rect 46846 281551 46848 281560
rect 46900 281551 46902 281560
rect 46848 281522 46900 281528
rect 46846 277808 46902 277817
rect 46846 277743 46902 277752
rect 46860 277438 46888 277743
rect 46848 277432 46900 277438
rect 46848 277374 46900 277380
rect 46952 274922 46980 285223
rect 46940 274916 46992 274922
rect 46940 274858 46992 274864
rect 46846 268288 46902 268297
rect 46846 268223 46902 268232
rect 46860 267850 46888 268223
rect 46848 267844 46900 267850
rect 46848 267786 46900 267792
rect 46940 263628 46992 263634
rect 46940 263570 46992 263576
rect 46952 259486 46980 263570
rect 46940 259480 46992 259486
rect 46940 259422 46992 259428
rect 46754 247616 46810 247625
rect 46754 247551 46810 247560
rect 46754 247480 46810 247489
rect 46754 247415 46810 247424
rect 46768 247110 46796 247415
rect 46756 247104 46808 247110
rect 46756 247046 46808 247052
rect 46754 245848 46810 245857
rect 46754 245783 46810 245792
rect 46662 244352 46718 244361
rect 46662 244287 46718 244296
rect 46664 233232 46716 233238
rect 46664 233174 46716 233180
rect 46570 226672 46626 226681
rect 46570 226607 46626 226616
rect 46676 225554 46704 233174
rect 46664 225548 46716 225554
rect 46664 225490 46716 225496
rect 46662 221368 46718 221377
rect 46662 221303 46718 221312
rect 46570 218648 46626 218657
rect 46570 218583 46626 218592
rect 46584 218142 46612 218583
rect 46572 218136 46624 218142
rect 46572 218078 46624 218084
rect 46572 213172 46624 213178
rect 46572 213114 46624 213120
rect 46584 198558 46612 213114
rect 46676 199986 46704 221303
rect 46664 199980 46716 199986
rect 46664 199922 46716 199928
rect 46572 198552 46624 198558
rect 46572 198494 46624 198500
rect 46768 195294 46796 245783
rect 46848 238740 46900 238746
rect 46848 238682 46900 238688
rect 46860 238241 46888 238682
rect 46846 238232 46902 238241
rect 46846 238167 46902 238176
rect 46846 237552 46902 237561
rect 46846 237487 46902 237496
rect 46860 237454 46888 237487
rect 46848 237448 46900 237454
rect 46848 237390 46900 237396
rect 46940 236700 46992 236706
rect 46940 236642 46992 236648
rect 46846 236056 46902 236065
rect 46846 235991 46902 236000
rect 46860 232626 46888 235991
rect 46848 232620 46900 232626
rect 46848 232562 46900 232568
rect 46846 232384 46902 232393
rect 46846 232319 46902 232328
rect 46860 231878 46888 232319
rect 46848 231872 46900 231878
rect 46848 231814 46900 231820
rect 46846 230616 46902 230625
rect 46846 230551 46902 230560
rect 46860 230518 46888 230551
rect 46848 230512 46900 230518
rect 46848 230454 46900 230460
rect 46846 227896 46902 227905
rect 46846 227831 46902 227840
rect 46860 227798 46888 227831
rect 46848 227792 46900 227798
rect 46848 227734 46900 227740
rect 46952 227050 46980 236642
rect 47044 233481 47072 566510
rect 47124 561604 47176 561610
rect 47124 561546 47176 561552
rect 47136 270201 47164 561546
rect 47228 376281 47256 585958
rect 47400 562352 47452 562358
rect 47400 562294 47452 562300
rect 47308 561400 47360 561406
rect 47308 561342 47360 561348
rect 47214 376272 47270 376281
rect 47214 376207 47270 376216
rect 47216 374740 47268 374746
rect 47216 374682 47268 374688
rect 47228 348430 47256 374682
rect 47216 348424 47268 348430
rect 47216 348366 47268 348372
rect 47214 335472 47270 335481
rect 47214 335407 47270 335416
rect 47122 270192 47178 270201
rect 47122 270127 47178 270136
rect 47124 242208 47176 242214
rect 47124 242150 47176 242156
rect 47030 233472 47086 233481
rect 47030 233407 47086 233416
rect 47136 233238 47164 242150
rect 47124 233232 47176 233238
rect 47124 233174 47176 233180
rect 47030 230888 47086 230897
rect 47030 230823 47086 230832
rect 46940 227044 46992 227050
rect 46940 226986 46992 226992
rect 46846 224088 46902 224097
rect 46846 224023 46902 224032
rect 46860 223650 46888 224023
rect 46848 223644 46900 223650
rect 46848 223586 46900 223592
rect 46846 222456 46902 222465
rect 46846 222391 46902 222400
rect 46860 222222 46888 222391
rect 46848 222216 46900 222222
rect 46848 222158 46900 222164
rect 46846 221096 46902 221105
rect 46846 221031 46902 221040
rect 46860 220862 46888 221031
rect 46848 220856 46900 220862
rect 46848 220798 46900 220804
rect 46846 218104 46902 218113
rect 46846 218039 46848 218048
rect 46900 218039 46902 218048
rect 46848 218010 46900 218016
rect 46846 215384 46902 215393
rect 46846 215319 46848 215328
rect 46900 215319 46902 215328
rect 46848 215290 46900 215296
rect 46846 214024 46902 214033
rect 46846 213959 46848 213968
rect 46900 213959 46902 213968
rect 46848 213930 46900 213936
rect 46846 211304 46902 211313
rect 46846 211239 46902 211248
rect 46860 211206 46888 211239
rect 46848 211200 46900 211206
rect 46848 211142 46900 211148
rect 46848 208344 46900 208350
rect 46848 208286 46900 208292
rect 46860 207641 46888 208286
rect 46846 207632 46902 207641
rect 46846 207567 46902 207576
rect 46848 206984 46900 206990
rect 46846 206952 46848 206961
rect 46900 206952 46902 206961
rect 46846 206887 46902 206896
rect 46846 205728 46902 205737
rect 46846 205663 46848 205672
rect 46900 205663 46902 205672
rect 46848 205634 46900 205640
rect 46848 204332 46900 204338
rect 46848 204274 46900 204280
rect 46756 195288 46808 195294
rect 46756 195230 46808 195236
rect 46860 192370 46888 204274
rect 47044 199510 47072 230823
rect 47124 227860 47176 227866
rect 47124 227802 47176 227808
rect 47136 215422 47164 227802
rect 47124 215416 47176 215422
rect 47124 215358 47176 215364
rect 47124 214600 47176 214606
rect 47124 214542 47176 214548
rect 47136 204338 47164 214542
rect 47124 204332 47176 204338
rect 47124 204274 47176 204280
rect 47032 199504 47084 199510
rect 47032 199446 47084 199452
rect 46848 192364 46900 192370
rect 46848 192306 46900 192312
rect 46848 191208 46900 191214
rect 46848 191150 46900 191156
rect 46662 178800 46718 178809
rect 46662 178735 46718 178744
rect 46572 169380 46624 169386
rect 46572 169322 46624 169328
rect 46478 156768 46534 156777
rect 46478 156703 46534 156712
rect 46386 155952 46442 155961
rect 46386 155887 46442 155896
rect 46388 155304 46440 155310
rect 46388 155246 46440 155252
rect 46296 21752 46348 21758
rect 46296 21694 46348 21700
rect 46400 21214 46428 155246
rect 46584 21486 46612 169322
rect 46676 23390 46704 178735
rect 46756 174888 46808 174894
rect 46756 174830 46808 174836
rect 46664 23384 46716 23390
rect 46664 23326 46716 23332
rect 46572 21480 46624 21486
rect 46572 21422 46624 21428
rect 46388 21208 46440 21214
rect 46388 21150 46440 21156
rect 46204 20324 46256 20330
rect 46204 20266 46256 20272
rect 46112 18556 46164 18562
rect 46112 18498 46164 18504
rect 45928 18420 45980 18426
rect 45928 18362 45980 18368
rect 45468 17332 45520 17338
rect 45468 17274 45520 17280
rect 46662 11656 46718 11665
rect 46662 11591 46718 11600
rect 42248 3800 42300 3806
rect 42248 3742 42300 3748
rect 39764 3528 39816 3534
rect 39764 3470 39816 3476
rect 43074 3496 43130 3505
rect 43074 3431 43130 3440
rect 43088 480 43116 3431
rect 46676 480 46704 11591
rect 46768 4010 46796 174830
rect 46860 18358 46888 191150
rect 47228 49026 47256 335407
rect 47320 298081 47348 561342
rect 47412 504121 47440 562294
rect 47492 560924 47544 560930
rect 47492 560866 47544 560872
rect 47504 521801 47532 560866
rect 47490 521792 47546 521801
rect 47490 521727 47546 521736
rect 47398 504112 47454 504121
rect 47398 504047 47454 504056
rect 47306 298072 47362 298081
rect 47306 298007 47362 298016
rect 47398 281888 47454 281897
rect 47398 281823 47454 281832
rect 47306 273320 47362 273329
rect 47306 273255 47362 273264
rect 47216 49020 47268 49026
rect 47216 48962 47268 48968
rect 47320 29374 47348 273255
rect 47412 132462 47440 281823
rect 47490 259584 47546 259593
rect 47490 259519 47546 259528
rect 47504 241505 47532 259519
rect 47490 241496 47546 241505
rect 47490 241431 47546 241440
rect 47490 216744 47546 216753
rect 47490 216679 47546 216688
rect 47400 132456 47452 132462
rect 47400 132398 47452 132404
rect 47308 29368 47360 29374
rect 47308 29310 47360 29316
rect 47504 28966 47532 216679
rect 47596 213178 47624 589222
rect 78864 589076 78916 589082
rect 78864 589018 78916 589024
rect 52458 587888 52514 587897
rect 52458 587823 52514 587832
rect 53838 587888 53894 587897
rect 53838 587823 53894 587832
rect 56598 587888 56654 587897
rect 56598 587823 56654 587832
rect 57886 587888 57942 587897
rect 57886 587823 57942 587832
rect 58070 587888 58126 587897
rect 58070 587823 58126 587832
rect 59358 587888 59414 587897
rect 59358 587823 59414 587832
rect 62118 587888 62174 587897
rect 62118 587823 62174 587832
rect 63498 587888 63554 587897
rect 63498 587823 63554 587832
rect 63682 587888 63738 587897
rect 63682 587823 63738 587832
rect 64970 587888 65026 587897
rect 64970 587823 65026 587832
rect 66350 587888 66406 587897
rect 66350 587823 66406 587832
rect 67638 587888 67694 587897
rect 67638 587823 67694 587832
rect 69018 587888 69074 587897
rect 69018 587823 69074 587832
rect 70398 587888 70454 587897
rect 70398 587823 70454 587832
rect 71778 587888 71834 587897
rect 71778 587823 71834 587832
rect 72422 587888 72478 587897
rect 72422 587823 72478 587832
rect 74630 587888 74686 587897
rect 74630 587823 74686 587832
rect 77298 587888 77354 587897
rect 77298 587823 77354 587832
rect 78678 587888 78734 587897
rect 78678 587823 78734 587832
rect 49056 587376 49108 587382
rect 49056 587318 49108 587324
rect 48964 586628 49016 586634
rect 48964 586570 49016 586576
rect 47768 570716 47820 570722
rect 47768 570658 47820 570664
rect 47676 232620 47728 232626
rect 47676 232562 47728 232568
rect 47584 213172 47636 213178
rect 47584 213114 47636 213120
rect 47584 211812 47636 211818
rect 47584 211754 47636 211760
rect 47596 156942 47624 211754
rect 47584 156936 47636 156942
rect 47584 156878 47636 156884
rect 47688 82754 47716 232562
rect 47780 229401 47808 570658
rect 48976 567194 49004 586570
rect 48884 567166 49004 567194
rect 48228 563032 48280 563038
rect 48228 562974 48280 562980
rect 48240 559994 48268 562974
rect 48884 560182 48912 567166
rect 48962 561776 49018 561785
rect 48962 561711 49018 561720
rect 48872 560176 48924 560182
rect 48872 560118 48924 560124
rect 48070 559966 48268 559994
rect 48976 559994 49004 561711
rect 49068 560250 49096 587318
rect 49148 576224 49200 576230
rect 49148 576166 49200 576172
rect 49160 563038 49188 576166
rect 49148 563032 49200 563038
rect 49148 562974 49200 562980
rect 51540 562080 51592 562086
rect 51540 562022 51592 562028
rect 51632 562080 51684 562086
rect 51632 562022 51684 562028
rect 51080 561876 51132 561882
rect 51080 561818 51132 561824
rect 50252 561740 50304 561746
rect 50252 561682 50304 561688
rect 49606 560280 49662 560289
rect 49056 560244 49108 560250
rect 49606 560215 49608 560224
rect 49056 560186 49108 560192
rect 49660 560215 49662 560224
rect 49608 560186 49660 560192
rect 50264 559994 50292 561682
rect 51092 560017 51120 561818
rect 51078 560008 51134 560017
rect 48976 559966 49358 559994
rect 50264 559966 50600 559994
rect 51552 559994 51580 562022
rect 51644 560153 51672 562022
rect 52472 561542 52500 587823
rect 53852 577522 53880 587823
rect 56506 587752 56562 587761
rect 56506 587687 56562 587696
rect 56520 578921 56548 587687
rect 56506 578912 56562 578921
rect 56506 578847 56562 578856
rect 53840 577516 53892 577522
rect 53840 577458 53892 577464
rect 52644 573368 52696 573374
rect 52644 573310 52696 573316
rect 52460 561536 52512 561542
rect 52460 561478 52512 561484
rect 51630 560144 51686 560153
rect 51630 560079 51686 560088
rect 52656 559994 52684 573310
rect 56612 563990 56640 587823
rect 57900 587450 57928 587823
rect 57888 587444 57940 587450
rect 57888 587386 57940 587392
rect 56600 563984 56652 563990
rect 56600 563926 56652 563932
rect 57426 562184 57482 562193
rect 57426 562119 57482 562128
rect 51552 559966 51934 559994
rect 52578 559966 52684 559994
rect 57440 559994 57468 562119
rect 57978 562048 58034 562057
rect 57978 561983 58034 561992
rect 57992 559994 58020 561983
rect 58084 560969 58112 587823
rect 59174 562184 59230 562193
rect 59174 562119 59230 562128
rect 58070 560960 58126 560969
rect 58070 560895 58126 560904
rect 59188 560250 59216 562119
rect 59266 562048 59322 562057
rect 59266 561983 59322 561992
rect 59280 561241 59308 561983
rect 59372 561270 59400 587823
rect 62026 587752 62082 587761
rect 62026 587687 62082 587696
rect 62040 574870 62068 587687
rect 62028 574864 62080 574870
rect 62028 574806 62080 574812
rect 59818 564496 59874 564505
rect 59818 564431 59874 564440
rect 59360 561264 59412 561270
rect 59266 561232 59322 561241
rect 59360 561206 59412 561212
rect 59266 561167 59322 561176
rect 59176 560244 59228 560250
rect 59176 560186 59228 560192
rect 59832 559994 59860 564431
rect 59910 561912 59966 561921
rect 59910 561847 59966 561856
rect 57440 559966 57730 559994
rect 57992 559966 58374 559994
rect 59662 559966 59860 559994
rect 59924 559994 59952 561847
rect 62132 560930 62160 587823
rect 63512 561134 63540 587823
rect 63590 587752 63646 587761
rect 63590 587687 63646 587696
rect 63604 576162 63632 587687
rect 63592 576156 63644 576162
rect 63592 576098 63644 576104
rect 63696 561474 63724 587823
rect 64788 565208 64840 565214
rect 64788 565150 64840 565156
rect 63684 561468 63736 561474
rect 63684 561410 63736 561416
rect 63500 561128 63552 561134
rect 63500 561070 63552 561076
rect 62120 560924 62172 560930
rect 62120 560866 62172 560872
rect 63222 560552 63278 560561
rect 62488 560516 62540 560522
rect 63222 560487 63278 560496
rect 62488 560458 62540 560464
rect 62500 559994 62528 560458
rect 63236 559994 63264 560487
rect 64800 560266 64828 565150
rect 64984 561105 65012 587823
rect 66364 585886 66392 587823
rect 67546 586392 67602 586401
rect 67546 586327 67602 586336
rect 66352 585880 66404 585886
rect 66352 585822 66404 585828
rect 67560 570654 67588 586327
rect 67548 570648 67600 570654
rect 67548 570590 67600 570596
rect 65708 562624 65760 562630
rect 65708 562566 65760 562572
rect 64970 561096 65026 561105
rect 64970 561031 65026 561040
rect 59924 559966 60260 559994
rect 62238 559966 62528 559994
rect 62882 559966 63264 559994
rect 64754 560238 64828 560266
rect 64754 559980 64782 560238
rect 65720 559994 65748 562566
rect 67652 561610 67680 587823
rect 67640 561604 67692 561610
rect 67640 561546 67692 561552
rect 69032 561338 69060 587823
rect 70306 587752 70362 587761
rect 70306 587687 70362 587696
rect 70320 571985 70348 587687
rect 70306 571976 70362 571985
rect 70306 571911 70362 571920
rect 69020 561332 69072 561338
rect 69020 561274 69072 561280
rect 70412 561202 70440 587823
rect 71792 587314 71820 587823
rect 71780 587308 71832 587314
rect 71780 587250 71832 587256
rect 72436 581641 72464 587823
rect 73066 587752 73122 587761
rect 73066 587687 73122 587696
rect 74538 587752 74594 587761
rect 74538 587687 74594 587696
rect 72422 581632 72478 581641
rect 72422 581567 72478 581576
rect 73080 562630 73108 587687
rect 74446 587616 74502 587625
rect 74446 587551 74502 587560
rect 74460 577522 74488 587551
rect 74448 577516 74500 577522
rect 74448 577458 74500 577464
rect 73068 562624 73120 562630
rect 73068 562566 73120 562572
rect 74552 562358 74580 587687
rect 74644 563922 74672 587823
rect 77206 587752 77262 587761
rect 77206 587687 77262 587696
rect 77220 586770 77248 587687
rect 77208 586764 77260 586770
rect 77208 586706 77260 586712
rect 77114 586392 77170 586401
rect 77114 586327 77170 586336
rect 77128 565146 77156 586327
rect 77116 565140 77168 565146
rect 77116 565082 77168 565088
rect 74632 563916 74684 563922
rect 74632 563858 74684 563864
rect 75828 562556 75880 562562
rect 75828 562498 75880 562504
rect 74540 562352 74592 562358
rect 74540 562294 74592 562300
rect 70400 561196 70452 561202
rect 70400 561138 70452 561144
rect 75840 559994 75868 562498
rect 76656 562352 76708 562358
rect 76656 562294 76708 562300
rect 76668 559994 76696 562294
rect 77312 561406 77340 587823
rect 78692 587382 78720 587823
rect 78770 587752 78826 587761
rect 78770 587687 78826 587696
rect 78680 587376 78732 587382
rect 78680 587318 78732 587324
rect 77758 568712 77814 568721
rect 77758 568647 77814 568656
rect 77300 561400 77352 561406
rect 77300 561342 77352 561348
rect 77772 559994 77800 568647
rect 78784 565282 78812 587687
rect 78772 565276 78824 565282
rect 78772 565218 78824 565224
rect 78876 560266 78904 589018
rect 79782 587888 79838 587897
rect 79782 587823 79838 587832
rect 81162 587888 81218 587897
rect 81162 587823 81218 587832
rect 81806 587888 81862 587897
rect 81806 587823 81862 587832
rect 82910 587888 82966 587897
rect 82910 587823 82966 587832
rect 79796 584526 79824 587823
rect 81176 586566 81204 587823
rect 81164 586560 81216 586566
rect 81164 586502 81216 586508
rect 81820 585954 81848 587823
rect 81898 587752 81954 587761
rect 81898 587687 81954 587696
rect 81912 587246 81940 587687
rect 82084 587444 82136 587450
rect 82084 587386 82136 587392
rect 81900 587240 81952 587246
rect 81900 587182 81952 587188
rect 81808 585948 81860 585954
rect 81808 585890 81860 585896
rect 79784 584520 79836 584526
rect 79784 584462 79836 584468
rect 82096 566642 82124 587386
rect 82924 576854 82952 587823
rect 84396 583030 84424 589455
rect 140780 589144 140832 589150
rect 140780 589086 140832 589092
rect 86040 589076 86092 589082
rect 86040 589018 86092 589024
rect 85486 586392 85542 586401
rect 85486 586327 85542 586336
rect 84384 583024 84436 583030
rect 84384 582966 84436 582972
rect 82924 576826 83044 576854
rect 82084 566636 82136 566642
rect 82084 566578 82136 566584
rect 82820 565004 82872 565010
rect 82820 564946 82872 564952
rect 82832 562494 82860 564946
rect 81624 562488 81676 562494
rect 81624 562430 81676 562436
rect 82820 562488 82872 562494
rect 82820 562430 82872 562436
rect 78876 560238 78950 560266
rect 65720 559966 66102 559994
rect 75762 559966 75868 559994
rect 76406 559966 76696 559994
rect 77694 559966 77800 559994
rect 78922 559980 78950 560238
rect 81636 559994 81664 562430
rect 83016 561066 83044 576826
rect 85500 573646 85528 586327
rect 86052 576854 86080 589018
rect 87142 587888 87198 587897
rect 87142 587823 87198 587832
rect 88338 587888 88394 587897
rect 88338 587823 88394 587832
rect 91098 587888 91154 587897
rect 91098 587823 91154 587832
rect 93122 587888 93178 587897
rect 93122 587823 93178 587832
rect 93858 587888 93914 587897
rect 93858 587823 93914 587832
rect 95146 587888 95202 587897
rect 95146 587823 95202 587832
rect 99470 587888 99526 587897
rect 99470 587823 99526 587832
rect 101954 587888 102010 587897
rect 101954 587823 102010 587832
rect 106922 587888 106978 587897
rect 106922 587823 106978 587832
rect 109038 587888 109094 587897
rect 109038 587823 109094 587832
rect 111798 587888 111854 587897
rect 111798 587823 111854 587832
rect 115202 587888 115258 587897
rect 115202 587823 115258 587832
rect 118698 587888 118754 587897
rect 118698 587823 118754 587832
rect 124402 587888 124458 587897
rect 124402 587823 124458 587832
rect 128358 587888 128414 587897
rect 128358 587823 128414 587832
rect 131762 587888 131818 587897
rect 131762 587823 131818 587832
rect 133970 587888 134026 587897
rect 133970 587823 134026 587832
rect 136638 587888 136694 587897
rect 136638 587823 136694 587832
rect 139398 587888 139454 587897
rect 139398 587823 139454 587832
rect 86958 587752 87014 587761
rect 86958 587687 87014 587696
rect 86866 586392 86922 586401
rect 86866 586327 86922 586336
rect 86052 576826 86172 576854
rect 85488 573640 85540 573646
rect 85488 573582 85540 573588
rect 85486 567216 85542 567225
rect 85486 567151 85542 567160
rect 83094 563272 83150 563281
rect 83094 563207 83150 563216
rect 83004 561060 83056 561066
rect 83004 561002 83056 561008
rect 83108 559994 83136 563207
rect 83740 562420 83792 562426
rect 83740 562362 83792 562368
rect 81558 559966 81664 559994
rect 82846 559966 83136 559994
rect 83752 559994 83780 562362
rect 85500 559994 85528 567151
rect 86144 559994 86172 576826
rect 86880 572082 86908 586327
rect 86868 572076 86920 572082
rect 86868 572018 86920 572024
rect 86314 562456 86370 562465
rect 86314 562391 86370 562400
rect 83752 559966 84088 559994
rect 85422 559966 85528 559994
rect 86066 559966 86172 559994
rect 86328 559994 86356 562391
rect 86972 560998 87000 587687
rect 87050 586392 87106 586401
rect 87050 586327 87106 586336
rect 87064 563786 87092 586327
rect 87156 583098 87184 587823
rect 87144 583092 87196 583098
rect 87144 583034 87196 583040
rect 87328 581800 87380 581806
rect 87328 581742 87380 581748
rect 87340 576854 87368 581742
rect 87340 576826 87460 576854
rect 87052 563780 87104 563786
rect 87052 563722 87104 563728
rect 86960 560992 87012 560998
rect 86960 560934 87012 560940
rect 87432 559994 87460 576826
rect 88352 563854 88380 587823
rect 89626 586392 89682 586401
rect 89626 586327 89682 586336
rect 91006 586392 91062 586401
rect 91006 586327 91062 586336
rect 89640 576162 89668 586327
rect 89628 576156 89680 576162
rect 89628 576098 89680 576104
rect 91020 565282 91048 586327
rect 91112 572150 91140 587823
rect 92386 586392 92442 586401
rect 92386 586327 92442 586336
rect 92400 576065 92428 586327
rect 93136 583001 93164 587823
rect 93122 582992 93178 583001
rect 93122 582927 93178 582936
rect 92386 576056 92442 576065
rect 92386 575991 92442 576000
rect 91100 572144 91152 572150
rect 91100 572086 91152 572092
rect 93872 565418 93900 587823
rect 93860 565412 93912 565418
rect 93860 565354 93912 565360
rect 91008 565276 91060 565282
rect 91008 565218 91060 565224
rect 88340 563848 88392 563854
rect 88340 563790 88392 563796
rect 95160 563786 95188 587823
rect 95238 587752 95294 587761
rect 95238 587687 95294 587696
rect 95252 587178 95280 587687
rect 95240 587172 95292 587178
rect 95240 587114 95292 587120
rect 97906 586392 97962 586401
rect 97906 586327 97962 586336
rect 97920 573510 97948 586327
rect 99484 580310 99512 587823
rect 101968 587110 101996 587823
rect 101956 587104 102008 587110
rect 101956 587046 102008 587052
rect 106936 587042 106964 587823
rect 106924 587036 106976 587042
rect 106924 586978 106976 586984
rect 104806 586392 104862 586401
rect 104806 586327 104862 586336
rect 100852 585812 100904 585818
rect 100852 585754 100904 585760
rect 99472 580304 99524 580310
rect 99472 580246 99524 580252
rect 100864 576854 100892 585754
rect 100864 576826 100984 576854
rect 97908 573504 97960 573510
rect 97908 573446 97960 573452
rect 95148 563780 95200 563786
rect 95148 563722 95200 563728
rect 91284 562624 91336 562630
rect 91284 562566 91336 562572
rect 90824 562420 90876 562426
rect 90824 562362 90876 562368
rect 89718 562320 89774 562329
rect 89718 562255 89774 562264
rect 86328 559966 86710 559994
rect 87354 559966 87460 559994
rect 89732 559994 89760 562255
rect 90836 559994 90864 562362
rect 91296 559994 91324 562566
rect 94780 562284 94832 562290
rect 94780 562226 94832 562232
rect 89732 559966 89930 559994
rect 90574 559966 90864 559994
rect 91218 559966 91324 559994
rect 94792 559994 94820 562226
rect 99380 562216 99432 562222
rect 99380 562158 99432 562164
rect 99392 559994 99420 562158
rect 100956 559994 100984 576826
rect 104820 566506 104848 586327
rect 109052 581670 109080 587823
rect 109040 581664 109092 581670
rect 109040 581606 109092 581612
rect 111812 577658 111840 587823
rect 115216 584594 115244 587823
rect 117226 586392 117282 586401
rect 117226 586327 117282 586336
rect 115204 584588 115256 584594
rect 115204 584530 115256 584536
rect 111800 577652 111852 577658
rect 111800 577594 111852 577600
rect 107660 577584 107712 577590
rect 107660 577526 107712 577532
rect 106094 567352 106150 567361
rect 106094 567287 106150 567296
rect 104808 566500 104860 566506
rect 104808 566442 104860 566448
rect 104348 564936 104400 564942
rect 104348 564878 104400 564884
rect 94792 559966 95082 559994
rect 99392 559966 99590 559994
rect 100878 559966 100984 559994
rect 104360 559994 104388 564878
rect 105084 562148 105136 562154
rect 105084 562090 105136 562096
rect 105096 559994 105124 562090
rect 106108 559994 106136 567287
rect 104360 559966 104742 559994
rect 105096 559966 105386 559994
rect 106030 559966 106136 559994
rect 107672 559994 107700 577526
rect 117240 569226 117268 586327
rect 117320 575000 117372 575006
rect 117320 574942 117372 574948
rect 117228 569220 117280 569226
rect 117228 569162 117280 569168
rect 116400 567248 116452 567254
rect 116400 567190 116452 567196
rect 109590 565992 109646 566001
rect 109590 565927 109646 565936
rect 109604 559994 109632 565927
rect 111892 564868 111944 564874
rect 111892 564810 111944 564816
rect 110144 561808 110196 561814
rect 110144 561750 110196 561756
rect 110156 559994 110184 561750
rect 111904 559994 111932 564810
rect 113456 562760 113508 562766
rect 113456 562702 113508 562708
rect 107672 559966 107916 559994
rect 109250 559966 109632 559994
rect 109894 559966 110184 559994
rect 111826 559966 111932 559994
rect 113468 559994 113496 562702
rect 116412 559994 116440 567190
rect 113468 559966 113758 559994
rect 116334 559966 116440 559994
rect 117332 559994 117360 574942
rect 118712 566574 118740 587823
rect 124416 586838 124444 587823
rect 128266 587752 128322 587761
rect 128266 587687 128322 587696
rect 124404 586832 124456 586838
rect 124404 586774 124456 586780
rect 124864 586832 124916 586838
rect 124864 586774 124916 586780
rect 122746 586392 122802 586401
rect 122746 586327 122802 586336
rect 122760 569294 122788 586327
rect 122748 569288 122800 569294
rect 122748 569230 122800 569236
rect 118700 566568 118752 566574
rect 118700 566510 118752 566516
rect 121552 566092 121604 566098
rect 121552 566034 121604 566040
rect 121564 559994 121592 566034
rect 124876 562562 124904 586774
rect 128280 566574 128308 587687
rect 128372 567866 128400 587823
rect 131776 586974 131804 587823
rect 131764 586968 131816 586974
rect 131764 586910 131816 586916
rect 133984 586838 134012 587823
rect 133972 586832 134024 586838
rect 133972 586774 134024 586780
rect 136652 574938 136680 587823
rect 139412 586906 139440 587823
rect 139400 586900 139452 586906
rect 139400 586842 139452 586848
rect 140792 576854 140820 589086
rect 141974 587888 142030 587897
rect 141974 587823 142030 587832
rect 159086 587888 159142 587897
rect 159086 587823 159142 587832
rect 141988 586906 142016 587823
rect 141976 586900 142028 586906
rect 141976 586842 142028 586848
rect 153844 586832 153896 586838
rect 153844 586774 153896 586780
rect 147220 581868 147272 581874
rect 147220 581810 147272 581816
rect 147232 576854 147260 581810
rect 140792 576826 140912 576854
rect 147232 576826 147352 576854
rect 136640 574932 136692 574938
rect 136640 574874 136692 574880
rect 128360 567860 128412 567866
rect 128360 567802 128412 567808
rect 140228 567452 140280 567458
rect 140228 567394 140280 567400
rect 131212 567384 131264 567390
rect 131212 567326 131264 567332
rect 128268 566568 128320 566574
rect 128268 566510 128320 566516
rect 130752 565548 130804 565554
rect 130752 565490 130804 565496
rect 124956 564596 125008 564602
rect 124956 564538 125008 564544
rect 124864 562556 124916 562562
rect 124864 562498 124916 562504
rect 117332 559966 117576 559994
rect 121486 559966 121592 559994
rect 124968 559994 124996 564538
rect 125690 562184 125746 562193
rect 125690 562119 125746 562128
rect 125704 559994 125732 562119
rect 130764 559994 130792 565490
rect 124968 559966 125350 559994
rect 125704 559966 125994 559994
rect 130502 559966 130792 559994
rect 131224 559994 131252 567326
rect 135904 565412 135956 565418
rect 135904 565354 135956 565360
rect 135916 559994 135944 565354
rect 138020 562080 138072 562086
rect 138020 562022 138072 562028
rect 131224 559966 131744 559994
rect 135654 559966 135944 559994
rect 138032 559994 138060 562022
rect 138572 562012 138624 562018
rect 138572 561954 138624 561960
rect 138584 559994 138612 561954
rect 140240 559994 140268 567394
rect 140884 559994 140912 576826
rect 143448 567316 143500 567322
rect 143448 567258 143500 567264
rect 143460 559994 143488 567258
rect 146208 560652 146260 560658
rect 146208 560594 146260 560600
rect 146220 559994 146248 560594
rect 147324 559994 147352 576826
rect 150532 576292 150584 576298
rect 150532 576234 150584 576240
rect 147956 573640 148008 573646
rect 147956 573582 148008 573588
rect 147968 559994 147996 573582
rect 148140 562488 148192 562494
rect 148140 562430 148192 562436
rect 138032 559966 138230 559994
rect 138584 559966 138874 559994
rect 140162 559966 140268 559994
rect 140806 559966 140912 559994
rect 143382 559966 143488 559994
rect 145958 559966 146248 559994
rect 147246 559966 147352 559994
rect 147890 559966 147996 559994
rect 148152 559994 148180 562430
rect 150544 559994 150572 576234
rect 153856 563689 153884 586774
rect 159100 583098 159128 587823
rect 163964 586900 164016 586906
rect 163964 586842 164016 586848
rect 160006 586392 160062 586401
rect 160006 586327 160062 586336
rect 159088 583092 159140 583098
rect 159088 583034 159140 583040
rect 160020 573646 160048 586327
rect 160100 580440 160152 580446
rect 160100 580382 160152 580388
rect 160112 576854 160140 580382
rect 163976 576854 164004 586842
rect 171692 579148 171744 579154
rect 171692 579090 171744 579096
rect 171704 576854 171732 579090
rect 160112 576826 160232 576854
rect 163976 576826 164096 576854
rect 171704 576826 171824 576854
rect 160008 573640 160060 573646
rect 160008 573582 160060 573588
rect 155224 572144 155276 572150
rect 155224 572086 155276 572092
rect 153936 563848 153988 563854
rect 153936 563790 153988 563796
rect 153842 563680 153898 563689
rect 153842 563615 153898 563624
rect 153948 559994 153976 563790
rect 148152 559966 148534 559994
rect 148888 559978 149178 559994
rect 148876 559972 149178 559978
rect 51078 559943 51134 559952
rect 148928 559966 149178 559972
rect 150466 559966 150572 559994
rect 153686 559966 153976 559994
rect 155236 559994 155264 572086
rect 157798 566128 157854 566137
rect 157798 566063 157854 566072
rect 157812 559994 157840 566063
rect 160204 559994 160232 576826
rect 163412 573708 163464 573714
rect 163412 573650 163464 573656
rect 162308 563576 162360 563582
rect 162308 563518 162360 563524
rect 155236 559966 155572 559994
rect 157550 559966 157840 559994
rect 160126 559966 160232 559994
rect 162320 559994 162348 563518
rect 163424 559994 163452 573650
rect 164068 559994 164096 576826
rect 168564 564800 168616 564806
rect 168564 564742 168616 564748
rect 164330 562592 164386 562601
rect 164330 562527 164386 562536
rect 162320 559966 162702 559994
rect 163346 559966 163452 559994
rect 163990 559966 164096 559994
rect 164344 559994 164372 562527
rect 168576 559994 168604 564742
rect 170770 562048 170826 562057
rect 170770 561983 170826 561992
rect 164344 559966 164634 559994
rect 168498 559966 168604 559994
rect 170784 559994 170812 561983
rect 171796 559994 171824 576826
rect 172624 576298 172652 668607
rect 172716 588538 172744 674834
rect 172704 588532 172756 588538
rect 172704 588474 172756 588480
rect 172612 576292 172664 576298
rect 172612 576234 172664 576240
rect 173176 562426 173204 685374
rect 347044 680944 347096 680950
rect 347044 680886 347096 680892
rect 173256 680468 173308 680474
rect 173256 680410 173308 680416
rect 173164 562420 173216 562426
rect 173164 562362 173216 562368
rect 173268 562358 173296 680410
rect 340880 676184 340932 676190
rect 340880 676126 340932 676132
rect 340892 675034 340920 676126
rect 340880 675028 340932 675034
rect 340880 674970 340932 674976
rect 328552 674960 328604 674966
rect 328550 674928 328552 674937
rect 340892 674937 340920 674970
rect 328604 674928 328606 674937
rect 328550 674863 328606 674872
rect 329746 674928 329802 674937
rect 329746 674863 329748 674872
rect 329800 674863 329802 674872
rect 340878 674928 340934 674937
rect 340878 674863 340934 674872
rect 329748 674834 329800 674840
rect 208306 626648 208362 626657
rect 208306 626583 208362 626592
rect 207662 625424 207718 625433
rect 207662 625359 207718 625368
rect 175278 608832 175334 608841
rect 175278 608767 175334 608776
rect 174544 599004 174596 599010
rect 174544 598946 174596 598952
rect 174556 566710 174584 598946
rect 174544 566704 174596 566710
rect 174544 566646 174596 566652
rect 175292 563718 175320 608767
rect 176566 607336 176622 607345
rect 176566 607271 176622 607280
rect 176580 607238 176608 607271
rect 176568 607232 176620 607238
rect 176568 607174 176620 607180
rect 176566 605976 176622 605985
rect 176566 605911 176622 605920
rect 176580 605878 176608 605911
rect 176568 605872 176620 605878
rect 176568 605814 176620 605820
rect 203524 605872 203576 605878
rect 203524 605814 203576 605820
rect 175370 604480 175426 604489
rect 175370 604415 175426 604424
rect 175384 565350 175412 604415
rect 175462 603120 175518 603129
rect 175462 603055 175518 603064
rect 175372 565344 175424 565350
rect 175372 565286 175424 565292
rect 175476 563854 175504 603055
rect 180064 586764 180116 586770
rect 180064 586706 180116 586712
rect 180076 565350 180104 586706
rect 200672 585200 200724 585206
rect 200672 585142 200724 585148
rect 200684 576854 200712 585142
rect 200684 576826 200804 576854
rect 190366 566264 190422 566273
rect 190366 566199 190422 566208
rect 180064 565344 180116 565350
rect 180064 565286 180116 565292
rect 175464 563848 175516 563854
rect 175464 563790 175516 563796
rect 179696 563848 179748 563854
rect 179696 563790 179748 563796
rect 175280 563712 175332 563718
rect 175280 563654 175332 563660
rect 179144 563508 179196 563514
rect 179144 563450 179196 563456
rect 173256 562352 173308 562358
rect 173256 562294 173308 562300
rect 174542 561912 174598 561921
rect 174542 561847 174598 561856
rect 174556 559994 174584 561847
rect 179156 559994 179184 563450
rect 179708 559994 179736 563790
rect 180708 563576 180760 563582
rect 180708 563518 180760 563524
rect 180720 560130 180748 563518
rect 181076 563440 181128 563446
rect 181076 563382 181128 563388
rect 188710 563408 188766 563417
rect 180720 560102 180840 560130
rect 180812 559994 180840 560102
rect 170784 559966 171074 559994
rect 171718 559966 171824 559994
rect 174294 559966 174584 559994
rect 178802 559966 179184 559994
rect 179446 559966 179736 559994
rect 180734 559966 180840 559994
rect 181088 559994 181116 563382
rect 188710 563343 188766 563352
rect 186872 562420 186924 562426
rect 186872 562362 186924 562368
rect 181628 561876 181680 561882
rect 181628 561818 181680 561824
rect 184848 561876 184900 561882
rect 184848 561818 184900 561824
rect 181640 559994 181668 561818
rect 183008 560584 183060 560590
rect 183008 560526 183060 560532
rect 183020 559994 183048 560526
rect 184860 559994 184888 561818
rect 186884 559994 186912 562362
rect 188724 559994 188752 563343
rect 189446 562048 189502 562057
rect 189446 561983 189502 561992
rect 189460 559994 189488 561983
rect 190380 560130 190408 566199
rect 198464 566160 198516 566166
rect 198464 566102 198516 566108
rect 191380 564732 191432 564738
rect 191380 564674 191432 564680
rect 190380 560102 190454 560130
rect 190426 559994 190454 560102
rect 181088 559966 181378 559994
rect 181640 559966 182022 559994
rect 182666 559966 183048 559994
rect 184598 559966 184888 559994
rect 186530 559966 186912 559994
rect 188462 559966 188752 559994
rect 189106 559966 189488 559994
rect 190394 559966 190454 559994
rect 191392 559994 191420 564674
rect 195886 564632 195942 564641
rect 195886 564567 195942 564576
rect 192574 562184 192630 562193
rect 192574 562119 192630 562128
rect 192588 559994 192616 562119
rect 193864 561944 193916 561950
rect 193864 561886 193916 561892
rect 191392 559966 191682 559994
rect 192326 559966 192616 559994
rect 193876 559994 193904 561886
rect 195900 559994 195928 564567
rect 198476 559994 198504 566102
rect 200776 559994 200804 576826
rect 203536 565486 203564 605814
rect 207018 599448 207074 599457
rect 207018 599383 207074 599392
rect 207032 599010 207060 599383
rect 207020 599004 207072 599010
rect 207020 598946 207072 598952
rect 207676 589218 207704 625359
rect 207754 623792 207810 623801
rect 207754 623727 207810 623736
rect 207768 589286 207796 623727
rect 208214 622432 208270 622441
rect 208214 622367 208270 622376
rect 208122 621072 208178 621081
rect 208122 621007 208178 621016
rect 208030 617672 208086 617681
rect 208030 617607 208086 617616
rect 207938 597680 207994 597689
rect 207938 597615 207994 597624
rect 207756 589280 207808 589286
rect 207756 589222 207808 589228
rect 207664 589212 207716 589218
rect 207664 589154 207716 589160
rect 207952 570926 207980 597615
rect 208044 579086 208072 617607
rect 208032 579080 208084 579086
rect 208032 579022 208084 579028
rect 207940 570920 207992 570926
rect 207940 570862 207992 570868
rect 208136 570858 208164 621007
rect 208124 570852 208176 570858
rect 208124 570794 208176 570800
rect 208228 567866 208256 622367
rect 208320 570790 208348 626583
rect 209686 619984 209742 619993
rect 209686 619919 209742 619928
rect 209044 607232 209096 607238
rect 209044 607174 209096 607180
rect 209056 574938 209084 607174
rect 209134 598360 209190 598369
rect 209134 598295 209190 598304
rect 209148 590034 209176 598295
rect 209136 590028 209188 590034
rect 209136 589970 209188 589976
rect 209148 580514 209176 589970
rect 209136 580508 209188 580514
rect 209136 580450 209188 580456
rect 209044 574932 209096 574938
rect 209044 574874 209096 574880
rect 209700 572218 209728 619919
rect 239312 589280 239364 589286
rect 239312 589222 239364 589228
rect 225144 589212 225196 589218
rect 225144 589154 225196 589160
rect 224958 587888 225014 587897
rect 224958 587823 225014 587832
rect 209780 586764 209832 586770
rect 209780 586706 209832 586712
rect 209792 580378 209820 586706
rect 215484 584656 215536 584662
rect 215484 584598 215536 584604
rect 211620 584588 211672 584594
rect 211620 584530 211672 584536
rect 209780 580372 209832 580378
rect 209780 580314 209832 580320
rect 211632 576854 211660 584530
rect 215496 576854 215524 584598
rect 219992 577652 220044 577658
rect 219992 577594 220044 577600
rect 220004 576854 220032 577594
rect 211632 576826 211752 576854
rect 215496 576826 215616 576854
rect 220004 576826 220124 576854
rect 209688 572212 209740 572218
rect 209688 572154 209740 572160
rect 208308 570784 208360 570790
rect 208308 570726 208360 570732
rect 208216 567860 208268 567866
rect 208216 567802 208268 567808
rect 203524 565480 203576 565486
rect 203524 565422 203576 565428
rect 204168 563916 204220 563922
rect 204168 563858 204220 563864
rect 203616 562760 203668 562766
rect 203616 562702 203668 562708
rect 201408 561944 201460 561950
rect 201408 561886 201460 561892
rect 201420 559994 201448 561886
rect 203628 559994 203656 562702
rect 204180 559994 204208 563858
rect 208032 563712 208084 563718
rect 208032 563654 208084 563660
rect 207478 560960 207534 560969
rect 207478 560895 207534 560904
rect 207492 559994 207520 560895
rect 208044 559994 208072 563654
rect 208768 562488 208820 562494
rect 208768 562430 208820 562436
rect 208780 559994 208808 562430
rect 211724 559994 211752 576826
rect 214472 562556 214524 562562
rect 214472 562498 214524 562504
rect 214484 559994 214512 562498
rect 215588 559994 215616 576826
rect 217508 568676 217560 568682
rect 217508 568618 217560 568624
rect 217048 566092 217100 566098
rect 217048 566034 217100 566040
rect 217060 559994 217088 566034
rect 217520 559994 217548 568618
rect 220096 559994 220124 576826
rect 224972 576230 225000 587823
rect 225156 576854 225184 589154
rect 227810 587888 227866 587897
rect 227810 587823 227866 587832
rect 231674 587888 231730 587897
rect 231674 587823 231730 587832
rect 234526 587888 234582 587897
rect 234526 587823 234582 587832
rect 235998 587888 236054 587897
rect 235998 587823 236054 587832
rect 237378 587888 237434 587897
rect 237378 587823 237434 587832
rect 238666 587888 238722 587897
rect 238666 587823 238722 587832
rect 238850 587888 238906 587897
rect 238850 587823 238906 587832
rect 227824 586838 227852 587823
rect 227812 586832 227864 586838
rect 227812 586774 227864 586780
rect 231688 577658 231716 587823
rect 231766 586392 231822 586401
rect 231766 586327 231822 586336
rect 233146 586392 233202 586401
rect 233146 586327 233202 586336
rect 231676 577652 231728 577658
rect 231676 577594 231728 577600
rect 225156 576826 225276 576854
rect 224960 576224 225012 576230
rect 224960 576166 225012 576172
rect 222016 568744 222068 568750
rect 222016 568686 222068 568692
rect 222028 559994 222056 568686
rect 222200 563780 222252 563786
rect 222200 563722 222252 563728
rect 224776 563780 224828 563786
rect 224776 563722 224828 563728
rect 193876 559966 194212 559994
rect 195546 559966 195928 559994
rect 198122 559966 198504 559994
rect 200698 559966 200804 559994
rect 201342 559966 201448 559994
rect 203274 559966 203656 559994
rect 203918 559966 204208 559994
rect 207138 559966 207520 559994
rect 207782 559966 208072 559994
rect 208426 559966 208808 559994
rect 211646 559966 211752 559994
rect 214222 559966 214512 559994
rect 215510 559966 215616 559994
rect 216798 559966 217088 559994
rect 217442 559966 217548 559994
rect 220018 559966 220124 559994
rect 221950 559966 222056 559994
rect 222212 559994 222240 563722
rect 224224 563644 224276 563650
rect 224224 563586 224276 563592
rect 224236 559994 224264 563586
rect 224788 559994 224816 563722
rect 225248 559994 225276 576826
rect 231780 569362 231808 586327
rect 231768 569356 231820 569362
rect 231768 569298 231820 569304
rect 233160 567934 233188 586327
rect 234540 569430 234568 587823
rect 234618 587752 234674 587761
rect 234618 587687 234674 587696
rect 234632 577590 234660 587687
rect 234620 577584 234672 577590
rect 234620 577526 234672 577532
rect 236012 573714 236040 587823
rect 237392 575006 237420 587823
rect 238680 576230 238708 587823
rect 238758 586800 238814 586809
rect 238758 586735 238760 586744
rect 238812 586735 238814 586744
rect 238760 586706 238812 586712
rect 238864 579154 238892 587823
rect 238852 579148 238904 579154
rect 238852 579090 238904 579096
rect 239324 576854 239352 589222
rect 257342 588976 257398 588985
rect 257342 588911 257398 588920
rect 240506 587888 240562 587897
rect 240506 587823 240562 587832
rect 242438 587888 242494 587897
rect 242438 587823 242494 587832
rect 243542 587888 243598 587897
rect 243542 587823 243598 587832
rect 245566 587888 245622 587897
rect 245566 587823 245622 587832
rect 245842 587888 245898 587897
rect 245842 587823 245898 587832
rect 247038 587888 247094 587897
rect 247038 587823 247094 587832
rect 248142 587888 248198 587897
rect 248142 587823 248198 587832
rect 248418 587888 248474 587897
rect 248418 587823 248474 587832
rect 249706 587888 249762 587897
rect 249706 587823 249762 587832
rect 252650 587888 252706 587897
rect 252650 587823 252706 587832
rect 253938 587888 253994 587897
rect 253938 587823 253994 587832
rect 255318 587888 255374 587897
rect 255318 587823 255374 587832
rect 256606 587888 256662 587897
rect 256606 587823 256662 587832
rect 240520 586022 240548 587823
rect 240782 587752 240838 587761
rect 240782 587687 240838 587696
rect 240796 586838 240824 587687
rect 240784 586832 240836 586838
rect 240784 586774 240836 586780
rect 242452 586770 242480 587823
rect 242440 586764 242492 586770
rect 242440 586706 242492 586712
rect 240508 586016 240560 586022
rect 240508 585958 240560 585964
rect 243556 581942 243584 587823
rect 245580 586702 245608 587823
rect 245568 586696 245620 586702
rect 245568 586638 245620 586644
rect 245856 586634 245884 587823
rect 246946 587752 247002 587761
rect 246946 587687 247002 587696
rect 245844 586628 245896 586634
rect 245844 586570 245896 586576
rect 244186 586392 244242 586401
rect 244186 586327 244242 586336
rect 243544 581936 243596 581942
rect 243544 581878 243596 581884
rect 239324 576826 239444 576854
rect 238668 576224 238720 576230
rect 238668 576166 238720 576172
rect 237380 575000 237432 575006
rect 237380 574942 237432 574948
rect 236000 573708 236052 573714
rect 236000 573650 236052 573656
rect 237380 572076 237432 572082
rect 237380 572018 237432 572024
rect 234528 569424 234580 569430
rect 234528 569366 234580 569372
rect 234896 568880 234948 568886
rect 234896 568822 234948 568828
rect 233148 567928 233200 567934
rect 233148 567870 233200 567876
rect 226892 566636 226944 566642
rect 226892 566578 226944 566584
rect 225420 565344 225472 565350
rect 225420 565286 225472 565292
rect 222212 559966 222548 559994
rect 223882 559966 224264 559994
rect 224526 559966 224816 559994
rect 225170 559966 225276 559994
rect 225432 559994 225460 565286
rect 226800 562352 226852 562358
rect 226800 562294 226852 562300
rect 226812 559994 226840 562294
rect 225432 559966 225814 559994
rect 226458 559966 226840 559994
rect 226904 559994 226932 566578
rect 230388 565344 230440 565350
rect 230388 565286 230440 565292
rect 230400 559994 230428 565286
rect 232504 564732 232556 564738
rect 232504 564674 232556 564680
rect 232516 559994 232544 564674
rect 233792 560788 233844 560794
rect 233792 560730 233844 560736
rect 233804 559994 233832 560730
rect 234908 559994 234936 568822
rect 236368 562216 236420 562222
rect 236368 562158 236420 562164
rect 235816 560720 235868 560726
rect 235816 560662 235868 560668
rect 235828 559994 235856 560662
rect 236380 559994 236408 562158
rect 237392 560266 237420 572018
rect 238668 564936 238720 564942
rect 238668 564878 238720 564884
rect 226904 559966 227102 559994
rect 230322 559966 230428 559994
rect 232254 559966 232544 559994
rect 233542 559966 233832 559994
rect 234830 559966 234936 559994
rect 235474 559966 235856 559994
rect 236118 559966 236408 559994
rect 237346 560238 237420 560266
rect 237346 559980 237374 560238
rect 238680 560130 238708 564878
rect 238680 560102 238800 560130
rect 238772 559994 238800 560102
rect 239416 559994 239444 576826
rect 244200 576298 244228 586327
rect 245752 580372 245804 580378
rect 245752 580314 245804 580320
rect 245764 576854 245792 580314
rect 246960 577590 246988 587687
rect 246948 577584 247000 577590
rect 246948 577526 247000 577532
rect 245764 576826 245884 576854
rect 244188 576292 244240 576298
rect 244188 576234 244240 576240
rect 244556 568812 244608 568818
rect 244556 568754 244608 568760
rect 243268 567520 243320 567526
rect 243268 567462 243320 567468
rect 241426 566400 241482 566409
rect 241426 566335 241482 566344
rect 240968 566228 241020 566234
rect 240968 566170 241020 566176
rect 240046 562320 240102 562329
rect 240046 562255 240102 562264
rect 240060 559994 240088 562255
rect 240980 559994 241008 566170
rect 241440 559994 241468 566335
rect 243280 559994 243308 567462
rect 243452 565480 243504 565486
rect 243452 565422 243504 565428
rect 238694 559966 238800 559994
rect 239338 559966 239444 559994
rect 239982 559966 240088 559994
rect 240626 559966 241008 559994
rect 241270 559966 241468 559994
rect 243202 559966 243308 559994
rect 243464 559994 243492 565422
rect 244568 559994 244596 568754
rect 244740 564664 244792 564670
rect 244740 564606 244792 564612
rect 243464 559966 243846 559994
rect 244490 559966 244596 559994
rect 244752 559994 244780 564606
rect 245856 559994 245884 576826
rect 247052 563922 247080 587823
rect 248156 586974 248184 587823
rect 248144 586968 248196 586974
rect 248144 586910 248196 586916
rect 248432 581806 248460 587823
rect 248420 581800 248472 581806
rect 248420 581742 248472 581748
rect 249720 568070 249748 587823
rect 249798 587752 249854 587761
rect 249798 587687 249854 587696
rect 252558 587752 252614 587761
rect 252558 587687 252614 587696
rect 249708 568064 249760 568070
rect 249708 568006 249760 568012
rect 249812 565214 249840 587687
rect 252466 586392 252522 586401
rect 252466 586327 252522 586336
rect 250444 580508 250496 580514
rect 250444 580450 250496 580456
rect 249800 565208 249852 565214
rect 249800 565150 249852 565156
rect 248328 564664 248380 564670
rect 248328 564606 248380 564612
rect 247040 563916 247092 563922
rect 247040 563858 247092 563864
rect 248340 560130 248368 564606
rect 249708 563440 249760 563446
rect 249708 563382 249760 563388
rect 249720 562562 249748 563382
rect 249708 562556 249760 562562
rect 249708 562498 249760 562504
rect 250456 562086 250484 580450
rect 252480 569498 252508 586327
rect 252468 569492 252520 569498
rect 252468 569434 252520 569440
rect 252572 565418 252600 587687
rect 252664 569265 252692 587823
rect 253952 581738 253980 587823
rect 253940 581732 253992 581738
rect 253940 581674 253992 581680
rect 255332 572150 255360 587823
rect 256620 586906 256648 587823
rect 256608 586900 256660 586906
rect 256608 586842 256660 586848
rect 257356 576854 257384 588911
rect 292764 588532 292816 588538
rect 292764 588474 292816 588480
rect 257986 587888 258042 587897
rect 257986 587823 258042 587832
rect 260654 587888 260710 587897
rect 260654 587823 260710 587832
rect 261022 587888 261078 587897
rect 261022 587823 261078 587832
rect 262034 587888 262090 587897
rect 262034 587823 262090 587832
rect 262218 587888 262274 587897
rect 262218 587823 262274 587832
rect 264886 587888 264942 587897
rect 264886 587823 264942 587832
rect 266266 587888 266322 587897
rect 266266 587823 266322 587832
rect 268934 587888 268990 587897
rect 268934 587823 268990 587832
rect 269762 587888 269818 587897
rect 269762 587823 269818 587832
rect 270498 587888 270554 587897
rect 270498 587823 270554 587832
rect 273534 587888 273590 587897
rect 273534 587823 273590 587832
rect 274638 587888 274694 587897
rect 274638 587823 274694 587832
rect 281078 587888 281134 587897
rect 281078 587823 281134 587832
rect 282918 587888 282974 587897
rect 282918 587823 282974 587832
rect 286322 587888 286378 587897
rect 286322 587823 286378 587832
rect 288438 587888 288494 587897
rect 288438 587823 288494 587832
rect 291014 587888 291070 587897
rect 291014 587823 291070 587832
rect 257356 576826 257476 576854
rect 255320 572144 255372 572150
rect 255320 572086 255372 572092
rect 252650 569256 252706 569265
rect 252650 569191 252706 569200
rect 254860 567588 254912 567594
rect 254860 567530 254912 567536
rect 252560 565412 252612 565418
rect 252560 565354 252612 565360
rect 253940 565276 253992 565282
rect 253940 565218 253992 565224
rect 251824 564868 251876 564874
rect 251824 564810 251876 564816
rect 250444 562080 250496 562086
rect 250444 562022 250496 562028
rect 248340 560102 248414 560130
rect 248386 559994 248414 560102
rect 250456 559994 250484 562022
rect 251836 559994 251864 564810
rect 244752 559966 245134 559994
rect 245778 559966 245884 559994
rect 248354 559966 248414 559994
rect 250286 559966 250484 559994
rect 251574 559966 251864 559994
rect 253952 559994 253980 565218
rect 254872 559994 254900 567530
rect 255780 564052 255832 564058
rect 255780 563994 255832 564000
rect 255688 560856 255740 560862
rect 255688 560798 255740 560804
rect 255700 559994 255728 560798
rect 253952 559966 254150 559994
rect 254794 559966 254900 559994
rect 255438 559966 255728 559994
rect 255792 559994 255820 563994
rect 257448 559994 257476 576826
rect 258000 566642 258028 587823
rect 258170 586800 258226 586809
rect 258170 586735 258226 586744
rect 258078 586392 258134 586401
rect 258078 586327 258134 586336
rect 258092 570722 258120 586327
rect 258184 580446 258212 586735
rect 260668 586634 260696 587823
rect 261036 587042 261064 587823
rect 261024 587036 261076 587042
rect 261024 586978 261076 586984
rect 260656 586628 260708 586634
rect 260656 586570 260708 586576
rect 258172 580440 258224 580446
rect 258172 580382 258224 580388
rect 258080 570716 258132 570722
rect 258080 570658 258132 570664
rect 262048 566710 262076 587823
rect 262036 566704 262088 566710
rect 262036 566646 262088 566652
rect 257988 566636 258040 566642
rect 257988 566578 258040 566584
rect 262232 563854 262260 587823
rect 264426 587752 264482 587761
rect 264426 587687 264482 587696
rect 264440 587586 264468 587687
rect 264428 587580 264480 587586
rect 264428 587522 264480 587528
rect 263506 586392 263562 586401
rect 263506 586327 263562 586336
rect 263520 570722 263548 586327
rect 263508 570716 263560 570722
rect 263508 570658 263560 570664
rect 263416 565004 263468 565010
rect 263416 564946 263468 564952
rect 262220 563848 262272 563854
rect 262220 563790 262272 563796
rect 260746 563544 260802 563553
rect 260746 563479 260802 563488
rect 260288 562148 260340 562154
rect 260288 562090 260340 562096
rect 260300 559994 260328 562090
rect 260760 559994 260788 563479
rect 263428 559994 263456 564946
rect 264900 563922 264928 587823
rect 264978 587752 265034 587761
rect 264978 587687 265034 587696
rect 264992 573578 265020 587687
rect 265072 586016 265124 586022
rect 265072 585958 265124 585964
rect 265084 576854 265112 585958
rect 265084 576826 265204 576854
rect 264980 573572 265032 573578
rect 264980 573514 265032 573520
rect 264888 563916 264940 563922
rect 264888 563858 264940 563864
rect 265176 559994 265204 576826
rect 266280 569566 266308 587823
rect 267646 586392 267702 586401
rect 267646 586327 267702 586336
rect 266268 569560 266320 569566
rect 266268 569502 266320 569508
rect 267660 568002 267688 586327
rect 268948 572082 268976 587823
rect 269026 586392 269082 586401
rect 269026 586327 269082 586336
rect 268936 572076 268988 572082
rect 268936 572018 268988 572024
rect 269040 568138 269068 586327
rect 269776 584594 269804 587823
rect 269764 584588 269816 584594
rect 269764 584530 269816 584536
rect 270224 583092 270276 583098
rect 270224 583034 270276 583040
rect 270236 576854 270264 583034
rect 270512 577561 270540 587823
rect 273548 586090 273576 587823
rect 273536 586084 273588 586090
rect 273536 586026 273588 586032
rect 274652 581874 274680 587823
rect 281092 587110 281120 587823
rect 281080 587104 281132 587110
rect 281080 587046 281132 587052
rect 277490 586528 277546 586537
rect 277490 586463 277546 586472
rect 274640 581868 274692 581874
rect 274640 581810 274692 581816
rect 270498 577552 270554 577561
rect 270498 577487 270554 577496
rect 270236 576826 270356 576854
rect 269028 568132 269080 568138
rect 269028 568074 269080 568080
rect 267648 567996 267700 568002
rect 267648 567938 267700 567944
rect 265992 565072 266044 565078
rect 265992 565014 266044 565020
rect 266004 559994 266032 565014
rect 269856 564800 269908 564806
rect 269856 564742 269908 564748
rect 268014 560824 268070 560833
rect 268014 560759 268070 560768
rect 255792 559966 256036 559994
rect 257370 559966 257476 559994
rect 259946 559966 260328 559994
rect 260590 559966 260788 559994
rect 263166 559966 263456 559994
rect 265098 559966 265204 559994
rect 265742 559966 266032 559994
rect 268028 559994 268056 560759
rect 269868 559994 269896 564742
rect 270328 559994 270356 576826
rect 277504 570761 277532 586463
rect 282932 584662 282960 587823
rect 286336 587178 286364 587823
rect 286324 587172 286376 587178
rect 286324 587114 286376 587120
rect 282920 584656 282972 584662
rect 282920 584598 282972 584604
rect 288452 583137 288480 587823
rect 291028 587246 291056 587823
rect 291016 587240 291068 587246
rect 291016 587182 291068 587188
rect 288438 583128 288494 583137
rect 288438 583063 288494 583072
rect 281816 577584 281868 577590
rect 281816 577526 281868 577532
rect 281828 576854 281856 577526
rect 292776 576854 292804 588474
rect 317420 588464 317472 588470
rect 317420 588406 317472 588412
rect 298098 587888 298154 587897
rect 298098 587823 298154 587832
rect 300858 587888 300914 587897
rect 300858 587823 300914 587832
rect 302238 587888 302294 587897
rect 302238 587823 302294 587832
rect 305090 587888 305146 587897
rect 305090 587823 305146 587832
rect 308494 587888 308550 587897
rect 308494 587823 308550 587832
rect 310518 587888 310574 587897
rect 310518 587823 310574 587832
rect 313278 587888 313334 587897
rect 313278 587823 313334 587832
rect 316038 587888 316094 587897
rect 316038 587823 316094 587832
rect 293866 586392 293922 586401
rect 293866 586327 293922 586336
rect 296626 586392 296682 586401
rect 296626 586327 296682 586336
rect 281828 576826 281948 576854
rect 292776 576826 292896 576854
rect 278688 572212 278740 572218
rect 278688 572154 278740 572160
rect 277490 570752 277546 570761
rect 277490 570687 277546 570696
rect 272892 568948 272944 568954
rect 272892 568890 272944 568896
rect 272904 559994 272932 568890
rect 275008 566296 275060 566302
rect 275008 566238 275060 566244
rect 274454 562592 274510 562601
rect 274454 562527 274510 562536
rect 274468 559994 274496 562527
rect 275020 559994 275048 566238
rect 278320 562284 278372 562290
rect 278320 562226 278372 562232
rect 278332 559994 278360 562226
rect 278700 559994 278728 572154
rect 281920 559994 281948 576826
rect 289174 568848 289230 568857
rect 289174 568783 289230 568792
rect 287888 560924 287940 560930
rect 287888 560866 287940 560872
rect 287900 559994 287928 560866
rect 268028 559966 268318 559994
rect 269606 559966 269896 559994
rect 270250 559966 270356 559994
rect 272826 559966 272932 559994
rect 274114 559966 274496 559994
rect 274758 559966 275048 559994
rect 276690 559978 277072 559994
rect 276690 559972 277084 559978
rect 276690 559966 277032 559972
rect 148876 559914 148928 559920
rect 277978 559966 278360 559994
rect 278622 559966 278728 559994
rect 281842 559966 281948 559994
rect 287638 559966 287928 559994
rect 289188 559994 289216 568783
rect 291200 560992 291252 560998
rect 291200 560934 291252 560940
rect 291212 559994 291240 560934
rect 292868 559994 292896 576826
rect 293880 566778 293908 586327
rect 296640 568206 296668 586327
rect 298112 586022 298140 587823
rect 298100 586016 298152 586022
rect 298100 585958 298152 585964
rect 297916 580440 297968 580446
rect 297916 580382 297968 580388
rect 297928 576854 297956 580382
rect 297928 576826 298048 576854
rect 296628 568200 296680 568206
rect 296628 568142 296680 568148
rect 293868 566772 293920 566778
rect 293868 566714 293920 566720
rect 295708 565140 295760 565146
rect 295708 565082 295760 565088
rect 294326 562728 294382 562737
rect 294326 562663 294382 562672
rect 289188 559966 289524 559994
rect 290858 559966 291240 559994
rect 292790 559966 292896 559994
rect 294340 559994 294368 562663
rect 294788 560108 294840 560114
rect 294788 560050 294840 560056
rect 294340 559966 294676 559994
rect 294800 559978 294828 560050
rect 295720 559994 295748 565082
rect 297638 564768 297694 564777
rect 297638 564703 297694 564712
rect 297652 559994 297680 564703
rect 298020 559994 298048 576826
rect 300872 572014 300900 587823
rect 302252 579018 302280 587823
rect 302240 579012 302292 579018
rect 302240 578954 302292 578960
rect 305104 574705 305132 587823
rect 308508 587314 308536 587823
rect 308496 587308 308548 587314
rect 308496 587250 308548 587256
rect 306932 586084 306984 586090
rect 306932 586026 306984 586032
rect 306288 578944 306340 578950
rect 306288 578886 306340 578892
rect 305090 574696 305146 574705
rect 305090 574631 305146 574640
rect 300860 572008 300912 572014
rect 300860 571950 300912 571956
rect 298928 564528 298980 564534
rect 298928 564470 298980 564476
rect 298940 559994 298968 564470
rect 299388 563848 299440 563854
rect 299388 563790 299440 563796
rect 299400 559994 299428 563790
rect 301412 563372 301464 563378
rect 301412 563314 301464 563320
rect 294788 559972 294840 559978
rect 277032 559914 277084 559920
rect 295720 559966 296010 559994
rect 297298 559966 297680 559994
rect 297942 559966 298048 559994
rect 298586 559966 298968 559994
rect 299230 559966 299428 559994
rect 301424 559994 301452 563314
rect 306300 563054 306328 578886
rect 306944 576854 306972 586026
rect 307760 584656 307812 584662
rect 307760 584598 307812 584604
rect 307772 576854 307800 584598
rect 306944 576826 307064 576854
rect 307772 576826 308352 576854
rect 306300 563026 306420 563054
rect 304080 562556 304132 562562
rect 304080 562498 304132 562504
rect 304092 559994 304120 562498
rect 305920 561060 305972 561066
rect 305920 561002 305972 561008
rect 305932 559994 305960 561002
rect 306392 559994 306420 563026
rect 307036 559994 307064 576826
rect 307668 563372 307720 563378
rect 307668 563314 307720 563320
rect 307680 559994 307708 563314
rect 308034 562456 308090 562465
rect 308034 562391 308090 562400
rect 301424 559966 301806 559994
rect 303738 559966 304120 559994
rect 305670 559966 305960 559994
rect 306314 559966 306420 559994
rect 306958 559966 307064 559994
rect 307602 559966 307708 559994
rect 308048 559994 308076 562391
rect 308324 559994 308352 576826
rect 310532 565350 310560 587823
rect 313292 567905 313320 587823
rect 316052 587382 316080 587823
rect 316040 587376 316092 587382
rect 316040 587318 316092 587324
rect 317432 576854 317460 588406
rect 333886 587888 333942 587897
rect 333886 587823 333942 587832
rect 333900 586566 333928 587823
rect 333888 586560 333940 586566
rect 333888 586502 333940 586508
rect 333794 586392 333850 586401
rect 333794 586327 333850 586336
rect 320456 586016 320508 586022
rect 320456 585958 320508 585964
rect 320468 576854 320496 585958
rect 330116 581664 330168 581670
rect 330116 581606 330168 581612
rect 330128 576854 330156 581606
rect 317432 576826 318012 576854
rect 320468 576826 320588 576854
rect 330128 576826 330248 576854
rect 313278 567896 313334 567905
rect 313278 567831 313334 567840
rect 317788 566432 317840 566438
rect 317788 566374 317840 566380
rect 314936 566364 314988 566370
rect 314936 566306 314988 566312
rect 311164 565616 311216 565622
rect 311164 565558 311216 565564
rect 310520 565344 310572 565350
rect 310520 565286 310572 565292
rect 311176 559994 311204 565558
rect 313096 561128 313148 561134
rect 313096 561070 313148 561076
rect 313108 559994 313136 561070
rect 314948 559994 314976 566306
rect 315948 565140 316000 565146
rect 315948 565082 316000 565088
rect 315960 560130 315988 565082
rect 317800 560294 317828 566374
rect 317984 560294 318012 576826
rect 317800 560266 317920 560294
rect 317984 560266 318104 560294
rect 317892 560130 317920 560266
rect 315960 560102 316080 560130
rect 317892 560102 318012 560130
rect 315578 560008 315634 560017
rect 308048 559966 308246 559994
rect 308324 559966 308844 559994
rect 311176 559966 311466 559994
rect 312754 559966 313136 559994
rect 314686 559966 314976 559994
rect 315330 559966 315578 559994
rect 316052 559994 316080 560102
rect 317984 559994 318012 560102
rect 315974 559966 316080 559994
rect 317906 559966 318012 559994
rect 318076 559994 318104 560266
rect 320560 559994 320588 576826
rect 324688 565208 324740 565214
rect 324688 565150 324740 565156
rect 322110 564904 322166 564913
rect 322110 564839 322166 564848
rect 322124 559994 322152 564839
rect 324700 559994 324728 565150
rect 327816 563984 327868 563990
rect 327816 563926 327868 563932
rect 325976 563304 326028 563310
rect 325976 563246 326028 563252
rect 325608 560312 325660 560318
rect 325608 560254 325660 560260
rect 325620 560130 325648 560254
rect 325620 560102 325694 560130
rect 325666 559994 325694 560102
rect 318076 559966 318504 559994
rect 320482 559966 320588 559994
rect 321770 559966 322152 559994
rect 324346 559966 324728 559994
rect 325634 559966 325694 559994
rect 325988 559994 326016 563246
rect 327828 559994 327856 563926
rect 328366 563680 328422 563689
rect 328366 563615 328422 563624
rect 328380 559994 328408 563615
rect 330220 559994 330248 576826
rect 331496 573504 331548 573510
rect 331496 573446 331548 573452
rect 330482 560688 330538 560697
rect 330482 560623 330538 560632
rect 325988 559966 326278 559994
rect 327566 559966 327856 559994
rect 328210 559966 328408 559994
rect 330142 559966 330248 559994
rect 330496 559994 330524 560623
rect 331508 559994 331536 573446
rect 333808 565282 333836 586327
rect 346860 584588 346912 584594
rect 346860 584530 346912 584536
rect 346872 576854 346900 584530
rect 346872 576826 346992 576854
rect 335358 567488 335414 567497
rect 335358 567423 335414 567432
rect 333796 565276 333848 565282
rect 333796 565218 333848 565224
rect 335372 562426 335400 567423
rect 340144 564596 340196 564602
rect 340144 564538 340196 564544
rect 339132 564120 339184 564126
rect 339132 564062 339184 564068
rect 338764 563304 338816 563310
rect 338764 563246 338816 563252
rect 336648 563236 336700 563242
rect 336648 563178 336700 563184
rect 335360 562420 335412 562426
rect 335360 562362 335412 562368
rect 336372 562216 336424 562222
rect 336372 562158 336424 562164
rect 336280 562012 336332 562018
rect 336280 561954 336332 561960
rect 336292 559994 336320 561954
rect 336384 561105 336412 562158
rect 336370 561096 336426 561105
rect 336370 561031 336426 561040
rect 336660 559994 336688 563178
rect 338028 562624 338080 562630
rect 338028 562566 338080 562572
rect 337568 561740 337620 561746
rect 337568 561682 337620 561688
rect 337580 559994 337608 561682
rect 338040 559994 338068 562566
rect 338776 562494 338804 563246
rect 338764 562488 338816 562494
rect 338764 562430 338816 562436
rect 339144 562426 339172 564062
rect 339132 562420 339184 562426
rect 339132 562362 339184 562368
rect 339406 560416 339462 560425
rect 339406 560351 339462 560360
rect 330496 559966 330786 559994
rect 331430 559966 331536 559994
rect 334650 559978 335032 559994
rect 334650 559972 335044 559978
rect 334650 559966 334992 559972
rect 315578 559943 315634 559952
rect 294788 559914 294840 559920
rect 335938 559966 336320 559994
rect 336582 559966 336688 559994
rect 337226 559966 337608 559994
rect 337870 559966 338068 559994
rect 339420 559978 339448 560351
rect 340156 559994 340184 564538
rect 343732 563916 343784 563922
rect 343732 563858 343784 563864
rect 340788 562760 340840 562766
rect 340788 562702 340840 562708
rect 339408 559972 339460 559978
rect 334992 559914 335044 559920
rect 339802 559966 340184 559994
rect 340446 559978 340736 559994
rect 340800 559978 340828 562702
rect 341982 561776 342038 561785
rect 341982 561711 342038 561720
rect 341996 559994 342024 561711
rect 343744 559994 343772 563858
rect 346492 562284 346544 562290
rect 346492 562226 346544 562232
rect 346400 561740 346452 561746
rect 346400 561682 346452 561688
rect 340446 559972 340748 559978
rect 340446 559966 340696 559972
rect 339408 559914 339460 559920
rect 340696 559914 340748 559920
rect 340788 559972 340840 559978
rect 341734 559966 342024 559994
rect 343666 559966 343772 559994
rect 346412 559978 346440 561682
rect 346504 560046 346532 562226
rect 346492 560040 346544 560046
rect 346964 559994 346992 576826
rect 347056 562630 347084 680886
rect 347148 655518 347176 700470
rect 347240 670682 347268 700538
rect 347792 686594 347820 702406
rect 364352 689314 364380 702406
rect 381544 700664 381596 700670
rect 381544 700606 381596 700612
rect 374828 698964 374880 698970
rect 374828 698906 374880 698912
rect 364340 689308 364392 689314
rect 364340 689250 364392 689256
rect 347780 686588 347832 686594
rect 347780 686530 347832 686536
rect 363604 685976 363656 685982
rect 363604 685918 363656 685924
rect 362224 685024 362276 685030
rect 362224 684966 362276 684972
rect 359464 684956 359516 684962
rect 359464 684898 359516 684904
rect 351184 675028 351236 675034
rect 351184 674970 351236 674976
rect 347780 674960 347832 674966
rect 347780 674902 347832 674908
rect 347228 670676 347280 670682
rect 347228 670618 347280 670624
rect 347136 655512 347188 655518
rect 347136 655454 347188 655460
rect 347136 641776 347188 641782
rect 347136 641718 347188 641724
rect 347148 580378 347176 641718
rect 347792 588470 347820 674902
rect 349158 669216 349214 669225
rect 349158 669151 349214 669160
rect 348792 661088 348844 661094
rect 348792 661030 348844 661036
rect 347780 588464 347832 588470
rect 347780 588406 347832 588412
rect 348424 587172 348476 587178
rect 348424 587114 348476 587120
rect 347136 580372 347188 580378
rect 347136 580314 347188 580320
rect 347964 579080 348016 579086
rect 347964 579022 348016 579028
rect 347780 569560 347832 569566
rect 347780 569502 347832 569508
rect 347044 562624 347096 562630
rect 347044 562566 347096 562572
rect 347688 562216 347740 562222
rect 347688 562158 347740 562164
rect 347700 559994 347728 562158
rect 346492 559982 346544 559988
rect 346400 559972 346452 559978
rect 340788 559914 340840 559920
rect 346886 559966 346992 559994
rect 347530 559966 347728 559994
rect 346400 559914 346452 559920
rect 347688 559904 347740 559910
rect 347688 559846 347740 559852
rect 347700 559638 347728 559846
rect 347688 559632 347740 559638
rect 347688 559574 347740 559580
rect 347688 559496 347740 559502
rect 347688 559438 347740 559444
rect 347700 559026 347728 559438
rect 347688 559020 347740 559026
rect 347688 558962 347740 558968
rect 347792 478009 347820 569502
rect 347872 565276 347924 565282
rect 347872 565218 347924 565224
rect 347884 522889 347912 565218
rect 347870 522880 347926 522889
rect 347870 522815 347926 522824
rect 347778 478000 347834 478009
rect 347778 477935 347834 477944
rect 347778 475008 347834 475017
rect 347778 474943 347834 474952
rect 47766 229392 47822 229401
rect 47766 229327 47822 229336
rect 47766 226400 47822 226409
rect 47766 226335 47822 226344
rect 47780 220289 47808 226335
rect 47766 220280 47822 220289
rect 47766 220215 47822 220224
rect 47860 202360 47912 202366
rect 47860 202302 47912 202308
rect 47872 199617 47900 202302
rect 347686 200968 347742 200977
rect 347686 200903 347742 200912
rect 347700 200394 347728 200903
rect 347688 200388 347740 200394
rect 347688 200330 347740 200336
rect 347686 200288 347742 200297
rect 347686 200223 347742 200232
rect 47858 199608 47914 199617
rect 47858 199543 47914 199552
rect 48056 198014 48084 200124
rect 48700 198694 48728 200124
rect 48688 198688 48740 198694
rect 48688 198630 48740 198636
rect 48044 198008 48096 198014
rect 48044 197950 48096 197956
rect 49344 197470 49372 200124
rect 49988 198150 50016 200124
rect 50344 199980 50396 199986
rect 50344 199922 50396 199928
rect 49976 198144 50028 198150
rect 49976 198086 50028 198092
rect 50068 198008 50120 198014
rect 50068 197950 50120 197956
rect 49516 197872 49568 197878
rect 49516 197814 49568 197820
rect 49332 197464 49384 197470
rect 49332 197406 49384 197412
rect 48964 192704 49016 192710
rect 48964 192646 49016 192652
rect 48686 187096 48742 187105
rect 48686 187031 48742 187040
rect 47860 182844 47912 182850
rect 47860 182786 47912 182792
rect 47872 142118 47900 182786
rect 48228 177336 48280 177342
rect 48228 177278 48280 177284
rect 48136 176180 48188 176186
rect 48136 176122 48188 176128
rect 47952 155780 48004 155786
rect 47952 155722 48004 155728
rect 47860 142112 47912 142118
rect 47860 142054 47912 142060
rect 47860 139460 47912 139466
rect 47860 139402 47912 139408
rect 47872 107642 47900 139402
rect 47860 107636 47912 107642
rect 47860 107578 47912 107584
rect 47676 82748 47728 82754
rect 47676 82690 47728 82696
rect 47492 28960 47544 28966
rect 47492 28902 47544 28908
rect 47964 22030 47992 155722
rect 48044 151360 48096 151366
rect 48044 151302 48096 151308
rect 47952 22024 48004 22030
rect 47952 21966 48004 21972
rect 46848 18352 46900 18358
rect 46848 18294 46900 18300
rect 48056 16590 48084 151302
rect 48044 16584 48096 16590
rect 48044 16526 48096 16532
rect 48148 16522 48176 176122
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48240 4146 48268 177278
rect 48700 149161 48728 187031
rect 48872 181484 48924 181490
rect 48872 181426 48924 181432
rect 48780 150136 48832 150142
rect 48780 150078 48832 150084
rect 48686 149152 48742 149161
rect 48686 149087 48742 149096
rect 48792 139466 48820 150078
rect 48780 139460 48832 139466
rect 48780 139402 48832 139408
rect 48884 108866 48912 181426
rect 48976 108934 49004 192646
rect 49424 191140 49476 191146
rect 49424 191082 49476 191088
rect 49332 178968 49384 178974
rect 49332 178910 49384 178916
rect 49056 177472 49108 177478
rect 49056 177414 49108 177420
rect 48964 108928 49016 108934
rect 48964 108870 49016 108876
rect 48872 108860 48924 108866
rect 48872 108802 48924 108808
rect 48964 107636 49016 107642
rect 48964 107578 49016 107584
rect 48976 11014 49004 107578
rect 49068 63510 49096 177414
rect 49148 151020 49200 151026
rect 49148 150962 49200 150968
rect 49056 63504 49108 63510
rect 49056 63446 49108 63452
rect 49160 27062 49188 150962
rect 49240 150884 49292 150890
rect 49240 150826 49292 150832
rect 49148 27056 49200 27062
rect 49148 26998 49200 27004
rect 49252 26178 49280 150826
rect 49344 41342 49372 178910
rect 49332 41336 49384 41342
rect 49332 41278 49384 41284
rect 49240 26172 49292 26178
rect 49240 26114 49292 26120
rect 49436 22778 49464 191082
rect 49528 28830 49556 197814
rect 50080 195242 50108 197950
rect 49804 195214 50108 195242
rect 49608 193112 49660 193118
rect 49608 193054 49660 193060
rect 49516 28824 49568 28830
rect 49516 28766 49568 28772
rect 49424 22772 49476 22778
rect 49424 22714 49476 22720
rect 49620 21350 49648 193054
rect 49804 175982 49832 195214
rect 49976 192432 50028 192438
rect 49976 192374 50028 192380
rect 49792 175976 49844 175982
rect 49792 175918 49844 175924
rect 49608 21344 49660 21350
rect 49608 21286 49660 21292
rect 49988 18766 50016 192374
rect 50252 180124 50304 180130
rect 50252 180066 50304 180072
rect 50068 174548 50120 174554
rect 50068 174490 50120 174496
rect 50080 129742 50108 174490
rect 50160 149796 50212 149802
rect 50160 149738 50212 149744
rect 50068 129736 50120 129742
rect 50068 129678 50120 129684
rect 50172 102270 50200 149738
rect 50160 102264 50212 102270
rect 50160 102206 50212 102212
rect 50264 93838 50292 180066
rect 50356 152726 50384 199922
rect 50632 198014 50660 200124
rect 50620 198008 50672 198014
rect 50620 197950 50672 197956
rect 51276 197402 51304 200124
rect 51908 198144 51960 198150
rect 53208 198098 53236 200124
rect 53852 198257 53880 200124
rect 55784 198422 55812 200124
rect 55772 198416 55824 198422
rect 55772 198358 55824 198364
rect 53838 198248 53894 198257
rect 53838 198183 53894 198192
rect 51908 198086 51960 198092
rect 51264 197396 51316 197402
rect 51264 197338 51316 197344
rect 50896 195424 50948 195430
rect 50896 195366 50948 195372
rect 50804 192568 50856 192574
rect 50804 192510 50856 192516
rect 50434 177576 50490 177585
rect 50434 177511 50490 177520
rect 50344 152720 50396 152726
rect 50344 152662 50396 152668
rect 50448 124982 50476 177511
rect 50712 171828 50764 171834
rect 50712 171770 50764 171776
rect 50620 151768 50672 151774
rect 50620 151710 50672 151716
rect 50528 151156 50580 151162
rect 50528 151098 50580 151104
rect 50436 124976 50488 124982
rect 50436 124918 50488 124924
rect 50342 124128 50398 124137
rect 50342 124063 50398 124072
rect 50252 93832 50304 93838
rect 50252 93774 50304 93780
rect 49976 18760 50028 18766
rect 49976 18702 50028 18708
rect 50356 18698 50384 124063
rect 50436 117632 50488 117638
rect 50436 117574 50488 117580
rect 50344 18692 50396 18698
rect 50344 18634 50396 18640
rect 48964 11008 49016 11014
rect 48964 10950 49016 10956
rect 48228 4140 48280 4146
rect 48228 4082 48280 4088
rect 46756 4004 46808 4010
rect 46756 3946 46808 3952
rect 50448 3942 50476 117574
rect 50540 24342 50568 151098
rect 50632 24750 50660 151710
rect 50724 28762 50752 171770
rect 50712 28756 50764 28762
rect 50712 28698 50764 28704
rect 50816 27538 50844 192510
rect 50908 28354 50936 195366
rect 51448 192840 51500 192846
rect 51448 192782 51500 192788
rect 51356 152924 51408 152930
rect 51356 152866 51408 152872
rect 51264 149864 51316 149870
rect 51264 149806 51316 149812
rect 51276 140826 51304 149806
rect 51264 140820 51316 140826
rect 51264 140762 51316 140768
rect 50988 126948 51040 126954
rect 50988 126890 51040 126896
rect 51000 119474 51028 126890
rect 50988 119468 51040 119474
rect 50988 119410 51040 119416
rect 50896 28348 50948 28354
rect 50896 28290 50948 28296
rect 50804 27532 50856 27538
rect 50804 27474 50856 27480
rect 50620 24744 50672 24750
rect 50620 24686 50672 24692
rect 50528 24336 50580 24342
rect 50528 24278 50580 24284
rect 51368 21622 51396 152866
rect 51460 23934 51488 192782
rect 51722 155544 51778 155553
rect 51722 155479 51778 155488
rect 51736 147801 51764 155479
rect 51722 147792 51778 147801
rect 51722 147727 51778 147736
rect 51814 147656 51870 147665
rect 51814 147591 51870 147600
rect 51632 143540 51684 143546
rect 51632 143482 51684 143488
rect 51538 142080 51594 142089
rect 51538 142015 51594 142024
rect 51552 124137 51580 142015
rect 51538 124128 51594 124137
rect 51538 124063 51594 124072
rect 51644 110430 51672 143482
rect 51724 138780 51776 138786
rect 51724 138722 51776 138728
rect 51736 126954 51764 138722
rect 51724 126948 51776 126954
rect 51724 126890 51776 126896
rect 51724 125112 51776 125118
rect 51724 125054 51776 125060
rect 51632 110424 51684 110430
rect 51632 110366 51684 110372
rect 51448 23928 51500 23934
rect 51448 23870 51500 23876
rect 51736 21826 51764 125054
rect 51828 118046 51856 147591
rect 51816 118040 51868 118046
rect 51816 117982 51868 117988
rect 51920 75886 51948 198086
rect 52564 198070 53236 198098
rect 52276 195764 52328 195770
rect 52276 195706 52328 195712
rect 52184 183456 52236 183462
rect 52184 183398 52236 183404
rect 52000 152448 52052 152454
rect 52000 152390 52052 152396
rect 51908 75880 51960 75886
rect 51908 75822 51960 75828
rect 52012 25906 52040 152390
rect 52092 151564 52144 151570
rect 52092 151506 52144 151512
rect 52000 25900 52052 25906
rect 52000 25842 52052 25848
rect 52104 21894 52132 151506
rect 52196 142225 52224 183398
rect 52182 142216 52238 142225
rect 52182 142151 52238 142160
rect 52288 28898 52316 195706
rect 52366 146568 52422 146577
rect 52366 146503 52422 146512
rect 52380 142202 52408 146503
rect 52380 142174 52500 142202
rect 52472 138786 52500 142174
rect 52460 138780 52512 138786
rect 52460 138722 52512 138728
rect 52368 123480 52420 123486
rect 52368 123422 52420 123428
rect 52276 28892 52328 28898
rect 52276 28834 52328 28840
rect 52092 21888 52144 21894
rect 52092 21830 52144 21836
rect 51724 21820 51776 21826
rect 51724 21762 51776 21768
rect 51356 21616 51408 21622
rect 51356 21558 51408 21564
rect 52380 17202 52408 123422
rect 52460 102264 52512 102270
rect 52460 102206 52512 102212
rect 52472 97918 52500 102206
rect 52460 97912 52512 97918
rect 52460 97854 52512 97860
rect 52564 27334 52592 198070
rect 53012 198008 53064 198014
rect 53012 197950 53064 197956
rect 52644 177404 52696 177410
rect 52644 177346 52696 177352
rect 52552 27328 52604 27334
rect 52552 27270 52604 27276
rect 52368 17196 52420 17202
rect 52368 17138 52420 17144
rect 52656 16574 52684 177346
rect 52828 169176 52880 169182
rect 52828 169118 52880 169124
rect 52736 151700 52788 151706
rect 52736 151642 52788 151648
rect 52748 24070 52776 151642
rect 52840 25634 52868 169118
rect 52920 149932 52972 149938
rect 52920 149874 52972 149880
rect 52828 25628 52880 25634
rect 52828 25570 52880 25576
rect 52736 24064 52788 24070
rect 52736 24006 52788 24012
rect 52932 23322 52960 149874
rect 52920 23316 52972 23322
rect 52920 23258 52972 23264
rect 52656 16546 52960 16574
rect 50436 3936 50488 3942
rect 50436 3878 50488 3884
rect 50158 3496 50214 3505
rect 50158 3431 50214 3440
rect 50172 480 50200 3431
rect 52932 490 52960 16546
rect 53024 3398 53052 197950
rect 54484 197464 54536 197470
rect 54484 197406 54536 197412
rect 53196 197396 53248 197402
rect 53196 197338 53248 197344
rect 53208 180794 53236 197338
rect 54208 192636 54260 192642
rect 54208 192578 54260 192584
rect 53472 187604 53524 187610
rect 53472 187546 53524 187552
rect 53380 185904 53432 185910
rect 53380 185846 53432 185852
rect 53116 180766 53236 180794
rect 53116 180266 53144 180766
rect 53104 180260 53156 180266
rect 53104 180202 53156 180208
rect 53288 175024 53340 175030
rect 53288 174966 53340 174972
rect 53300 123554 53328 174966
rect 53288 123548 53340 123554
rect 53288 123490 53340 123496
rect 53196 117700 53248 117706
rect 53196 117642 53248 117648
rect 53208 95130 53236 117642
rect 53392 104786 53420 185846
rect 53484 146130 53512 187546
rect 53564 187400 53616 187406
rect 53564 187342 53616 187348
rect 53472 146124 53524 146130
rect 53472 146066 53524 146072
rect 53576 135930 53604 187342
rect 53840 142180 53892 142186
rect 53840 142122 53892 142128
rect 53746 135960 53802 135969
rect 53564 135924 53616 135930
rect 53746 135895 53802 135904
rect 53564 135866 53616 135872
rect 53760 124817 53788 135895
rect 53746 124808 53802 124817
rect 53746 124743 53802 124752
rect 53656 123616 53708 123622
rect 53656 123558 53708 123564
rect 53668 111178 53696 123558
rect 53748 123276 53800 123282
rect 53748 123218 53800 123224
rect 53760 116618 53788 123218
rect 53852 117638 53880 142122
rect 53932 118040 53984 118046
rect 53932 117982 53984 117988
rect 53840 117632 53892 117638
rect 53840 117574 53892 117580
rect 53748 116612 53800 116618
rect 53748 116554 53800 116560
rect 53748 111240 53800 111246
rect 53748 111182 53800 111188
rect 53656 111172 53708 111178
rect 53656 111114 53708 111120
rect 53380 104780 53432 104786
rect 53380 104722 53432 104728
rect 53760 103514 53788 111182
rect 53760 103486 53880 103514
rect 53288 102196 53340 102202
rect 53288 102138 53340 102144
rect 53196 95124 53248 95130
rect 53196 95066 53248 95072
rect 53300 68882 53328 102138
rect 53852 96626 53880 103486
rect 53944 102202 53972 117982
rect 53932 102196 53984 102202
rect 53932 102138 53984 102144
rect 53380 96620 53432 96626
rect 53380 96562 53432 96568
rect 53840 96620 53892 96626
rect 53840 96562 53892 96568
rect 53288 68876 53340 68882
rect 53288 68818 53340 68824
rect 53392 19106 53420 96562
rect 54220 29714 54248 192578
rect 54392 150204 54444 150210
rect 54392 150146 54444 150152
rect 54404 117706 54432 150146
rect 54392 117700 54444 117706
rect 54392 117642 54444 117648
rect 54208 29708 54260 29714
rect 54208 29650 54260 29656
rect 53654 25528 53710 25537
rect 53654 25463 53710 25472
rect 53668 24886 53696 25463
rect 53656 24880 53708 24886
rect 53656 24822 53708 24828
rect 54496 21962 54524 197406
rect 56138 195528 56194 195537
rect 54760 195492 54812 195498
rect 56138 195463 56194 195472
rect 54760 195434 54812 195440
rect 54668 183184 54720 183190
rect 54668 183126 54720 183132
rect 54576 177608 54628 177614
rect 54576 177550 54628 177556
rect 54588 140690 54616 177550
rect 54576 140684 54628 140690
rect 54576 140626 54628 140632
rect 54576 137284 54628 137290
rect 54576 137226 54628 137232
rect 54588 123282 54616 137226
rect 54680 126954 54708 183126
rect 54668 126948 54720 126954
rect 54668 126890 54720 126896
rect 54576 123276 54628 123282
rect 54576 123218 54628 123224
rect 54666 122088 54722 122097
rect 54666 122023 54722 122032
rect 54576 119468 54628 119474
rect 54576 119410 54628 119416
rect 54588 112470 54616 119410
rect 54576 112464 54628 112470
rect 54576 112406 54628 112412
rect 54576 95124 54628 95130
rect 54576 95066 54628 95072
rect 54484 21956 54536 21962
rect 54484 21898 54536 21904
rect 54588 21554 54616 95066
rect 54680 83706 54708 122023
rect 54772 120018 54800 195434
rect 55588 195356 55640 195362
rect 55588 195298 55640 195304
rect 55036 190052 55088 190058
rect 55036 189994 55088 190000
rect 54944 181960 54996 181966
rect 54944 181902 54996 181908
rect 54852 166388 54904 166394
rect 54852 166330 54904 166336
rect 54760 120012 54812 120018
rect 54760 119954 54812 119960
rect 54760 111104 54812 111110
rect 54760 111046 54812 111052
rect 54668 83700 54720 83706
rect 54668 83642 54720 83648
rect 54576 21548 54628 21554
rect 54576 21490 54628 21496
rect 54772 19242 54800 111046
rect 54864 25566 54892 166330
rect 54852 25560 54904 25566
rect 54852 25502 54904 25508
rect 54956 25498 54984 181902
rect 55048 29753 55076 189994
rect 55128 146396 55180 146402
rect 55128 146338 55180 146344
rect 55140 143614 55168 146338
rect 55128 143608 55180 143614
rect 55128 143550 55180 143556
rect 55220 140820 55272 140826
rect 55220 140762 55272 140768
rect 55232 137290 55260 140762
rect 55220 137284 55272 137290
rect 55220 137226 55272 137232
rect 55128 126404 55180 126410
rect 55128 126346 55180 126352
rect 55140 120086 55168 126346
rect 55128 120080 55180 120086
rect 55128 120022 55180 120028
rect 55128 84244 55180 84250
rect 55128 84186 55180 84192
rect 55034 29744 55090 29753
rect 55034 29679 55090 29688
rect 54944 25492 54996 25498
rect 54944 25434 54996 25440
rect 55140 20262 55168 84186
rect 55600 45354 55628 195298
rect 55956 190256 56008 190262
rect 55956 190198 56008 190204
rect 55864 185632 55916 185638
rect 55864 185574 55916 185580
rect 55680 174820 55732 174826
rect 55680 174762 55732 174768
rect 55692 142186 55720 174762
rect 55770 151192 55826 151201
rect 55770 151127 55826 151136
rect 55680 142180 55732 142186
rect 55680 142122 55732 142128
rect 55784 109002 55812 151127
rect 55772 108996 55824 109002
rect 55772 108938 55824 108944
rect 55876 98161 55904 185574
rect 55862 98152 55918 98161
rect 55862 98087 55918 98096
rect 55864 97912 55916 97918
rect 55864 97854 55916 97860
rect 55772 75812 55824 75818
rect 55772 75754 55824 75760
rect 55588 45348 55640 45354
rect 55588 45290 55640 45296
rect 55128 20256 55180 20262
rect 55128 20198 55180 20204
rect 55784 20194 55812 75754
rect 55772 20188 55824 20194
rect 55772 20130 55824 20136
rect 55876 19922 55904 97854
rect 55968 77081 55996 190198
rect 56048 155712 56100 155718
rect 56048 155654 56100 155660
rect 55954 77072 56010 77081
rect 55954 77007 56010 77016
rect 55956 68876 56008 68882
rect 55956 68818 56008 68824
rect 55864 19916 55916 19922
rect 55864 19858 55916 19864
rect 54760 19236 54812 19242
rect 54760 19178 54812 19184
rect 53380 19100 53432 19106
rect 53380 19042 53432 19048
rect 55968 18494 55996 68818
rect 56060 41721 56088 155654
rect 56152 70281 56180 195463
rect 58360 190454 58388 200124
rect 58624 198416 58676 198422
rect 58624 198358 58676 198364
rect 57992 190426 58388 190454
rect 56322 184376 56378 184385
rect 56322 184311 56378 184320
rect 56230 149016 56286 149025
rect 56230 148951 56286 148960
rect 56138 70272 56194 70281
rect 56138 70207 56194 70216
rect 56046 41712 56102 41721
rect 56046 41647 56102 41656
rect 56244 21690 56272 148951
rect 56336 54641 56364 184311
rect 56416 170536 56468 170542
rect 56416 170478 56468 170484
rect 56322 54632 56378 54641
rect 56322 54567 56378 54576
rect 56428 32201 56456 170478
rect 57888 170400 57940 170406
rect 57888 170342 57940 170348
rect 56784 160948 56836 160954
rect 56784 160890 56836 160896
rect 56600 153060 56652 153066
rect 56600 153002 56652 153008
rect 56612 125118 56640 153002
rect 56692 142112 56744 142118
rect 56692 142054 56744 142060
rect 56704 141681 56732 142054
rect 56690 141672 56746 141681
rect 56690 141607 56746 141616
rect 56692 140752 56744 140758
rect 56692 140694 56744 140700
rect 56704 140321 56732 140694
rect 56690 140312 56746 140321
rect 56690 140247 56746 140256
rect 56692 128852 56744 128858
rect 56692 128794 56744 128800
rect 56704 126410 56732 128794
rect 56692 126404 56744 126410
rect 56692 126346 56744 126352
rect 56690 125352 56746 125361
rect 56690 125287 56746 125296
rect 56600 125112 56652 125118
rect 56600 125054 56652 125060
rect 56704 124982 56732 125287
rect 56692 124976 56744 124982
rect 56692 124918 56744 124924
rect 56692 120080 56744 120086
rect 56692 120022 56744 120028
rect 56704 111110 56732 120022
rect 56692 111104 56744 111110
rect 56692 111046 56744 111052
rect 56600 108996 56652 109002
rect 56600 108938 56652 108944
rect 56612 107681 56640 108938
rect 56598 107672 56654 107681
rect 56598 107607 56654 107616
rect 56796 56001 56824 160890
rect 56874 159624 56930 159633
rect 56874 159559 56930 159568
rect 56888 113121 56916 159559
rect 57794 159352 57850 159361
rect 57794 159287 57850 159296
rect 56966 158536 57022 158545
rect 56966 158471 57022 158480
rect 56980 119921 57008 158471
rect 57612 155576 57664 155582
rect 57612 155518 57664 155524
rect 57518 154048 57574 154057
rect 57518 153983 57574 153992
rect 57336 150068 57388 150074
rect 57336 150010 57388 150016
rect 57244 140684 57296 140690
rect 57244 140626 57296 140632
rect 57256 139641 57284 140626
rect 57242 139632 57298 139641
rect 57242 139567 57298 139576
rect 57152 124636 57204 124642
rect 57152 124578 57204 124584
rect 56966 119912 57022 119921
rect 56966 119847 57022 119856
rect 56966 118008 57022 118017
rect 56966 117943 57022 117952
rect 56980 113174 57008 117943
rect 57060 117292 57112 117298
rect 57060 117234 57112 117240
rect 57072 117201 57100 117234
rect 57058 117192 57114 117201
rect 57058 117127 57114 117136
rect 56980 113146 57100 113174
rect 56874 113112 56930 113121
rect 56874 113047 56930 113056
rect 56876 104780 56928 104786
rect 56876 104722 56928 104728
rect 56888 104281 56916 104722
rect 56874 104272 56930 104281
rect 56874 104207 56930 104216
rect 57072 84250 57100 113146
rect 57164 90681 57192 124578
rect 57348 120222 57376 150010
rect 57428 145036 57480 145042
rect 57428 144978 57480 144984
rect 57440 121582 57468 144978
rect 57428 121576 57480 121582
rect 57428 121518 57480 121524
rect 57428 121440 57480 121446
rect 57428 121382 57480 121388
rect 57440 120601 57468 121382
rect 57426 120592 57482 120601
rect 57426 120527 57482 120536
rect 57336 120216 57388 120222
rect 57336 120158 57388 120164
rect 57428 120012 57480 120018
rect 57428 119954 57480 119960
rect 57440 119241 57468 119954
rect 57426 119232 57482 119241
rect 57426 119167 57482 119176
rect 57428 115932 57480 115938
rect 57428 115874 57480 115880
rect 57440 115161 57468 115874
rect 57426 115152 57482 115161
rect 57426 115087 57482 115096
rect 57428 114504 57480 114510
rect 57426 114472 57428 114481
rect 57480 114472 57482 114481
rect 57426 114407 57482 114416
rect 57244 112464 57296 112470
rect 57244 112406 57296 112412
rect 57150 90672 57206 90681
rect 57150 90607 57206 90616
rect 57060 84244 57112 84250
rect 57060 84186 57112 84192
rect 57152 84176 57204 84182
rect 57152 84118 57204 84124
rect 57164 75818 57192 84118
rect 57152 75812 57204 75818
rect 57152 75754 57204 75760
rect 57060 69692 57112 69698
rect 57060 69634 57112 69640
rect 57072 64874 57100 69634
rect 57152 68944 57204 68950
rect 57152 68886 57204 68892
rect 57164 68241 57192 68886
rect 57150 68232 57206 68241
rect 57150 68167 57206 68176
rect 57072 64846 57192 64874
rect 57060 60036 57112 60042
rect 57060 59978 57112 59984
rect 56782 55992 56838 56001
rect 56782 55927 56838 55936
rect 57072 46481 57100 59978
rect 57164 47161 57192 64846
rect 57150 47152 57206 47161
rect 57150 47087 57206 47096
rect 57058 46472 57114 46481
rect 57058 46407 57114 46416
rect 57152 45348 57204 45354
rect 57152 45290 57204 45296
rect 57164 45121 57192 45290
rect 57150 45112 57206 45121
rect 57150 45047 57206 45056
rect 56692 41336 56744 41342
rect 56692 41278 56744 41284
rect 56704 41041 56732 41278
rect 56690 41032 56746 41041
rect 56690 40967 56746 40976
rect 56414 32192 56470 32201
rect 56414 32127 56470 32136
rect 56232 21684 56284 21690
rect 56232 21626 56284 21632
rect 57256 19281 57284 112406
rect 57336 110424 57388 110430
rect 57532 110401 57560 153983
rect 57624 143585 57652 155518
rect 57704 155440 57756 155446
rect 57704 155382 57756 155388
rect 57610 143576 57666 143585
rect 57610 143511 57666 143520
rect 57612 137964 57664 137970
rect 57612 137906 57664 137912
rect 57624 137601 57652 137906
rect 57610 137592 57666 137601
rect 57610 137527 57666 137536
rect 57612 135244 57664 135250
rect 57612 135186 57664 135192
rect 57624 134881 57652 135186
rect 57610 134872 57666 134881
rect 57610 134807 57666 134816
rect 57612 133884 57664 133890
rect 57612 133826 57664 133832
rect 57624 132841 57652 133826
rect 57610 132832 57666 132841
rect 57610 132767 57666 132776
rect 57612 132456 57664 132462
rect 57612 132398 57664 132404
rect 57624 131481 57652 132398
rect 57610 131472 57666 131481
rect 57610 131407 57666 131416
rect 57612 131096 57664 131102
rect 57612 131038 57664 131044
rect 57624 130801 57652 131038
rect 57610 130792 57666 130801
rect 57610 130727 57666 130736
rect 57612 129736 57664 129742
rect 57612 129678 57664 129684
rect 57624 129441 57652 129678
rect 57610 129432 57666 129441
rect 57610 129367 57666 129376
rect 57612 128308 57664 128314
rect 57612 128250 57664 128256
rect 57624 128081 57652 128250
rect 57610 128072 57666 128081
rect 57610 128007 57666 128016
rect 57612 126948 57664 126954
rect 57612 126890 57664 126896
rect 57624 126721 57652 126890
rect 57610 126712 57666 126721
rect 57610 126647 57666 126656
rect 57612 124160 57664 124166
rect 57612 124102 57664 124108
rect 57624 123321 57652 124102
rect 57610 123312 57666 123321
rect 57610 123247 57666 123256
rect 57612 123208 57664 123214
rect 57612 123150 57664 123156
rect 57336 110366 57388 110372
rect 57518 110392 57574 110401
rect 57242 19272 57298 19281
rect 57242 19207 57298 19216
rect 55956 18488 56008 18494
rect 55956 18430 56008 18436
rect 57348 17406 57376 110366
rect 57518 110327 57574 110336
rect 57520 108928 57572 108934
rect 57520 108870 57572 108876
rect 57428 108860 57480 108866
rect 57428 108802 57480 108808
rect 57440 18834 57468 108802
rect 57532 108361 57560 108870
rect 57518 108352 57574 108361
rect 57518 108287 57574 108296
rect 57520 104848 57572 104854
rect 57520 104790 57572 104796
rect 57532 103601 57560 104790
rect 57518 103592 57574 103601
rect 57518 103527 57574 103536
rect 57520 103488 57572 103494
rect 57520 103430 57572 103436
rect 57532 102921 57560 103430
rect 57518 102912 57574 102921
rect 57518 102847 57574 102856
rect 57520 102128 57572 102134
rect 57520 102070 57572 102076
rect 57532 101561 57560 102070
rect 57518 101552 57574 101561
rect 57518 101487 57574 101496
rect 57520 100700 57572 100706
rect 57520 100642 57572 100648
rect 57532 99521 57560 100642
rect 57518 99512 57574 99521
rect 57518 99447 57574 99456
rect 57520 95192 57572 95198
rect 57520 95134 57572 95140
rect 57532 94081 57560 95134
rect 57518 94072 57574 94081
rect 57518 94007 57574 94016
rect 57520 93832 57572 93838
rect 57520 93774 57572 93780
rect 57532 92721 57560 93774
rect 57518 92712 57574 92721
rect 57518 92647 57574 92656
rect 57624 89842 57652 123150
rect 57532 89814 57652 89842
rect 57532 85474 57560 89814
rect 57612 89684 57664 89690
rect 57612 89626 57664 89632
rect 57624 89321 57652 89626
rect 57610 89312 57666 89321
rect 57610 89247 57666 89256
rect 57612 86964 57664 86970
rect 57612 86906 57664 86912
rect 57624 86601 57652 86906
rect 57610 86592 57666 86601
rect 57610 86527 57666 86536
rect 57520 85468 57572 85474
rect 57520 85410 57572 85416
rect 57716 83858 57744 155382
rect 57808 143041 57836 159287
rect 57900 145761 57928 170342
rect 57992 152454 58020 190426
rect 58256 185972 58308 185978
rect 58256 185914 58308 185920
rect 57980 152448 58032 152454
rect 57980 152390 58032 152396
rect 58164 152448 58216 152454
rect 58164 152390 58216 152396
rect 57886 145752 57942 145761
rect 57886 145687 57942 145696
rect 57794 143032 57850 143041
rect 57794 142967 57850 142976
rect 57796 142112 57848 142118
rect 57796 142054 57848 142060
rect 57808 132494 57836 142054
rect 57980 135924 58032 135930
rect 57980 135866 58032 135872
rect 57808 132466 57928 132494
rect 57796 126948 57848 126954
rect 57796 126890 57848 126896
rect 57808 123214 57836 126890
rect 57900 123486 57928 132466
rect 57992 123622 58020 135866
rect 58070 124128 58126 124137
rect 58070 124063 58126 124072
rect 57980 123616 58032 123622
rect 57980 123558 58032 123564
rect 57888 123480 57940 123486
rect 57888 123422 57940 123428
rect 57796 123208 57848 123214
rect 57796 123150 57848 123156
rect 57888 121440 57940 121446
rect 57888 121382 57940 121388
rect 57796 120148 57848 120154
rect 57796 120090 57848 120096
rect 57808 83978 57836 120090
rect 57900 117094 57928 121382
rect 57888 117088 57940 117094
rect 57888 117030 57940 117036
rect 57980 116612 58032 116618
rect 57980 116554 58032 116560
rect 57888 103420 57940 103426
rect 57888 103362 57940 103368
rect 57900 102241 57928 103362
rect 57886 102232 57942 102241
rect 57886 102167 57942 102176
rect 57796 83972 57848 83978
rect 57796 83914 57848 83920
rect 57716 83830 57928 83858
rect 57796 83768 57848 83774
rect 57796 83710 57848 83716
rect 57704 83700 57756 83706
rect 57704 83642 57756 83648
rect 57612 82816 57664 82822
rect 57612 82758 57664 82764
rect 57520 82748 57572 82754
rect 57520 82690 57572 82696
rect 57532 81841 57560 82690
rect 57624 82521 57652 82758
rect 57610 82512 57666 82521
rect 57610 82447 57666 82456
rect 57518 81832 57574 81841
rect 57518 81767 57574 81776
rect 57716 81682 57744 83642
rect 57532 81654 57744 81682
rect 57532 21729 57560 81654
rect 57704 79348 57756 79354
rect 57704 79290 57756 79296
rect 57612 75880 57664 75886
rect 57612 75822 57664 75828
rect 57624 75721 57652 75822
rect 57610 75712 57666 75721
rect 57610 75647 57666 75656
rect 57612 75608 57664 75614
rect 57612 75550 57664 75556
rect 57518 21720 57574 21729
rect 57518 21655 57574 21664
rect 57624 21282 57652 75550
rect 57612 21276 57664 21282
rect 57612 21218 57664 21224
rect 57428 18828 57480 18834
rect 57428 18770 57480 18776
rect 57716 17542 57744 79290
rect 57808 19854 57836 83710
rect 57900 81161 57928 83830
rect 57886 81152 57942 81161
rect 57886 81087 57942 81096
rect 57888 79416 57940 79422
rect 57888 79358 57940 79364
rect 57900 75614 57928 79358
rect 57992 79354 58020 116554
rect 57980 79348 58032 79354
rect 57980 79290 58032 79296
rect 57888 75608 57940 75614
rect 57888 75550 57940 75556
rect 57888 69012 57940 69018
rect 57888 68954 57940 68960
rect 57900 68921 57928 68954
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57888 67584 57940 67590
rect 57886 67552 57888 67561
rect 57940 67552 57942 67561
rect 57886 67487 57942 67496
rect 57888 64864 57940 64870
rect 57888 64806 57940 64812
rect 57900 64161 57928 64806
rect 57886 64152 57942 64161
rect 57886 64087 57942 64096
rect 57888 63504 57940 63510
rect 57886 63472 57888 63481
rect 57940 63472 57942 63481
rect 57886 63407 57942 63416
rect 57886 62112 57942 62121
rect 57886 62047 57888 62056
rect 57940 62047 57942 62056
rect 57888 62018 57940 62024
rect 57888 59356 57940 59362
rect 57888 59298 57940 59304
rect 57900 58721 57928 59298
rect 57886 58712 57942 58721
rect 57886 58647 57942 58656
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57900 57361 57928 57870
rect 57886 57352 57942 57361
rect 57886 57287 57942 57296
rect 57888 56568 57940 56574
rect 57888 56510 57940 56516
rect 57900 55321 57928 56510
rect 57886 55312 57942 55321
rect 57886 55247 57942 55256
rect 57888 49020 57940 49026
rect 57888 48962 57940 48968
rect 57900 41562 57928 48962
rect 57900 41534 58020 41562
rect 57888 41404 57940 41410
rect 57888 41346 57940 41352
rect 57900 40361 57928 41346
rect 57886 40352 57942 40361
rect 57886 40287 57942 40296
rect 57992 40202 58020 41534
rect 57900 40174 58020 40202
rect 57900 39681 57928 40174
rect 57886 39672 57942 39681
rect 57886 39607 57942 39616
rect 57888 34468 57940 34474
rect 57888 34410 57940 34416
rect 57900 33561 57928 34410
rect 57886 33552 57942 33561
rect 57886 33487 57942 33496
rect 57888 33040 57940 33046
rect 57888 32982 57940 32988
rect 57900 32881 57928 32982
rect 57886 32872 57942 32881
rect 57886 32807 57942 32816
rect 57796 19848 57848 19854
rect 57796 19790 57848 19796
rect 58084 17678 58112 124063
rect 58176 45801 58204 152390
rect 58268 115841 58296 185914
rect 58532 146328 58584 146334
rect 58532 146270 58584 146276
rect 58440 146124 58492 146130
rect 58440 146066 58492 146072
rect 58452 135250 58480 146066
rect 58440 135244 58492 135250
rect 58440 135186 58492 135192
rect 58544 128858 58572 146270
rect 58532 128852 58584 128858
rect 58532 128794 58584 128800
rect 58348 127628 58400 127634
rect 58348 127570 58400 127576
rect 58254 115832 58310 115841
rect 58254 115767 58310 115776
rect 58256 85536 58308 85542
rect 58256 85478 58308 85484
rect 58268 84182 58296 85478
rect 58256 84176 58308 84182
rect 58256 84118 58308 84124
rect 58162 45792 58218 45801
rect 58162 45727 58218 45736
rect 58360 20126 58388 127570
rect 58636 124642 58664 198358
rect 59004 197169 59032 200124
rect 58990 197160 59046 197169
rect 58990 197095 59046 197104
rect 60292 195809 60320 200124
rect 60278 195800 60334 195809
rect 60278 195735 60334 195744
rect 58808 190324 58860 190330
rect 58808 190266 58860 190272
rect 58716 187468 58768 187474
rect 58716 187410 58768 187416
rect 58728 136542 58756 187410
rect 58716 136536 58768 136542
rect 58716 136478 58768 136484
rect 58716 134428 58768 134434
rect 58716 134370 58768 134376
rect 58728 126954 58756 134370
rect 58716 126948 58768 126954
rect 58716 126890 58768 126896
rect 58716 125316 58768 125322
rect 58716 125258 58768 125264
rect 58624 124636 58676 124642
rect 58624 124578 58676 124584
rect 58624 123548 58676 123554
rect 58624 123490 58676 123496
rect 58440 98660 58492 98666
rect 58440 98602 58492 98608
rect 58452 85542 58480 98602
rect 58440 85536 58492 85542
rect 58440 85478 58492 85484
rect 58532 85468 58584 85474
rect 58532 85410 58584 85416
rect 58544 22098 58572 85410
rect 58636 26858 58664 123490
rect 58728 98682 58756 125258
rect 58820 100162 58848 190266
rect 59452 189644 59504 189650
rect 59452 189586 59504 189592
rect 59084 184408 59136 184414
rect 59084 184350 59136 184356
rect 58900 182096 58952 182102
rect 58900 182038 58952 182044
rect 58912 143698 58940 182038
rect 58992 150952 59044 150958
rect 58992 150894 59044 150900
rect 59004 143834 59032 150894
rect 59096 144945 59124 184350
rect 59360 156664 59412 156670
rect 59360 156606 59412 156612
rect 59268 150000 59320 150006
rect 59268 149942 59320 149948
rect 59082 144936 59138 144945
rect 59280 144922 59308 149942
rect 59372 145042 59400 156606
rect 59464 151745 59492 189586
rect 59728 187332 59780 187338
rect 59728 187274 59780 187280
rect 59636 184476 59688 184482
rect 59636 184418 59688 184424
rect 59544 174956 59596 174962
rect 59544 174898 59596 174904
rect 59450 151736 59506 151745
rect 59450 151671 59506 151680
rect 59452 151632 59504 151638
rect 59452 151574 59504 151580
rect 59464 146334 59492 151574
rect 59556 150210 59584 174898
rect 59648 156670 59676 184418
rect 59636 156664 59688 156670
rect 59636 156606 59688 156612
rect 59634 151736 59690 151745
rect 59634 151671 59690 151680
rect 59544 150204 59596 150210
rect 59544 150146 59596 150152
rect 59542 150104 59598 150113
rect 59542 150039 59598 150048
rect 59556 146402 59584 150039
rect 59648 147665 59676 151671
rect 59740 151473 59768 187274
rect 59820 184544 59872 184550
rect 59820 184486 59872 184492
rect 59726 151464 59782 151473
rect 59726 151399 59782 151408
rect 59726 151328 59782 151337
rect 59726 151263 59782 151272
rect 59740 149025 59768 151263
rect 59726 149016 59782 149025
rect 59726 148951 59782 148960
rect 59634 147656 59690 147665
rect 59634 147591 59690 147600
rect 59544 146396 59596 146402
rect 59544 146338 59596 146344
rect 59452 146328 59504 146334
rect 59452 146270 59504 146276
rect 59360 145036 59412 145042
rect 59360 144978 59412 144984
rect 59280 144894 59400 144922
rect 59082 144871 59138 144880
rect 59004 143806 59216 143834
rect 58912 143670 59124 143698
rect 58898 143576 58954 143585
rect 58898 143511 58954 143520
rect 58912 136649 58940 143511
rect 59096 142118 59124 143670
rect 59084 142112 59136 142118
rect 59084 142054 59136 142060
rect 59188 138014 59216 143806
rect 59372 142066 59400 144894
rect 59280 142038 59400 142066
rect 59280 139346 59308 142038
rect 59280 139318 59400 139346
rect 59266 139224 59322 139233
rect 59266 139159 59322 139168
rect 59004 137986 59216 138014
rect 58898 136640 58954 136649
rect 58898 136575 58954 136584
rect 58900 136536 58952 136542
rect 58900 136478 58952 136484
rect 58912 121446 58940 136478
rect 58900 121440 58952 121446
rect 58900 121382 58952 121388
rect 58898 111888 58954 111897
rect 58898 111823 58954 111832
rect 58808 100156 58860 100162
rect 58808 100098 58860 100104
rect 58728 98654 58848 98682
rect 58716 98592 58768 98598
rect 58716 98534 58768 98540
rect 58624 26852 58676 26858
rect 58624 26794 58676 26800
rect 58728 25838 58756 98534
rect 58716 25832 58768 25838
rect 58716 25774 58768 25780
rect 58532 22092 58584 22098
rect 58532 22034 58584 22040
rect 58348 20120 58400 20126
rect 58348 20062 58400 20068
rect 58072 17672 58124 17678
rect 58072 17614 58124 17620
rect 57704 17536 57756 17542
rect 57704 17478 57756 17484
rect 57336 17400 57388 17406
rect 57336 17342 57388 17348
rect 58820 16454 58848 98654
rect 58912 20670 58940 111823
rect 59004 53281 59032 137986
rect 59082 137320 59138 137329
rect 59082 137255 59138 137264
rect 59096 124166 59124 137255
rect 59280 136762 59308 139159
rect 59372 137306 59400 139318
rect 59372 137278 59492 137306
rect 59280 136734 59400 136762
rect 59372 135402 59400 136734
rect 59280 135374 59400 135402
rect 59280 134434 59308 135374
rect 59360 135244 59412 135250
rect 59360 135186 59412 135192
rect 59268 134428 59320 134434
rect 59268 134370 59320 134376
rect 59372 127634 59400 135186
rect 59360 127628 59412 127634
rect 59360 127570 59412 127576
rect 59266 125488 59322 125497
rect 59266 125423 59322 125432
rect 59084 124160 59136 124166
rect 59084 124102 59136 124108
rect 59280 120193 59308 125423
rect 59464 125322 59492 137278
rect 59452 125316 59504 125322
rect 59452 125258 59504 125264
rect 59360 124160 59412 124166
rect 59360 124102 59412 124108
rect 59266 120184 59322 120193
rect 59266 120119 59322 120128
rect 59372 120068 59400 124102
rect 59452 121372 59504 121378
rect 59452 121314 59504 121320
rect 59280 120040 59400 120068
rect 59280 117298 59308 120040
rect 59464 120000 59492 121314
rect 59636 120216 59688 120222
rect 59636 120158 59688 120164
rect 59372 119972 59492 120000
rect 59268 117292 59320 117298
rect 59268 117234 59320 117240
rect 59268 117020 59320 117026
rect 59268 116962 59320 116968
rect 59084 100156 59136 100162
rect 59084 100098 59136 100104
rect 59096 96801 59124 100098
rect 59280 98734 59308 116962
rect 59372 111246 59400 119972
rect 59544 117292 59596 117298
rect 59544 117234 59596 117240
rect 59452 117088 59504 117094
rect 59452 117030 59504 117036
rect 59360 111240 59412 111246
rect 59360 111182 59412 111188
rect 59268 98728 59320 98734
rect 59268 98670 59320 98676
rect 59464 98666 59492 117030
rect 59452 98660 59504 98666
rect 59452 98602 59504 98608
rect 59556 98598 59584 117234
rect 59648 117026 59676 120158
rect 59832 120154 59860 184486
rect 60936 180794 60964 200124
rect 61534 199866 61562 200124
rect 61534 199838 61608 199866
rect 61580 191350 61608 199838
rect 64156 198286 64184 200124
rect 67376 198490 67404 200124
rect 67364 198484 67416 198490
rect 67364 198426 67416 198432
rect 64144 198280 64196 198286
rect 64144 198222 64196 198228
rect 63500 197940 63552 197946
rect 63500 197882 63552 197888
rect 61568 191344 61620 191350
rect 61568 191286 61620 191292
rect 60752 180766 60964 180794
rect 59912 180192 59964 180198
rect 59912 180134 59964 180140
rect 59924 150142 59952 180134
rect 60002 151464 60058 151473
rect 60002 151399 60058 151408
rect 59912 150136 59964 150142
rect 60016 150113 60044 151399
rect 60752 150890 60780 180766
rect 61934 153096 61990 153105
rect 61934 153031 61990 153040
rect 61292 152312 61344 152318
rect 61292 152254 61344 152260
rect 60740 150884 60792 150890
rect 60740 150826 60792 150832
rect 59912 150078 59964 150084
rect 60002 150104 60058 150113
rect 60002 150039 60058 150048
rect 59910 149968 59966 149977
rect 61304 149940 61332 152254
rect 61948 149940 61976 153031
rect 63512 149954 63540 197882
rect 68020 186969 68048 200124
rect 68284 197396 68336 197402
rect 68284 197338 68336 197344
rect 68006 186960 68062 186969
rect 68006 186895 68062 186904
rect 65800 180260 65852 180266
rect 65800 180202 65852 180208
rect 64512 169108 64564 169114
rect 64512 169050 64564 169056
rect 63512 149926 63894 149954
rect 64524 149940 64552 169050
rect 65812 149940 65840 180202
rect 66444 170468 66496 170474
rect 66444 170410 66496 170416
rect 66456 149940 66484 170410
rect 67088 152516 67140 152522
rect 67088 152458 67140 152464
rect 67100 149940 67128 152458
rect 68296 152318 68324 197338
rect 69020 195152 69072 195158
rect 69020 195094 69072 195100
rect 68284 152312 68336 152318
rect 68284 152254 68336 152260
rect 68744 152244 68796 152250
rect 68744 152186 68796 152192
rect 68756 149954 68784 152186
rect 68418 149926 68784 149954
rect 69032 149940 69060 195094
rect 70596 180794 70624 200124
rect 71194 200002 71222 200124
rect 71148 199974 71222 200002
rect 71148 197402 71176 199974
rect 72528 197878 72556 200124
rect 72516 197872 72568 197878
rect 72516 197814 72568 197820
rect 71136 197396 71188 197402
rect 71136 197338 71188 197344
rect 73172 190454 73200 200124
rect 73816 197334 73844 200124
rect 73804 197328 73856 197334
rect 73804 197270 73856 197276
rect 74460 195242 74488 200124
rect 75702 200002 75730 200124
rect 75656 199974 75730 200002
rect 75460 199708 75512 199714
rect 75460 199650 75512 199656
rect 73356 195214 74488 195242
rect 73172 190426 73292 190454
rect 70504 180766 70624 180794
rect 69664 180328 69716 180334
rect 69664 180270 69716 180276
rect 69676 152250 69704 180270
rect 69664 152244 69716 152250
rect 69664 152186 69716 152192
rect 70504 151026 70532 180766
rect 73264 154086 73292 190426
rect 73356 177313 73384 195214
rect 73528 195084 73580 195090
rect 73528 195026 73580 195032
rect 73342 177304 73398 177313
rect 73342 177239 73398 177248
rect 73252 154080 73304 154086
rect 73252 154022 73304 154028
rect 72882 152416 72938 152425
rect 72882 152351 72938 152360
rect 70492 151020 70544 151026
rect 70492 150962 70544 150968
rect 72896 149940 72924 152351
rect 73540 149940 73568 195026
rect 74816 177744 74868 177750
rect 74816 177686 74868 177692
rect 74828 149940 74856 177686
rect 75472 149940 75500 199650
rect 75656 196654 75684 199974
rect 75644 196648 75696 196654
rect 75644 196590 75696 196596
rect 77036 180794 77064 200124
rect 77680 198422 77708 200124
rect 77668 198416 77720 198422
rect 77668 198358 77720 198364
rect 78324 180794 78352 200124
rect 78680 195152 78732 195158
rect 78680 195094 78732 195100
rect 75932 180766 77064 180794
rect 77404 180766 78352 180794
rect 75932 151162 75960 180766
rect 77404 180033 77432 180766
rect 77390 180024 77446 180033
rect 77390 179959 77446 179968
rect 78036 169244 78088 169250
rect 78036 169186 78088 169192
rect 77390 167648 77446 167657
rect 77390 167583 77446 167592
rect 76748 152380 76800 152386
rect 76748 152322 76800 152328
rect 75920 151156 75972 151162
rect 75920 151098 75972 151104
rect 76760 149940 76788 152322
rect 77404 149940 77432 167583
rect 78048 149940 78076 169186
rect 78692 150958 78720 195094
rect 78968 180794 78996 200124
rect 79612 195158 79640 200124
rect 80152 196648 80204 196654
rect 80152 196590 80204 196596
rect 79600 195152 79652 195158
rect 79600 195094 79652 195100
rect 80060 195152 80112 195158
rect 80060 195094 80112 195100
rect 78784 180766 78996 180794
rect 78784 156738 78812 180766
rect 79324 171896 79376 171902
rect 79324 171838 79376 171844
rect 78772 156732 78824 156738
rect 78772 156674 78824 156680
rect 78680 150952 78732 150958
rect 78680 150894 78732 150900
rect 79336 149940 79364 171838
rect 80072 151162 80100 195094
rect 80060 151156 80112 151162
rect 80060 151098 80112 151104
rect 80164 149954 80192 196590
rect 80256 156806 80284 200124
rect 80854 200002 80882 200124
rect 80808 199974 80882 200002
rect 80808 195158 80836 199974
rect 82188 196994 82216 200124
rect 82832 198393 82860 200124
rect 83476 198801 83504 200124
rect 84120 199034 84148 200124
rect 85362 200002 85390 200124
rect 85316 199974 85390 200002
rect 84108 199028 84160 199034
rect 84108 198970 84160 198976
rect 83462 198792 83518 198801
rect 83462 198727 83518 198736
rect 82818 198384 82874 198393
rect 82818 198319 82874 198328
rect 82176 196988 82228 196994
rect 82176 196930 82228 196936
rect 80796 195152 80848 195158
rect 80796 195094 80848 195100
rect 85316 192302 85344 199974
rect 86696 197810 86724 200124
rect 88628 198506 88656 200124
rect 88444 198478 88656 198506
rect 86684 197804 86736 197810
rect 86684 197746 86736 197752
rect 86408 195560 86460 195566
rect 86408 195502 86460 195508
rect 85304 192296 85356 192302
rect 85304 192238 85356 192244
rect 85764 189916 85816 189922
rect 85764 189858 85816 189864
rect 84200 166592 84252 166598
rect 84200 166534 84252 166540
rect 81900 165096 81952 165102
rect 81900 165038 81952 165044
rect 80244 156800 80296 156806
rect 80244 156742 80296 156748
rect 81256 152516 81308 152522
rect 81256 152458 81308 152464
rect 80164 149926 80638 149954
rect 81268 149940 81296 152458
rect 81912 149940 81940 165038
rect 82544 152720 82596 152726
rect 82544 152662 82596 152668
rect 82556 149940 82584 152662
rect 84212 149954 84240 166534
rect 84212 149926 85146 149954
rect 85776 149940 85804 189858
rect 86420 149940 86448 195502
rect 87696 192976 87748 192982
rect 87696 192918 87748 192924
rect 87708 149940 87736 192918
rect 88444 173194 88472 198478
rect 88616 198348 88668 198354
rect 88616 198290 88668 198296
rect 88628 180794 88656 198290
rect 89272 197266 89300 200124
rect 89870 200002 89898 200124
rect 89824 199974 89898 200002
rect 89260 197260 89312 197266
rect 89260 197202 89312 197208
rect 88536 180766 88656 180794
rect 88432 173188 88484 173194
rect 88432 173130 88484 173136
rect 88536 149954 88564 180766
rect 89824 177546 89852 199974
rect 90916 199640 90968 199646
rect 90916 199582 90968 199588
rect 89812 177540 89864 177546
rect 89812 177482 89864 177488
rect 88536 149926 89010 149954
rect 90928 149940 90956 199582
rect 91204 180794 91232 200124
rect 92492 190454 92520 200124
rect 92664 199572 92716 199578
rect 92664 199514 92716 199520
rect 92492 190426 92612 190454
rect 91112 180766 91232 180794
rect 91112 154018 91140 180766
rect 92584 158506 92612 190426
rect 92572 158500 92624 158506
rect 92572 158442 92624 158448
rect 91100 154012 91152 154018
rect 91100 153954 91152 153960
rect 92676 149954 92704 199514
rect 93136 197985 93164 200124
rect 94424 198393 94452 200124
rect 94410 198384 94466 198393
rect 94410 198319 94466 198328
rect 93122 197976 93178 197985
rect 93122 197911 93178 197920
rect 96356 180794 96384 200124
rect 97000 195242 97028 200124
rect 95252 180766 96384 180794
rect 96632 195214 97028 195242
rect 95252 176050 95280 180766
rect 95240 176044 95292 176050
rect 95240 175986 95292 175992
rect 94780 152380 94832 152386
rect 94780 152322 94832 152328
rect 92676 149926 93518 149954
rect 94792 149940 94820 152322
rect 96632 151774 96660 195214
rect 97644 180794 97672 200124
rect 100864 198762 100892 200124
rect 100852 198756 100904 198762
rect 100852 198698 100904 198704
rect 101508 198626 101536 200124
rect 101496 198620 101548 198626
rect 101496 198562 101548 198568
rect 102152 194138 102180 200124
rect 104084 199646 104112 200124
rect 104682 200002 104710 200124
rect 104636 199974 104710 200002
rect 104072 199640 104124 199646
rect 104072 199582 104124 199588
rect 104636 199102 104664 199974
rect 104716 199640 104768 199646
rect 104716 199582 104768 199588
rect 104728 199102 104756 199582
rect 106016 199306 106044 200124
rect 106004 199300 106056 199306
rect 106004 199242 106056 199248
rect 104624 199096 104676 199102
rect 104624 199038 104676 199044
rect 104716 199096 104768 199102
rect 104716 199038 104768 199044
rect 102140 194132 102192 194138
rect 102140 194074 102192 194080
rect 98644 191276 98696 191282
rect 98644 191218 98696 191224
rect 96724 180766 97672 180794
rect 96724 172038 96752 180766
rect 96712 172032 96764 172038
rect 96712 171974 96764 171980
rect 96712 159724 96764 159730
rect 96712 159666 96764 159672
rect 96620 151768 96672 151774
rect 96620 151710 96672 151716
rect 96724 149954 96752 159666
rect 96724 149926 97382 149954
rect 98656 149940 98684 191218
rect 99932 187536 99984 187542
rect 99932 187478 99984 187484
rect 99288 177540 99340 177546
rect 99288 177482 99340 177488
rect 99300 149940 99328 177482
rect 99944 149940 99972 187478
rect 106660 180794 106688 200124
rect 108592 197402 108620 200124
rect 108948 199504 109000 199510
rect 108948 199446 109000 199452
rect 108580 197396 108632 197402
rect 108580 197338 108632 197344
rect 106292 180766 106688 180794
rect 103796 180260 103848 180266
rect 103796 180202 103848 180208
rect 103808 149940 103836 180202
rect 106292 154154 106320 180766
rect 108302 180704 108358 180713
rect 108302 180639 108358 180648
rect 106280 154148 106332 154154
rect 106280 154090 106332 154096
rect 107660 152788 107712 152794
rect 107660 152730 107712 152736
rect 106372 152720 106424 152726
rect 106372 152662 106424 152668
rect 106384 149940 106412 152662
rect 107672 149940 107700 152730
rect 108316 149940 108344 180639
rect 108960 149940 108988 199446
rect 109684 197396 109736 197402
rect 109684 197338 109736 197344
rect 109696 155854 109724 197338
rect 111168 180794 111196 200124
rect 111812 195242 111840 200124
rect 111812 195214 111932 195242
rect 111800 195152 111852 195158
rect 111800 195094 111852 195100
rect 110432 180766 111196 180794
rect 110432 160857 110460 180766
rect 110880 163872 110932 163878
rect 110880 163814 110932 163820
rect 110418 160848 110474 160857
rect 110418 160783 110474 160792
rect 109684 155848 109736 155854
rect 109684 155790 109736 155796
rect 110892 149940 110920 163814
rect 111812 152454 111840 195094
rect 111904 153921 111932 195214
rect 112456 180794 112484 200124
rect 113100 195158 113128 200124
rect 113088 195152 113140 195158
rect 113088 195094 113140 195100
rect 113180 195152 113232 195158
rect 113180 195094 113232 195100
rect 111996 180766 112484 180794
rect 111996 179110 112024 180766
rect 111984 179104 112036 179110
rect 111984 179046 112036 179052
rect 112168 172100 112220 172106
rect 112168 172042 112220 172048
rect 111890 153912 111946 153921
rect 111890 153847 111946 153856
rect 111800 152448 111852 152454
rect 111800 152390 111852 152396
rect 112180 149940 112208 172042
rect 113192 151706 113220 195094
rect 113744 180794 113772 200124
rect 114342 200002 114370 200124
rect 114296 199974 114370 200002
rect 114296 195158 114324 199974
rect 114284 195152 114336 195158
rect 114284 195094 114336 195100
rect 116320 190454 116348 200124
rect 116964 195566 116992 200124
rect 116952 195560 117004 195566
rect 116952 195502 117004 195508
rect 113284 180766 113772 180794
rect 115952 190426 116348 190454
rect 113180 151700 113232 151706
rect 113180 151642 113232 151648
rect 113284 151570 113312 180766
rect 113364 176248 113416 176254
rect 113364 176190 113416 176196
rect 113272 151564 113324 151570
rect 113272 151506 113324 151512
rect 113376 149954 113404 176190
rect 115952 171970 115980 190426
rect 116676 186040 116728 186046
rect 116676 185982 116728 185988
rect 116032 182980 116084 182986
rect 116032 182922 116084 182928
rect 115940 171964 115992 171970
rect 115940 171906 115992 171912
rect 113376 149926 114126 149954
rect 116044 149940 116072 182922
rect 116688 149940 116716 185982
rect 118252 180794 118280 200124
rect 118850 199866 118878 200124
rect 118804 199838 118878 199866
rect 118804 199238 118832 199838
rect 118792 199232 118844 199238
rect 118792 199174 118844 199180
rect 120184 197033 120212 200124
rect 120170 197024 120226 197033
rect 120170 196959 120226 196968
rect 121472 195838 121500 200124
rect 122760 198257 122788 200124
rect 123358 199866 123386 200124
rect 123358 199838 123432 199866
rect 123404 198626 123432 199838
rect 123392 198620 123444 198626
rect 123392 198562 123444 198568
rect 122746 198248 122802 198257
rect 122746 198183 122802 198192
rect 121460 195832 121512 195838
rect 121460 195774 121512 195780
rect 124692 180794 124720 200124
rect 127268 199170 127296 200124
rect 127256 199164 127308 199170
rect 127256 199106 127308 199112
rect 125048 196512 125100 196518
rect 125048 196454 125100 196460
rect 117332 180766 118280 180794
rect 124324 180766 124720 180794
rect 117332 151337 117360 180766
rect 121460 159520 121512 159526
rect 121460 159462 121512 159468
rect 121472 152386 121500 159462
rect 124324 156670 124352 180766
rect 124404 169448 124456 169454
rect 124404 169390 124456 169396
rect 124312 156664 124364 156670
rect 124312 156606 124364 156612
rect 122748 152788 122800 152794
rect 122748 152730 122800 152736
rect 121460 152380 121512 152386
rect 121460 152322 121512 152328
rect 119896 151564 119948 151570
rect 119896 151506 119948 151512
rect 117318 151328 117374 151337
rect 117318 151263 117374 151272
rect 119908 149940 119936 151506
rect 122760 149954 122788 152730
rect 122514 149926 122788 149954
rect 124416 149940 124444 169390
rect 125060 149940 125088 196454
rect 127912 180794 127940 200124
rect 128510 199866 128538 200124
rect 128464 199838 128538 199866
rect 128464 195770 128492 199838
rect 128452 195764 128504 195770
rect 128452 195706 128504 195712
rect 126992 180766 127940 180794
rect 126992 152930 127020 180766
rect 129844 172106 129872 200124
rect 133018 199866 133046 200124
rect 133018 199838 133092 199866
rect 133064 194177 133092 199838
rect 133050 194168 133106 194177
rect 133050 194103 133106 194112
rect 134352 192982 134380 200124
rect 135260 196580 135312 196586
rect 135260 196522 135312 196528
rect 134340 192976 134392 192982
rect 134340 192918 134392 192924
rect 130200 179104 130252 179110
rect 130200 179046 130252 179052
rect 129832 172100 129884 172106
rect 129832 172042 129884 172048
rect 127072 162172 127124 162178
rect 127072 162114 127124 162120
rect 126980 152924 127032 152930
rect 126980 152866 127032 152872
rect 127084 149954 127112 162114
rect 129556 153196 129608 153202
rect 129556 153138 129608 153144
rect 127624 152924 127676 152930
rect 127624 152866 127676 152872
rect 127022 149926 127112 149954
rect 127636 149940 127664 152866
rect 129568 149940 129596 153138
rect 130212 149940 130240 179046
rect 135272 149954 135300 196522
rect 137572 180794 137600 200124
rect 138170 199866 138198 200124
rect 138170 199838 138244 199866
rect 138216 195838 138244 199838
rect 138204 195832 138256 195838
rect 138204 195774 138256 195780
rect 142080 194342 142108 200124
rect 147830 199866 147858 200124
rect 147830 199838 147904 199866
rect 147876 198354 147904 199838
rect 147864 198348 147916 198354
rect 147864 198290 147916 198296
rect 145656 198212 145708 198218
rect 145656 198154 145708 198160
rect 142068 194336 142120 194342
rect 142068 194278 142120 194284
rect 141792 193860 141844 193866
rect 141792 193802 141844 193808
rect 139398 192944 139454 192953
rect 139398 192879 139454 192888
rect 136652 180766 137600 180794
rect 136652 155786 136680 180766
rect 137284 163940 137336 163946
rect 137284 163882 137336 163888
rect 136640 155780 136692 155786
rect 136640 155722 136692 155728
rect 135996 153196 136048 153202
rect 135996 153138 136048 153144
rect 135272 149926 135378 149954
rect 136008 149940 136036 153138
rect 137296 149940 137324 163882
rect 139412 149954 139440 192879
rect 141148 153128 141200 153134
rect 141148 153070 141200 153076
rect 139412 149926 139886 149954
rect 141160 149940 141188 153070
rect 141804 149940 141832 193802
rect 142436 161084 142488 161090
rect 142436 161026 142488 161032
rect 142448 149940 142476 161026
rect 145012 153128 145064 153134
rect 145012 153070 145064 153076
rect 145024 149940 145052 153070
rect 145668 149940 145696 198154
rect 146298 192944 146354 192953
rect 146298 192879 146354 192888
rect 146312 149940 146340 192879
rect 146944 184680 146996 184686
rect 146944 184622 146996 184628
rect 146956 149940 146984 184622
rect 147678 181656 147734 181665
rect 147678 181591 147734 181600
rect 147692 149954 147720 181591
rect 150452 166326 150480 200124
rect 151740 195158 151768 200124
rect 153672 198121 153700 200124
rect 153658 198112 153714 198121
rect 153658 198047 153714 198056
rect 150532 195152 150584 195158
rect 150532 195094 150584 195100
rect 151728 195152 151780 195158
rect 151728 195094 151780 195100
rect 150544 166462 150572 195094
rect 154316 192914 154344 200124
rect 154304 192908 154356 192914
rect 154304 192850 154356 192856
rect 151820 192364 151872 192370
rect 151820 192306 151872 192312
rect 150532 166456 150584 166462
rect 150532 166398 150584 166404
rect 150440 166320 150492 166326
rect 150440 166262 150492 166268
rect 150164 158568 150216 158574
rect 150164 158510 150216 158516
rect 147692 149926 148258 149954
rect 150176 149940 150204 158510
rect 151832 149954 151860 192306
rect 155604 180794 155632 200124
rect 156846 199866 156874 200124
rect 156340 199838 156874 199866
rect 156340 180794 156368 199838
rect 158180 191729 158208 200124
rect 158536 199436 158588 199442
rect 158536 199378 158588 199384
rect 158166 191720 158222 191729
rect 158166 191655 158222 191664
rect 154592 180766 155632 180794
rect 155972 180766 156368 180794
rect 154592 155718 154620 180766
rect 155316 159792 155368 159798
rect 155316 159734 155368 159740
rect 154580 155712 154632 155718
rect 154580 155654 154632 155660
rect 153382 152688 153438 152697
rect 153382 152623 153438 152632
rect 151832 149926 152122 149954
rect 153396 149940 153424 152623
rect 155328 149940 155356 159734
rect 155972 158166 156000 180766
rect 157890 170368 157946 170377
rect 157890 170303 157946 170312
rect 155960 158160 156012 158166
rect 155960 158102 156012 158108
rect 157904 149940 157932 170303
rect 158548 149940 158576 199378
rect 158824 180794 158852 200124
rect 160112 198830 160140 200124
rect 160100 198824 160152 198830
rect 160100 198766 160152 198772
rect 160756 198218 160784 200124
rect 160744 198212 160796 198218
rect 160744 198154 160796 198160
rect 161400 195158 161428 200124
rect 160100 195152 160152 195158
rect 160100 195094 160152 195100
rect 161388 195152 161440 195158
rect 161388 195094 161440 195100
rect 159180 184748 159232 184754
rect 159180 184690 159232 184696
rect 158732 180766 158852 180794
rect 158732 158098 158760 180766
rect 158720 158092 158772 158098
rect 158720 158034 158772 158040
rect 159192 149940 159220 184690
rect 160112 152862 160140 195094
rect 163332 190454 163360 200124
rect 165264 198150 165292 200124
rect 167840 198966 167868 200124
rect 167828 198960 167880 198966
rect 167828 198902 167880 198908
rect 168484 198558 168512 200124
rect 168472 198552 168524 198558
rect 168472 198494 168524 198500
rect 166264 198212 166316 198218
rect 166264 198154 166316 198160
rect 165252 198144 165304 198150
rect 165252 198086 165304 198092
rect 162872 190426 163360 190454
rect 161756 155848 161808 155854
rect 161756 155790 161808 155796
rect 160100 152856 160152 152862
rect 160100 152798 160152 152804
rect 161768 149940 161796 155790
rect 162872 155310 162900 190426
rect 163044 183524 163096 183530
rect 163044 183466 163096 183472
rect 162860 155304 162912 155310
rect 162860 155246 162912 155252
rect 163056 149940 163084 183466
rect 166276 157010 166304 198154
rect 169128 189990 169156 200124
rect 169116 189984 169168 189990
rect 169116 189926 169168 189932
rect 169772 188902 169800 200124
rect 170416 198121 170444 200124
rect 170402 198112 170458 198121
rect 170402 198047 170458 198056
rect 172992 192438 173020 200124
rect 173636 192914 173664 200124
rect 174280 195770 174308 200124
rect 174924 199073 174952 200124
rect 174910 199064 174966 199073
rect 174910 198999 174966 199008
rect 174268 195764 174320 195770
rect 174268 195706 174320 195712
rect 175924 195220 175976 195226
rect 175924 195162 175976 195168
rect 173624 192908 173676 192914
rect 173624 192850 173676 192856
rect 172980 192432 173032 192438
rect 172980 192374 173032 192380
rect 174636 189984 174688 189990
rect 174636 189926 174688 189932
rect 169760 188896 169812 188902
rect 169760 188838 169812 188844
rect 172058 179888 172114 179897
rect 172058 179823 172114 179832
rect 170772 169516 170824 169522
rect 170772 169458 170824 169464
rect 168380 159588 168432 159594
rect 168380 159530 168432 159536
rect 166264 157004 166316 157010
rect 166264 156946 166316 156952
rect 166908 154012 166960 154018
rect 166908 153954 166960 153960
rect 166920 149940 166948 153954
rect 168392 153105 168420 159530
rect 168378 153096 168434 153105
rect 168378 153031 168434 153040
rect 170126 152824 170182 152833
rect 170126 152759 170182 152768
rect 170140 149940 170168 152759
rect 170784 149940 170812 169458
rect 172072 149940 172100 179823
rect 174648 149940 174676 189926
rect 175280 154216 175332 154222
rect 175280 154158 175332 154164
rect 175292 149940 175320 154158
rect 175936 149940 175964 195162
rect 178788 180794 178816 200124
rect 180076 195242 180104 200124
rect 178052 180766 178816 180794
rect 179432 195214 180104 195242
rect 176660 169584 176712 169590
rect 176660 169526 176712 169532
rect 176672 149954 176700 169526
rect 178052 154018 178080 180766
rect 178132 160744 178184 160750
rect 178132 160686 178184 160692
rect 178040 154012 178092 154018
rect 178040 153954 178092 153960
rect 178144 153134 178172 160686
rect 179432 155786 179460 195214
rect 180720 195158 180748 200124
rect 181318 199866 181346 200124
rect 181318 199838 181392 199866
rect 179512 195152 179564 195158
rect 179512 195094 179564 195100
rect 180708 195152 180760 195158
rect 180708 195094 180760 195100
rect 179524 187678 179552 195094
rect 181364 194274 181392 199838
rect 182652 196586 182680 200124
rect 182640 196580 182692 196586
rect 182640 196522 182692 196528
rect 181352 194268 181404 194274
rect 181352 194210 181404 194216
rect 183940 189038 183968 200124
rect 184584 191690 184612 200124
rect 185826 199866 185854 200124
rect 185320 199838 185854 199866
rect 184572 191684 184624 191690
rect 184572 191626 184624 191632
rect 183928 189032 183980 189038
rect 183928 188974 183980 188980
rect 179512 187672 179564 187678
rect 179512 187614 179564 187620
rect 183008 184340 183060 184346
rect 183008 184282 183060 184288
rect 180800 172100 180852 172106
rect 180800 172042 180852 172048
rect 179420 155780 179472 155786
rect 179420 155722 179472 155728
rect 178132 153128 178184 153134
rect 178132 153070 178184 153076
rect 179788 153128 179840 153134
rect 179788 153070 179840 153076
rect 179142 152824 179198 152833
rect 179142 152759 179198 152768
rect 176672 149926 177238 149954
rect 179156 149940 179184 152759
rect 179800 149940 179828 153070
rect 180812 149954 180840 172042
rect 180812 149926 181746 149954
rect 183020 149940 183048 184282
rect 185320 180794 185348 199838
rect 187804 196761 187832 200124
rect 187790 196752 187846 196761
rect 187790 196687 187846 196696
rect 189092 193118 189120 200124
rect 190334 199866 190362 200124
rect 190334 199838 190408 199866
rect 190380 198218 190408 199838
rect 190368 198212 190420 198218
rect 190368 198154 190420 198160
rect 189080 193112 189132 193118
rect 189080 193054 189132 193060
rect 192956 190454 192984 200124
rect 194244 198830 194272 200124
rect 194232 198824 194284 198830
rect 194232 198766 194284 198772
rect 194888 192846 194916 200124
rect 195486 199866 195514 200124
rect 194980 199838 195514 199866
rect 194876 192840 194928 192846
rect 194876 192782 194928 192788
rect 191852 190426 192984 190454
rect 187516 186108 187568 186114
rect 187516 186050 187568 186056
rect 184952 180766 185348 180794
rect 184952 163606 184980 180766
rect 184940 163600 184992 163606
rect 184940 163542 184992 163548
rect 187528 149940 187556 186050
rect 191852 180470 191880 190426
rect 192024 187672 192076 187678
rect 192024 187614 192076 187620
rect 191840 180464 191892 180470
rect 191840 180406 191892 180412
rect 188160 176316 188212 176322
rect 188160 176258 188212 176264
rect 188172 149940 188200 176258
rect 188804 157004 188856 157010
rect 188804 156946 188856 156952
rect 188816 149940 188844 156946
rect 192036 149940 192064 187614
rect 194980 184890 195008 199838
rect 196820 194041 196848 200124
rect 197464 195242 197492 200124
rect 197372 195214 197492 195242
rect 196806 194032 196862 194041
rect 196806 193967 196862 193976
rect 194968 184884 195020 184890
rect 194968 184826 195020 184832
rect 197372 180334 197400 195214
rect 198108 182170 198136 200124
rect 198096 182164 198148 182170
rect 198096 182106 198148 182112
rect 197360 180328 197412 180334
rect 197360 180270 197412 180276
rect 195242 172408 195298 172417
rect 195242 172343 195298 172352
rect 193220 170604 193272 170610
rect 193220 170546 193272 170552
rect 193232 149954 193260 170546
rect 193232 149926 193982 149954
rect 195256 149940 195284 172343
rect 197176 164892 197228 164898
rect 197176 164834 197228 164840
rect 197188 149940 197216 164834
rect 198752 151638 198780 200124
rect 199994 199866 200022 200124
rect 199994 199838 200068 199866
rect 200040 199073 200068 199838
rect 200026 199064 200082 199073
rect 200026 198999 200082 199008
rect 201328 198150 201356 200124
rect 201972 198422 202000 200124
rect 201960 198416 202012 198422
rect 201960 198358 202012 198364
rect 201316 198144 201368 198150
rect 201316 198086 201368 198092
rect 204548 195226 204576 200124
rect 205146 199866 205174 200124
rect 205146 199838 205220 199866
rect 204536 195220 204588 195226
rect 204536 195162 204588 195168
rect 205192 193118 205220 199838
rect 208412 199238 208440 200124
rect 209654 200002 209682 200124
rect 209148 199974 209682 200002
rect 208400 199232 208452 199238
rect 208400 199174 208452 199180
rect 209148 198234 209176 199974
rect 208504 198206 209176 198234
rect 208122 197976 208178 197985
rect 208122 197911 208178 197920
rect 205180 193112 205232 193118
rect 205180 193054 205232 193060
rect 202972 191412 203024 191418
rect 202972 191354 203024 191360
rect 201500 184884 201552 184890
rect 201500 184826 201552 184832
rect 199752 166728 199804 166734
rect 199752 166670 199804 166676
rect 199106 152688 199162 152697
rect 199106 152623 199162 152632
rect 198740 151632 198792 151638
rect 198740 151574 198792 151580
rect 199120 149940 199148 152623
rect 199764 149940 199792 166670
rect 200396 152856 200448 152862
rect 200396 152798 200448 152804
rect 200408 149940 200436 152798
rect 201512 149954 201540 184826
rect 201512 149926 202354 149954
rect 202984 149940 203012 191354
rect 207480 167748 207532 167754
rect 207480 167690 207532 167696
rect 204260 156936 204312 156942
rect 204260 156878 204312 156884
rect 204272 149940 204300 156878
rect 205640 155712 205692 155718
rect 205640 155654 205692 155660
rect 204902 152960 204958 152969
rect 204902 152895 204958 152904
rect 204916 149940 204944 152895
rect 205652 149954 205680 155654
rect 205652 149926 206862 149954
rect 207492 149940 207520 167690
rect 208136 149940 208164 197911
rect 208504 153066 208532 198206
rect 208768 198076 208820 198082
rect 208768 198018 208820 198024
rect 208492 153060 208544 153066
rect 208492 153002 208544 153008
rect 208780 149940 208808 198018
rect 210988 195158 211016 200124
rect 209780 195152 209832 195158
rect 209780 195094 209832 195100
rect 210976 195152 211028 195158
rect 210976 195094 211028 195100
rect 209412 153060 209464 153066
rect 209412 153002 209464 153008
rect 209424 149940 209452 153002
rect 209792 152998 209820 195094
rect 211986 190360 212042 190369
rect 211986 190295 212042 190304
rect 209872 184816 209924 184822
rect 209872 184758 209924 184764
rect 209780 152992 209832 152998
rect 209780 152934 209832 152940
rect 209884 149954 209912 184758
rect 209884 149926 210726 149954
rect 212000 149940 212028 190295
rect 213564 180794 213592 200124
rect 214806 200002 214834 200124
rect 214484 199974 214834 200002
rect 214484 180794 214512 199974
rect 216140 189718 216168 200124
rect 216128 189712 216180 189718
rect 216128 189654 216180 189660
rect 216496 184884 216548 184890
rect 216496 184826 216548 184832
rect 212552 180766 213592 180794
rect 213932 180766 214512 180794
rect 212552 163674 212580 180766
rect 213932 179110 213960 180766
rect 213920 179104 213972 179110
rect 213920 179046 213972 179052
rect 213276 176384 213328 176390
rect 213276 176326 213328 176332
rect 212540 163668 212592 163674
rect 212540 163610 212592 163616
rect 213288 149940 213316 176326
rect 214104 163736 214156 163742
rect 214104 163678 214156 163684
rect 213920 152992 213972 152998
rect 213920 152934 213972 152940
rect 213932 149940 213960 152934
rect 214116 149954 214144 163678
rect 214116 149926 215234 149954
rect 216508 149940 216536 184826
rect 216784 180794 216812 200124
rect 220360 196716 220412 196722
rect 220360 196658 220412 196664
rect 217784 192840 217836 192846
rect 217784 192782 217836 192788
rect 216692 180766 216812 180794
rect 216692 155310 216720 180766
rect 216772 159452 216824 159458
rect 216772 159394 216824 159400
rect 216680 155304 216732 155310
rect 216680 155246 216732 155252
rect 216784 153134 216812 159394
rect 216772 153128 216824 153134
rect 216772 153070 216824 153076
rect 217796 149940 217824 192782
rect 219716 160812 219768 160818
rect 219716 160754 219768 160760
rect 219728 149940 219756 160754
rect 220372 149940 220400 196658
rect 221292 188358 221320 200124
rect 221936 198898 221964 200124
rect 221924 198892 221976 198898
rect 221924 198834 221976 198840
rect 222580 190454 222608 200124
rect 223868 198558 223896 200124
rect 223856 198552 223908 198558
rect 223856 198494 223908 198500
rect 222212 190426 222608 190454
rect 221280 188352 221332 188358
rect 221280 188294 221332 188300
rect 222212 163742 222240 190426
rect 226444 189650 226472 200124
rect 227732 196722 227760 200124
rect 227720 196716 227772 196722
rect 227720 196658 227772 196664
rect 228376 195634 228404 200124
rect 228364 195628 228416 195634
rect 228364 195570 228416 195576
rect 226432 189644 226484 189650
rect 226432 189586 226484 189592
rect 222292 185700 222344 185706
rect 222292 185642 222344 185648
rect 222200 163736 222252 163742
rect 222200 163678 222252 163684
rect 221648 161152 221700 161158
rect 221648 161094 221700 161100
rect 221660 149940 221688 161094
rect 222304 149940 222332 185642
rect 224224 183252 224276 183258
rect 224224 183194 224276 183200
rect 223948 154080 224000 154086
rect 223948 154022 224000 154028
rect 223960 149954 223988 154022
rect 224236 153202 224264 183194
rect 230952 180794 230980 200124
rect 232240 195242 232268 200124
rect 230492 180766 230980 180794
rect 231872 195214 232268 195242
rect 226800 180396 226852 180402
rect 226800 180338 226852 180344
rect 225512 169652 225564 169658
rect 225512 169594 225564 169600
rect 224868 154080 224920 154086
rect 224868 154022 224920 154028
rect 224224 153196 224276 153202
rect 224224 153138 224276 153144
rect 223960 149926 224250 149954
rect 224880 149940 224908 154022
rect 225524 149940 225552 169594
rect 226156 164008 226208 164014
rect 226156 163950 226208 163956
rect 226168 149940 226196 163950
rect 226812 149940 226840 180338
rect 227720 177812 227772 177818
rect 227720 177754 227772 177760
rect 227732 149954 227760 177754
rect 230492 170542 230520 180766
rect 230480 170536 230532 170542
rect 230480 170478 230532 170484
rect 228732 165164 228784 165170
rect 228732 165106 228784 165112
rect 227732 149926 228114 149954
rect 228744 149940 228772 165106
rect 231872 158234 231900 195214
rect 232884 180794 232912 200124
rect 233482 199866 233510 200124
rect 233482 199838 233556 199866
rect 233528 198966 233556 199838
rect 233516 198960 233568 198966
rect 233516 198902 233568 198908
rect 235170 196616 235226 196625
rect 235170 196551 235226 196560
rect 234528 184340 234580 184346
rect 234528 184282 234580 184288
rect 231964 180766 232912 180794
rect 231964 165102 231992 180766
rect 233884 170536 233936 170542
rect 233884 170478 233936 170484
rect 231952 165096 232004 165102
rect 231952 165038 232004 165044
rect 231860 158228 231912 158234
rect 231860 158170 231912 158176
rect 232596 155848 232648 155854
rect 232596 155790 232648 155796
rect 229376 155780 229428 155786
rect 229376 155722 229428 155728
rect 230020 155780 230072 155786
rect 230020 155722 230072 155728
rect 229388 149940 229416 155722
rect 230032 149940 230060 155722
rect 232608 149940 232636 155790
rect 233896 149940 233924 170478
rect 234540 149940 234568 184282
rect 235184 149940 235212 196551
rect 236748 187610 236776 200124
rect 238634 200002 238662 200124
rect 238588 199974 238662 200002
rect 238588 194954 238616 199974
rect 239968 195158 239996 200124
rect 238760 195152 238812 195158
rect 238760 195094 238812 195100
rect 239956 195152 240008 195158
rect 239956 195094 240008 195100
rect 237380 194948 237432 194954
rect 237380 194890 237432 194896
rect 238576 194948 238628 194954
rect 238576 194890 238628 194896
rect 236736 187604 236788 187610
rect 236736 187546 236788 187552
rect 237392 165102 237420 194890
rect 237380 165096 237432 165102
rect 237380 165038 237432 165044
rect 237748 164076 237800 164082
rect 237748 164018 237800 164024
rect 237760 149940 237788 164018
rect 238772 155650 238800 195094
rect 241256 194002 241284 200124
rect 243142 200002 243170 200124
rect 243096 199974 243170 200002
rect 241244 193996 241296 194002
rect 241244 193938 241296 193944
rect 242992 193928 243044 193934
rect 242992 193870 243044 193876
rect 239036 186924 239088 186930
rect 239036 186866 239088 186872
rect 238760 155644 238812 155650
rect 238760 155586 238812 155592
rect 239048 149940 239076 186866
rect 241612 177880 241664 177886
rect 241612 177822 241664 177828
rect 240140 160880 240192 160886
rect 240140 160822 240192 160828
rect 240152 149954 240180 160822
rect 240966 152552 241022 152561
rect 240966 152487 241022 152496
rect 240152 149926 240350 149954
rect 240980 149940 241008 152487
rect 241624 149940 241652 177822
rect 242256 172032 242308 172038
rect 242256 171974 242308 171980
rect 242268 149940 242296 171974
rect 243004 149954 243032 193870
rect 243096 192778 243124 199974
rect 244476 198490 244504 200124
rect 244464 198484 244516 198490
rect 244464 198426 244516 198432
rect 246408 196790 246436 200124
rect 247052 198898 247080 200124
rect 247040 198892 247092 198898
rect 247040 198834 247092 198840
rect 246396 196784 246448 196790
rect 246396 196726 246448 196732
rect 247696 195498 247724 200124
rect 247684 195492 247736 195498
rect 247684 195434 247736 195440
rect 249628 194070 249656 200124
rect 252802 200002 252830 200124
rect 252572 199974 252830 200002
rect 249616 194064 249668 194070
rect 249616 194006 249668 194012
rect 243084 192772 243136 192778
rect 243084 192714 243136 192720
rect 245476 184612 245528 184618
rect 245476 184554 245528 184560
rect 242926 149926 243032 149954
rect 245488 149940 245516 184554
rect 249984 184136 250036 184142
rect 249984 184078 250036 184084
rect 246120 182776 246172 182782
rect 246120 182718 246172 182724
rect 246132 149940 246160 182718
rect 249340 173392 249392 173398
rect 249340 173334 249392 173340
rect 248420 161220 248472 161226
rect 248420 161162 248472 161168
rect 248432 149954 248460 161162
rect 248432 149926 248722 149954
rect 249352 149940 249380 173334
rect 249996 149940 250024 184078
rect 250628 177540 250680 177546
rect 250628 177482 250680 177488
rect 250640 149940 250668 177482
rect 251270 162072 251326 162081
rect 251270 162007 251326 162016
rect 251284 149940 251312 162007
rect 252572 159662 252600 199974
rect 254780 198098 254808 200124
rect 254860 198348 254912 198354
rect 254860 198290 254912 198296
rect 253952 198070 254808 198098
rect 252652 188352 252704 188358
rect 252652 188294 252704 188300
rect 252560 159656 252612 159662
rect 252560 159598 252612 159604
rect 251916 153264 251968 153270
rect 251916 153206 251968 153212
rect 251928 149940 251956 153206
rect 252664 149954 252692 188294
rect 253952 160886 253980 198070
rect 254872 195974 254900 198290
rect 254780 195946 254900 195974
rect 254780 180794 254808 195946
rect 256068 190454 256096 200124
rect 257954 199866 257982 200124
rect 257908 199838 257982 199866
rect 257908 198937 257936 199838
rect 257894 198928 257950 198937
rect 257894 198863 257950 198872
rect 259460 195424 259512 195430
rect 259460 195366 259512 195372
rect 254596 180766 254808 180794
rect 255332 190426 256096 190454
rect 253940 160880 253992 160886
rect 253940 160822 253992 160828
rect 254596 155922 254624 180766
rect 254584 155916 254636 155922
rect 254584 155858 254636 155864
rect 254492 153128 254544 153134
rect 254492 153070 254544 153076
rect 252664 149926 253230 149954
rect 254504 149940 254532 153070
rect 255332 150074 255360 190426
rect 255780 182028 255832 182034
rect 255780 181970 255832 181976
rect 255320 150068 255372 150074
rect 255320 150010 255372 150016
rect 255792 149940 255820 181970
rect 259000 166796 259052 166802
rect 259000 166738 259052 166744
rect 259012 149940 259040 166738
rect 259472 153270 259500 195366
rect 259932 180794 259960 200124
rect 260576 195430 260604 200124
rect 262462 199866 262490 200124
rect 262462 199838 262536 199866
rect 262508 197402 262536 199838
rect 262496 197396 262548 197402
rect 262496 197338 262548 197344
rect 260564 195424 260616 195430
rect 260564 195366 260616 195372
rect 263796 192710 263824 200124
rect 264244 197396 264296 197402
rect 264244 197338 264296 197344
rect 263784 192704 263836 192710
rect 263784 192646 263836 192652
rect 259564 180766 259960 180794
rect 259564 158302 259592 180766
rect 264152 172168 264204 172174
rect 264152 172110 264204 172116
rect 260840 163804 260892 163810
rect 260840 163746 260892 163752
rect 259552 158296 259604 158302
rect 259552 158238 259604 158244
rect 259644 157004 259696 157010
rect 259644 156946 259696 156952
rect 259460 153264 259512 153270
rect 259460 153206 259512 153212
rect 259656 149940 259684 156946
rect 260288 154284 260340 154290
rect 260288 154226 260340 154232
rect 260300 149940 260328 154226
rect 260852 149954 260880 163746
rect 260852 149926 261602 149954
rect 264164 149940 264192 172110
rect 264256 157894 264284 197338
rect 266084 196784 266136 196790
rect 266084 196726 266136 196732
rect 264244 157888 264296 157894
rect 264244 157830 264296 157836
rect 266096 149940 266124 196726
rect 266372 162314 266400 200124
rect 266970 199866 266998 200124
rect 266924 199838 266998 199866
rect 266924 195498 266952 199838
rect 268384 198144 268436 198150
rect 268384 198086 268436 198092
rect 266912 195492 266964 195498
rect 266912 195434 266964 195440
rect 268396 173330 268424 198086
rect 270236 180794 270264 200124
rect 271524 199306 271552 200124
rect 272122 199866 272150 200124
rect 272122 199838 272196 199866
rect 271512 199300 271564 199306
rect 271512 199242 271564 199248
rect 272168 198082 272196 199838
rect 272156 198076 272208 198082
rect 272156 198018 272208 198024
rect 270590 196616 270646 196625
rect 270590 196551 270646 196560
rect 269132 180766 270264 180794
rect 268660 177676 268712 177682
rect 268660 177618 268712 177624
rect 268384 173324 268436 173330
rect 268384 173266 268436 173272
rect 266360 162308 266412 162314
rect 266360 162250 266412 162256
rect 268016 158636 268068 158642
rect 268016 158578 268068 158584
rect 268028 149940 268056 158578
rect 268672 149940 268700 177618
rect 269132 155106 269160 180766
rect 269120 155100 269172 155106
rect 269120 155042 269172 155048
rect 270604 149940 270632 196551
rect 272524 184612 272576 184618
rect 272524 184554 272576 184560
rect 271234 163432 271290 163441
rect 271234 163367 271290 163376
rect 271248 149940 271276 163367
rect 271880 156936 271932 156942
rect 271880 156878 271932 156884
rect 271892 149940 271920 156878
rect 272536 149940 272564 184554
rect 273456 180794 273484 200124
rect 275388 198150 275416 200124
rect 275836 199572 275888 199578
rect 275836 199514 275888 199520
rect 275376 198144 275428 198150
rect 275376 198086 275428 198092
rect 275848 196858 275876 199514
rect 275836 196852 275888 196858
rect 275836 196794 275888 196800
rect 276032 193798 276060 200124
rect 276630 199866 276658 200124
rect 276630 199838 276704 199866
rect 276676 196858 276704 199838
rect 276664 196852 276716 196858
rect 276664 196794 276716 196800
rect 276020 193792 276072 193798
rect 276020 193734 276072 193740
rect 278608 191593 278636 200124
rect 278594 191584 278650 191593
rect 278594 191519 278650 191528
rect 279252 190454 279280 200124
rect 280540 193730 280568 200124
rect 281184 195498 281212 200124
rect 281782 199866 281810 200124
rect 281736 199838 281810 199866
rect 281172 195492 281224 195498
rect 281172 195434 281224 195440
rect 281736 194206 281764 199838
rect 281724 194200 281776 194206
rect 281724 194142 281776 194148
rect 280528 193724 280580 193730
rect 280528 193666 280580 193672
rect 278792 190426 279280 190454
rect 275744 190392 275796 190398
rect 275744 190334 275796 190340
rect 273364 180766 273484 180794
rect 273364 176390 273392 180766
rect 274456 180464 274508 180470
rect 274456 180406 274508 180412
rect 273352 176384 273404 176390
rect 273352 176326 273404 176332
rect 274468 149940 274496 180406
rect 275756 149940 275784 190334
rect 277400 166864 277452 166870
rect 277400 166806 277452 166812
rect 277412 149954 277440 166806
rect 278792 163878 278820 190426
rect 278964 186176 279016 186182
rect 278964 186118 279016 186124
rect 278780 163872 278832 163878
rect 278780 163814 278832 163820
rect 277412 149926 278346 149954
rect 278976 149940 279004 186118
rect 283116 180794 283144 200124
rect 287624 198354 287652 200124
rect 287612 198348 287664 198354
rect 287612 198290 287664 198296
rect 284760 194200 284812 194206
rect 284760 194142 284812 194148
rect 283472 184068 283524 184074
rect 283472 184010 283524 184016
rect 282932 180766 283144 180794
rect 279608 180464 279660 180470
rect 279608 180406 279660 180412
rect 279620 149940 279648 180406
rect 282828 160676 282880 160682
rect 282828 160618 282880 160624
rect 281540 156800 281592 156806
rect 281540 156742 281592 156748
rect 281552 149954 281580 156742
rect 281552 149926 282210 149954
rect 282840 149940 282868 160618
rect 282932 158438 282960 180766
rect 282920 158432 282972 158438
rect 282920 158374 282972 158380
rect 283484 149940 283512 184010
rect 284116 155508 284168 155514
rect 284116 155450 284168 155456
rect 284128 149940 284156 155450
rect 284772 149940 284800 194142
rect 287980 193656 288032 193662
rect 287980 193598 288032 193604
rect 285404 191412 285456 191418
rect 285404 191354 285456 191360
rect 285416 149940 285444 191354
rect 285680 162240 285732 162246
rect 285680 162182 285732 162188
rect 285692 149954 285720 162182
rect 285692 149926 286718 149954
rect 287992 149940 288020 193598
rect 290844 180794 290872 200124
rect 291442 200002 291470 200124
rect 289832 180766 290872 180794
rect 291212 199974 291470 200002
rect 289832 154222 289860 180766
rect 291212 154222 291240 199974
rect 292776 180794 292804 200124
rect 293960 195424 294012 195430
rect 293960 195366 294012 195372
rect 293132 188420 293184 188426
rect 293132 188362 293184 188368
rect 292592 180766 292804 180794
rect 292592 158710 292620 180766
rect 292580 158704 292632 158710
rect 292580 158646 292632 158652
rect 292488 155644 292540 155650
rect 292488 155586 292540 155592
rect 289820 154216 289872 154222
rect 289820 154158 289872 154164
rect 291200 154216 291252 154222
rect 291200 154158 291252 154164
rect 291200 153196 291252 153202
rect 291200 153138 291252 153144
rect 291212 149940 291240 153138
rect 292500 149940 292528 155586
rect 293144 149940 293172 188362
rect 293972 150006 294000 195366
rect 294064 169590 294092 200124
rect 294708 195430 294736 200124
rect 295352 196926 295380 200124
rect 295340 196920 295392 196926
rect 295340 196862 295392 196868
rect 297928 195430 297956 200124
rect 294696 195424 294748 195430
rect 294696 195366 294748 195372
rect 297916 195424 297968 195430
rect 297916 195366 297968 195372
rect 296352 188352 296404 188358
rect 296352 188294 296404 188300
rect 294052 169584 294104 169590
rect 294052 169526 294104 169532
rect 295708 155168 295760 155174
rect 295708 155110 295760 155116
rect 293960 150000 294012 150006
rect 293960 149942 294012 149948
rect 295720 149940 295748 155110
rect 296364 149940 296392 188294
rect 299860 180794 299888 200124
rect 300458 199866 300486 200124
rect 300458 199838 300532 199866
rect 300504 199170 300532 199838
rect 300492 199164 300544 199170
rect 300492 199106 300544 199112
rect 300860 191480 300912 191486
rect 300860 191422 300912 191428
rect 299492 180766 299888 180794
rect 299492 154290 299520 180766
rect 299480 154284 299532 154290
rect 299480 154226 299532 154232
rect 297640 152652 297692 152658
rect 297640 152594 297692 152600
rect 297652 149940 297680 152594
rect 300872 149940 300900 191422
rect 301792 180794 301820 200124
rect 302148 182164 302200 182170
rect 302148 182106 302200 182112
rect 301056 180766 301820 180794
rect 301056 172038 301084 180766
rect 301044 172032 301096 172038
rect 301044 171974 301096 171980
rect 302160 149940 302188 182106
rect 303080 180794 303108 200124
rect 303724 185978 303752 200124
rect 304368 196926 304396 200124
rect 304356 196920 304408 196926
rect 304356 196862 304408 196868
rect 303712 185972 303764 185978
rect 303712 185914 303764 185920
rect 302252 180766 303108 180794
rect 302252 163810 302280 180766
rect 302240 163804 302292 163810
rect 302240 163746 302292 163752
rect 305012 158370 305040 200124
rect 305610 200002 305638 200124
rect 305104 199974 305638 200002
rect 305104 163878 305132 199974
rect 306944 180794 306972 200124
rect 310118 200002 310146 200124
rect 309612 199974 310146 200002
rect 307024 198076 307076 198082
rect 307024 198018 307076 198024
rect 306392 180766 306972 180794
rect 305092 163872 305144 163878
rect 305092 163814 305144 163820
rect 305000 158364 305052 158370
rect 305000 158306 305052 158312
rect 306392 151638 306420 180766
rect 306472 169720 306524 169726
rect 306472 169662 306524 169668
rect 306380 151632 306432 151638
rect 306380 151574 306432 151580
rect 306484 149954 306512 169662
rect 307036 164218 307064 198018
rect 307944 191344 307996 191350
rect 307944 191286 307996 191292
rect 307024 164212 307076 164218
rect 307024 164154 307076 164160
rect 306484 149926 307326 149954
rect 307956 149940 307984 191286
rect 309612 180794 309640 199974
rect 312740 195634 312768 200124
rect 312728 195628 312780 195634
rect 312728 195570 312780 195576
rect 314028 180794 314056 200124
rect 315270 199866 315298 200124
rect 315270 199838 315344 199866
rect 315316 197878 315344 199838
rect 317248 199442 317276 200124
rect 317236 199436 317288 199442
rect 317236 199378 317288 199384
rect 317892 197946 317920 200124
rect 319778 199866 319806 200124
rect 319778 199838 319852 199866
rect 319824 199374 319852 199838
rect 319812 199368 319864 199374
rect 319812 199310 319864 199316
rect 317880 197940 317932 197946
rect 317880 197882 317932 197888
rect 315304 197872 315356 197878
rect 315304 197814 315356 197820
rect 318892 193860 318944 193866
rect 318892 193802 318944 193808
rect 309152 180766 309640 180794
rect 313292 180766 314056 180794
rect 309152 157010 309180 180766
rect 313096 176384 313148 176390
rect 313096 176326 313148 176332
rect 312452 175092 312504 175098
rect 312452 175034 312504 175040
rect 309876 164212 309928 164218
rect 309876 164154 309928 164160
rect 309140 157004 309192 157010
rect 309140 156946 309192 156952
rect 309232 155032 309284 155038
rect 309232 154974 309284 154980
rect 308588 154148 308640 154154
rect 308588 154090 308640 154096
rect 308600 149940 308628 154090
rect 309244 149940 309272 154974
rect 309888 149940 309916 164154
rect 310520 152652 310572 152658
rect 310520 152594 310572 152600
rect 310532 149940 310560 152594
rect 312464 149940 312492 175034
rect 313108 149940 313136 176326
rect 313292 149938 313320 180766
rect 315304 169584 315356 169590
rect 315304 169526 315356 169532
rect 314384 167680 314436 167686
rect 314384 167622 314436 167628
rect 313740 154148 313792 154154
rect 313740 154090 313792 154096
rect 313752 149940 313780 154090
rect 314396 149940 314424 167622
rect 315316 152930 315344 169526
rect 318248 156800 318300 156806
rect 318248 156742 318300 156748
rect 317602 155816 317658 155825
rect 317602 155751 317658 155760
rect 315304 152924 315356 152930
rect 315304 152866 315356 152872
rect 316592 152924 316644 152930
rect 316592 152866 316644 152872
rect 315028 152448 315080 152454
rect 315028 152390 315080 152396
rect 315040 149940 315068 152390
rect 316604 149954 316632 152866
rect 313280 149932 313332 149938
rect 59910 149903 59966 149912
rect 59820 120148 59872 120154
rect 59820 120090 59872 120096
rect 59636 117020 59688 117026
rect 59636 116962 59688 116968
rect 59636 111172 59688 111178
rect 59636 111114 59688 111120
rect 59544 98592 59596 98598
rect 59544 98534 59596 98540
rect 59082 96792 59138 96801
rect 59082 96727 59138 96736
rect 59648 79422 59676 111114
rect 59820 98728 59872 98734
rect 59820 98670 59872 98676
rect 59636 79416 59688 79422
rect 59636 79358 59688 79364
rect 58990 53272 59046 53281
rect 58990 53207 59046 53216
rect 58900 20664 58952 20670
rect 58900 20606 58952 20612
rect 59832 17474 59860 98670
rect 59924 17610 59952 149903
rect 316358 149926 316632 149954
rect 317616 149940 317644 155751
rect 318260 149940 318288 156742
rect 318904 149940 318932 193802
rect 321112 180794 321140 200124
rect 324332 195242 324360 200124
rect 324930 200002 324958 200124
rect 324884 199974 324958 200002
rect 324332 195214 324452 195242
rect 324320 195152 324372 195158
rect 324320 195094 324372 195100
rect 322112 187604 322164 187610
rect 322112 187546 322164 187552
rect 320192 180766 321140 180794
rect 320192 161022 320220 180766
rect 321466 163704 321522 163713
rect 321466 163639 321522 163648
rect 320180 161016 320232 161022
rect 320180 160958 320232 160964
rect 320824 158500 320876 158506
rect 320824 158442 320876 158448
rect 320836 149940 320864 158442
rect 321480 149940 321508 163639
rect 322124 149940 322152 187546
rect 324332 164014 324360 195094
rect 324424 166666 324452 195214
rect 324884 195158 324912 199974
rect 326908 195158 326936 200124
rect 324872 195152 324924 195158
rect 324872 195094 324924 195100
rect 325700 195152 325752 195158
rect 325700 195094 325752 195100
rect 326896 195152 326948 195158
rect 326896 195094 326948 195100
rect 325712 169386 325740 195094
rect 327552 180794 327580 200124
rect 328196 199510 328224 200124
rect 328184 199504 328236 199510
rect 328184 199446 328236 199452
rect 328840 195242 328868 200124
rect 329438 200002 329466 200124
rect 327092 180766 327580 180794
rect 328472 195214 328868 195242
rect 328932 199974 329466 200002
rect 327092 172106 327120 180766
rect 327080 172100 327132 172106
rect 327080 172042 327132 172048
rect 325700 169380 325752 169386
rect 325700 169322 325752 169328
rect 324412 166660 324464 166666
rect 324412 166602 324464 166608
rect 324320 164008 324372 164014
rect 324320 163950 324372 163956
rect 328472 156806 328500 195214
rect 328932 180794 328960 199974
rect 330772 194313 330800 200124
rect 332060 198082 332088 200124
rect 332048 198076 332100 198082
rect 332048 198018 332100 198024
rect 330758 194304 330814 194313
rect 330758 194239 330814 194248
rect 333348 191214 333376 200124
rect 333946 199866 333974 200124
rect 333946 199838 334112 199866
rect 333980 195152 334032 195158
rect 333980 195094 334032 195100
rect 333336 191208 333388 191214
rect 333336 191150 333388 191156
rect 328564 180766 328960 180794
rect 328460 156800 328512 156806
rect 328460 156742 328512 156748
rect 328564 156738 328592 180766
rect 329194 180568 329250 180577
rect 329194 180503 329250 180512
rect 328736 169380 328788 169386
rect 328736 169322 328788 169328
rect 323400 156732 323452 156738
rect 323400 156674 323452 156680
rect 328552 156732 328604 156738
rect 328552 156674 328604 156680
rect 322756 155100 322808 155106
rect 322756 155042 322808 155048
rect 322768 149940 322796 155042
rect 323412 149940 323440 156674
rect 326620 152584 326672 152590
rect 325054 152552 325110 152561
rect 326620 152526 326672 152532
rect 327264 152584 327316 152590
rect 327264 152526 327316 152532
rect 325054 152487 325110 152496
rect 325068 149954 325096 152487
rect 324730 149926 325096 149954
rect 326632 149940 326660 152526
rect 327276 149940 327304 152526
rect 328748 149954 328776 169322
rect 328594 149926 328776 149954
rect 329208 149940 329236 180503
rect 330484 180328 330536 180334
rect 330484 180270 330536 180276
rect 330496 152794 330524 180270
rect 333992 156806 334020 195094
rect 334084 158681 334112 199838
rect 335280 195158 335308 200124
rect 335268 195152 335320 195158
rect 335268 195094 335320 195100
rect 337856 193050 337884 200124
rect 339098 200002 339126 200124
rect 338592 199974 339126 200002
rect 337844 193044 337896 193050
rect 337844 192986 337896 192992
rect 338592 180794 338620 199974
rect 340432 197334 340460 200124
rect 340880 199572 340932 199578
rect 340880 199514 340932 199520
rect 340420 197328 340472 197334
rect 340420 197270 340472 197276
rect 340892 197266 340920 199514
rect 340880 197260 340932 197266
rect 340880 197202 340932 197208
rect 339500 191208 339552 191214
rect 339500 191150 339552 191156
rect 338132 180766 338620 180794
rect 335636 169312 335688 169318
rect 335636 169254 335688 169260
rect 334070 158672 334126 158681
rect 334070 158607 334126 158616
rect 333980 156800 334032 156806
rect 333980 156742 334032 156748
rect 330484 152788 330536 152794
rect 330484 152730 330536 152736
rect 334992 152788 335044 152794
rect 334992 152730 335044 152736
rect 335004 149940 335032 152730
rect 335648 149940 335676 169254
rect 338132 155514 338160 180766
rect 338120 155508 338172 155514
rect 338120 155450 338172 155456
rect 339512 149940 339540 191150
rect 341076 190330 341104 200124
rect 342364 196897 342392 200124
rect 343008 198286 343036 200124
rect 346122 199336 346178 199345
rect 346122 199271 346178 199280
rect 342996 198280 343048 198286
rect 342996 198222 343048 198228
rect 346136 197810 346164 199271
rect 346228 198694 346256 200124
rect 347516 199730 347544 200124
rect 347700 200002 347728 200223
rect 346412 199702 347544 199730
rect 347608 199974 347728 200002
rect 346308 199640 346360 199646
rect 346308 199582 346360 199588
rect 346216 198688 346268 198694
rect 346216 198630 346268 198636
rect 346124 197804 346176 197810
rect 346124 197746 346176 197752
rect 342350 196888 342406 196897
rect 342350 196823 342406 196832
rect 342720 195152 342772 195158
rect 342720 195094 342772 195100
rect 341064 190324 341116 190330
rect 341064 190266 341116 190272
rect 340144 154216 340196 154222
rect 340144 154158 340196 154164
rect 340156 149940 340184 154158
rect 341798 152960 341854 152969
rect 341798 152895 341854 152904
rect 341812 149954 341840 152895
rect 342076 152244 342128 152250
rect 342076 152186 342128 152192
rect 341474 149926 341840 149954
rect 342088 149940 342116 152186
rect 342732 149940 342760 195094
rect 346320 192982 346348 199582
rect 346308 192976 346360 192982
rect 346308 192918 346360 192924
rect 345020 179036 345072 179042
rect 345020 178978 345072 178984
rect 343364 171964 343416 171970
rect 343364 171906 343416 171912
rect 343376 149940 343404 171906
rect 344008 152380 344060 152386
rect 344008 152322 344060 152328
rect 344020 149940 344048 152322
rect 345032 149954 345060 178978
rect 346412 164014 346440 199702
rect 347608 199617 347636 199974
rect 347688 199912 347740 199918
rect 347688 199854 347740 199860
rect 347594 199608 347650 199617
rect 347504 199572 347556 199578
rect 347594 199543 347650 199552
rect 347504 199514 347556 199520
rect 347516 184074 347544 199514
rect 347700 198529 347728 199854
rect 347686 198520 347742 198529
rect 347686 198455 347742 198464
rect 347792 184890 347820 474943
rect 347976 377097 348004 579022
rect 348240 576224 348292 576230
rect 348240 576166 348292 576172
rect 348148 568200 348200 568206
rect 348148 568142 348200 568148
rect 348056 566704 348108 566710
rect 348056 566646 348108 566652
rect 348068 402974 348096 566646
rect 348160 433401 348188 568142
rect 348252 456521 348280 576166
rect 348332 560040 348384 560046
rect 348332 559982 348384 559988
rect 348344 559570 348372 559982
rect 348332 559564 348384 559570
rect 348332 559506 348384 559512
rect 348330 523560 348386 523569
rect 348330 523495 348386 523504
rect 348238 456512 348294 456521
rect 348238 456447 348294 456456
rect 348146 433392 348202 433401
rect 348146 433327 348202 433336
rect 348068 402946 348188 402974
rect 348160 396681 348188 402946
rect 348146 396672 348202 396681
rect 348146 396607 348202 396616
rect 348054 390688 348110 390697
rect 348054 390623 348110 390632
rect 347962 377088 348018 377097
rect 347962 377023 348018 377032
rect 347962 368520 348018 368529
rect 347962 368455 348018 368464
rect 347870 276040 347926 276049
rect 347870 275975 347926 275984
rect 347780 184884 347832 184890
rect 347780 184826 347832 184832
rect 347504 184068 347556 184074
rect 347504 184010 347556 184016
rect 347884 180266 347912 275975
rect 347872 180260 347924 180266
rect 347872 180202 347924 180208
rect 346584 179104 346636 179110
rect 346584 179046 346636 179052
rect 346400 164008 346452 164014
rect 346400 163950 346452 163956
rect 345032 149926 345322 149954
rect 346596 149940 346624 179046
rect 347976 170474 348004 368455
rect 348068 191486 348096 390623
rect 348344 296041 348372 523495
rect 348330 296032 348386 296041
rect 348330 295967 348386 295976
rect 348436 295390 348464 587114
rect 348700 586968 348752 586974
rect 348700 586910 348752 586916
rect 348516 586832 348568 586838
rect 348516 586774 348568 586780
rect 348528 488918 348556 586774
rect 348608 586560 348660 586566
rect 348608 586502 348660 586508
rect 348620 494018 348648 586502
rect 348712 498574 348740 586910
rect 348804 586022 348832 661030
rect 348792 586016 348844 586022
rect 348792 585958 348844 585964
rect 349172 584662 349200 669151
rect 351196 650690 351224 674970
rect 351184 650684 351236 650690
rect 351184 650626 351236 650632
rect 358084 640348 358136 640354
rect 358084 640290 358136 640296
rect 350446 609376 350502 609385
rect 350446 609311 350502 609320
rect 350460 608666 350488 609311
rect 350448 608660 350500 608666
rect 350448 608602 350500 608608
rect 349250 607744 349306 607753
rect 349250 607679 349306 607688
rect 349160 584656 349212 584662
rect 349160 584598 349212 584604
rect 349264 584458 349292 607679
rect 350446 606384 350502 606393
rect 350446 606319 350502 606328
rect 350460 605878 350488 606319
rect 350448 605872 350500 605878
rect 350448 605814 350500 605820
rect 350446 604888 350502 604897
rect 350446 604823 350502 604832
rect 350460 604518 350488 604823
rect 350448 604512 350500 604518
rect 350448 604454 350500 604460
rect 349342 603664 349398 603673
rect 349342 603599 349398 603608
rect 349356 589150 349384 603599
rect 349344 589144 349396 589150
rect 349344 589086 349396 589092
rect 350540 587376 350592 587382
rect 350540 587318 350592 587324
rect 349712 585948 349764 585954
rect 349712 585890 349764 585896
rect 349252 584452 349304 584458
rect 349252 584394 349304 584400
rect 349620 583024 349672 583030
rect 349620 582966 349672 582972
rect 349252 581936 349304 581942
rect 349252 581878 349304 581884
rect 349160 573436 349212 573442
rect 349160 573378 349212 573384
rect 349172 541521 349200 573378
rect 349158 541512 349214 541521
rect 349158 541447 349214 541456
rect 348700 498568 348752 498574
rect 348700 498510 348752 498516
rect 349160 498568 349212 498574
rect 349160 498510 349212 498516
rect 348608 494012 348660 494018
rect 348608 493954 348660 493960
rect 348976 491700 349028 491706
rect 348976 491642 349028 491648
rect 348516 488912 348568 488918
rect 348516 488854 348568 488860
rect 348882 433256 348938 433265
rect 348882 433191 348938 433200
rect 348516 397316 348568 397322
rect 348516 397258 348568 397264
rect 348424 295384 348476 295390
rect 348424 295326 348476 295332
rect 348424 282056 348476 282062
rect 348424 281998 348476 282004
rect 348056 191480 348108 191486
rect 348056 191422 348108 191428
rect 347964 170468 348016 170474
rect 347964 170410 348016 170416
rect 348436 155854 348464 281998
rect 348528 199442 348556 397258
rect 348896 389434 348924 433191
rect 348884 389428 348936 389434
rect 348884 389370 348936 389376
rect 348884 388476 348936 388482
rect 348884 388418 348936 388424
rect 348792 358556 348844 358562
rect 348792 358498 348844 358504
rect 348804 249762 348832 358498
rect 348896 276078 348924 388418
rect 348988 349858 349016 491642
rect 349172 489841 349200 498510
rect 349158 489832 349214 489841
rect 349158 489767 349214 489776
rect 349068 456136 349120 456142
rect 349068 456078 349120 456084
rect 348976 349852 349028 349858
rect 348976 349794 349028 349800
rect 348976 294092 349028 294098
rect 348976 294034 349028 294040
rect 348884 276072 348936 276078
rect 348884 276014 348936 276020
rect 348884 269068 348936 269074
rect 348884 269010 348936 269016
rect 348792 249756 348844 249762
rect 348792 249698 348844 249704
rect 348608 247104 348660 247110
rect 348608 247046 348660 247052
rect 348620 199510 348648 247046
rect 348896 244934 348924 269010
rect 348988 269006 349016 294034
rect 348976 269000 349028 269006
rect 348976 268942 349028 268948
rect 348976 268864 349028 268870
rect 348976 268806 349028 268812
rect 348988 262206 349016 268806
rect 348976 262200 349028 262206
rect 348976 262142 349028 262148
rect 348976 260840 349028 260846
rect 348976 260782 349028 260788
rect 348884 244928 348936 244934
rect 348884 244870 348936 244876
rect 348792 223916 348844 223922
rect 348792 223858 348844 223864
rect 348700 218068 348752 218074
rect 348700 218010 348752 218016
rect 348712 200297 348740 218010
rect 348698 200288 348754 200297
rect 348698 200223 348754 200232
rect 348804 199646 348832 223858
rect 348988 218142 349016 260782
rect 349080 233918 349108 456078
rect 349264 347041 349292 581878
rect 349344 573640 349396 573646
rect 349344 573582 349396 573588
rect 349356 451761 349384 573582
rect 349528 566636 349580 566642
rect 349528 566578 349580 566584
rect 349436 566500 349488 566506
rect 349436 566442 349488 566448
rect 349448 558210 349476 566442
rect 349436 558204 349488 558210
rect 349436 558146 349488 558152
rect 349436 554736 349488 554742
rect 349436 554678 349488 554684
rect 349448 554441 349476 554678
rect 349434 554432 349490 554441
rect 349434 554367 349490 554376
rect 349434 532128 349490 532137
rect 349434 532063 349490 532072
rect 349448 531350 349476 532063
rect 349436 531344 349488 531350
rect 349436 531286 349488 531292
rect 349436 494012 349488 494018
rect 349436 493954 349488 493960
rect 349342 451752 349398 451761
rect 349342 451687 349398 451696
rect 349250 347032 349306 347041
rect 349250 346967 349306 346976
rect 349158 299432 349214 299441
rect 349158 299367 349214 299376
rect 349172 282062 349200 299367
rect 349448 296721 349476 493954
rect 349540 409601 349568 566578
rect 349632 500041 349660 582966
rect 349618 500032 349674 500041
rect 349618 499967 349674 499976
rect 349620 488912 349672 488918
rect 349620 488854 349672 488860
rect 349526 409592 349582 409601
rect 349526 409527 349582 409536
rect 349528 389428 349580 389434
rect 349528 389370 349580 389376
rect 349434 296712 349490 296721
rect 349434 296647 349490 296656
rect 349252 295384 349304 295390
rect 349252 295326 349304 295332
rect 349160 282056 349212 282062
rect 349160 281998 349212 282004
rect 349160 269000 349212 269006
rect 349160 268942 349212 268948
rect 349172 260846 349200 268942
rect 349264 262721 349292 295326
rect 349344 286272 349396 286278
rect 349344 286214 349396 286220
rect 349356 279721 349384 286214
rect 349342 279712 349398 279721
rect 349342 279647 349398 279656
rect 349540 268870 349568 389370
rect 349632 336161 349660 488854
rect 349724 470801 349752 585890
rect 350356 576156 350408 576162
rect 350356 576098 350408 576104
rect 349896 574932 349948 574938
rect 349896 574874 349948 574880
rect 349804 558204 349856 558210
rect 349804 558146 349856 558152
rect 349710 470792 349766 470801
rect 349710 470727 349766 470736
rect 349710 456920 349766 456929
rect 349710 456855 349766 456864
rect 349618 336152 349674 336161
rect 349618 336087 349674 336096
rect 349618 280528 349674 280537
rect 349618 280463 349674 280472
rect 349528 268864 349580 268870
rect 349528 268806 349580 268812
rect 349434 262848 349490 262857
rect 349434 262783 349490 262792
rect 349250 262712 349306 262721
rect 349250 262647 349306 262656
rect 349448 262274 349476 262783
rect 349436 262268 349488 262274
rect 349436 262210 349488 262216
rect 349252 262200 349304 262206
rect 349252 262142 349304 262148
rect 349160 260840 349212 260846
rect 349160 260782 349212 260788
rect 349068 233912 349120 233918
rect 349068 233854 349120 233860
rect 349158 233880 349214 233889
rect 349158 233815 349214 233824
rect 349068 233776 349120 233782
rect 349068 233718 349120 233724
rect 348976 218136 349028 218142
rect 348976 218078 349028 218084
rect 348976 212492 349028 212498
rect 348976 212434 349028 212440
rect 348988 206174 349016 212434
rect 349080 212430 349108 233718
rect 349172 223922 349200 233815
rect 349160 223916 349212 223922
rect 349160 223858 349212 223864
rect 349160 218136 349212 218142
rect 349160 218078 349212 218084
rect 349068 212424 349120 212430
rect 349068 212366 349120 212372
rect 348976 206168 349028 206174
rect 348976 206110 349028 206116
rect 349172 204898 349200 218078
rect 348896 204870 349200 204898
rect 348792 199640 348844 199646
rect 348792 199582 348844 199588
rect 348608 199504 348660 199510
rect 348608 199446 348660 199452
rect 348516 199436 348568 199442
rect 348516 199378 348568 199384
rect 348698 198928 348754 198937
rect 348698 198863 348754 198872
rect 348424 155848 348476 155854
rect 348424 155790 348476 155796
rect 348712 153202 348740 198863
rect 348896 183530 348924 204870
rect 349068 200796 349120 200802
rect 349068 200738 349120 200744
rect 348976 199436 349028 199442
rect 348976 199378 349028 199384
rect 348988 195498 349016 199378
rect 349080 197878 349108 200738
rect 349068 197872 349120 197878
rect 349068 197814 349120 197820
rect 348976 195492 349028 195498
rect 348976 195434 349028 195440
rect 349264 192846 349292 262142
rect 349526 258768 349582 258777
rect 349526 258703 349582 258712
rect 349540 258126 349568 258703
rect 349528 258120 349580 258126
rect 349528 258062 349580 258068
rect 349344 249756 349396 249762
rect 349344 249698 349396 249704
rect 349356 212498 349384 249698
rect 349436 233912 349488 233918
rect 349436 233854 349488 233860
rect 349448 218074 349476 233854
rect 349436 218068 349488 218074
rect 349436 218010 349488 218016
rect 349344 212492 349396 212498
rect 349344 212434 349396 212440
rect 349526 210080 349582 210089
rect 349526 210015 349582 210024
rect 349342 202328 349398 202337
rect 349342 202263 349398 202272
rect 349252 192840 349304 192846
rect 349252 192782 349304 192788
rect 348884 183524 348936 183530
rect 348884 183466 348936 183472
rect 349356 175030 349384 202263
rect 349540 187270 349568 210015
rect 349632 190262 349660 280463
rect 349724 257961 349752 456855
rect 349816 455841 349844 558146
rect 349908 521801 349936 574874
rect 350264 566772 350316 566778
rect 350264 566714 350316 566720
rect 350170 547088 350226 547097
rect 350170 547023 350226 547032
rect 350184 546582 350212 547023
rect 350172 546576 350224 546582
rect 350172 546518 350224 546524
rect 350170 533488 350226 533497
rect 350170 533423 350226 533432
rect 350184 532846 350212 533423
rect 350172 532840 350224 532846
rect 350172 532782 350224 532788
rect 349894 521792 349950 521801
rect 349894 521727 349950 521736
rect 350080 521212 350132 521218
rect 350080 521154 350132 521160
rect 350092 518894 350120 521154
rect 350092 518866 350212 518894
rect 350078 516624 350134 516633
rect 350078 516559 350134 516568
rect 350092 516254 350120 516559
rect 350080 516248 350132 516254
rect 350080 516190 350132 516196
rect 350078 513496 350134 513505
rect 350078 513431 350080 513440
rect 350132 513431 350134 513440
rect 350080 513402 350132 513408
rect 349986 506968 350042 506977
rect 349986 506903 350042 506912
rect 350000 506598 350028 506903
rect 349988 506592 350040 506598
rect 349988 506534 350040 506540
rect 349896 506524 349948 506530
rect 349896 506466 349948 506472
rect 349908 491706 349936 506466
rect 350078 505608 350134 505617
rect 350078 505543 350134 505552
rect 350092 505170 350120 505543
rect 350080 505164 350132 505170
rect 350080 505106 350132 505112
rect 349896 491700 349948 491706
rect 349896 491642 349948 491648
rect 349986 485208 350042 485217
rect 349986 485143 350042 485152
rect 350000 484430 350028 485143
rect 349988 484424 350040 484430
rect 349988 484366 350040 484372
rect 350078 480720 350134 480729
rect 350078 480655 350134 480664
rect 350092 480350 350120 480655
rect 350080 480344 350132 480350
rect 350080 480286 350132 480292
rect 350078 476504 350134 476513
rect 350078 476439 350134 476448
rect 350092 476202 350120 476439
rect 350080 476196 350132 476202
rect 350080 476138 350132 476144
rect 350080 466404 350132 466410
rect 350080 466346 350132 466352
rect 350092 466041 350120 466346
rect 350078 466032 350134 466041
rect 350078 465967 350134 465976
rect 350078 462904 350134 462913
rect 350078 462839 350134 462848
rect 350092 462466 350120 462839
rect 350080 462460 350132 462466
rect 350080 462402 350132 462408
rect 350078 461408 350134 461417
rect 350078 461343 350134 461352
rect 350092 460970 350120 461343
rect 350080 460964 350132 460970
rect 350080 460906 350132 460912
rect 349802 455832 349858 455841
rect 349802 455767 349858 455776
rect 350078 445904 350134 445913
rect 350078 445839 350134 445848
rect 350092 445806 350120 445839
rect 350080 445800 350132 445806
rect 350080 445742 350132 445748
rect 350078 437880 350134 437889
rect 350078 437815 350134 437824
rect 350092 437510 350120 437815
rect 350080 437504 350132 437510
rect 350080 437446 350132 437452
rect 350078 430944 350134 430953
rect 350078 430879 350134 430888
rect 350092 430642 350120 430879
rect 350080 430636 350132 430642
rect 350080 430578 350132 430584
rect 350078 421288 350134 421297
rect 350078 421223 350134 421232
rect 350092 421054 350120 421223
rect 350080 421048 350132 421054
rect 350080 420990 350132 420996
rect 350078 404968 350134 404977
rect 350078 404903 350134 404912
rect 350092 404394 350120 404903
rect 350080 404388 350132 404394
rect 350080 404330 350132 404336
rect 350078 395448 350134 395457
rect 350078 395383 350134 395392
rect 349802 394904 349858 394913
rect 349802 394839 349858 394848
rect 349816 394806 349844 394839
rect 349804 394800 349856 394806
rect 349804 394742 349856 394748
rect 350092 394738 350120 395383
rect 350080 394732 350132 394738
rect 350080 394674 350132 394680
rect 350078 391368 350134 391377
rect 350078 391303 350134 391312
rect 350092 390590 350120 391303
rect 350080 390584 350132 390590
rect 350080 390526 350132 390532
rect 350080 390108 350132 390114
rect 350080 390050 350132 390056
rect 350092 385014 350120 390050
rect 350080 385008 350132 385014
rect 350080 384950 350132 384956
rect 349986 356688 350042 356697
rect 349986 356623 350042 356632
rect 350000 356114 350028 356623
rect 349988 356108 350040 356114
rect 349988 356050 350040 356056
rect 350184 350674 350212 518866
rect 350172 350668 350224 350674
rect 350172 350610 350224 350616
rect 349804 349852 349856 349858
rect 349804 349794 349856 349800
rect 349816 302258 349844 349794
rect 350170 344040 350226 344049
rect 350170 343975 350226 343984
rect 350184 343670 350212 343975
rect 350172 343664 350224 343670
rect 350172 343606 350224 343612
rect 349894 331256 349950 331265
rect 349894 331191 349950 331200
rect 349908 305046 349936 331191
rect 350172 320136 350224 320142
rect 350172 320078 350224 320084
rect 350184 319161 350212 320078
rect 350170 319152 350226 319161
rect 350170 319087 350226 319096
rect 350170 315208 350226 315217
rect 350170 315143 350226 315152
rect 350184 314702 350212 315143
rect 350172 314696 350224 314702
rect 350172 314638 350224 314644
rect 350172 309800 350224 309806
rect 350172 309742 350224 309748
rect 349896 305040 349948 305046
rect 349896 304982 349948 304988
rect 349894 302968 349950 302977
rect 349894 302903 349950 302912
rect 349804 302252 349856 302258
rect 349804 302194 349856 302200
rect 349804 285728 349856 285734
rect 349804 285670 349856 285676
rect 349710 257952 349766 257961
rect 349710 257887 349766 257896
rect 349712 212424 349764 212430
rect 349712 212366 349764 212372
rect 349724 200569 349752 212366
rect 349710 200560 349766 200569
rect 349710 200495 349766 200504
rect 349816 197266 349844 285670
rect 349908 238066 349936 302903
rect 350080 300824 350132 300830
rect 350080 300766 350132 300772
rect 350092 298042 350120 300766
rect 350080 298036 350132 298042
rect 350080 297978 350132 297984
rect 350080 295520 350132 295526
rect 350080 295462 350132 295468
rect 350092 288561 350120 295462
rect 350078 288552 350134 288561
rect 350078 288487 350134 288496
rect 350184 277394 350212 309742
rect 350276 295526 350304 566714
rect 350368 493921 350396 576098
rect 350446 551168 350502 551177
rect 350446 551103 350502 551112
rect 350460 550662 350488 551103
rect 350448 550656 350500 550662
rect 350448 550598 350500 550604
rect 350446 546544 350502 546553
rect 350446 546479 350448 546488
rect 350500 546479 350502 546488
rect 350448 546450 350500 546456
rect 350446 543008 350502 543017
rect 350446 542943 350502 542952
rect 350460 542434 350488 542943
rect 350448 542428 350500 542434
rect 350448 542370 350500 542376
rect 350446 538384 350502 538393
rect 350446 538319 350502 538328
rect 350460 538286 350488 538319
rect 350448 538280 350500 538286
rect 350448 538222 350500 538228
rect 350446 536888 350502 536897
rect 350446 536823 350448 536832
rect 350500 536823 350502 536832
rect 350448 536794 350500 536800
rect 350446 534712 350502 534721
rect 350446 534647 350502 534656
rect 350460 534138 350488 534647
rect 350448 534132 350500 534138
rect 350448 534074 350500 534080
rect 350446 532808 350502 532817
rect 350446 532743 350448 532752
rect 350500 532743 350502 532752
rect 350448 532714 350500 532720
rect 350446 530768 350502 530777
rect 350446 530703 350502 530712
rect 350460 529990 350488 530703
rect 350448 529984 350500 529990
rect 350448 529926 350500 529932
rect 350446 527232 350502 527241
rect 350446 527167 350448 527176
rect 350500 527167 350502 527176
rect 350448 527138 350500 527144
rect 350446 526008 350502 526017
rect 350446 525943 350448 525952
rect 350500 525943 350502 525952
rect 350448 525914 350500 525920
rect 350446 523288 350502 523297
rect 350446 523223 350502 523232
rect 350460 523054 350488 523223
rect 350448 523048 350500 523054
rect 350552 523025 350580 587318
rect 354772 587308 354824 587314
rect 354772 587250 354824 587256
rect 352012 587240 352064 587246
rect 352012 587182 352064 587188
rect 350632 587104 350684 587110
rect 350632 587046 350684 587052
rect 350448 522990 350500 522996
rect 350538 523016 350594 523025
rect 350538 522951 350594 522960
rect 350446 517576 350502 517585
rect 350446 517511 350448 517520
rect 350500 517511 350502 517520
rect 350448 517482 350500 517488
rect 350446 516352 350502 516361
rect 350446 516287 350448 516296
rect 350500 516287 350502 516296
rect 350448 516258 350500 516264
rect 350446 513768 350502 513777
rect 350446 513703 350502 513712
rect 350460 513398 350488 513703
rect 350448 513392 350500 513398
rect 350448 513334 350500 513340
rect 350448 511964 350500 511970
rect 350448 511906 350500 511912
rect 350460 511601 350488 511906
rect 350446 511592 350502 511601
rect 350446 511527 350502 511536
rect 350448 509244 350500 509250
rect 350448 509186 350500 509192
rect 350460 508881 350488 509186
rect 350446 508872 350502 508881
rect 350446 508807 350502 508816
rect 350448 506456 350500 506462
rect 350448 506398 350500 506404
rect 350460 505481 350488 506398
rect 350446 505472 350502 505481
rect 350446 505407 350502 505416
rect 350446 503840 350502 503849
rect 350446 503775 350502 503784
rect 350460 503742 350488 503775
rect 350448 503736 350500 503742
rect 350448 503678 350500 503684
rect 350446 500168 350502 500177
rect 350446 500103 350502 500112
rect 350460 499594 350488 500103
rect 350448 499588 350500 499594
rect 350448 499530 350500 499536
rect 350446 498264 350502 498273
rect 350446 498199 350448 498208
rect 350500 498199 350502 498208
rect 350448 498170 350500 498176
rect 350446 495544 350502 495553
rect 350446 495479 350448 495488
rect 350500 495479 350502 495488
rect 350448 495450 350500 495456
rect 350446 494592 350502 494601
rect 350446 494527 350448 494536
rect 350500 494527 350502 494536
rect 350448 494498 350500 494504
rect 350354 493912 350410 493921
rect 350354 493847 350410 493856
rect 350354 492008 350410 492017
rect 350354 491943 350410 491952
rect 350368 491434 350396 491943
rect 350446 491464 350502 491473
rect 350356 491428 350408 491434
rect 350446 491399 350502 491408
rect 350356 491370 350408 491376
rect 350460 491366 350488 491399
rect 350448 491360 350500 491366
rect 350448 491302 350500 491308
rect 350356 491292 350408 491298
rect 350356 491234 350408 491240
rect 350368 390114 350396 491234
rect 350446 490104 350502 490113
rect 350446 490039 350502 490048
rect 350460 490006 350488 490039
rect 350448 490000 350500 490006
rect 350448 489942 350500 489948
rect 350448 488504 350500 488510
rect 350448 488446 350500 488452
rect 350460 487801 350488 488446
rect 350446 487792 350502 487801
rect 350446 487727 350502 487736
rect 350446 483168 350502 483177
rect 350446 483103 350502 483112
rect 350460 483070 350488 483103
rect 350448 483064 350500 483070
rect 350448 483006 350500 483012
rect 350448 481704 350500 481710
rect 350446 481672 350448 481681
rect 350500 481672 350502 481681
rect 350446 481607 350502 481616
rect 350446 480312 350502 480321
rect 350446 480247 350448 480256
rect 350500 480247 350502 480256
rect 350448 480218 350500 480224
rect 350446 476232 350502 476241
rect 350446 476167 350502 476176
rect 350460 476134 350488 476167
rect 350448 476128 350500 476134
rect 350448 476070 350500 476076
rect 350446 473512 350502 473521
rect 350446 473447 350502 473456
rect 350460 473414 350488 473447
rect 350448 473408 350500 473414
rect 350448 473350 350500 473356
rect 350446 466576 350502 466585
rect 350446 466511 350502 466520
rect 350460 466478 350488 466511
rect 350448 466472 350500 466478
rect 350448 466414 350500 466420
rect 350446 465216 350502 465225
rect 350446 465151 350502 465160
rect 350460 465118 350488 465151
rect 350448 465112 350500 465118
rect 350448 465054 350500 465060
rect 350446 462496 350502 462505
rect 350446 462431 350502 462440
rect 350460 462398 350488 462431
rect 350448 462392 350500 462398
rect 350448 462334 350500 462340
rect 350446 461136 350502 461145
rect 350446 461071 350502 461080
rect 350460 461038 350488 461071
rect 350448 461032 350500 461038
rect 350448 460974 350500 460980
rect 350446 459640 350502 459649
rect 350446 459575 350448 459584
rect 350500 459575 350502 459584
rect 350448 459546 350500 459552
rect 350446 457328 350502 457337
rect 350446 457263 350448 457272
rect 350500 457263 350502 457272
rect 350448 457234 350500 457240
rect 350446 454200 350502 454209
rect 350446 454135 350448 454144
rect 350500 454135 350502 454144
rect 350448 454106 350500 454112
rect 350446 451888 350502 451897
rect 350446 451823 350502 451832
rect 350460 451314 350488 451823
rect 350448 451308 350500 451314
rect 350448 451250 350500 451256
rect 350448 451172 350500 451178
rect 350448 451114 350500 451120
rect 350460 451081 350488 451114
rect 350446 451072 350502 451081
rect 350446 451007 350502 451016
rect 350446 449984 350502 449993
rect 350446 449919 350448 449928
rect 350500 449919 350502 449928
rect 350448 449890 350500 449896
rect 350446 447808 350502 447817
rect 350446 447743 350502 447752
rect 350460 447166 350488 447743
rect 350448 447160 350500 447166
rect 350448 447102 350500 447108
rect 350446 446448 350502 446457
rect 350446 446383 350502 446392
rect 350460 445874 350488 446383
rect 350448 445868 350500 445874
rect 350448 445810 350500 445816
rect 350448 445732 350500 445738
rect 350448 445674 350500 445680
rect 350460 445641 350488 445674
rect 350446 445632 350502 445641
rect 350446 445567 350502 445576
rect 350446 441688 350502 441697
rect 350446 441623 350448 441632
rect 350500 441623 350502 441632
rect 350448 441594 350500 441600
rect 350446 440328 350502 440337
rect 350446 440263 350448 440272
rect 350500 440263 350502 440272
rect 350448 440234 350500 440240
rect 350448 437436 350500 437442
rect 350448 437378 350500 437384
rect 350460 436801 350488 437378
rect 350446 436792 350502 436801
rect 350446 436727 350502 436736
rect 350448 434784 350500 434790
rect 350446 434752 350448 434761
rect 350500 434752 350502 434761
rect 350446 434687 350502 434696
rect 350448 430704 350500 430710
rect 350446 430672 350448 430681
rect 350500 430672 350502 430681
rect 350446 430607 350502 430616
rect 350446 427952 350502 427961
rect 350446 427887 350502 427896
rect 350460 427854 350488 427887
rect 350448 427848 350500 427854
rect 350448 427790 350500 427796
rect 350446 426592 350502 426601
rect 350446 426527 350502 426536
rect 350460 426494 350488 426527
rect 350448 426488 350500 426494
rect 350448 426430 350500 426436
rect 350446 425368 350502 425377
rect 350446 425303 350502 425312
rect 350460 425134 350488 425303
rect 350448 425128 350500 425134
rect 350448 425070 350500 425076
rect 350446 422376 350502 422385
rect 350446 422311 350448 422320
rect 350500 422311 350502 422320
rect 350448 422282 350500 422288
rect 350446 421016 350502 421025
rect 350446 420951 350448 420960
rect 350500 420951 350502 420960
rect 350448 420922 350500 420928
rect 350446 419656 350502 419665
rect 350446 419591 350502 419600
rect 350460 419558 350488 419591
rect 350448 419552 350500 419558
rect 350448 419494 350500 419500
rect 350446 418432 350502 418441
rect 350446 418367 350502 418376
rect 350460 418198 350488 418367
rect 350448 418192 350500 418198
rect 350448 418134 350500 418140
rect 350446 416936 350502 416945
rect 350446 416871 350502 416880
rect 350460 416838 350488 416871
rect 350448 416832 350500 416838
rect 350448 416774 350500 416780
rect 350446 414488 350502 414497
rect 350446 414423 350448 414432
rect 350500 414423 350502 414432
rect 350448 414394 350500 414400
rect 350446 414080 350502 414089
rect 350446 414015 350448 414024
rect 350500 414015 350502 414024
rect 350448 413986 350500 413992
rect 350446 411360 350502 411369
rect 350446 411295 350448 411304
rect 350500 411295 350502 411304
rect 350448 411266 350500 411272
rect 350446 407280 350502 407289
rect 350446 407215 350448 407224
rect 350500 407215 350502 407224
rect 350448 407186 350500 407192
rect 350446 404560 350502 404569
rect 350446 404495 350502 404504
rect 350460 404462 350488 404495
rect 350448 404456 350500 404462
rect 350448 404398 350500 404404
rect 350446 400344 350502 400353
rect 350446 400279 350502 400288
rect 350460 400246 350488 400279
rect 350448 400240 350500 400246
rect 350448 400182 350500 400188
rect 350446 399528 350502 399537
rect 350446 399463 350502 399472
rect 350460 398886 350488 399463
rect 350448 398880 350500 398886
rect 350448 398822 350500 398828
rect 350446 397624 350502 397633
rect 350446 397559 350502 397568
rect 350460 397526 350488 397559
rect 350448 397520 350500 397526
rect 350448 397462 350500 397468
rect 350446 396808 350502 396817
rect 350446 396743 350502 396752
rect 350460 396098 350488 396743
rect 350448 396092 350500 396098
rect 350448 396034 350500 396040
rect 350448 394664 350500 394670
rect 350446 394632 350448 394641
rect 350500 394632 350502 394641
rect 350446 394567 350502 394576
rect 350446 392048 350502 392057
rect 350446 391983 350448 391992
rect 350500 391983 350502 391992
rect 350448 391954 350500 391960
rect 350448 390516 350500 390522
rect 350448 390458 350500 390464
rect 350356 390108 350408 390114
rect 350356 390050 350408 390056
rect 350354 390008 350410 390017
rect 350354 389943 350410 389952
rect 350368 389230 350396 389943
rect 350460 389881 350488 390458
rect 350446 389872 350502 389881
rect 350446 389807 350502 389816
rect 350356 389224 350408 389230
rect 350356 389166 350408 389172
rect 350448 387864 350500 387870
rect 350446 387832 350448 387841
rect 350500 387832 350502 387841
rect 350356 387796 350408 387802
rect 350446 387767 350502 387776
rect 350356 387738 350408 387744
rect 350368 387161 350396 387738
rect 350354 387152 350410 387161
rect 350354 387087 350410 387096
rect 350446 382392 350502 382401
rect 350446 382327 350502 382336
rect 350460 382294 350488 382327
rect 350448 382288 350500 382294
rect 350448 382230 350500 382236
rect 350354 381440 350410 381449
rect 350354 381375 350410 381384
rect 350368 381002 350396 381375
rect 350446 381032 350502 381041
rect 350356 380996 350408 381002
rect 350446 380967 350502 380976
rect 350356 380938 350408 380944
rect 350460 380934 350488 380967
rect 350448 380928 350500 380934
rect 350448 380870 350500 380876
rect 350446 377224 350502 377233
rect 350446 377159 350502 377168
rect 350460 376786 350488 377159
rect 350448 376780 350500 376786
rect 350448 376722 350500 376728
rect 350354 375864 350410 375873
rect 350354 375799 350410 375808
rect 350368 375426 350396 375799
rect 350356 375420 350408 375426
rect 350356 375362 350408 375368
rect 350448 375352 350500 375358
rect 350448 375294 350500 375300
rect 350460 374921 350488 375294
rect 350446 374912 350502 374921
rect 350446 374847 350502 374856
rect 350446 372872 350502 372881
rect 350446 372807 350502 372816
rect 350460 372638 350488 372807
rect 350448 372632 350500 372638
rect 350448 372574 350500 372580
rect 350446 371376 350502 371385
rect 350446 371311 350502 371320
rect 350460 371278 350488 371311
rect 350448 371272 350500 371278
rect 350448 371214 350500 371220
rect 350448 365696 350500 365702
rect 350448 365638 350500 365644
rect 350460 365401 350488 365638
rect 350446 365392 350502 365401
rect 350446 365327 350502 365336
rect 350446 364440 350502 364449
rect 350446 364375 350448 364384
rect 350500 364375 350502 364384
rect 350448 364346 350500 364352
rect 350446 358048 350502 358057
rect 350446 357983 350448 357992
rect 350500 357983 350502 357992
rect 350448 357954 350500 357960
rect 350448 356040 350500 356046
rect 350448 355982 350500 355988
rect 350460 355881 350488 355982
rect 350446 355872 350502 355881
rect 350446 355807 350502 355816
rect 350446 354784 350502 354793
rect 350446 354719 350448 354728
rect 350500 354719 350502 354728
rect 350448 354690 350500 354696
rect 350356 351960 350408 351966
rect 350356 351902 350408 351908
rect 350368 350010 350396 351902
rect 350446 350704 350502 350713
rect 350446 350639 350502 350648
rect 350460 350606 350488 350639
rect 350448 350600 350500 350606
rect 350448 350542 350500 350548
rect 350368 349982 350488 350010
rect 350354 349888 350410 349897
rect 350354 349823 350410 349832
rect 350368 349178 350396 349823
rect 350460 349466 350488 349982
rect 350460 349438 350580 349466
rect 350446 349344 350502 349353
rect 350446 349279 350502 349288
rect 350460 349246 350488 349279
rect 350448 349240 350500 349246
rect 350448 349182 350500 349188
rect 350356 349172 350408 349178
rect 350356 349114 350408 349120
rect 350552 349058 350580 349438
rect 350460 349030 350580 349058
rect 350354 345808 350410 345817
rect 350354 345743 350410 345752
rect 350368 345506 350396 345743
rect 350356 345500 350408 345506
rect 350356 345442 350408 345448
rect 350354 344448 350410 344457
rect 350354 344383 350410 344392
rect 350368 343738 350396 344383
rect 350356 343732 350408 343738
rect 350356 343674 350408 343680
rect 350356 343596 350408 343602
rect 350356 343538 350408 343544
rect 350368 342281 350396 343538
rect 350354 342272 350410 342281
rect 350354 342207 350410 342216
rect 350354 338192 350410 338201
rect 350354 338127 350356 338136
rect 350408 338127 350410 338136
rect 350356 338098 350408 338104
rect 350354 334112 350410 334121
rect 350354 334047 350410 334056
rect 350368 334014 350396 334047
rect 350356 334008 350408 334014
rect 350356 333950 350408 333956
rect 350354 332752 350410 332761
rect 350354 332687 350410 332696
rect 350368 332654 350396 332687
rect 350356 332648 350408 332654
rect 350356 332590 350408 332596
rect 350354 329896 350410 329905
rect 350354 329831 350356 329840
rect 350408 329831 350410 329840
rect 350356 329802 350408 329808
rect 350354 328944 350410 328953
rect 350354 328879 350410 328888
rect 350368 328506 350396 328879
rect 350356 328500 350408 328506
rect 350356 328442 350408 328448
rect 350354 325816 350410 325825
rect 350354 325751 350410 325760
rect 350368 325718 350396 325751
rect 350356 325712 350408 325718
rect 350356 325654 350408 325660
rect 350354 321736 350410 321745
rect 350354 321671 350410 321680
rect 350368 321638 350396 321671
rect 350356 321632 350408 321638
rect 350356 321574 350408 321580
rect 350354 320648 350410 320657
rect 350354 320583 350410 320592
rect 350368 320210 350396 320583
rect 350356 320204 350408 320210
rect 350356 320146 350408 320152
rect 350354 319288 350410 319297
rect 350354 319223 350410 319232
rect 350368 318850 350396 319223
rect 350356 318844 350408 318850
rect 350356 318786 350408 318792
rect 350354 317792 350410 317801
rect 350354 317727 350410 317736
rect 350368 317490 350396 317727
rect 350356 317484 350408 317490
rect 350356 317426 350408 317432
rect 350356 315988 350408 315994
rect 350356 315930 350408 315936
rect 350368 315081 350396 315930
rect 350354 315072 350410 315081
rect 350354 315007 350410 315016
rect 350354 312352 350410 312361
rect 350354 312287 350410 312296
rect 350368 311914 350396 312287
rect 350356 311908 350408 311914
rect 350356 311850 350408 311856
rect 350354 311128 350410 311137
rect 350354 311063 350410 311072
rect 350368 310554 350396 311063
rect 350356 310548 350408 310554
rect 350356 310490 350408 310496
rect 350354 308408 350410 308417
rect 350354 308343 350410 308352
rect 350368 307834 350396 308343
rect 350356 307828 350408 307834
rect 350356 307770 350408 307776
rect 350354 304328 350410 304337
rect 350354 304263 350410 304272
rect 350368 303754 350396 304263
rect 350356 303748 350408 303754
rect 350356 303690 350408 303696
rect 350354 302424 350410 302433
rect 350354 302359 350410 302368
rect 350368 302326 350396 302359
rect 350356 302320 350408 302326
rect 350356 302262 350408 302268
rect 350354 300928 350410 300937
rect 350354 300863 350356 300872
rect 350408 300863 350410 300872
rect 350356 300834 350408 300840
rect 350354 300248 350410 300257
rect 350354 300183 350410 300192
rect 350368 299606 350396 300183
rect 350356 299600 350408 299606
rect 350356 299542 350408 299548
rect 350354 298888 350410 298897
rect 350354 298823 350410 298832
rect 350368 298178 350396 298823
rect 350356 298172 350408 298178
rect 350356 298114 350408 298120
rect 350356 298036 350408 298042
rect 350356 297978 350408 297984
rect 350264 295520 350316 295526
rect 350264 295462 350316 295468
rect 350264 295384 350316 295390
rect 350262 295352 350264 295361
rect 350316 295352 350318 295361
rect 350262 295287 350318 295296
rect 350264 294024 350316 294030
rect 350262 293992 350264 294001
rect 350316 293992 350318 294001
rect 350262 293927 350318 293936
rect 350262 288688 350318 288697
rect 350262 288623 350318 288632
rect 350276 288454 350304 288623
rect 350264 288448 350316 288454
rect 350264 288390 350316 288396
rect 350262 287192 350318 287201
rect 350262 287127 350264 287136
rect 350316 287127 350318 287136
rect 350264 287098 350316 287104
rect 350264 287020 350316 287026
rect 350264 286962 350316 286968
rect 350276 286521 350304 286962
rect 350262 286512 350318 286521
rect 350262 286447 350318 286456
rect 350264 285660 350316 285666
rect 350264 285602 350316 285608
rect 350276 285161 350304 285602
rect 350262 285152 350318 285161
rect 350262 285087 350318 285096
rect 350262 277536 350318 277545
rect 350262 277471 350318 277480
rect 350276 277438 350304 277471
rect 350092 277366 350212 277394
rect 350264 277432 350316 277438
rect 350264 277374 350316 277380
rect 349988 273352 350040 273358
rect 349988 273294 350040 273300
rect 350000 258074 350028 273294
rect 350092 270434 350120 277366
rect 350264 275936 350316 275942
rect 350264 275878 350316 275884
rect 350276 275641 350304 275878
rect 350262 275632 350318 275641
rect 350262 275567 350318 275576
rect 350170 273864 350226 273873
rect 350170 273799 350226 273808
rect 350184 273290 350212 273799
rect 350262 273456 350318 273465
rect 350262 273391 350264 273400
rect 350316 273391 350318 273400
rect 350264 273362 350316 273368
rect 350172 273284 350224 273290
rect 350172 273226 350224 273232
rect 350262 272232 350318 272241
rect 350262 272167 350318 272176
rect 350276 271930 350304 272167
rect 350264 271924 350316 271930
rect 350264 271866 350316 271872
rect 350264 270496 350316 270502
rect 350264 270438 350316 270444
rect 350080 270428 350132 270434
rect 350080 270370 350132 270376
rect 350276 270201 350304 270438
rect 350262 270192 350318 270201
rect 350262 270127 350318 270136
rect 350264 269000 350316 269006
rect 350264 268942 350316 268948
rect 350276 268841 350304 268942
rect 350262 268832 350318 268841
rect 350262 268767 350318 268776
rect 350262 266792 350318 266801
rect 350262 266727 350318 266736
rect 350276 266422 350304 266727
rect 350264 266416 350316 266422
rect 350264 266358 350316 266364
rect 350262 263936 350318 263945
rect 350262 263871 350318 263880
rect 350276 263702 350304 263871
rect 350264 263696 350316 263702
rect 350264 263638 350316 263644
rect 350264 262200 350316 262206
rect 350264 262142 350316 262148
rect 350276 261361 350304 262142
rect 350262 261352 350318 261361
rect 350262 261287 350318 261296
rect 350000 258046 350304 258074
rect 349986 256048 350042 256057
rect 349986 255983 350042 255992
rect 349896 238060 349948 238066
rect 349896 238002 349948 238008
rect 349896 236020 349948 236026
rect 349896 235962 349948 235968
rect 349804 197260 349856 197266
rect 349804 197202 349856 197208
rect 349620 190256 349672 190262
rect 349620 190198 349672 190204
rect 349528 187264 349580 187270
rect 349528 187206 349580 187212
rect 349344 175024 349396 175030
rect 349344 174966 349396 174972
rect 349908 158642 349936 235962
rect 350000 233918 350028 255983
rect 350172 255468 350224 255474
rect 350172 255410 350224 255416
rect 350080 248396 350132 248402
rect 350080 248338 350132 248344
rect 350092 247761 350120 248338
rect 350078 247752 350134 247761
rect 350078 247687 350134 247696
rect 350184 244662 350212 255410
rect 350172 244656 350224 244662
rect 350172 244598 350224 244604
rect 350078 244352 350134 244361
rect 350078 244287 350134 244296
rect 349988 233912 350040 233918
rect 349988 233854 350040 233860
rect 349988 204468 350040 204474
rect 349988 204410 350040 204416
rect 349896 158636 349948 158642
rect 349896 158578 349948 158584
rect 350000 155650 350028 204410
rect 350092 203590 350120 244287
rect 350170 242992 350226 243001
rect 350170 242927 350226 242936
rect 350184 235278 350212 242927
rect 350172 235272 350224 235278
rect 350172 235214 350224 235220
rect 350172 222624 350224 222630
rect 350172 222566 350224 222572
rect 350080 203584 350132 203590
rect 350080 203526 350132 203532
rect 350184 199578 350212 222566
rect 350276 222154 350304 258046
rect 350368 246242 350396 297978
rect 350460 255474 350488 349030
rect 350540 302252 350592 302258
rect 350540 302194 350592 302200
rect 350552 294098 350580 302194
rect 350540 294092 350592 294098
rect 350540 294034 350592 294040
rect 350644 286278 350672 587046
rect 350724 584520 350776 584526
rect 350724 584462 350776 584468
rect 350736 330721 350764 584462
rect 351092 577516 351144 577522
rect 351092 577458 351144 577464
rect 350816 576292 350868 576298
rect 350816 576234 350868 576240
rect 350722 330712 350778 330721
rect 350722 330647 350778 330656
rect 350828 324601 350856 576234
rect 350908 574864 350960 574870
rect 350908 574806 350960 574812
rect 350920 385121 350948 574806
rect 351000 570920 351052 570926
rect 351000 570862 351052 570868
rect 350906 385112 350962 385121
rect 350906 385047 350962 385056
rect 351012 370161 351040 570862
rect 351104 383761 351132 577458
rect 351184 568132 351236 568138
rect 351184 568074 351236 568080
rect 351196 397322 351224 568074
rect 351920 568064 351972 568070
rect 351920 568006 351972 568012
rect 351276 560788 351328 560794
rect 351276 560730 351328 560736
rect 351288 506530 351316 560730
rect 351932 554742 351960 568006
rect 351920 554736 351972 554742
rect 351920 554678 351972 554684
rect 351368 531344 351420 531350
rect 351368 531286 351420 531292
rect 351276 506524 351328 506530
rect 351276 506466 351328 506472
rect 351184 397316 351236 397322
rect 351184 397258 351236 397264
rect 351184 385008 351236 385014
rect 351184 384950 351236 384956
rect 351090 383752 351146 383761
rect 351090 383687 351146 383696
rect 351090 379808 351146 379817
rect 351090 379743 351146 379752
rect 350998 370152 351054 370161
rect 350998 370087 351054 370096
rect 350998 363352 351054 363361
rect 350998 363287 351054 363296
rect 350814 324592 350870 324601
rect 350814 324527 350870 324536
rect 350724 305040 350776 305046
rect 350724 304982 350776 304988
rect 350632 286272 350684 286278
rect 350632 286214 350684 286220
rect 350630 284336 350686 284345
rect 350630 284271 350686 284280
rect 350540 276072 350592 276078
rect 350540 276014 350592 276020
rect 350552 269074 350580 276014
rect 350540 269068 350592 269074
rect 350540 269010 350592 269016
rect 350448 255468 350500 255474
rect 350448 255410 350500 255416
rect 350446 255368 350502 255377
rect 350446 255303 350448 255312
rect 350500 255303 350502 255312
rect 350448 255274 350500 255280
rect 350446 254008 350502 254017
rect 350446 253943 350448 253952
rect 350500 253943 350502 253952
rect 350448 253914 350500 253920
rect 350446 249928 350502 249937
rect 350446 249863 350502 249872
rect 350460 249830 350488 249863
rect 350448 249824 350500 249830
rect 350448 249766 350500 249772
rect 350446 248568 350502 248577
rect 350446 248503 350502 248512
rect 350460 248470 350488 248503
rect 350448 248464 350500 248470
rect 350448 248406 350500 248412
rect 350368 246214 350488 246242
rect 350354 246120 350410 246129
rect 350354 246055 350410 246064
rect 350368 245682 350396 246055
rect 350460 245857 350488 246214
rect 350446 245848 350502 245857
rect 350446 245783 350502 245792
rect 350448 245744 350500 245750
rect 350446 245712 350448 245721
rect 350500 245712 350502 245721
rect 350356 245676 350408 245682
rect 350446 245647 350502 245656
rect 350356 245618 350408 245624
rect 350538 244488 350594 244497
rect 350538 244423 350594 244432
rect 350446 243264 350502 243273
rect 350446 243199 350502 243208
rect 350460 242962 350488 243199
rect 350448 242956 350500 242962
rect 350448 242898 350500 242904
rect 350354 239320 350410 239329
rect 350354 239255 350410 239264
rect 350368 238950 350396 239255
rect 350356 238944 350408 238950
rect 350356 238886 350408 238892
rect 350446 238912 350502 238921
rect 350446 238847 350448 238856
rect 350500 238847 350502 238856
rect 350448 238818 350500 238824
rect 350448 237312 350500 237318
rect 350448 237254 350500 237260
rect 350460 236201 350488 237254
rect 350446 236192 350502 236201
rect 350446 236127 350502 236136
rect 350446 234968 350502 234977
rect 350446 234903 350448 234912
rect 350500 234903 350502 234912
rect 350448 234874 350500 234880
rect 350446 232248 350502 232257
rect 350446 232183 350502 232192
rect 350460 231878 350488 232183
rect 350448 231872 350500 231878
rect 350448 231814 350500 231820
rect 350446 230616 350502 230625
rect 350446 230551 350502 230560
rect 350460 230518 350488 230551
rect 350448 230512 350500 230518
rect 350448 230454 350500 230460
rect 350446 229256 350502 229265
rect 350446 229191 350502 229200
rect 350460 229158 350488 229191
rect 350448 229152 350500 229158
rect 350448 229094 350500 229100
rect 350446 225040 350502 225049
rect 350446 224975 350448 224984
rect 350500 224975 350502 224984
rect 350448 224946 350500 224952
rect 350448 223576 350500 223582
rect 350448 223518 350500 223524
rect 350460 222601 350488 223518
rect 350446 222592 350502 222601
rect 350446 222527 350502 222536
rect 350264 222148 350316 222154
rect 350264 222090 350316 222096
rect 350446 221232 350502 221241
rect 350446 221167 350448 221176
rect 350500 221167 350502 221176
rect 350448 221138 350500 221144
rect 350354 220008 350410 220017
rect 350354 219943 350410 219952
rect 350264 218000 350316 218006
rect 350264 217942 350316 217948
rect 350276 217161 350304 217942
rect 350262 217152 350318 217161
rect 350262 217087 350318 217096
rect 350262 207768 350318 207777
rect 350262 207703 350318 207712
rect 350276 207058 350304 207703
rect 350264 207052 350316 207058
rect 350264 206994 350316 207000
rect 350262 205048 350318 205057
rect 350262 204983 350318 204992
rect 350276 204338 350304 204983
rect 350264 204332 350316 204338
rect 350264 204274 350316 204280
rect 350172 199572 350224 199578
rect 350172 199514 350224 199520
rect 350368 195362 350396 219943
rect 350446 218104 350502 218113
rect 350446 218039 350448 218048
rect 350500 218039 350502 218048
rect 350448 218010 350500 218016
rect 350446 217560 350502 217569
rect 350446 217495 350502 217504
rect 350460 217258 350488 217495
rect 350448 217252 350500 217258
rect 350448 217194 350500 217200
rect 350446 215384 350502 215393
rect 350446 215319 350448 215328
rect 350500 215319 350502 215328
rect 350448 215290 350500 215296
rect 350446 213208 350502 213217
rect 350446 213143 350502 213152
rect 350460 212566 350488 213143
rect 350448 212560 350500 212566
rect 350448 212502 350500 212508
rect 350446 209128 350502 209137
rect 350446 209063 350502 209072
rect 350460 208418 350488 209063
rect 350448 208412 350500 208418
rect 350448 208354 350500 208360
rect 350446 207224 350502 207233
rect 350446 207159 350502 207168
rect 350460 207126 350488 207159
rect 350448 207120 350500 207126
rect 350448 207062 350500 207068
rect 350448 206984 350500 206990
rect 350446 206952 350448 206961
rect 350500 206952 350502 206961
rect 350446 206887 350502 206896
rect 350448 204264 350500 204270
rect 350446 204232 350448 204241
rect 350500 204232 350502 204241
rect 350446 204167 350502 204176
rect 350446 203144 350502 203153
rect 350446 203079 350502 203088
rect 350460 202910 350488 203079
rect 350448 202904 350500 202910
rect 350448 202846 350500 202852
rect 350446 201784 350502 201793
rect 350446 201719 350502 201728
rect 350460 201550 350488 201719
rect 350448 201544 350500 201550
rect 350448 201486 350500 201492
rect 350356 195356 350408 195362
rect 350356 195298 350408 195304
rect 350448 165028 350500 165034
rect 350448 164970 350500 164976
rect 349988 155644 350040 155650
rect 349988 155586 350040 155592
rect 348700 153196 348752 153202
rect 348700 153138 348752 153144
rect 347872 152312 347924 152318
rect 347872 152254 347924 152260
rect 347884 149940 347912 152254
rect 350460 149940 350488 164970
rect 350552 155174 350580 244423
rect 350644 166802 350672 284271
rect 350632 166796 350684 166802
rect 350632 166738 350684 166744
rect 350540 155168 350592 155174
rect 350540 155110 350592 155116
rect 350736 152250 350764 304982
rect 350816 270428 350868 270434
rect 350816 270370 350868 270376
rect 350828 236026 350856 270370
rect 350816 236020 350868 236026
rect 350816 235962 350868 235968
rect 351012 191214 351040 363287
rect 351000 191208 351052 191214
rect 351000 191150 351052 191156
rect 351104 184686 351132 379743
rect 351196 304366 351224 384950
rect 351184 304360 351236 304366
rect 351184 304302 351236 304308
rect 351184 288516 351236 288522
rect 351184 288458 351236 288464
rect 351196 193730 351224 288458
rect 351276 262268 351328 262274
rect 351276 262210 351328 262216
rect 351288 196790 351316 262210
rect 351276 196784 351328 196790
rect 351276 196726 351328 196732
rect 351184 193724 351236 193730
rect 351184 193666 351236 193672
rect 351092 184680 351144 184686
rect 351092 184622 351144 184628
rect 351380 182782 351408 531286
rect 352024 456142 352052 587182
rect 353300 570716 353352 570722
rect 353300 570658 353352 570664
rect 352380 569424 352432 569430
rect 352380 569366 352432 569372
rect 352196 567928 352248 567934
rect 352196 567870 352248 567876
rect 352104 558952 352156 558958
rect 352104 558894 352156 558900
rect 352116 521218 352144 558894
rect 352104 521212 352156 521218
rect 352104 521154 352156 521160
rect 352104 506592 352156 506598
rect 352104 506534 352156 506540
rect 352012 456136 352064 456142
rect 352012 456078 352064 456084
rect 352012 394800 352064 394806
rect 352012 394742 352064 394748
rect 351460 394732 351512 394738
rect 351460 394674 351512 394680
rect 351472 186046 351500 394674
rect 351920 222148 351972 222154
rect 351920 222090 351972 222096
rect 351932 204474 351960 222090
rect 351920 204468 351972 204474
rect 351920 204410 351972 204416
rect 351460 186040 351512 186046
rect 351460 185982 351512 185988
rect 351368 182776 351420 182782
rect 351368 182718 351420 182724
rect 351092 162376 351144 162382
rect 351092 162318 351144 162324
rect 350724 152244 350776 152250
rect 350724 152186 350776 152192
rect 351104 149940 351132 162318
rect 352024 149954 352052 394742
rect 352116 175098 352144 506534
rect 352208 247110 352236 567870
rect 352288 560992 352340 560998
rect 352288 560934 352340 560940
rect 352300 491298 352328 560934
rect 352288 491292 352340 491298
rect 352288 491234 352340 491240
rect 352288 484424 352340 484430
rect 352288 484366 352340 484372
rect 352196 247104 352248 247110
rect 352196 247046 352248 247052
rect 352196 244656 352248 244662
rect 352196 244598 352248 244604
rect 352208 193798 352236 244598
rect 352196 193792 352248 193798
rect 352196 193734 352248 193740
rect 352300 184142 352328 484366
rect 352392 351966 352420 569366
rect 352472 569288 352524 569294
rect 352472 569230 352524 569236
rect 352484 358562 352512 569230
rect 352840 563984 352892 563990
rect 352840 563926 352892 563932
rect 352564 561128 352616 561134
rect 352564 561070 352616 561076
rect 352472 358556 352524 358562
rect 352472 358498 352524 358504
rect 352472 356108 352524 356114
rect 352472 356050 352524 356056
rect 352380 351960 352432 351966
rect 352380 351902 352432 351908
rect 352380 350668 352432 350674
rect 352380 350610 352432 350616
rect 352392 184754 352420 350610
rect 352380 184748 352432 184754
rect 352380 184690 352432 184696
rect 352288 184136 352340 184142
rect 352288 184078 352340 184084
rect 352104 175092 352156 175098
rect 352104 175034 352156 175040
rect 352484 173398 352512 356050
rect 352576 275330 352604 561070
rect 352656 560652 352708 560658
rect 352656 560594 352708 560600
rect 352668 305017 352696 560594
rect 352748 390584 352800 390590
rect 352748 390526 352800 390532
rect 352654 305008 352710 305017
rect 352654 304943 352710 304952
rect 352656 304360 352708 304366
rect 352656 304302 352708 304308
rect 352564 275324 352616 275330
rect 352564 275266 352616 275272
rect 352564 247104 352616 247110
rect 352564 247046 352616 247052
rect 352576 233782 352604 247046
rect 352564 233776 352616 233782
rect 352564 233718 352616 233724
rect 352668 222630 352696 304302
rect 352656 222624 352708 222630
rect 352656 222566 352708 222572
rect 352564 206168 352616 206174
rect 352564 206110 352616 206116
rect 352576 196858 352604 206110
rect 352564 196852 352616 196858
rect 352564 196794 352616 196800
rect 352760 188426 352788 390526
rect 352748 188420 352800 188426
rect 352748 188362 352800 188368
rect 352852 184822 352880 563926
rect 353312 511970 353340 570658
rect 353852 570648 353904 570654
rect 353852 570590 353904 570596
rect 353760 569492 353812 569498
rect 353760 569434 353812 569440
rect 353392 569220 353444 569226
rect 353392 569162 353444 569168
rect 353300 511964 353352 511970
rect 353300 511906 353352 511912
rect 353404 247110 353432 569162
rect 353576 565548 353628 565554
rect 353576 565490 353628 565496
rect 353484 491428 353536 491434
rect 353484 491370 353536 491376
rect 353392 247104 353444 247110
rect 353392 247046 353444 247052
rect 353392 231872 353444 231878
rect 353392 231814 353444 231820
rect 353300 215348 353352 215354
rect 353300 215290 353352 215296
rect 353312 201113 353340 215290
rect 353298 201104 353354 201113
rect 353298 201039 353354 201048
rect 352840 184816 352892 184822
rect 352840 184758 352892 184764
rect 353404 183394 353432 231814
rect 353496 191418 353524 491370
rect 353588 273358 353616 565490
rect 353668 563712 353720 563718
rect 353668 563654 353720 563660
rect 353680 300830 353708 563654
rect 353772 451178 353800 569434
rect 353760 451172 353812 451178
rect 353760 451114 353812 451120
rect 353760 421048 353812 421054
rect 353760 420990 353812 420996
rect 353668 300824 353720 300830
rect 353668 300766 353720 300772
rect 353576 273352 353628 273358
rect 353576 273294 353628 273300
rect 353576 271924 353628 271930
rect 353576 271866 353628 271872
rect 353484 191412 353536 191418
rect 353484 191354 353536 191360
rect 353392 183388 353444 183394
rect 353392 183330 353444 183336
rect 352472 173392 352524 173398
rect 352472 173334 352524 173340
rect 353588 172174 353616 271866
rect 353772 186930 353800 420990
rect 353864 365702 353892 570590
rect 353944 567384 353996 567390
rect 353944 567326 353996 567332
rect 353956 542366 353984 567326
rect 354680 565208 354732 565214
rect 354680 565150 354732 565156
rect 353944 542360 353996 542366
rect 353944 542302 353996 542308
rect 354128 513460 354180 513466
rect 354128 513402 354180 513408
rect 353852 365696 353904 365702
rect 353852 365638 353904 365644
rect 353852 345500 353904 345506
rect 353852 345442 353904 345448
rect 353760 186924 353812 186930
rect 353760 186866 353812 186872
rect 353864 176186 353892 345442
rect 353944 307828 353996 307834
rect 353944 307770 353996 307776
rect 353852 176180 353904 176186
rect 353852 176122 353904 176128
rect 353576 172168 353628 172174
rect 353576 172110 353628 172116
rect 353956 155650 353984 307770
rect 354036 298172 354088 298178
rect 354036 298114 354088 298120
rect 354048 220114 354076 298114
rect 354036 220108 354088 220114
rect 354036 220050 354088 220056
rect 354140 186114 354168 513402
rect 354220 302320 354272 302326
rect 354220 302262 354272 302268
rect 354232 187406 354260 302262
rect 354588 219496 354640 219502
rect 354588 219438 354640 219444
rect 354600 215286 354628 219438
rect 354588 215280 354640 215286
rect 354588 215222 354640 215228
rect 354220 187400 354272 187406
rect 354220 187342 354272 187348
rect 354128 186108 354180 186114
rect 354128 186050 354180 186056
rect 354312 175024 354364 175030
rect 354312 174966 354364 174972
rect 353944 155644 353996 155650
rect 353944 155586 353996 155592
rect 352024 149926 352406 149954
rect 354324 149940 354352 174966
rect 354692 153066 354720 565150
rect 354784 196586 354812 587250
rect 356520 587036 356572 587042
rect 356520 586978 356572 586984
rect 356428 585880 356480 585886
rect 356428 585822 356480 585828
rect 355140 580304 355192 580310
rect 355140 580246 355192 580252
rect 355048 577652 355100 577658
rect 355048 577594 355100 577600
rect 354956 572076 355008 572082
rect 354956 572018 355008 572024
rect 354864 569356 354916 569362
rect 354864 569298 354916 569304
rect 354876 199442 354904 569298
rect 354968 218006 354996 572018
rect 355060 248402 355088 577594
rect 355152 269006 355180 580246
rect 356152 570852 356204 570858
rect 356152 570794 356204 570800
rect 355324 563780 355376 563786
rect 355324 563722 355376 563728
rect 355232 498228 355284 498234
rect 355232 498170 355284 498176
rect 355140 269000 355192 269006
rect 355140 268942 355192 268948
rect 355140 253972 355192 253978
rect 355140 253914 355192 253920
rect 355048 248396 355100 248402
rect 355048 248338 355100 248344
rect 354956 218000 355008 218006
rect 354956 217942 355008 217948
rect 355048 217252 355100 217258
rect 355048 217194 355100 217200
rect 354864 199436 354916 199442
rect 354864 199378 354916 199384
rect 354772 196580 354824 196586
rect 354772 196522 354824 196528
rect 355060 184550 355088 217194
rect 355152 192642 355180 253914
rect 355244 195158 355272 498170
rect 355336 238134 355364 563722
rect 355416 494556 355468 494562
rect 355416 494498 355468 494504
rect 355428 456793 355456 494498
rect 355414 456784 355470 456793
rect 355414 456719 355470 456728
rect 355416 358012 355468 358018
rect 355416 357954 355468 357960
rect 355324 238128 355376 238134
rect 355324 238070 355376 238076
rect 355324 226364 355376 226370
rect 355324 226306 355376 226312
rect 355232 195152 355284 195158
rect 355232 195094 355284 195100
rect 355140 192636 355192 192642
rect 355140 192578 355192 192584
rect 355048 184544 355100 184550
rect 355048 184486 355100 184492
rect 355336 155786 355364 226306
rect 355428 169522 355456 357954
rect 355506 285832 355562 285841
rect 355506 285767 355508 285776
rect 355560 285767 355562 285776
rect 355508 285738 355560 285744
rect 355508 273420 355560 273426
rect 355508 273362 355560 273368
rect 355520 234734 355548 273362
rect 355876 245676 355928 245682
rect 355876 245618 355928 245624
rect 355508 234728 355560 234734
rect 355508 234670 355560 234676
rect 355600 233980 355652 233986
rect 355600 233922 355652 233928
rect 355508 218068 355560 218074
rect 355508 218010 355560 218016
rect 355520 171902 355548 218010
rect 355508 171896 355560 171902
rect 355508 171838 355560 171844
rect 355416 169516 355468 169522
rect 355416 169458 355468 169464
rect 355324 155780 355376 155786
rect 355324 155722 355376 155728
rect 354680 153060 354732 153066
rect 354680 153002 354732 153008
rect 354772 153060 354824 153066
rect 354772 153002 354824 153008
rect 354784 152794 354812 153002
rect 354772 152788 354824 152794
rect 354772 152730 354824 152736
rect 354864 152788 354916 152794
rect 354864 152730 354916 152736
rect 354876 152658 354904 152730
rect 354864 152652 354916 152658
rect 354864 152594 354916 152600
rect 354956 152652 355008 152658
rect 354956 152594 355008 152600
rect 354968 149940 354996 152594
rect 355612 149940 355640 233922
rect 355888 233238 355916 245618
rect 356164 238754 356192 570794
rect 356244 473408 356296 473414
rect 356244 473350 356296 473356
rect 356072 238726 356192 238754
rect 356072 236042 356100 238726
rect 355980 236014 356100 236042
rect 355876 233232 355928 233238
rect 355876 233174 355928 233180
rect 355980 220794 356008 236014
rect 356152 234932 356204 234938
rect 356152 234874 356204 234880
rect 356060 233232 356112 233238
rect 356060 233174 356112 233180
rect 355968 220788 356020 220794
rect 355968 220730 356020 220736
rect 356072 219502 356100 233174
rect 356060 219496 356112 219502
rect 356060 219438 356112 219444
rect 356164 192574 356192 234874
rect 356152 192568 356204 192574
rect 356152 192510 356204 192516
rect 356060 162308 356112 162314
rect 356060 162250 356112 162256
rect 356072 149954 356100 162250
rect 356256 161158 356284 473350
rect 356336 457292 356388 457298
rect 356336 457234 356388 457240
rect 356244 161152 356296 161158
rect 356244 161094 356296 161100
rect 356348 151502 356376 457234
rect 356440 287026 356468 585822
rect 356532 288522 356560 586978
rect 357716 586764 357768 586770
rect 357716 586706 357768 586712
rect 357624 568880 357676 568886
rect 357624 568822 357676 568828
rect 357440 568676 357492 568682
rect 357440 568618 357492 568624
rect 357164 566160 357216 566166
rect 357164 566102 357216 566108
rect 356704 525972 356756 525978
rect 356704 525914 356756 525920
rect 356520 288516 356572 288522
rect 356520 288458 356572 288464
rect 356428 287020 356480 287026
rect 356428 286962 356480 286968
rect 356428 221196 356480 221202
rect 356428 221138 356480 221144
rect 356440 185910 356468 221138
rect 356612 220788 356664 220794
rect 356612 220730 356664 220736
rect 356520 215280 356572 215286
rect 356520 215222 356572 215228
rect 356532 188902 356560 215222
rect 356624 195430 356652 220730
rect 356716 217326 356744 525914
rect 356796 414452 356848 414458
rect 356796 414394 356848 414400
rect 356808 228954 356836 414394
rect 356888 392012 356940 392018
rect 356888 391954 356940 391960
rect 356796 228948 356848 228954
rect 356796 228890 356848 228896
rect 356704 217320 356756 217326
rect 356704 217262 356756 217268
rect 356900 213246 356928 391954
rect 357072 287156 357124 287162
rect 357072 287098 357124 287104
rect 356980 256760 357032 256766
rect 356980 256702 357032 256708
rect 356888 213240 356940 213246
rect 356888 213182 356940 213188
rect 356612 195424 356664 195430
rect 356612 195366 356664 195372
rect 356520 188896 356572 188902
rect 356520 188838 356572 188844
rect 356428 185904 356480 185910
rect 356428 185846 356480 185852
rect 356992 166870 357020 256702
rect 357084 227254 357112 287098
rect 357072 227248 357124 227254
rect 357072 227190 357124 227196
rect 356980 166864 357032 166870
rect 356980 166806 357032 166812
rect 357176 155038 357204 566102
rect 357452 184482 357480 568618
rect 357532 560312 357584 560318
rect 357532 560254 357584 560260
rect 357440 184476 357492 184482
rect 357440 184418 357492 184424
rect 357544 180470 357572 560254
rect 357636 309806 357664 568822
rect 357728 388482 357756 586706
rect 357716 388476 357768 388482
rect 357716 388418 357768 388424
rect 357624 309800 357676 309806
rect 357624 309742 357676 309748
rect 357624 275324 357676 275330
rect 357624 275266 357676 275272
rect 357532 180464 357584 180470
rect 357532 180406 357584 180412
rect 357164 155032 357216 155038
rect 357164 154974 357216 154980
rect 357636 152590 357664 275266
rect 357716 245812 357768 245818
rect 357716 245754 357768 245760
rect 357728 187474 357756 245754
rect 357716 187468 357768 187474
rect 357716 187410 357768 187416
rect 358096 180402 358124 640290
rect 359280 586900 359332 586906
rect 359280 586842 359332 586848
rect 359188 566568 359240 566574
rect 359188 566510 359240 566516
rect 358820 566228 358872 566234
rect 358820 566170 358872 566176
rect 358268 549296 358320 549302
rect 358268 549238 358320 549244
rect 358176 516180 358228 516186
rect 358176 516122 358228 516128
rect 358084 180396 358136 180402
rect 358084 180338 358136 180344
rect 358188 152726 358216 516122
rect 358280 199306 358308 549238
rect 358452 404456 358504 404462
rect 358452 404398 358504 404404
rect 358360 390584 358412 390590
rect 358360 390526 358412 390532
rect 358268 199300 358320 199306
rect 358268 199242 358320 199248
rect 358372 193662 358400 390526
rect 358464 232558 358492 404398
rect 358544 307828 358596 307834
rect 358544 307770 358596 307776
rect 358452 232552 358504 232558
rect 358452 232494 358504 232500
rect 358360 193656 358412 193662
rect 358360 193598 358412 193604
rect 358556 160954 358584 307770
rect 358544 160948 358596 160954
rect 358544 160890 358596 160896
rect 358176 152720 358228 152726
rect 358176 152662 358228 152668
rect 357624 152584 357676 152590
rect 357624 152526 357676 152532
rect 358832 152318 358860 566170
rect 358912 565072 358964 565078
rect 358912 565014 358964 565020
rect 358924 152794 358952 565014
rect 359004 560856 359056 560862
rect 359004 560798 359056 560804
rect 359016 183462 359044 560798
rect 359096 532840 359148 532846
rect 359096 532782 359148 532788
rect 359004 183456 359056 183462
rect 359004 183398 359056 183404
rect 359108 158574 359136 532782
rect 359200 200802 359228 566510
rect 359292 245682 359320 586842
rect 359372 398880 359424 398886
rect 359372 398822 359424 398828
rect 359280 245676 359332 245682
rect 359280 245618 359332 245624
rect 359280 244928 359332 244934
rect 359280 244870 359332 244876
rect 359188 200796 359240 200802
rect 359188 200738 359240 200744
rect 359292 191690 359320 244870
rect 359280 191684 359332 191690
rect 359280 191626 359332 191632
rect 359384 185842 359412 398822
rect 359372 185836 359424 185842
rect 359372 185778 359424 185784
rect 359096 158568 359148 158574
rect 359096 158510 359148 158516
rect 358912 152788 358964 152794
rect 358912 152730 358964 152736
rect 359476 152454 359504 684898
rect 361580 674892 361632 674898
rect 361580 674834 361632 674840
rect 360844 632120 360896 632126
rect 360844 632062 360896 632068
rect 360384 567860 360436 567866
rect 360384 567802 360436 567808
rect 359556 567452 359608 567458
rect 359556 567394 359608 567400
rect 359568 509182 359596 567394
rect 360200 565004 360252 565010
rect 360200 564946 360252 564952
rect 359556 509176 359608 509182
rect 359556 509118 359608 509124
rect 359556 506524 359608 506530
rect 359556 506466 359608 506472
rect 359568 159497 359596 506466
rect 359648 303680 359700 303686
rect 359648 303622 359700 303628
rect 359554 159488 359610 159497
rect 359554 159423 359610 159432
rect 359660 159390 359688 303622
rect 360108 176112 360160 176118
rect 360108 176054 360160 176060
rect 359648 159384 359700 159390
rect 359648 159326 359700 159332
rect 359464 152448 359516 152454
rect 359464 152390 359516 152396
rect 358820 152312 358872 152318
rect 358820 152254 358872 152260
rect 356336 151496 356388 151502
rect 356336 151438 356388 151444
rect 356072 149926 356270 149954
rect 360120 149940 360148 176054
rect 360212 152386 360240 564946
rect 360292 564936 360344 564942
rect 360292 564878 360344 564884
rect 360304 152930 360332 564878
rect 360396 198694 360424 567802
rect 360568 559700 360620 559706
rect 360568 559642 360620 559648
rect 360476 503736 360528 503742
rect 360476 503678 360528 503684
rect 360384 198688 360436 198694
rect 360384 198630 360436 198636
rect 360488 163946 360516 503678
rect 360580 226370 360608 559642
rect 360660 425128 360712 425134
rect 360660 425070 360712 425076
rect 360568 226364 360620 226370
rect 360568 226306 360620 226312
rect 360568 225004 360620 225010
rect 360568 224946 360620 224952
rect 360580 183326 360608 224946
rect 360672 187678 360700 425070
rect 360856 199374 360884 632062
rect 360936 492720 360988 492726
rect 360936 492662 360988 492668
rect 360844 199368 360896 199374
rect 360844 199310 360896 199316
rect 360660 187672 360712 187678
rect 360660 187614 360712 187620
rect 360568 183320 360620 183326
rect 360568 183262 360620 183268
rect 360476 163940 360528 163946
rect 360476 163882 360528 163888
rect 360948 155718 360976 492662
rect 361028 430704 361080 430710
rect 361028 430646 361080 430652
rect 361040 224330 361068 430646
rect 361120 249892 361172 249898
rect 361120 249834 361172 249840
rect 361028 224324 361080 224330
rect 361028 224266 361080 224272
rect 361132 161090 361160 249834
rect 361592 196722 361620 674834
rect 361856 586696 361908 586702
rect 361856 586638 361908 586644
rect 361764 586628 361816 586634
rect 361764 586570 361816 586576
rect 361672 568744 361724 568750
rect 361672 568686 361724 568692
rect 361580 196716 361632 196722
rect 361580 196658 361632 196664
rect 361120 161084 361172 161090
rect 361120 161026 361172 161032
rect 360936 155712 360988 155718
rect 360936 155654 360988 155660
rect 361684 155582 361712 568686
rect 361776 192914 361804 586570
rect 361868 195226 361896 586638
rect 361948 419552 362000 419558
rect 361948 419494 362000 419500
rect 361856 195220 361908 195226
rect 361856 195162 361908 195168
rect 361764 192908 361816 192914
rect 361764 192850 361816 192856
rect 361960 156874 361988 419494
rect 361948 156868 362000 156874
rect 361948 156810 362000 156816
rect 361672 155576 361724 155582
rect 361672 155518 361724 155524
rect 360292 152924 360344 152930
rect 360292 152866 360344 152872
rect 362236 152658 362264 684966
rect 363144 570784 363196 570790
rect 363144 570726 363196 570732
rect 362316 489932 362368 489938
rect 362316 489874 362368 489880
rect 362328 176322 362356 489874
rect 362960 480344 363012 480350
rect 362960 480286 363012 480292
rect 362408 419552 362460 419558
rect 362408 419494 362460 419500
rect 362420 199753 362448 419494
rect 362500 350600 362552 350606
rect 362500 350542 362552 350548
rect 362512 232694 362540 350542
rect 362500 232688 362552 232694
rect 362500 232630 362552 232636
rect 362406 199744 362462 199753
rect 362406 199679 362462 199688
rect 362972 177857 363000 480286
rect 363052 461032 363104 461038
rect 363052 460974 363104 460980
rect 363064 187338 363092 460974
rect 363156 343602 363184 570726
rect 363144 343596 363196 343602
rect 363144 343538 363196 343544
rect 363144 329860 363196 329866
rect 363144 329802 363196 329808
rect 363052 187332 363104 187338
rect 363052 187274 363104 187280
rect 362958 177848 363014 177857
rect 362958 177783 363014 177792
rect 362316 176316 362368 176322
rect 362316 176258 362368 176264
rect 363156 169454 363184 329802
rect 363236 325712 363288 325718
rect 363236 325654 363288 325660
rect 363248 322930 363276 325654
rect 363236 322924 363288 322930
rect 363236 322866 363288 322872
rect 363236 245744 363288 245750
rect 363236 245686 363288 245692
rect 363248 187649 363276 245686
rect 363420 234728 363472 234734
rect 363420 234670 363472 234676
rect 363328 200796 363380 200802
rect 363328 200738 363380 200744
rect 363234 187640 363290 187649
rect 363234 187575 363290 187584
rect 363144 169448 363196 169454
rect 363144 169390 363196 169396
rect 362224 152652 362276 152658
rect 362224 152594 362276 152600
rect 360200 152380 360252 152386
rect 360200 152322 360252 152328
rect 363340 149940 363368 200738
rect 363432 184414 363460 234670
rect 363420 184408 363472 184414
rect 363420 184350 363472 184356
rect 363616 153066 363644 685918
rect 373908 682168 373960 682174
rect 373908 682110 373960 682116
rect 363694 680912 363750 680921
rect 363694 680847 363750 680856
rect 363708 199073 363736 680847
rect 369858 680504 369914 680513
rect 369858 680439 369914 680448
rect 367836 648644 367888 648650
rect 367836 648586 367888 648592
rect 367744 633480 367796 633486
rect 367744 633422 367796 633428
rect 364340 604512 364392 604518
rect 364340 604454 364392 604460
rect 363788 542428 363840 542434
rect 363788 542370 363840 542376
rect 363800 237386 363828 542370
rect 363880 474836 363932 474842
rect 363880 474778 363932 474784
rect 363788 237380 363840 237386
rect 363788 237322 363840 237328
rect 363694 199064 363750 199073
rect 363694 198999 363750 199008
rect 363892 195566 363920 474778
rect 363972 430636 364024 430642
rect 363972 430578 364024 430584
rect 363984 234122 364012 430578
rect 364064 360256 364116 360262
rect 364064 360198 364116 360204
rect 363972 234116 364024 234122
rect 363972 234058 364024 234064
rect 363880 195560 363932 195566
rect 363880 195502 363932 195508
rect 364076 194138 364104 360198
rect 364352 198150 364380 604454
rect 366364 601724 366416 601730
rect 366364 601666 366416 601672
rect 365076 574796 365128 574802
rect 365076 574738 365128 574744
rect 364432 563236 364484 563242
rect 364432 563178 364484 563184
rect 364340 198144 364392 198150
rect 364340 198086 364392 198092
rect 364444 194206 364472 563178
rect 364984 561060 365036 561066
rect 364984 561002 365036 561008
rect 364524 476196 364576 476202
rect 364524 476138 364576 476144
rect 364432 194200 364484 194206
rect 364432 194142 364484 194148
rect 364064 194132 364116 194138
rect 364064 194074 364116 194080
rect 364536 182102 364564 476138
rect 364524 182096 364576 182102
rect 364524 182038 364576 182044
rect 363604 153060 363656 153066
rect 363604 153002 363656 153008
rect 364996 152930 365024 561002
rect 365088 276010 365116 574738
rect 365168 567588 365220 567594
rect 365168 567530 365220 567536
rect 365180 294642 365208 567530
rect 365720 563304 365772 563310
rect 365720 563246 365772 563252
rect 365260 469260 365312 469266
rect 365260 469202 365312 469208
rect 365168 294636 365220 294642
rect 365168 294578 365220 294584
rect 365168 292596 365220 292602
rect 365168 292538 365220 292544
rect 365076 276004 365128 276010
rect 365076 275946 365128 275952
rect 365180 169658 365208 292538
rect 365272 198286 365300 469202
rect 365444 422340 365496 422346
rect 365444 422282 365496 422288
rect 365352 400240 365404 400246
rect 365352 400182 365404 400188
rect 365260 198280 365312 198286
rect 365260 198222 365312 198228
rect 365168 169652 365220 169658
rect 365168 169594 365220 169600
rect 365364 161090 365392 400182
rect 365456 345030 365484 422282
rect 365444 345024 365496 345030
rect 365444 344966 365496 344972
rect 365536 329860 365588 329866
rect 365536 329802 365588 329808
rect 365444 300892 365496 300898
rect 365444 300834 365496 300840
rect 365456 232626 365484 300834
rect 365548 285666 365576 329802
rect 365536 285660 365588 285666
rect 365536 285602 365588 285608
rect 365628 263628 365680 263634
rect 365628 263570 365680 263576
rect 365536 262948 365588 262954
rect 365536 262890 365588 262896
rect 365548 258074 365576 262890
rect 365640 262206 365668 263570
rect 365628 262200 365680 262206
rect 365628 262142 365680 262148
rect 365548 258046 365668 258074
rect 365640 240106 365668 258046
rect 365628 240100 365680 240106
rect 365628 240042 365680 240048
rect 365444 232620 365496 232626
rect 365444 232562 365496 232568
rect 365352 161084 365404 161090
rect 365352 161026 365404 161032
rect 365732 155689 365760 563246
rect 365812 559088 365864 559094
rect 365812 559030 365864 559036
rect 365824 193934 365852 559030
rect 365904 447160 365956 447166
rect 365904 447102 365956 447108
rect 365812 193928 365864 193934
rect 365812 193870 365864 193876
rect 365916 190233 365944 447102
rect 366088 338156 366140 338162
rect 366088 338098 366140 338104
rect 366100 191282 366128 338098
rect 366180 229152 366232 229158
rect 366180 229094 366232 229100
rect 366088 191276 366140 191282
rect 366088 191218 366140 191224
rect 365902 190224 365958 190233
rect 365902 190159 365958 190168
rect 365718 155680 365774 155689
rect 365718 155615 365774 155624
rect 364984 152924 365036 152930
rect 364984 152866 365036 152872
rect 366192 151570 366220 229094
rect 366376 159730 366404 601666
rect 366456 571396 366508 571402
rect 366456 571338 366508 571344
rect 366468 199238 366496 571338
rect 367192 566432 367244 566438
rect 367192 566374 367244 566380
rect 366548 561944 366600 561950
rect 366548 561886 366600 561892
rect 366560 240145 366588 561886
rect 366640 546576 366692 546582
rect 366640 546518 366692 546524
rect 366546 240136 366602 240145
rect 366546 240071 366602 240080
rect 366652 232529 366680 546518
rect 367100 516316 367152 516322
rect 367100 516258 367152 516264
rect 366732 445868 366784 445874
rect 366732 445810 366784 445816
rect 366744 361554 366772 445810
rect 366732 361548 366784 361554
rect 366732 361490 366784 361496
rect 366824 332648 366876 332654
rect 366824 332590 366876 332596
rect 366732 300892 366784 300898
rect 366732 300834 366784 300840
rect 366638 232520 366694 232529
rect 366638 232455 366694 232464
rect 366456 199232 366508 199238
rect 366456 199174 366508 199180
rect 366744 186182 366772 300834
rect 366732 186176 366784 186182
rect 366732 186118 366784 186124
rect 366364 159724 366416 159730
rect 366364 159666 366416 159672
rect 366180 151564 366232 151570
rect 366180 151506 366232 151512
rect 366836 149938 366864 332590
rect 367112 187513 367140 516258
rect 367204 262954 367232 566374
rect 367284 481704 367336 481710
rect 367284 481646 367336 481652
rect 367192 262948 367244 262954
rect 367192 262890 367244 262896
rect 367098 187504 367154 187513
rect 367098 187439 367154 187448
rect 367296 184278 367324 481646
rect 367376 404388 367428 404394
rect 367376 404330 367428 404336
rect 367284 184272 367336 184278
rect 367284 184214 367336 184220
rect 367388 178974 367416 404330
rect 367468 263696 367520 263702
rect 367468 263638 367520 263644
rect 367376 178968 367428 178974
rect 367376 178910 367428 178916
rect 367480 166598 367508 263638
rect 367756 169726 367784 633422
rect 367848 580446 367876 648586
rect 368480 608660 368532 608666
rect 368480 608602 368532 608608
rect 367836 580440 367888 580446
rect 367836 580382 367888 580388
rect 367928 562148 367980 562154
rect 367928 562090 367980 562096
rect 367836 538280 367888 538286
rect 367836 538222 367888 538228
rect 367848 225622 367876 538222
rect 367940 265674 367968 562090
rect 368020 513392 368072 513398
rect 368020 513334 368072 513340
rect 368032 310486 368060 513334
rect 368296 349240 368348 349246
rect 368296 349182 368348 349188
rect 368112 310548 368164 310554
rect 368112 310490 368164 310496
rect 368020 310480 368072 310486
rect 368020 310422 368072 310428
rect 368020 299532 368072 299538
rect 368020 299474 368072 299480
rect 367928 265668 367980 265674
rect 367928 265610 367980 265616
rect 367836 225616 367888 225622
rect 367836 225558 367888 225564
rect 368032 173262 368060 299474
rect 368020 173256 368072 173262
rect 368020 173198 368072 173204
rect 367744 169720 367796 169726
rect 367744 169662 367796 169668
rect 367468 166592 367520 166598
rect 367468 166534 367520 166540
rect 368124 158574 368152 310490
rect 368308 284306 368336 349182
rect 368296 284300 368348 284306
rect 368296 284242 368348 284248
rect 368204 282940 368256 282946
rect 368204 282882 368256 282888
rect 368112 158568 368164 158574
rect 368112 158510 368164 158516
rect 368216 156942 368244 282882
rect 368492 194177 368520 608602
rect 368664 564732 368716 564738
rect 368664 564674 368716 564680
rect 368572 561876 368624 561882
rect 368572 561818 368624 561824
rect 368478 194168 368534 194177
rect 368478 194103 368534 194112
rect 368204 156936 368256 156942
rect 368204 156878 368256 156884
rect 368584 155378 368612 561818
rect 368676 187377 368704 564674
rect 368938 563680 368994 563689
rect 368938 563615 368994 563624
rect 368756 480276 368808 480282
rect 368756 480218 368808 480224
rect 368662 187368 368718 187377
rect 368662 187303 368718 187312
rect 368572 155372 368624 155378
rect 368572 155314 368624 155320
rect 368768 151434 368796 480218
rect 368848 441652 368900 441658
rect 368848 441594 368900 441600
rect 368860 177614 368888 441594
rect 368952 341465 368980 563615
rect 369124 562556 369176 562562
rect 369124 562498 369176 562504
rect 368938 341456 368994 341465
rect 368938 341391 368994 341400
rect 368940 294024 368992 294030
rect 368940 293966 368992 293972
rect 368952 181898 368980 293966
rect 369136 218754 369164 562498
rect 369216 462460 369268 462466
rect 369216 462402 369268 462408
rect 369228 232898 369256 462402
rect 369308 420980 369360 420986
rect 369308 420922 369360 420928
rect 369216 232892 369268 232898
rect 369216 232834 369268 232840
rect 369320 227050 369348 420922
rect 369400 328500 369452 328506
rect 369400 328442 369452 328448
rect 369412 228478 369440 328442
rect 369400 228472 369452 228478
rect 369400 228414 369452 228420
rect 369308 227044 369360 227050
rect 369308 226986 369360 226992
rect 369124 218748 369176 218754
rect 369124 218690 369176 218696
rect 368940 181892 368992 181898
rect 368940 181834 368992 181840
rect 368848 177608 368900 177614
rect 368848 177550 368900 177556
rect 369124 155916 369176 155922
rect 369124 155858 369176 155864
rect 368756 151428 368808 151434
rect 368756 151370 368808 151376
rect 369136 149940 369164 155858
rect 369872 149954 369900 680439
rect 371884 615528 371936 615534
rect 371884 615470 371936 615476
rect 371240 605872 371292 605878
rect 371240 605814 371292 605820
rect 370504 568948 370556 568954
rect 370504 568890 370556 568896
rect 369952 567996 370004 568002
rect 369952 567938 370004 567944
rect 369964 197334 369992 567938
rect 369952 197328 370004 197334
rect 369952 197270 370004 197276
rect 370516 155378 370544 568890
rect 370596 528624 370648 528630
rect 370596 528566 370648 528572
rect 370608 187202 370636 528566
rect 370688 484424 370740 484430
rect 370688 484366 370740 484372
rect 370700 187542 370728 484366
rect 370780 441652 370832 441658
rect 370780 441594 370832 441600
rect 370792 194002 370820 441594
rect 370872 426556 370924 426562
rect 370872 426498 370924 426504
rect 370884 199102 370912 426498
rect 370964 407176 371016 407182
rect 370964 407118 371016 407124
rect 370872 199096 370924 199102
rect 370872 199038 370924 199044
rect 370780 193996 370832 194002
rect 370780 193938 370832 193944
rect 370976 191321 371004 407118
rect 371148 320204 371200 320210
rect 371148 320146 371200 320152
rect 371056 292664 371108 292670
rect 371056 292606 371108 292612
rect 370962 191312 371018 191321
rect 370962 191247 371018 191256
rect 370688 187536 370740 187542
rect 370688 187478 370740 187484
rect 370596 187196 370648 187202
rect 370596 187138 370648 187144
rect 371068 169182 371096 292606
rect 371160 233034 371188 320146
rect 371148 233028 371200 233034
rect 371148 232970 371200 232976
rect 371252 196926 371280 605814
rect 371332 465112 371384 465118
rect 371332 465054 371384 465060
rect 371240 196920 371292 196926
rect 371240 196862 371292 196868
rect 371344 187134 371372 465054
rect 371424 460964 371476 460970
rect 371424 460906 371476 460912
rect 371332 187128 371384 187134
rect 371332 187070 371384 187076
rect 371436 184210 371464 460906
rect 371896 199034 371924 615470
rect 373264 566364 373316 566370
rect 373264 566306 373316 566312
rect 371974 562456 372030 562465
rect 371974 562391 372030 562400
rect 371884 199028 371936 199034
rect 371884 198970 371936 198976
rect 371424 184204 371476 184210
rect 371424 184146 371476 184152
rect 371238 173360 371294 173369
rect 371238 173295 371294 173304
rect 371056 169176 371108 169182
rect 371056 169118 371108 169124
rect 370504 155372 370556 155378
rect 370504 155314 370556 155320
rect 371252 151814 371280 173295
rect 371988 161294 372016 562391
rect 372068 562080 372120 562086
rect 372068 562022 372120 562028
rect 372158 562048 372214 562057
rect 372080 237930 372108 562022
rect 372158 561983 372214 561992
rect 372068 237924 372120 237930
rect 372068 237866 372120 237872
rect 372172 210361 372200 561983
rect 372620 536852 372672 536858
rect 372620 536794 372672 536800
rect 372436 491360 372488 491366
rect 372436 491302 372488 491308
rect 372252 473408 372304 473414
rect 372252 473350 372304 473356
rect 372158 210352 372214 210361
rect 372158 210287 372214 210296
rect 372264 166734 372292 473350
rect 372344 456816 372396 456822
rect 372344 456758 372396 456764
rect 372252 166728 372304 166734
rect 372252 166670 372304 166676
rect 371976 161288 372028 161294
rect 371976 161230 372028 161236
rect 372356 155446 372384 456758
rect 372448 233170 372476 491302
rect 372436 233164 372488 233170
rect 372436 233106 372488 233112
rect 372632 175001 372660 536794
rect 372712 434784 372764 434790
rect 372712 434726 372764 434732
rect 372724 180198 372752 434726
rect 372804 302932 372856 302938
rect 372804 302874 372856 302880
rect 372712 180192 372764 180198
rect 372712 180134 372764 180140
rect 372618 174992 372674 175001
rect 372618 174927 372674 174936
rect 372816 171134 372844 302874
rect 372816 171106 373212 171134
rect 372344 155440 372396 155446
rect 372344 155382 372396 155388
rect 373184 151814 373212 171106
rect 373276 154290 373304 566306
rect 373354 564632 373410 564641
rect 373354 564567 373410 564576
rect 373368 158545 373396 564567
rect 373540 520328 373592 520334
rect 373540 520270 373592 520276
rect 373448 512032 373500 512038
rect 373448 511974 373500 511980
rect 373354 158536 373410 158545
rect 373354 158471 373410 158480
rect 373264 154284 373316 154290
rect 373264 154226 373316 154232
rect 373460 153134 373488 511974
rect 373552 185745 373580 520270
rect 373816 459604 373868 459610
rect 373816 459546 373868 459552
rect 373632 436144 373684 436150
rect 373632 436086 373684 436092
rect 373538 185736 373594 185745
rect 373538 185671 373594 185680
rect 373644 181830 373672 436086
rect 373724 426624 373776 426630
rect 373724 426566 373776 426572
rect 373736 190097 373764 426566
rect 373828 240038 373856 459546
rect 373920 302297 373948 682110
rect 374644 599004 374696 599010
rect 374644 598946 374696 598952
rect 374000 568812 374052 568818
rect 374000 568754 374052 568760
rect 373906 302288 373962 302297
rect 373906 302223 373962 302232
rect 373816 240032 373868 240038
rect 373816 239974 373868 239980
rect 373722 190088 373778 190097
rect 373722 190023 373778 190032
rect 373632 181824 373684 181830
rect 373632 181766 373684 181772
rect 374012 158409 374040 568754
rect 374552 449948 374604 449954
rect 374552 449890 374604 449896
rect 374564 371210 374592 449890
rect 374552 371204 374604 371210
rect 374552 371146 374604 371152
rect 374552 303748 374604 303754
rect 374552 303690 374604 303696
rect 374564 232830 374592 303690
rect 374552 232824 374604 232830
rect 374552 232766 374604 232772
rect 374656 165170 374684 598946
rect 374736 565140 374788 565146
rect 374736 565082 374788 565088
rect 374644 165164 374696 165170
rect 374644 165106 374696 165112
rect 374748 163441 374776 565082
rect 374840 513330 374868 698906
rect 380164 681964 380216 681970
rect 380164 681906 380216 681912
rect 377404 681216 377456 681222
rect 377404 681158 377456 681164
rect 376024 652792 376076 652798
rect 376024 652734 376076 652740
rect 375104 567384 375156 567390
rect 375104 567326 375156 567332
rect 374828 513324 374880 513330
rect 374828 513266 374880 513272
rect 374828 490000 374880 490006
rect 374828 489942 374880 489948
rect 374840 236570 374868 489942
rect 374920 438932 374972 438938
rect 374920 438874 374972 438880
rect 374828 236564 374880 236570
rect 374828 236506 374880 236512
rect 374932 187241 374960 438874
rect 375012 376780 375064 376786
rect 375012 376722 375064 376728
rect 374918 187232 374974 187241
rect 374918 187167 374974 187176
rect 374734 163432 374790 163441
rect 374734 163367 374790 163376
rect 373998 158400 374054 158409
rect 373998 158335 374054 158344
rect 375024 156874 375052 376722
rect 375116 375358 375144 567326
rect 375288 454096 375340 454102
rect 375288 454038 375340 454044
rect 375104 375352 375156 375358
rect 375104 375294 375156 375300
rect 375196 371272 375248 371278
rect 375196 371214 375248 371220
rect 375104 354748 375156 354754
rect 375104 354690 375156 354696
rect 375116 160954 375144 354690
rect 375208 228818 375236 371214
rect 375196 228812 375248 228818
rect 375196 228754 375248 228760
rect 375104 160948 375156 160954
rect 375104 160890 375156 160896
rect 375012 156868 375064 156874
rect 375012 156810 375064 156816
rect 375300 155417 375328 454038
rect 375380 445800 375432 445806
rect 375380 445742 375432 445748
rect 375392 177886 375420 445742
rect 375472 407244 375524 407250
rect 375472 407186 375524 407192
rect 375380 177880 375432 177886
rect 375380 177822 375432 177828
rect 375484 171834 375512 407186
rect 376036 174865 376064 652734
rect 376116 585200 376168 585206
rect 376116 585142 376168 585148
rect 376022 174856 376078 174865
rect 376022 174791 376078 174800
rect 375472 171828 375524 171834
rect 375472 171770 375524 171776
rect 375286 155408 375342 155417
rect 375286 155343 375342 155352
rect 373448 153128 373500 153134
rect 373448 153070 373500 153076
rect 376128 152425 376156 585142
rect 376484 566024 376536 566030
rect 376484 565966 376536 565972
rect 376206 561096 376262 561105
rect 376206 561031 376262 561040
rect 376220 251841 376248 561031
rect 376300 527196 376352 527202
rect 376300 527138 376352 527144
rect 376312 259418 376340 527138
rect 376392 419620 376444 419626
rect 376392 419562 376444 419568
rect 376300 259412 376352 259418
rect 376300 259354 376352 259360
rect 376300 256828 376352 256834
rect 376300 256770 376352 256776
rect 376206 251832 376262 251841
rect 376206 251767 376262 251776
rect 376312 206990 376340 256770
rect 376300 206984 376352 206990
rect 376300 206926 376352 206932
rect 376404 178673 376432 419562
rect 376496 325650 376524 565966
rect 376668 339516 376720 339522
rect 376668 339458 376720 339464
rect 376576 331288 376628 331294
rect 376576 331230 376628 331236
rect 376484 325644 376536 325650
rect 376484 325586 376536 325592
rect 376484 269136 376536 269142
rect 376484 269078 376536 269084
rect 376390 178664 376446 178673
rect 376390 178599 376446 178608
rect 376496 161226 376524 269078
rect 376588 181966 376616 331230
rect 376680 237318 376708 339458
rect 377312 322992 377364 322998
rect 377312 322934 377364 322940
rect 377220 259412 377272 259418
rect 377220 259354 377272 259360
rect 376668 237312 376720 237318
rect 376668 237254 376720 237260
rect 377232 236609 377260 259354
rect 377218 236600 377274 236609
rect 377218 236535 377274 236544
rect 376760 234048 376812 234054
rect 376760 233990 376812 233996
rect 376576 181960 376628 181966
rect 376576 181902 376628 181908
rect 376484 161220 376536 161226
rect 376484 161162 376536 161168
rect 376772 156602 376800 233990
rect 376852 164960 376904 164966
rect 376852 164902 376904 164908
rect 376760 156596 376812 156602
rect 376760 156538 376812 156544
rect 376114 152416 376170 152425
rect 376114 152351 376170 152360
rect 371252 151786 372016 151814
rect 373184 151786 373304 151814
rect 371988 149954 372016 151786
rect 373276 149954 373304 151786
rect 366824 149932 366876 149938
rect 313280 149874 313332 149880
rect 369872 149926 370438 149954
rect 371988 149926 372370 149954
rect 373276 149926 373658 149954
rect 376864 149940 376892 164902
rect 377220 156596 377272 156602
rect 377220 156538 377272 156544
rect 377232 149954 377260 156538
rect 377324 154154 377352 322934
rect 377312 154148 377364 154154
rect 377312 154090 377364 154096
rect 377416 152833 377444 681158
rect 377496 583772 377548 583778
rect 377496 583714 377548 583720
rect 377402 152824 377458 152833
rect 377402 152759 377458 152768
rect 377508 152522 377536 583714
rect 379152 564868 379204 564874
rect 379152 564810 379204 564816
rect 378784 563576 378836 563582
rect 378784 563518 378836 563524
rect 377588 546576 377640 546582
rect 377588 546518 377640 546524
rect 377600 166530 377628 546518
rect 377680 543788 377732 543794
rect 377680 543730 377732 543736
rect 377692 187066 377720 543730
rect 377772 476128 377824 476134
rect 377772 476070 377824 476076
rect 377784 229838 377812 476070
rect 377864 451376 377916 451382
rect 377864 451318 377916 451324
rect 377876 387802 377904 451318
rect 377956 416832 378008 416838
rect 377956 416774 378008 416780
rect 377864 387796 377916 387802
rect 377864 387738 377916 387744
rect 377864 378208 377916 378214
rect 377864 378150 377916 378156
rect 377772 229832 377824 229838
rect 377772 229774 377824 229780
rect 377680 187060 377732 187066
rect 377680 187002 377732 187008
rect 377588 166524 377640 166530
rect 377588 166466 377640 166472
rect 377876 162382 377904 378150
rect 377968 220182 377996 416774
rect 378048 353320 378100 353326
rect 378048 353262 378100 353268
rect 377956 220176 378008 220182
rect 377956 220118 378008 220124
rect 378060 177750 378088 353262
rect 378692 321632 378744 321638
rect 378692 321574 378744 321580
rect 378140 235340 378192 235346
rect 378140 235282 378192 235288
rect 378048 177744 378100 177750
rect 378048 177686 378100 177692
rect 377864 162376 377916 162382
rect 377864 162318 377916 162324
rect 377496 152516 377548 152522
rect 377496 152458 377548 152464
rect 378152 149954 378180 235282
rect 378704 233102 378732 321574
rect 378692 233096 378744 233102
rect 378692 233038 378744 233044
rect 378796 153134 378824 563518
rect 378876 562216 378928 562222
rect 378876 562158 378928 562164
rect 378888 161362 378916 562158
rect 378968 523048 379020 523054
rect 378968 522990 379020 522996
rect 378980 229770 379008 522990
rect 379060 483132 379112 483138
rect 379060 483074 379112 483080
rect 378968 229764 379020 229770
rect 378968 229706 379020 229712
rect 379072 196994 379100 483074
rect 379164 455394 379192 564810
rect 379152 455388 379204 455394
rect 379152 455330 379204 455336
rect 379428 447160 379480 447166
rect 379428 447102 379480 447108
rect 379152 372632 379204 372638
rect 379152 372574 379204 372580
rect 379060 196988 379112 196994
rect 379060 196930 379112 196936
rect 378876 161356 378928 161362
rect 378876 161298 378928 161304
rect 379164 159390 379192 372574
rect 379336 351960 379388 351966
rect 379336 351902 379388 351908
rect 379244 349240 379296 349246
rect 379244 349182 379296 349188
rect 379256 176254 379284 349182
rect 379348 188358 379376 351902
rect 379440 302938 379468 447102
rect 380072 381064 380124 381070
rect 380072 381006 380124 381012
rect 379428 302932 379480 302938
rect 379428 302874 379480 302880
rect 379428 299600 379480 299606
rect 379428 299542 379480 299548
rect 379440 232490 379468 299542
rect 379980 295384 380032 295390
rect 379980 295326 380032 295332
rect 379428 232484 379480 232490
rect 379428 232426 379480 232432
rect 379992 228750 380020 295326
rect 379980 228744 380032 228750
rect 379980 228686 380032 228692
rect 379336 188352 379388 188358
rect 379336 188294 379388 188300
rect 379244 176248 379296 176254
rect 379244 176190 379296 176196
rect 380084 174962 380112 381006
rect 380176 176390 380204 681906
rect 380256 534132 380308 534138
rect 380256 534074 380308 534080
rect 380268 224398 380296 534074
rect 380440 529984 380492 529990
rect 380440 529926 380492 529932
rect 380348 451308 380400 451314
rect 380348 451250 380400 451256
rect 380256 224392 380308 224398
rect 380256 224334 380308 224340
rect 380164 176384 380216 176390
rect 380164 176326 380216 176332
rect 380072 174956 380124 174962
rect 380072 174898 380124 174904
rect 379152 159384 379204 159390
rect 379152 159326 379204 159332
rect 378784 153128 378836 153134
rect 378784 153070 378836 153076
rect 380360 151298 380388 451250
rect 380452 235385 380480 529926
rect 380624 505164 380676 505170
rect 380624 505106 380676 505112
rect 380532 499588 380584 499594
rect 380532 499530 380584 499536
rect 380438 235376 380494 235385
rect 380438 235311 380494 235320
rect 380544 228886 380572 499530
rect 380636 234394 380664 505106
rect 380808 454164 380860 454170
rect 380808 454106 380860 454112
rect 380716 423700 380768 423706
rect 380716 423642 380768 423648
rect 380624 234388 380676 234394
rect 380624 234330 380676 234336
rect 380532 228880 380584 228886
rect 380532 228822 380584 228828
rect 380728 190194 380756 423642
rect 380820 227186 380848 454106
rect 381452 343732 381504 343738
rect 381452 343674 381504 343680
rect 381360 328500 381412 328506
rect 381360 328442 381412 328448
rect 380808 227180 380860 227186
rect 380808 227122 380860 227128
rect 380716 190188 380768 190194
rect 380716 190130 380768 190136
rect 381372 181762 381400 328442
rect 381360 181756 381412 181762
rect 381360 181698 381412 181704
rect 381464 156942 381492 343674
rect 381556 238814 381584 700606
rect 396908 687404 396960 687410
rect 396908 687346 396960 687352
rect 384948 686180 385000 686186
rect 384948 686122 385000 686128
rect 384302 684856 384358 684865
rect 384302 684791 384358 684800
rect 382924 682372 382976 682378
rect 382924 682314 382976 682320
rect 381636 608660 381688 608666
rect 381636 608602 381688 608608
rect 381544 238808 381596 238814
rect 381544 238750 381596 238756
rect 381648 185774 381676 608602
rect 381728 566092 381780 566098
rect 381728 566034 381780 566040
rect 381636 185768 381688 185774
rect 381636 185710 381688 185716
rect 381452 156936 381504 156942
rect 381452 156878 381504 156884
rect 381740 154193 381768 566034
rect 382188 564460 382240 564466
rect 382188 564402 382240 564408
rect 382004 562420 382056 562426
rect 382004 562362 382056 562368
rect 381820 562012 381872 562018
rect 381820 561954 381872 561960
rect 381726 154184 381782 154193
rect 381726 154119 381782 154128
rect 381832 151502 381860 561954
rect 381912 532772 381964 532778
rect 381912 532714 381964 532720
rect 381924 151706 381952 532714
rect 382016 236910 382044 562362
rect 382096 440292 382148 440298
rect 382096 440234 382148 440240
rect 382004 236904 382056 236910
rect 382004 236846 382056 236852
rect 382108 154426 382136 440234
rect 382200 336734 382228 564402
rect 382280 560924 382332 560930
rect 382280 560866 382332 560872
rect 382188 336728 382240 336734
rect 382188 336670 382240 336676
rect 382188 334008 382240 334014
rect 382188 333950 382240 333956
rect 382200 162314 382228 333950
rect 382188 162308 382240 162314
rect 382188 162250 382240 162256
rect 382096 154420 382148 154426
rect 382096 154362 382148 154368
rect 381912 151700 381964 151706
rect 381912 151642 381964 151648
rect 381820 151496 381872 151502
rect 381820 151438 381872 151444
rect 380348 151292 380400 151298
rect 380348 151234 380400 151240
rect 380716 150816 380768 150822
rect 380716 150758 380768 150764
rect 377232 149926 377522 149954
rect 378152 149926 378810 149954
rect 380728 149940 380756 150758
rect 382292 149954 382320 560866
rect 382832 396092 382884 396098
rect 382832 396034 382884 396040
rect 382740 318844 382792 318850
rect 382740 318786 382792 318792
rect 382752 211886 382780 318786
rect 382844 237726 382872 396034
rect 382832 237720 382884 237726
rect 382832 237662 382884 237668
rect 382740 211880 382792 211886
rect 382740 211822 382792 211828
rect 382936 199345 382964 682314
rect 383016 667956 383068 667962
rect 383016 667898 383068 667904
rect 382922 199336 382978 199345
rect 382922 199271 382978 199280
rect 383028 198218 383056 667898
rect 383568 636268 383620 636274
rect 383568 636210 383620 636216
rect 383384 579692 383436 579698
rect 383384 579634 383436 579640
rect 383108 564596 383160 564602
rect 383108 564538 383160 564544
rect 383016 198212 383068 198218
rect 383016 198154 383068 198160
rect 383120 158642 383148 564538
rect 383200 517540 383252 517546
rect 383200 517482 383252 517488
rect 383108 158636 383160 158642
rect 383108 158578 383160 158584
rect 383212 150958 383240 517482
rect 383292 463752 383344 463758
rect 383292 463694 383344 463700
rect 383304 162178 383332 463694
rect 383396 320142 383424 579634
rect 383476 414044 383528 414050
rect 383476 413986 383528 413992
rect 383384 320136 383436 320142
rect 383384 320078 383436 320084
rect 383384 201544 383436 201550
rect 383384 201486 383436 201492
rect 383396 171834 383424 201486
rect 383384 171828 383436 171834
rect 383384 171770 383436 171776
rect 383292 162172 383344 162178
rect 383292 162114 383344 162120
rect 383488 155922 383516 413986
rect 383580 231441 383608 636210
rect 383660 364404 383712 364410
rect 383660 364346 383712 364352
rect 383566 231432 383622 231441
rect 383566 231367 383622 231376
rect 383672 184618 383700 364346
rect 384212 294636 384264 294642
rect 384212 294578 384264 294584
rect 383660 184612 383712 184618
rect 383660 184554 383712 184560
rect 383934 166288 383990 166297
rect 383934 166223 383990 166232
rect 383476 155916 383528 155922
rect 383476 155858 383528 155864
rect 383200 150952 383252 150958
rect 383200 150894 383252 150900
rect 382292 149926 383318 149954
rect 383948 149940 383976 166223
rect 384224 155553 384252 294578
rect 384210 155544 384266 155553
rect 384210 155479 384266 155488
rect 384316 152998 384344 684791
rect 384396 682032 384448 682038
rect 384396 681974 384448 681980
rect 384408 164082 384436 681974
rect 384488 567316 384540 567322
rect 384488 567258 384540 567264
rect 384396 164076 384448 164082
rect 384396 164018 384448 164024
rect 384500 163946 384528 567258
rect 384578 562592 384634 562601
rect 384578 562527 384634 562536
rect 384592 166569 384620 562527
rect 384672 516248 384724 516254
rect 384672 516190 384724 516196
rect 384578 166560 384634 166569
rect 384578 166495 384634 166504
rect 384488 163940 384540 163946
rect 384488 163882 384540 163888
rect 384578 157040 384634 157049
rect 384578 156975 384634 156984
rect 384304 152992 384356 152998
rect 384304 152934 384356 152940
rect 384592 149940 384620 156975
rect 384684 155689 384712 516190
rect 384856 481704 384908 481710
rect 384856 481646 384908 481652
rect 384764 472048 384816 472054
rect 384764 471990 384816 471996
rect 384776 234598 384804 471990
rect 384764 234592 384816 234598
rect 384764 234534 384816 234540
rect 384868 228410 384896 481646
rect 384960 240786 384988 686122
rect 388720 684616 388772 684622
rect 388720 684558 388772 684564
rect 385684 665236 385736 665242
rect 385684 665178 385736 665184
rect 385592 448588 385644 448594
rect 385592 448530 385644 448536
rect 385500 343664 385552 343670
rect 385500 343606 385552 343612
rect 385512 260846 385540 343606
rect 385500 260840 385552 260846
rect 385500 260782 385552 260788
rect 385500 258120 385552 258126
rect 385500 258062 385552 258068
rect 384948 240780 385000 240786
rect 384948 240722 385000 240728
rect 385040 235408 385092 235414
rect 385040 235350 385092 235356
rect 384856 228404 384908 228410
rect 384856 228346 384908 228352
rect 385052 171134 385080 235350
rect 385052 171106 385448 171134
rect 384670 155680 384726 155689
rect 384670 155615 384726 155624
rect 385420 149954 385448 171106
rect 385512 151774 385540 258062
rect 385604 235482 385632 448530
rect 385592 235476 385644 235482
rect 385592 235418 385644 235424
rect 385696 197946 385724 665178
rect 387248 661156 387300 661162
rect 387248 661098 387300 661104
rect 385960 567520 386012 567526
rect 385960 567462 386012 567468
rect 385776 563508 385828 563514
rect 385776 563450 385828 563456
rect 385684 197940 385736 197946
rect 385684 197882 385736 197888
rect 385788 153202 385816 563450
rect 385868 509312 385920 509318
rect 385868 509254 385920 509260
rect 385880 174894 385908 509254
rect 385972 237289 386000 567462
rect 387154 564768 387210 564777
rect 387154 564703 387210 564712
rect 387062 562320 387118 562329
rect 387062 562255 387118 562264
rect 386328 485852 386380 485858
rect 386328 485794 386380 485800
rect 386052 483064 386104 483070
rect 386052 483006 386104 483012
rect 385958 237280 386014 237289
rect 385958 237215 386014 237224
rect 385868 174888 385920 174894
rect 385868 174830 385920 174836
rect 386064 158506 386092 483006
rect 386236 467900 386288 467906
rect 386236 467842 386288 467848
rect 386144 462392 386196 462398
rect 386144 462334 386196 462340
rect 386156 236774 386184 462334
rect 386144 236768 386196 236774
rect 386144 236710 386196 236716
rect 386248 234190 386276 467842
rect 386236 234184 386288 234190
rect 386236 234126 386288 234132
rect 386052 158500 386104 158506
rect 386052 158442 386104 158448
rect 385776 153196 385828 153202
rect 385776 153138 385828 153144
rect 385500 151768 385552 151774
rect 385500 151710 385552 151716
rect 386340 149977 386368 485794
rect 386972 357468 387024 357474
rect 386972 357410 387024 357416
rect 386880 288448 386932 288454
rect 386880 288390 386932 288396
rect 386892 236842 386920 288390
rect 386880 236836 386932 236842
rect 386880 236778 386932 236784
rect 386984 228614 387012 357410
rect 386972 228608 387024 228614
rect 386972 228550 387024 228556
rect 386420 171828 386472 171834
rect 386420 171770 386472 171776
rect 386326 149968 386382 149977
rect 385420 149926 385894 149954
rect 386432 149954 386460 171770
rect 387076 154154 387104 562255
rect 387168 161129 387196 564703
rect 387260 275942 387288 661098
rect 387432 618316 387484 618322
rect 387432 618258 387484 618264
rect 387340 523116 387392 523122
rect 387340 523058 387392 523064
rect 387248 275936 387300 275942
rect 387248 275878 387300 275884
rect 387248 260840 387300 260846
rect 387248 260782 387300 260788
rect 387260 241330 387288 260782
rect 387248 241324 387300 241330
rect 387248 241266 387300 241272
rect 387352 181694 387380 523058
rect 387444 488510 387472 618258
rect 388444 576904 388496 576910
rect 388444 576846 388496 576852
rect 387524 495508 387576 495514
rect 387524 495450 387576 495456
rect 387432 488504 387484 488510
rect 387432 488446 387484 488452
rect 387536 456754 387564 495450
rect 387524 456748 387576 456754
rect 387524 456690 387576 456696
rect 387616 437504 387668 437510
rect 387616 437446 387668 437452
rect 387524 409896 387576 409902
rect 387524 409838 387576 409844
rect 387432 397588 387484 397594
rect 387432 397530 387484 397536
rect 387340 181688 387392 181694
rect 387340 181630 387392 181636
rect 387154 161120 387210 161129
rect 387154 161055 387210 161064
rect 387064 154148 387116 154154
rect 387064 154090 387116 154096
rect 386432 149926 387182 149954
rect 387444 149938 387472 397530
rect 387536 170406 387564 409838
rect 387628 224262 387656 437446
rect 387708 414044 387760 414050
rect 387708 413986 387760 413992
rect 387720 234326 387748 413986
rect 388352 394732 388404 394738
rect 388352 394674 388404 394680
rect 387800 380996 387852 381002
rect 387800 380938 387852 380944
rect 387708 234320 387760 234326
rect 387708 234262 387760 234268
rect 387616 224256 387668 224262
rect 387616 224198 387668 224204
rect 387524 170400 387576 170406
rect 387524 170342 387576 170348
rect 387812 151366 387840 380938
rect 388260 349172 388312 349178
rect 388260 349114 388312 349120
rect 388272 307766 388300 349114
rect 388260 307760 388312 307766
rect 388260 307702 388312 307708
rect 388364 231334 388392 394674
rect 388352 231328 388404 231334
rect 388352 231270 388404 231276
rect 388456 159798 388484 576846
rect 388536 550656 388588 550662
rect 388536 550598 388588 550604
rect 388548 211954 388576 550598
rect 388628 546508 388680 546514
rect 388628 546450 388680 546456
rect 388640 215966 388668 546450
rect 388732 356046 388760 684558
rect 392584 683732 392636 683738
rect 392584 683674 392636 683680
rect 389824 682304 389876 682310
rect 389824 682246 389876 682252
rect 389088 681760 389140 681766
rect 389088 681702 389140 681708
rect 388996 517540 389048 517546
rect 388996 517482 389048 517488
rect 388812 434784 388864 434790
rect 388812 434726 388864 434732
rect 388720 356040 388772 356046
rect 388720 355982 388772 355988
rect 388720 311908 388772 311914
rect 388720 311850 388772 311856
rect 388732 229974 388760 311850
rect 388720 229968 388772 229974
rect 388720 229910 388772 229916
rect 388628 215960 388680 215966
rect 388628 215902 388680 215908
rect 388536 211948 388588 211954
rect 388536 211890 388588 211896
rect 388824 169250 388852 434726
rect 388904 418260 388956 418266
rect 388904 418202 388956 418208
rect 388916 223582 388944 418202
rect 389008 233889 389036 517482
rect 389100 311953 389128 681702
rect 389180 563440 389232 563446
rect 389180 563382 389232 563388
rect 389086 311944 389142 311953
rect 389086 311879 389142 311888
rect 388994 233880 389050 233889
rect 388994 233815 389050 233824
rect 388904 223576 388956 223582
rect 388904 223518 388956 223524
rect 389088 204332 389140 204338
rect 389088 204274 389140 204280
rect 388812 169244 388864 169250
rect 388812 169186 388864 169192
rect 388444 159792 388496 159798
rect 388444 159734 388496 159740
rect 387800 151360 387852 151366
rect 387800 151302 387852 151308
rect 389100 149940 389128 204274
rect 389192 151814 389220 563382
rect 389732 266416 389784 266422
rect 389732 266358 389784 266364
rect 389744 161430 389772 266358
rect 389836 170542 389864 682246
rect 389916 563848 389968 563854
rect 389916 563790 389968 563796
rect 389824 170536 389876 170542
rect 389824 170478 389876 170484
rect 389732 161424 389784 161430
rect 389732 161366 389784 161372
rect 389928 152454 389956 563790
rect 390006 563272 390062 563281
rect 390006 563207 390062 563216
rect 390020 241262 390048 563207
rect 391480 561808 391532 561814
rect 391480 561750 391532 561756
rect 391296 559020 391348 559026
rect 391296 558962 391348 558968
rect 390376 524476 390428 524482
rect 390376 524418 390428 524424
rect 390284 422340 390336 422346
rect 390284 422282 390336 422288
rect 390192 411324 390244 411330
rect 390192 411266 390244 411272
rect 390100 390652 390152 390658
rect 390100 390594 390152 390600
rect 390008 241256 390060 241262
rect 390008 241198 390060 241204
rect 390112 194070 390140 390594
rect 390204 242894 390232 411266
rect 390192 242888 390244 242894
rect 390192 242830 390244 242836
rect 390296 228546 390324 422282
rect 390388 231266 390416 524418
rect 390468 473476 390520 473482
rect 390468 473418 390520 473424
rect 390376 231260 390428 231266
rect 390376 231202 390428 231208
rect 390284 228540 390336 228546
rect 390284 228482 390336 228488
rect 390100 194064 390152 194070
rect 390100 194006 390152 194012
rect 390480 155446 390508 473418
rect 391204 466472 391256 466478
rect 391204 466414 391256 466420
rect 391112 287224 391164 287230
rect 391112 287166 391164 287172
rect 391020 273284 391072 273290
rect 391020 273226 391072 273232
rect 391032 227118 391060 273226
rect 391020 227112 391072 227118
rect 391020 227054 391072 227060
rect 391124 191758 391152 287166
rect 391112 191752 391164 191758
rect 391112 191694 391164 191700
rect 391216 166598 391244 466414
rect 391308 277370 391336 558962
rect 391388 405748 391440 405754
rect 391388 405690 391440 405696
rect 391296 277364 391348 277370
rect 391296 277306 391348 277312
rect 391296 253972 391348 253978
rect 391296 253914 391348 253920
rect 391308 181626 391336 253914
rect 391296 181620 391348 181626
rect 391296 181562 391348 181568
rect 391400 174758 391428 405690
rect 391492 386374 391520 561750
rect 391848 495508 391900 495514
rect 391848 495450 391900 495456
rect 391756 488572 391808 488578
rect 391756 488514 391808 488520
rect 391664 411324 391716 411330
rect 391664 411266 391716 411272
rect 391572 401668 391624 401674
rect 391572 401610 391624 401616
rect 391480 386368 391532 386374
rect 391480 386310 391532 386316
rect 391480 350600 391532 350606
rect 391480 350542 391532 350548
rect 391492 177478 391520 350542
rect 391584 237114 391612 401610
rect 391572 237108 391624 237114
rect 391572 237050 391624 237056
rect 391480 177472 391532 177478
rect 391480 177414 391532 177420
rect 391388 174752 391440 174758
rect 391388 174694 391440 174700
rect 391204 166592 391256 166598
rect 391204 166534 391256 166540
rect 391676 161158 391704 411266
rect 391768 237318 391796 488514
rect 391756 237312 391808 237318
rect 391756 237254 391808 237260
rect 391860 166530 391888 495450
rect 392492 284368 392544 284374
rect 392492 284310 392544 284316
rect 392400 244316 392452 244322
rect 392400 244258 392452 244264
rect 392308 238876 392360 238882
rect 392308 238818 392360 238824
rect 392320 222970 392348 238818
rect 392308 222964 392360 222970
rect 392308 222906 392360 222912
rect 392412 190126 392440 244258
rect 392504 197062 392532 284310
rect 392492 197056 392544 197062
rect 392492 196998 392544 197004
rect 392400 190120 392452 190126
rect 392400 190062 392452 190068
rect 391848 166524 391900 166530
rect 391848 166466 391900 166472
rect 391664 161152 391716 161158
rect 391664 161094 391716 161100
rect 390468 155440 390520 155446
rect 390468 155382 390520 155388
rect 391664 153196 391716 153202
rect 391664 153138 391716 153144
rect 389916 152448 389968 152454
rect 389916 152390 389968 152396
rect 389192 151786 390048 151814
rect 390020 149954 390048 151786
rect 387432 149932 387484 149938
rect 386326 149903 386382 149912
rect 366824 149874 366876 149880
rect 390020 149926 390402 149954
rect 391676 149940 391704 153138
rect 392596 152862 392624 683674
rect 394238 680368 394294 680377
rect 394238 680303 394294 680312
rect 393964 661224 394016 661230
rect 393964 661166 394016 661172
rect 393228 637628 393280 637634
rect 393228 637570 393280 637576
rect 393136 587920 393188 587926
rect 393136 587862 393188 587868
rect 392676 566296 392728 566302
rect 392676 566238 392728 566244
rect 392584 152856 392636 152862
rect 392584 152798 392636 152804
rect 392688 151434 392716 566238
rect 392768 560516 392820 560522
rect 392768 560458 392820 560464
rect 392780 152318 392808 560458
rect 393044 437504 393096 437510
rect 393044 437446 393096 437452
rect 392952 380928 393004 380934
rect 392952 380870 393004 380876
rect 392860 314696 392912 314702
rect 392860 314638 392912 314644
rect 392872 166802 392900 314638
rect 392964 239630 392992 380870
rect 392952 239624 393004 239630
rect 392952 239566 393004 239572
rect 393056 239465 393084 437446
rect 393042 239456 393098 239465
rect 393042 239391 393098 239400
rect 393148 233782 393176 587862
rect 393136 233776 393188 233782
rect 393136 233718 393188 233724
rect 392860 166796 392912 166802
rect 392860 166738 392912 166744
rect 393240 159497 393268 637570
rect 393872 317484 393924 317490
rect 393872 317426 393924 317432
rect 393780 255332 393832 255338
rect 393780 255274 393832 255280
rect 393792 183326 393820 255274
rect 393884 235618 393912 317426
rect 393872 235612 393924 235618
rect 393872 235554 393924 235560
rect 393780 183320 393832 183326
rect 393780 183262 393832 183268
rect 393976 166433 394004 661166
rect 394054 564496 394110 564505
rect 394054 564431 394110 564440
rect 393962 166424 394018 166433
rect 393962 166359 394018 166368
rect 393226 159488 393282 159497
rect 393226 159423 393282 159432
rect 394068 152998 394096 564431
rect 394148 534132 394200 534138
rect 394148 534074 394200 534080
rect 394160 169386 394188 534074
rect 394148 169380 394200 169386
rect 394148 169322 394200 169328
rect 394056 152992 394108 152998
rect 394056 152934 394108 152940
rect 392768 152312 392820 152318
rect 392768 152254 392820 152260
rect 392676 151428 392728 151434
rect 392676 151370 392728 151376
rect 394252 149940 394280 680303
rect 395436 679040 395488 679046
rect 395436 678982 395488 678988
rect 395344 627972 395396 627978
rect 395344 627914 395396 627920
rect 394608 596216 394660 596222
rect 394608 596158 394660 596164
rect 394516 516248 394568 516254
rect 394516 516190 394568 516196
rect 394332 382288 394384 382294
rect 394332 382230 394384 382236
rect 394344 237250 394372 382230
rect 394424 380180 394476 380186
rect 394424 380122 394476 380128
rect 394332 237244 394384 237250
rect 394332 237186 394384 237192
rect 394436 155582 394464 380122
rect 394528 239902 394556 516190
rect 394516 239896 394568 239902
rect 394516 239838 394568 239844
rect 394620 157962 394648 596158
rect 395252 342304 395304 342310
rect 395252 342246 395304 342252
rect 395160 278792 395212 278798
rect 395160 278734 395212 278740
rect 395068 261112 395120 261118
rect 395068 261054 395120 261060
rect 395080 166734 395108 261054
rect 395172 234530 395200 278734
rect 395160 234524 395212 234530
rect 395160 234466 395212 234472
rect 395264 234258 395292 342246
rect 395356 270502 395384 627914
rect 395448 390522 395476 678982
rect 396724 618384 396776 618390
rect 396724 618326 396776 618332
rect 395528 563100 395580 563106
rect 395528 563042 395580 563048
rect 395540 447098 395568 563042
rect 395988 487212 396040 487218
rect 395988 487154 396040 487160
rect 395528 447092 395580 447098
rect 395528 447034 395580 447040
rect 395896 425128 395948 425134
rect 395896 425070 395948 425076
rect 395436 390516 395488 390522
rect 395436 390458 395488 390464
rect 395436 375420 395488 375426
rect 395436 375362 395488 375368
rect 395344 270496 395396 270502
rect 395344 270438 395396 270444
rect 395344 245676 395396 245682
rect 395344 245618 395396 245624
rect 395252 234252 395304 234258
rect 395252 234194 395304 234200
rect 395356 198014 395384 245618
rect 395344 198008 395396 198014
rect 395344 197950 395396 197956
rect 395068 166728 395120 166734
rect 395068 166670 395120 166676
rect 394608 157956 394660 157962
rect 394608 157898 394660 157904
rect 394424 155576 394476 155582
rect 394424 155518 394476 155524
rect 395448 152794 395476 375362
rect 395712 374060 395764 374066
rect 395712 374002 395764 374008
rect 395528 356108 395580 356114
rect 395528 356050 395580 356056
rect 395540 195702 395568 356050
rect 395620 288516 395672 288522
rect 395620 288458 395672 288464
rect 395528 195696 395580 195702
rect 395528 195638 395580 195644
rect 395632 163470 395660 288458
rect 395724 236978 395752 374002
rect 395804 320204 395856 320210
rect 395804 320146 395856 320152
rect 395712 236972 395764 236978
rect 395712 236914 395764 236920
rect 395620 163464 395672 163470
rect 395620 163406 395672 163412
rect 395436 152788 395488 152794
rect 395436 152730 395488 152736
rect 395816 151366 395844 320146
rect 395908 246362 395936 425070
rect 395896 246356 395948 246362
rect 395896 246298 395948 246304
rect 396000 166297 396028 487154
rect 396632 317484 396684 317490
rect 396632 317426 396684 317432
rect 396448 265668 396500 265674
rect 396448 265610 396500 265616
rect 396460 240009 396488 265610
rect 396540 259480 396592 259486
rect 396540 259422 396592 259428
rect 396446 240000 396502 240009
rect 396446 239935 396502 239944
rect 396552 198665 396580 259422
rect 396644 239290 396672 317426
rect 396736 261118 396764 618326
rect 396816 564664 396868 564670
rect 396816 564606 396868 564612
rect 396724 261112 396776 261118
rect 396724 261054 396776 261060
rect 396724 242956 396776 242962
rect 396724 242898 396776 242904
rect 396632 239284 396684 239290
rect 396632 239226 396684 239232
rect 396538 198656 396594 198665
rect 396538 198591 396594 198600
rect 395986 166288 396042 166297
rect 395986 166223 396042 166232
rect 396736 161226 396764 242898
rect 396828 237862 396856 564606
rect 396920 466410 396948 687346
rect 397368 682236 397420 682242
rect 397368 682178 397420 682184
rect 397000 676864 397052 676870
rect 397000 676806 397052 676812
rect 396908 466404 396960 466410
rect 396908 466346 396960 466352
rect 396908 462392 396960 462398
rect 396908 462334 396960 462340
rect 396816 237856 396868 237862
rect 396816 237798 396868 237804
rect 396920 188970 396948 462334
rect 397012 445670 397040 676806
rect 397276 501016 397328 501022
rect 397276 500958 397328 500964
rect 397000 445664 397052 445670
rect 397000 445606 397052 445612
rect 397184 427916 397236 427922
rect 397184 427858 397236 427864
rect 397000 397520 397052 397526
rect 397000 397462 397052 397468
rect 396908 188964 396960 188970
rect 396908 188906 396960 188912
rect 396724 161220 396776 161226
rect 396724 161162 396776 161168
rect 396172 155236 396224 155242
rect 396172 155178 396224 155184
rect 395804 151360 395856 151366
rect 395804 151302 395856 151308
rect 396184 149940 396212 155178
rect 397012 154494 397040 397462
rect 397092 387864 397144 387870
rect 397092 387806 397144 387812
rect 397000 154488 397052 154494
rect 397000 154430 397052 154436
rect 397104 154222 397132 387806
rect 397092 154216 397144 154222
rect 397092 154158 397144 154164
rect 397196 150414 397224 427858
rect 397288 164218 397316 500958
rect 397380 243545 397408 682178
rect 397472 663746 397500 703520
rect 400128 700664 400180 700670
rect 400128 700606 400180 700612
rect 399944 690668 399996 690674
rect 399944 690610 399996 690616
rect 398104 683596 398156 683602
rect 398104 683538 398156 683544
rect 397460 663740 397512 663746
rect 397460 663682 397512 663688
rect 398012 305040 398064 305046
rect 398012 304982 398064 304988
rect 397920 249824 397972 249830
rect 397920 249766 397972 249772
rect 397366 243536 397422 243545
rect 397366 243471 397422 243480
rect 397932 221474 397960 249766
rect 398024 233850 398052 304982
rect 398012 233844 398064 233850
rect 398012 233786 398064 233792
rect 397920 221468 397972 221474
rect 397920 221410 397972 221416
rect 397276 164212 397328 164218
rect 397276 164154 397328 164160
rect 398116 152697 398144 683538
rect 399484 679584 399536 679590
rect 399484 679526 399536 679532
rect 398748 594856 398800 594862
rect 398748 594798 398800 594804
rect 398288 563644 398340 563650
rect 398288 563586 398340 563592
rect 398194 560008 398250 560017
rect 398194 559943 398250 559952
rect 398208 152862 398236 559943
rect 398300 238513 398328 563586
rect 398564 552084 398616 552090
rect 398564 552026 398616 552032
rect 398472 517608 398524 517614
rect 398472 517550 398524 517556
rect 398380 393372 398432 393378
rect 398380 393314 398432 393320
rect 398392 315994 398420 393314
rect 398380 315988 398432 315994
rect 398380 315930 398432 315936
rect 398380 271924 398432 271930
rect 398380 271866 398432 271872
rect 398286 238504 398342 238513
rect 398286 238439 398342 238448
rect 398392 177410 398420 271866
rect 398484 234462 398512 517550
rect 398472 234456 398524 234462
rect 398472 234398 398524 234404
rect 398576 231130 398604 552026
rect 398656 550656 398708 550662
rect 398656 550598 398708 550604
rect 398564 231124 398616 231130
rect 398564 231066 398616 231072
rect 398380 177404 398432 177410
rect 398380 177346 398432 177352
rect 398668 157826 398696 550598
rect 398656 157820 398708 157826
rect 398656 157762 398708 157768
rect 398760 157010 398788 594798
rect 399496 588538 399524 679526
rect 399852 678292 399904 678298
rect 399852 678234 399904 678240
rect 399760 612808 399812 612814
rect 399760 612750 399812 612756
rect 399668 588600 399720 588606
rect 399668 588542 399720 588548
rect 399484 588532 399536 588538
rect 399484 588474 399536 588480
rect 399576 564800 399628 564806
rect 399576 564742 399628 564748
rect 399484 560720 399536 560726
rect 399484 560662 399536 560668
rect 399392 295384 399444 295390
rect 399392 295326 399444 295332
rect 399300 285796 399352 285802
rect 399300 285738 399352 285744
rect 399312 238610 399340 285738
rect 399300 238604 399352 238610
rect 399300 238546 399352 238552
rect 399404 231470 399432 295326
rect 399392 231464 399444 231470
rect 399392 231406 399444 231412
rect 398840 183456 398892 183462
rect 398840 183398 398892 183404
rect 398748 157004 398800 157010
rect 398748 156946 398800 156952
rect 398196 152856 398248 152862
rect 398196 152798 398248 152804
rect 398102 152688 398158 152697
rect 398102 152623 398158 152632
rect 397184 150408 397236 150414
rect 397184 150350 397236 150356
rect 398852 149954 398880 183398
rect 399496 152386 399524 560662
rect 399588 238649 399616 564742
rect 399680 292534 399708 588542
rect 399772 394670 399800 612750
rect 399864 509250 399892 678234
rect 399956 522986 399984 690610
rect 400036 683936 400088 683942
rect 400036 683878 400088 683884
rect 399944 522980 399996 522986
rect 399944 522922 399996 522928
rect 399852 509244 399904 509250
rect 399852 509186 399904 509192
rect 399760 394664 399812 394670
rect 399760 394606 399812 394612
rect 399944 372632 399996 372638
rect 399944 372574 399996 372580
rect 399852 311908 399904 311914
rect 399852 311850 399904 311856
rect 399760 310548 399812 310554
rect 399760 310490 399812 310496
rect 399668 292528 399720 292534
rect 399668 292470 399720 292476
rect 399668 245744 399720 245750
rect 399668 245686 399720 245692
rect 399574 238640 399630 238649
rect 399574 238575 399630 238584
rect 399680 177342 399708 245686
rect 399772 183190 399800 310490
rect 399760 183184 399812 183190
rect 399760 183126 399812 183132
rect 399668 177336 399720 177342
rect 399668 177278 399720 177284
rect 399484 152380 399536 152386
rect 399484 152322 399536 152328
rect 399864 151570 399892 311850
rect 399852 151564 399904 151570
rect 399852 151506 399904 151512
rect 399956 150113 399984 372574
rect 400048 238202 400076 683878
rect 400140 251190 400168 700606
rect 413664 700602 413692 703520
rect 413652 700596 413704 700602
rect 413652 700538 413704 700544
rect 405004 700528 405056 700534
rect 405004 700470 405056 700476
rect 400864 689376 400916 689382
rect 400864 689318 400916 689324
rect 400680 383716 400732 383722
rect 400680 383658 400732 383664
rect 400128 251184 400180 251190
rect 400128 251126 400180 251132
rect 400128 248464 400180 248470
rect 400128 248406 400180 248412
rect 400140 239766 400168 248406
rect 400128 239760 400180 239766
rect 400128 239702 400180 239708
rect 400036 238196 400088 238202
rect 400036 238138 400088 238144
rect 400692 231713 400720 383658
rect 400772 368552 400824 368558
rect 400772 368494 400824 368500
rect 400678 231704 400734 231713
rect 400678 231639 400734 231648
rect 400784 180130 400812 368494
rect 400876 238746 400904 689318
rect 403992 687472 404044 687478
rect 403992 687414 404044 687420
rect 402796 686044 402848 686050
rect 402796 685986 402848 685992
rect 402336 685568 402388 685574
rect 402336 685510 402388 685516
rect 402244 682440 402296 682446
rect 402244 682382 402296 682388
rect 400956 681012 401008 681018
rect 400956 680954 401008 680960
rect 400968 445738 400996 680954
rect 401508 590708 401560 590714
rect 401508 590650 401560 590656
rect 401048 567248 401100 567254
rect 401048 567190 401100 567196
rect 400956 445732 401008 445738
rect 400956 445674 401008 445680
rect 400956 418192 401008 418198
rect 400956 418134 401008 418140
rect 400864 238740 400916 238746
rect 400864 238682 400916 238688
rect 400772 180124 400824 180130
rect 400772 180066 400824 180072
rect 400680 162308 400732 162314
rect 400680 162250 400732 162256
rect 399942 150104 399998 150113
rect 399942 150039 399998 150048
rect 398852 149926 400062 149954
rect 400692 149940 400720 162250
rect 400968 157078 400996 418134
rect 401060 322862 401088 567190
rect 401140 563168 401192 563174
rect 401140 563110 401192 563116
rect 401152 441590 401180 563110
rect 401232 521756 401284 521762
rect 401232 521698 401284 521704
rect 401140 441584 401192 441590
rect 401140 441526 401192 441532
rect 401140 389224 401192 389230
rect 401140 389166 401192 389172
rect 401048 322856 401100 322862
rect 401048 322798 401100 322804
rect 401048 300960 401100 300966
rect 401048 300902 401100 300908
rect 401060 198082 401088 300902
rect 401048 198076 401100 198082
rect 401048 198018 401100 198024
rect 401152 159633 401180 389166
rect 401244 292466 401272 521698
rect 401416 477556 401468 477562
rect 401416 477498 401468 477504
rect 401324 465112 401376 465118
rect 401324 465054 401376 465060
rect 401232 292460 401284 292466
rect 401232 292402 401284 292408
rect 401232 260908 401284 260914
rect 401232 260850 401284 260856
rect 401244 174826 401272 260850
rect 401336 231198 401364 465054
rect 401324 231192 401376 231198
rect 401324 231134 401376 231140
rect 401324 229764 401376 229770
rect 401324 229706 401376 229712
rect 401232 174820 401284 174826
rect 401232 174762 401284 174768
rect 401138 159624 401194 159633
rect 401138 159559 401194 159568
rect 400956 157072 401008 157078
rect 400956 157014 401008 157020
rect 401336 149940 401364 229706
rect 401428 155786 401456 477498
rect 401416 155780 401468 155786
rect 401416 155722 401468 155728
rect 401520 152590 401548 590650
rect 402150 558240 402206 558249
rect 402150 558175 402206 558184
rect 402164 500954 402192 558175
rect 402152 500948 402204 500954
rect 402152 500890 402204 500896
rect 402152 323060 402204 323066
rect 402152 323002 402204 323008
rect 402060 278044 402112 278050
rect 402060 277986 402112 277992
rect 402072 237046 402100 277986
rect 402060 237040 402112 237046
rect 402060 236982 402112 236988
rect 402164 231402 402192 323002
rect 402152 231396 402204 231402
rect 402152 231338 402204 231344
rect 401968 178900 402020 178906
rect 401968 178842 402020 178848
rect 401508 152584 401560 152590
rect 401508 152526 401560 152532
rect 401980 149940 402008 178842
rect 402256 167754 402284 682382
rect 402348 589286 402376 685510
rect 402520 680536 402572 680542
rect 402520 680478 402572 680484
rect 402428 679652 402480 679658
rect 402428 679594 402480 679600
rect 402336 589280 402388 589286
rect 402336 589222 402388 589228
rect 402440 589014 402468 679594
rect 402428 589008 402480 589014
rect 402428 588950 402480 588956
rect 402428 564528 402480 564534
rect 402428 564470 402480 564476
rect 402336 563372 402388 563378
rect 402336 563314 402388 563320
rect 402244 167748 402296 167754
rect 402244 167690 402296 167696
rect 402348 151910 402376 563314
rect 402440 161265 402468 564470
rect 402532 405686 402560 680478
rect 402612 679176 402664 679182
rect 402612 679118 402664 679124
rect 402624 589082 402652 679118
rect 402704 650684 402756 650690
rect 402704 650626 402756 650632
rect 402612 589076 402664 589082
rect 402612 589018 402664 589024
rect 402716 528554 402744 650626
rect 402624 528526 402744 528554
rect 402624 525094 402652 528526
rect 402612 525088 402664 525094
rect 402612 525030 402664 525036
rect 402520 405680 402572 405686
rect 402520 405622 402572 405628
rect 402520 352028 402572 352034
rect 402520 351970 402572 351976
rect 402532 183462 402560 351970
rect 402624 244934 402652 525030
rect 402704 458244 402756 458250
rect 402704 458186 402756 458192
rect 402612 244928 402664 244934
rect 402612 244870 402664 244876
rect 402624 239698 402652 244870
rect 402612 239692 402664 239698
rect 402612 239634 402664 239640
rect 402520 183456 402572 183462
rect 402520 183398 402572 183404
rect 402426 161256 402482 161265
rect 402426 161191 402482 161200
rect 402716 153202 402744 458186
rect 402808 346390 402836 685986
rect 403716 681148 403768 681154
rect 403716 681090 403768 681096
rect 402888 644496 402940 644502
rect 402888 644438 402940 644444
rect 402796 346384 402848 346390
rect 402796 346326 402848 346332
rect 402796 267776 402848 267782
rect 402796 267718 402848 267724
rect 402808 159730 402836 267718
rect 402900 232354 402928 644438
rect 403624 560584 403676 560590
rect 403624 560526 403676 560532
rect 403532 310616 403584 310622
rect 403532 310558 403584 310564
rect 403440 277432 403492 277438
rect 403440 277374 403492 277380
rect 403452 238338 403480 277374
rect 403440 238332 403492 238338
rect 403440 238274 403492 238280
rect 402888 232348 402940 232354
rect 402888 232290 402940 232296
rect 402796 159724 402848 159730
rect 402796 159666 402848 159672
rect 402704 153196 402756 153202
rect 402704 153138 402756 153144
rect 403544 152522 403572 310558
rect 403636 153066 403664 560526
rect 403728 437442 403756 681090
rect 403808 680672 403860 680678
rect 403808 680614 403860 680620
rect 403820 506462 403848 680614
rect 403900 575544 403952 575550
rect 403900 575486 403952 575492
rect 403808 506456 403860 506462
rect 403808 506398 403860 506404
rect 403808 462460 403860 462466
rect 403808 462402 403860 462408
rect 403716 437436 403768 437442
rect 403716 437378 403768 437384
rect 403716 426488 403768 426494
rect 403716 426430 403768 426436
rect 403728 238678 403756 426430
rect 403716 238672 403768 238678
rect 403716 238614 403768 238620
rect 403820 232762 403848 462402
rect 403912 285666 403940 575486
rect 404004 574054 404032 687414
rect 404268 683528 404320 683534
rect 404268 683470 404320 683476
rect 404084 654220 404136 654226
rect 404084 654162 404136 654168
rect 403992 574048 404044 574054
rect 403992 573990 404044 573996
rect 403992 572756 404044 572762
rect 403992 572698 404044 572704
rect 403900 285660 403952 285666
rect 403900 285602 403952 285608
rect 404004 271862 404032 572698
rect 403992 271856 404044 271862
rect 403992 271798 404044 271804
rect 403900 262268 403952 262274
rect 403900 262210 403952 262216
rect 403808 232756 403860 232762
rect 403808 232698 403860 232704
rect 403912 162246 403940 262210
rect 403992 251252 404044 251258
rect 403992 251194 404044 251200
rect 403900 162240 403952 162246
rect 403900 162182 403952 162188
rect 404004 155106 404032 251194
rect 404096 240514 404124 654162
rect 404176 637696 404228 637702
rect 404176 637638 404228 637644
rect 404084 240508 404136 240514
rect 404084 240450 404136 240456
rect 404188 224466 404216 637638
rect 404280 603090 404308 683470
rect 404912 679244 404964 679250
rect 404912 679186 404964 679192
rect 404728 658300 404780 658306
rect 404728 658242 404780 658248
rect 404268 603084 404320 603090
rect 404268 603026 404320 603032
rect 404268 592068 404320 592074
rect 404268 592010 404320 592016
rect 404176 224460 404228 224466
rect 404176 224402 404228 224408
rect 404280 166433 404308 592010
rect 404266 166424 404322 166433
rect 404266 166359 404322 166368
rect 404740 164082 404768 658242
rect 404820 590912 404872 590918
rect 404820 590854 404872 590860
rect 404832 588849 404860 590854
rect 404924 589218 404952 679186
rect 404912 589212 404964 589218
rect 404912 589154 404964 589160
rect 404818 588840 404874 588849
rect 404818 588775 404874 588784
rect 405016 573374 405044 700470
rect 429856 698970 429884 703520
rect 429844 698964 429896 698970
rect 429844 698906 429896 698912
rect 462332 690674 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 690668 462372 690674
rect 462320 690610 462372 690616
rect 405096 687540 405148 687546
rect 405096 687482 405148 687488
rect 405108 588878 405136 687482
rect 407028 687336 407080 687342
rect 407028 687278 407080 687284
rect 405188 685908 405240 685914
rect 405188 685850 405240 685856
rect 405200 590918 405228 685850
rect 406660 684684 406712 684690
rect 406660 684626 406712 684632
rect 405280 684548 405332 684554
rect 405280 684490 405332 684496
rect 405188 590912 405240 590918
rect 405188 590854 405240 590860
rect 405188 590776 405240 590782
rect 405188 590718 405240 590724
rect 405096 588872 405148 588878
rect 405096 588814 405148 588820
rect 405200 588742 405228 590718
rect 405292 588946 405320 684490
rect 406568 681284 406620 681290
rect 406568 681226 406620 681232
rect 405464 680604 405516 680610
rect 405464 680546 405516 680552
rect 405370 679688 405426 679697
rect 405370 679623 405426 679632
rect 405280 588940 405332 588946
rect 405280 588882 405332 588888
rect 405188 588736 405240 588742
rect 405188 588678 405240 588684
rect 405384 585818 405412 679623
rect 405372 585812 405424 585818
rect 405372 585754 405424 585760
rect 405004 573368 405056 573374
rect 405004 573310 405056 573316
rect 405096 565956 405148 565962
rect 405096 565898 405148 565904
rect 405004 565888 405056 565894
rect 405004 565830 405056 565836
rect 405016 438870 405044 565830
rect 405004 438864 405056 438870
rect 405004 438806 405056 438812
rect 405004 427848 405056 427854
rect 405004 427790 405056 427796
rect 404912 287428 404964 287434
rect 404912 287370 404964 287376
rect 404924 228682 404952 287370
rect 405016 262206 405044 427790
rect 405108 416770 405136 565898
rect 405188 562692 405240 562698
rect 405188 562634 405240 562640
rect 405200 516118 405228 562634
rect 405280 560448 405332 560454
rect 405280 560390 405332 560396
rect 405292 552022 405320 560390
rect 405280 552016 405332 552022
rect 405280 551958 405332 551964
rect 405372 543856 405424 543862
rect 405372 543798 405424 543804
rect 405188 516112 405240 516118
rect 405188 516054 405240 516060
rect 405280 432540 405332 432546
rect 405280 432482 405332 432488
rect 405096 416764 405148 416770
rect 405096 416706 405148 416712
rect 405188 302252 405240 302258
rect 405188 302194 405240 302200
rect 405096 281444 405148 281450
rect 405096 281386 405148 281392
rect 405004 262200 405056 262206
rect 405004 262142 405056 262148
rect 405004 245812 405056 245818
rect 405004 245754 405056 245760
rect 405016 231538 405044 245754
rect 405004 231532 405056 231538
rect 405004 231474 405056 231480
rect 404912 228676 404964 228682
rect 404912 228618 404964 228624
rect 404728 164076 404780 164082
rect 404728 164018 404780 164024
rect 405108 160614 405136 281386
rect 405096 160608 405148 160614
rect 405096 160550 405148 160556
rect 403992 155100 404044 155106
rect 403992 155042 404044 155048
rect 405200 154562 405228 302194
rect 405292 167686 405320 432482
rect 405384 255270 405412 543798
rect 405476 485790 405504 680546
rect 406476 679380 406528 679386
rect 406476 679322 406528 679328
rect 405556 679312 405608 679318
rect 405556 679254 405608 679260
rect 405568 588810 405596 679254
rect 406382 642152 406438 642161
rect 406382 642087 406438 642096
rect 405556 588804 405608 588810
rect 405556 588746 405608 588752
rect 405556 564460 405608 564466
rect 405556 564402 405608 564408
rect 405464 485784 405516 485790
rect 405464 485726 405516 485732
rect 405464 452668 405516 452674
rect 405464 452610 405516 452616
rect 405372 255264 405424 255270
rect 405372 255206 405424 255212
rect 405372 251116 405424 251122
rect 405372 251058 405424 251064
rect 405280 167680 405332 167686
rect 405280 167622 405332 167628
rect 405384 155174 405412 251058
rect 405372 155168 405424 155174
rect 405372 155110 405424 155116
rect 405188 154556 405240 154562
rect 405188 154498 405240 154504
rect 403624 153060 403676 153066
rect 403624 153002 403676 153008
rect 405476 152658 405504 452610
rect 405568 238474 405596 564402
rect 406016 483064 406068 483070
rect 406016 483006 406068 483012
rect 405648 266416 405700 266422
rect 405648 266358 405700 266364
rect 405660 239834 405688 266358
rect 405648 239828 405700 239834
rect 405648 239770 405700 239776
rect 405556 238468 405608 238474
rect 405556 238410 405608 238416
rect 406028 152726 406056 483006
rect 406200 411392 406252 411398
rect 406200 411334 406252 411340
rect 406212 239494 406240 411334
rect 406292 408536 406344 408542
rect 406292 408478 406344 408484
rect 406200 239488 406252 239494
rect 406200 239430 406252 239436
rect 406304 232966 406332 408478
rect 406396 245818 406424 642087
rect 406488 459785 406516 679322
rect 406580 562358 406608 681226
rect 406568 562352 406620 562358
rect 406568 562294 406620 562300
rect 406566 531856 406622 531865
rect 406566 531791 406622 531800
rect 406474 459776 406530 459785
rect 406474 459711 406530 459720
rect 406474 429856 406530 429865
rect 406474 429791 406530 429800
rect 406384 245812 406436 245818
rect 406384 245754 406436 245760
rect 406292 232960 406344 232966
rect 406292 232902 406344 232908
rect 406488 203658 406516 429791
rect 406580 262993 406608 531791
rect 406672 372065 406700 684626
rect 406844 683324 406896 683330
rect 406844 683266 406896 683272
rect 406750 667856 406806 667865
rect 406750 667791 406806 667800
rect 406764 588674 406792 667791
rect 406752 588668 406804 588674
rect 406752 588610 406804 588616
rect 406750 556336 406806 556345
rect 406750 556271 406806 556280
rect 406658 372056 406714 372065
rect 406658 371991 406714 372000
rect 406658 356416 406714 356425
rect 406658 356351 406714 356360
rect 406566 262984 406622 262993
rect 406566 262919 406622 262928
rect 406568 262200 406620 262206
rect 406568 262142 406620 262148
rect 406580 237182 406608 262142
rect 406568 237176 406620 237182
rect 406568 237118 406620 237124
rect 406476 203652 406528 203658
rect 406476 203594 406528 203600
rect 406672 162178 406700 356351
rect 406764 239970 406792 556271
rect 406856 467945 406884 683266
rect 407040 644065 407068 687278
rect 413468 687268 413520 687274
rect 413468 687210 413520 687216
rect 407672 686112 407724 686118
rect 407672 686054 407724 686060
rect 407580 685500 407632 685506
rect 407580 685442 407632 685448
rect 407592 678230 407620 685442
rect 407580 678224 407632 678230
rect 407580 678166 407632 678172
rect 407118 678056 407174 678065
rect 407118 677991 407174 678000
rect 407132 677618 407160 677991
rect 407120 677612 407172 677618
rect 407120 677554 407172 677560
rect 407120 670676 407172 670682
rect 407120 670618 407172 670624
rect 407132 670585 407160 670618
rect 407118 670576 407174 670585
rect 407118 670511 407174 670520
rect 407118 669216 407174 669225
rect 407118 669151 407174 669160
rect 407132 667962 407160 669151
rect 407120 667956 407172 667962
rect 407120 667898 407172 667904
rect 407210 667176 407266 667185
rect 407210 667111 407266 667120
rect 407118 666496 407174 666505
rect 407118 666431 407174 666440
rect 407132 665242 407160 666431
rect 407120 665236 407172 665242
rect 407120 665178 407172 665184
rect 407224 665122 407252 667111
rect 407132 665094 407252 665122
rect 407026 644056 407082 644065
rect 407026 643991 407082 644000
rect 406934 631816 406990 631825
rect 406934 631751 406990 631760
rect 406842 467936 406898 467945
rect 406842 467871 406898 467880
rect 406844 246356 406896 246362
rect 406844 246298 406896 246304
rect 406752 239964 406804 239970
rect 406752 239906 406804 239912
rect 406856 239426 406884 246298
rect 406844 239420 406896 239426
rect 406844 239362 406896 239368
rect 406948 233238 406976 631751
rect 407026 625424 407082 625433
rect 407026 625359 407082 625368
rect 406936 233232 406988 233238
rect 406936 233174 406988 233180
rect 407040 213314 407068 625359
rect 407132 323202 407160 665094
rect 407210 663776 407266 663785
rect 407210 663711 407212 663720
rect 407264 663711 407266 663720
rect 407212 663682 407264 663688
rect 407394 662416 407450 662425
rect 407394 662351 407450 662360
rect 407210 661736 407266 661745
rect 407210 661671 407266 661680
rect 407224 661162 407252 661671
rect 407304 661224 407356 661230
rect 407304 661166 407356 661172
rect 407212 661156 407264 661162
rect 407212 661098 407264 661104
rect 407316 661065 407344 661166
rect 407408 661094 407436 662351
rect 407396 661088 407448 661094
rect 407302 661056 407358 661065
rect 407396 661030 407448 661036
rect 407302 660991 407358 661000
rect 407302 659016 407358 659025
rect 407302 658951 407358 658960
rect 407316 658306 407344 658951
rect 407304 658300 407356 658306
rect 407304 658242 407356 658248
rect 407212 655512 407264 655518
rect 407212 655454 407264 655460
rect 407224 654945 407252 655454
rect 407210 654936 407266 654945
rect 407210 654871 407266 654880
rect 407210 654256 407266 654265
rect 407210 654191 407212 654200
rect 407264 654191 407266 654200
rect 407212 654162 407264 654168
rect 407210 652896 407266 652905
rect 407210 652831 407266 652840
rect 407224 652798 407252 652831
rect 407212 652792 407264 652798
rect 407212 652734 407264 652740
rect 407212 650684 407264 650690
rect 407212 650626 407264 650632
rect 407224 650185 407252 650626
rect 407210 650176 407266 650185
rect 407210 650111 407266 650120
rect 407210 649496 407266 649505
rect 407210 649431 407266 649440
rect 407224 648650 407252 649431
rect 407486 648816 407542 648825
rect 407486 648751 407542 648760
rect 407212 648644 407264 648650
rect 407212 648586 407264 648592
rect 407210 644736 407266 644745
rect 407210 644671 407266 644680
rect 407224 644502 407252 644671
rect 407212 644496 407264 644502
rect 407212 644438 407264 644444
rect 407210 642016 407266 642025
rect 407210 641951 407266 641960
rect 407224 641782 407252 641951
rect 407212 641776 407264 641782
rect 407212 641718 407264 641724
rect 407210 641336 407266 641345
rect 407210 641271 407266 641280
rect 407224 640354 407252 641271
rect 407212 640348 407264 640354
rect 407212 640290 407264 640296
rect 407302 638072 407358 638081
rect 407302 638007 407358 638016
rect 407210 637936 407266 637945
rect 407210 637871 407266 637880
rect 407224 637634 407252 637871
rect 407316 637702 407344 638007
rect 407304 637696 407356 637702
rect 407304 637638 407356 637644
rect 407212 637628 407264 637634
rect 407212 637570 407264 637576
rect 407210 637256 407266 637265
rect 407210 637191 407266 637200
rect 407224 636274 407252 637191
rect 407212 636268 407264 636274
rect 407212 636210 407264 636216
rect 407210 633856 407266 633865
rect 407210 633791 407266 633800
rect 407224 633486 407252 633791
rect 407212 633480 407264 633486
rect 407212 633422 407264 633428
rect 407210 632496 407266 632505
rect 407210 632431 407266 632440
rect 407224 632126 407252 632431
rect 407212 632120 407264 632126
rect 407212 632062 407264 632068
rect 407210 629096 407266 629105
rect 407210 629031 407266 629040
rect 407224 627978 407252 629031
rect 407212 627972 407264 627978
rect 407212 627914 407264 627920
rect 407302 619576 407358 619585
rect 407302 619511 407358 619520
rect 407210 618896 407266 618905
rect 407210 618831 407266 618840
rect 407224 618322 407252 618831
rect 407316 618390 407344 619511
rect 407304 618384 407356 618390
rect 407304 618326 407356 618332
rect 407212 618316 407264 618322
rect 407212 618258 407264 618264
rect 407302 616856 407358 616865
rect 407302 616791 407358 616800
rect 407316 615534 407344 616791
rect 407304 615528 407356 615534
rect 407304 615470 407356 615476
rect 407302 614952 407358 614961
rect 407302 614887 407358 614896
rect 407212 612808 407264 612814
rect 407210 612776 407212 612785
rect 407264 612776 407266 612785
rect 407210 612711 407266 612720
rect 407210 608696 407266 608705
rect 407210 608631 407212 608640
rect 407264 608631 407266 608640
rect 407212 608602 407264 608608
rect 407316 605834 407344 614887
rect 407224 605806 407344 605834
rect 407224 440178 407252 605806
rect 407304 603084 407356 603090
rect 407304 603026 407356 603032
rect 407316 602585 407344 603026
rect 407302 602576 407358 602585
rect 407302 602511 407358 602520
rect 407302 601896 407358 601905
rect 407302 601831 407358 601840
rect 407316 601730 407344 601831
rect 407304 601724 407356 601730
rect 407304 601666 407356 601672
rect 407302 599176 407358 599185
rect 407302 599111 407358 599120
rect 407316 599010 407344 599111
rect 407304 599004 407356 599010
rect 407304 598946 407356 598952
rect 407302 597136 407358 597145
rect 407302 597071 407358 597080
rect 407316 596222 407344 597071
rect 407304 596216 407356 596222
rect 407304 596158 407356 596164
rect 407302 595096 407358 595105
rect 407302 595031 407358 595040
rect 407316 594862 407344 595031
rect 407304 594856 407356 594862
rect 407304 594798 407356 594804
rect 407302 593056 407358 593065
rect 407302 592991 407358 593000
rect 407316 592074 407344 592991
rect 407304 592068 407356 592074
rect 407304 592010 407356 592016
rect 407394 591152 407450 591161
rect 407394 591087 407450 591096
rect 407302 591016 407358 591025
rect 407302 590951 407358 590960
rect 407316 590714 407344 590951
rect 407408 590782 407436 591087
rect 407396 590776 407448 590782
rect 407396 590718 407448 590724
rect 407304 590708 407356 590714
rect 407304 590650 407356 590656
rect 407302 588976 407358 588985
rect 407302 588911 407358 588920
rect 407316 587926 407344 588911
rect 407500 588713 407528 648751
rect 407684 614825 407712 686054
rect 409696 685364 409748 685370
rect 409696 685306 409748 685312
rect 409052 685296 409104 685302
rect 409052 685238 409104 685244
rect 407764 685228 407816 685234
rect 407764 685170 407816 685176
rect 407776 678314 407804 685170
rect 407856 685160 407908 685166
rect 407856 685102 407908 685108
rect 407868 678434 407896 685102
rect 407948 683868 408000 683874
rect 407948 683810 408000 683816
rect 407856 678428 407908 678434
rect 407856 678370 407908 678376
rect 407776 678286 407896 678314
rect 407764 678224 407816 678230
rect 407764 678166 407816 678172
rect 407670 614816 407726 614825
rect 407670 614751 407726 614760
rect 407486 588704 407542 588713
rect 407486 588639 407542 588648
rect 407304 587920 407356 587926
rect 407304 587862 407356 587868
rect 407304 587512 407356 587518
rect 407304 587454 407356 587460
rect 407316 586945 407344 587454
rect 407302 586936 407358 586945
rect 407302 586871 407358 586880
rect 407776 586514 407804 678166
rect 407868 596174 407896 678286
rect 407960 605985 407988 683810
rect 408132 683664 408184 683670
rect 408132 683606 408184 683612
rect 408040 682100 408092 682106
rect 408040 682042 408092 682048
rect 408052 678570 408080 682042
rect 408040 678564 408092 678570
rect 408040 678506 408092 678512
rect 408040 678428 408092 678434
rect 408040 678370 408092 678376
rect 407946 605976 408002 605985
rect 407946 605911 408002 605920
rect 407868 596146 407988 596174
rect 407684 586486 407804 586514
rect 407684 585585 407712 586486
rect 407670 585576 407726 585585
rect 407670 585511 407726 585520
rect 407302 584896 407358 584905
rect 407302 584831 407358 584840
rect 407316 583778 407344 584831
rect 407304 583772 407356 583778
rect 407304 583714 407356 583720
rect 407302 580136 407358 580145
rect 407302 580071 407358 580080
rect 407316 579698 407344 580071
rect 407304 579692 407356 579698
rect 407304 579634 407356 579640
rect 407302 577416 407358 577425
rect 407302 577351 407358 577360
rect 407316 576910 407344 577351
rect 407304 576904 407356 576910
rect 407304 576846 407356 576852
rect 407302 576736 407358 576745
rect 407302 576671 407358 576680
rect 407316 575550 407344 576671
rect 407304 575544 407356 575550
rect 407304 575486 407356 575492
rect 407304 574048 407356 574054
rect 407302 574016 407304 574025
rect 407356 574016 407358 574025
rect 407302 573951 407358 573960
rect 407302 573336 407358 573345
rect 407302 573271 407358 573280
rect 407316 572762 407344 573271
rect 407304 572756 407356 572762
rect 407304 572698 407356 572704
rect 407302 572656 407358 572665
rect 407302 572591 407358 572600
rect 407316 571402 407344 572591
rect 407304 571396 407356 571402
rect 407304 571338 407356 571344
rect 407960 570625 407988 596146
rect 407946 570616 408002 570625
rect 407946 570551 408002 570560
rect 407302 569936 407358 569945
rect 407302 569871 407358 569880
rect 407316 568614 407344 569871
rect 407304 568608 407356 568614
rect 407304 568550 407356 568556
rect 407302 567896 407358 567905
rect 407302 567831 407358 567840
rect 407316 567390 407344 567831
rect 407304 567384 407356 567390
rect 407304 567326 407356 567332
rect 408052 565185 408080 678370
rect 408038 565176 408094 565185
rect 408038 565111 408094 565120
rect 407394 564496 407450 564505
rect 407394 564431 407396 564440
rect 407448 564431 407450 564440
rect 407396 564402 407448 564408
rect 407304 561672 407356 561678
rect 407304 561614 407356 561620
rect 407316 561105 407344 561614
rect 407854 561368 407910 561377
rect 407854 561303 407910 561312
rect 407302 561096 407358 561105
rect 407302 561031 407358 561040
rect 407764 560380 407816 560386
rect 407764 560322 407816 560328
rect 407580 559564 407632 559570
rect 407580 559506 407632 559512
rect 407592 555665 407620 559506
rect 407578 555656 407634 555665
rect 407578 555591 407634 555600
rect 407302 552936 407358 552945
rect 407302 552871 407358 552880
rect 407316 552090 407344 552871
rect 407304 552084 407356 552090
rect 407304 552026 407356 552032
rect 407396 552016 407448 552022
rect 407396 551958 407448 551964
rect 407408 551585 407436 551958
rect 407394 551576 407450 551585
rect 407394 551511 407450 551520
rect 407302 550896 407358 550905
rect 407302 550831 407358 550840
rect 407316 550662 407344 550831
rect 407304 550656 407356 550662
rect 407304 550598 407356 550604
rect 407302 550216 407358 550225
rect 407302 550151 407358 550160
rect 407316 549302 407344 550151
rect 407304 549296 407356 549302
rect 407304 549238 407356 549244
rect 407302 547496 407358 547505
rect 407302 547431 407358 547440
rect 407316 546582 407344 547431
rect 407304 546576 407356 546582
rect 407304 546518 407356 546524
rect 407776 546145 407804 560322
rect 407868 548865 407896 561303
rect 407948 559632 408000 559638
rect 407948 559574 408000 559580
rect 407960 557025 407988 559574
rect 408038 559056 408094 559065
rect 408038 558991 408094 559000
rect 407946 557016 408002 557025
rect 407946 556951 408002 556960
rect 407854 548856 407910 548865
rect 407854 548791 407910 548800
rect 407762 546136 407818 546145
rect 407762 546071 407818 546080
rect 407302 544776 407358 544785
rect 407302 544711 407358 544720
rect 407316 543794 407344 544711
rect 407394 544096 407450 544105
rect 407394 544031 407450 544040
rect 407408 543862 407436 544031
rect 407396 543856 407448 543862
rect 407396 543798 407448 543804
rect 407304 543788 407356 543794
rect 407304 543730 407356 543736
rect 407304 542360 407356 542366
rect 407304 542302 407356 542308
rect 407316 542065 407344 542302
rect 407302 542056 407358 542065
rect 407302 541991 407358 542000
rect 407762 537976 407818 537985
rect 407762 537911 407818 537920
rect 407302 535256 407358 535265
rect 407302 535191 407358 535200
rect 407316 534138 407344 535191
rect 407304 534132 407356 534138
rect 407304 534074 407356 534080
rect 407302 529136 407358 529145
rect 407302 529071 407358 529080
rect 407316 528630 407344 529071
rect 407304 528624 407356 528630
rect 407304 528566 407356 528572
rect 407394 525736 407450 525745
rect 407394 525671 407450 525680
rect 407304 525088 407356 525094
rect 407302 525056 407304 525065
rect 407356 525056 407358 525065
rect 407302 524991 407358 525000
rect 407408 524482 407436 525671
rect 407396 524476 407448 524482
rect 407396 524418 407448 524424
rect 407302 523696 407358 523705
rect 407302 523631 407358 523640
rect 407316 523122 407344 523631
rect 407304 523116 407356 523122
rect 407304 523058 407356 523064
rect 407394 523016 407450 523025
rect 407304 522980 407356 522986
rect 407394 522951 407450 522960
rect 407304 522922 407356 522928
rect 407316 522345 407344 522922
rect 407302 522336 407358 522345
rect 407302 522271 407358 522280
rect 407408 521762 407436 522951
rect 407396 521756 407448 521762
rect 407396 521698 407448 521704
rect 407302 521656 407358 521665
rect 407302 521591 407358 521600
rect 407316 520334 407344 521591
rect 407304 520328 407356 520334
rect 407304 520270 407356 520276
rect 407394 518256 407450 518265
rect 407394 518191 407450 518200
rect 407304 517608 407356 517614
rect 407302 517576 407304 517585
rect 407356 517576 407358 517585
rect 407408 517546 407436 518191
rect 407302 517511 407358 517520
rect 407396 517540 407448 517546
rect 407396 517482 407448 517488
rect 407394 516896 407450 516905
rect 407394 516831 407450 516840
rect 407304 516248 407356 516254
rect 407302 516216 407304 516225
rect 407356 516216 407358 516225
rect 407408 516186 407436 516831
rect 407302 516151 407358 516160
rect 407396 516180 407448 516186
rect 407396 516122 407448 516128
rect 407672 516112 407724 516118
rect 407672 516054 407724 516060
rect 407684 514865 407712 516054
rect 407670 514856 407726 514865
rect 407670 514791 407726 514800
rect 407304 513324 407356 513330
rect 407304 513266 407356 513272
rect 407316 512825 407344 513266
rect 407302 512816 407358 512825
rect 407302 512751 407358 512760
rect 407302 512136 407358 512145
rect 407302 512071 407358 512080
rect 407316 512038 407344 512071
rect 407304 512032 407356 512038
rect 407304 511974 407356 511980
rect 407302 509416 407358 509425
rect 407302 509351 407358 509360
rect 407316 509318 407344 509351
rect 407304 509312 407356 509318
rect 407304 509254 407356 509260
rect 407304 509176 407356 509182
rect 407304 509118 407356 509124
rect 407316 508065 407344 509118
rect 407302 508056 407358 508065
rect 407302 507991 407358 508000
rect 407302 506696 407358 506705
rect 407302 506631 407358 506640
rect 407316 506530 407344 506631
rect 407304 506524 407356 506530
rect 407304 506466 407356 506472
rect 407302 501256 407358 501265
rect 407302 501191 407358 501200
rect 407316 501022 407344 501191
rect 407304 501016 407356 501022
rect 407304 500958 407356 500964
rect 407396 500948 407448 500954
rect 407396 500890 407448 500896
rect 407408 500585 407436 500890
rect 407394 500576 407450 500585
rect 407394 500511 407450 500520
rect 407302 495816 407358 495825
rect 407302 495751 407358 495760
rect 407316 495514 407344 495751
rect 407304 495508 407356 495514
rect 407304 495450 407356 495456
rect 407302 493096 407358 493105
rect 407302 493031 407358 493040
rect 407316 492726 407344 493031
rect 407304 492720 407356 492726
rect 407304 492662 407356 492668
rect 407302 491056 407358 491065
rect 407302 490991 407358 491000
rect 407316 489938 407344 490991
rect 407304 489932 407356 489938
rect 407304 489874 407356 489880
rect 407302 489696 407358 489705
rect 407302 489631 407358 489640
rect 407316 488578 407344 489631
rect 407304 488572 407356 488578
rect 407304 488514 407356 488520
rect 407302 487656 407358 487665
rect 407302 487591 407358 487600
rect 407316 487218 407344 487591
rect 407304 487212 407356 487218
rect 407304 487154 407356 487160
rect 407302 486976 407358 486985
rect 407302 486911 407358 486920
rect 407316 485858 407344 486911
rect 407304 485852 407356 485858
rect 407304 485794 407356 485800
rect 407488 485784 407540 485790
rect 407488 485726 407540 485732
rect 407500 485625 407528 485726
rect 407486 485616 407542 485625
rect 407486 485551 407542 485560
rect 407302 484936 407358 484945
rect 407302 484871 407358 484880
rect 407316 484430 407344 484871
rect 407304 484424 407356 484430
rect 407304 484366 407356 484372
rect 407302 484256 407358 484265
rect 407302 484191 407358 484200
rect 407316 483138 407344 484191
rect 407304 483132 407356 483138
rect 407304 483074 407356 483080
rect 407302 482216 407358 482225
rect 407302 482151 407358 482160
rect 407316 481710 407344 482151
rect 407304 481704 407356 481710
rect 407304 481646 407356 481652
rect 407302 478136 407358 478145
rect 407302 478071 407358 478080
rect 407316 477562 407344 478071
rect 407304 477556 407356 477562
rect 407304 477498 407356 477504
rect 407302 475416 407358 475425
rect 407302 475351 407358 475360
rect 407316 474842 407344 475351
rect 407304 474836 407356 474842
rect 407304 474778 407356 474784
rect 407394 474736 407450 474745
rect 407394 474671 407450 474680
rect 407302 474056 407358 474065
rect 407302 473991 407358 474000
rect 407316 473482 407344 473991
rect 407304 473476 407356 473482
rect 407304 473418 407356 473424
rect 407408 473414 407436 474671
rect 407396 473408 407448 473414
rect 407396 473350 407448 473356
rect 407304 472048 407356 472054
rect 407302 472016 407304 472025
rect 407356 472016 407358 472025
rect 407302 471951 407358 471960
rect 407302 469976 407358 469985
rect 407302 469911 407358 469920
rect 407316 469266 407344 469911
rect 407304 469260 407356 469266
rect 407304 469202 407356 469208
rect 407302 468208 407358 468217
rect 407302 468143 407358 468152
rect 407316 467906 407344 468143
rect 407304 467900 407356 467906
rect 407304 467842 407356 467848
rect 407302 465896 407358 465905
rect 407302 465831 407358 465840
rect 407316 465118 407344 465831
rect 407304 465112 407356 465118
rect 407304 465054 407356 465060
rect 407302 463856 407358 463865
rect 407302 463791 407358 463800
rect 407316 463758 407344 463791
rect 407304 463752 407356 463758
rect 407304 463694 407356 463700
rect 407394 463176 407450 463185
rect 407394 463111 407450 463120
rect 407302 462496 407358 462505
rect 407408 462466 407436 463111
rect 407302 462431 407358 462440
rect 407396 462460 407448 462466
rect 407316 462398 407344 462431
rect 407396 462402 407448 462408
rect 407304 462392 407356 462398
rect 407304 462334 407356 462340
rect 407302 459096 407358 459105
rect 407302 459031 407358 459040
rect 407316 458250 407344 459031
rect 407304 458244 407356 458250
rect 407304 458186 407356 458192
rect 407302 457056 407358 457065
rect 407302 456991 407358 457000
rect 407316 456822 407344 456991
rect 407304 456816 407356 456822
rect 407304 456758 407356 456764
rect 407396 456748 407448 456754
rect 407396 456690 407448 456696
rect 407408 455705 407436 456690
rect 407394 455696 407450 455705
rect 407394 455631 407450 455640
rect 407396 455388 407448 455394
rect 407396 455330 407448 455336
rect 407302 455016 407358 455025
rect 407302 454951 407358 454960
rect 407316 454102 407344 454951
rect 407408 454345 407436 455330
rect 407394 454336 407450 454345
rect 407394 454271 407450 454280
rect 407304 454096 407356 454102
rect 407304 454038 407356 454044
rect 407670 452976 407726 452985
rect 407670 452911 407726 452920
rect 407684 452674 407712 452911
rect 407672 452668 407724 452674
rect 407672 452610 407724 452616
rect 407302 451616 407358 451625
rect 407302 451551 407358 451560
rect 407316 451382 407344 451551
rect 407304 451376 407356 451382
rect 407304 451318 407356 451324
rect 407302 449576 407358 449585
rect 407302 449511 407358 449520
rect 407316 448594 407344 449511
rect 407304 448588 407356 448594
rect 407304 448530 407356 448536
rect 407302 447264 407358 447273
rect 407302 447199 407358 447208
rect 407316 447166 407344 447199
rect 407304 447160 407356 447166
rect 407304 447102 407356 447108
rect 407396 447092 407448 447098
rect 407396 447034 407448 447040
rect 407408 446185 407436 447034
rect 407394 446176 407450 446185
rect 407394 446111 407450 446120
rect 407304 445664 407356 445670
rect 407304 445606 407356 445612
rect 407316 444825 407344 445606
rect 407302 444816 407358 444825
rect 407302 444751 407358 444760
rect 407302 442096 407358 442105
rect 407302 442031 407358 442040
rect 407316 441658 407344 442031
rect 407304 441652 407356 441658
rect 407304 441594 407356 441600
rect 407396 441584 407448 441590
rect 407396 441526 407448 441532
rect 407408 441425 407436 441526
rect 407394 441416 407450 441425
rect 407394 441351 407450 441360
rect 407224 440150 407344 440178
rect 407210 440056 407266 440065
rect 407210 439991 407266 440000
rect 407224 438938 407252 439991
rect 407212 438932 407264 438938
rect 407212 438874 407264 438880
rect 407210 438016 407266 438025
rect 407210 437951 407266 437960
rect 407224 437510 407252 437951
rect 407212 437504 407264 437510
rect 407212 437446 407264 437452
rect 407210 437336 407266 437345
rect 407210 437271 407266 437280
rect 407224 436150 407252 437271
rect 407212 436144 407264 436150
rect 407212 436086 407264 436092
rect 407210 435976 407266 435985
rect 407210 435911 407266 435920
rect 407224 434790 407252 435911
rect 407212 434784 407264 434790
rect 407212 434726 407264 434732
rect 407316 434625 407344 440150
rect 407488 438864 407540 438870
rect 407488 438806 407540 438812
rect 407500 438705 407528 438806
rect 407486 438696 407542 438705
rect 407486 438631 407542 438640
rect 407302 434616 407358 434625
rect 407302 434551 407358 434560
rect 407210 433256 407266 433265
rect 407210 433191 407266 433200
rect 407224 432546 407252 433191
rect 407212 432540 407264 432546
rect 407212 432482 407264 432488
rect 407210 429176 407266 429185
rect 407210 429111 407266 429120
rect 407224 427922 407252 429111
rect 407212 427916 407264 427922
rect 407212 427858 407264 427864
rect 407302 427816 407358 427825
rect 407302 427751 407358 427760
rect 407210 427136 407266 427145
rect 407210 427071 407266 427080
rect 407224 426562 407252 427071
rect 407316 426630 407344 427751
rect 407304 426624 407356 426630
rect 407304 426566 407356 426572
rect 407212 426556 407264 426562
rect 407212 426498 407264 426504
rect 407210 425776 407266 425785
rect 407210 425711 407266 425720
rect 407224 425134 407252 425711
rect 407212 425128 407264 425134
rect 407212 425070 407264 425076
rect 407210 423736 407266 423745
rect 407210 423671 407212 423680
rect 407264 423671 407266 423680
rect 407212 423642 407264 423648
rect 407210 423056 407266 423065
rect 407210 422991 407266 423000
rect 407224 422346 407252 422991
rect 407212 422340 407264 422346
rect 407212 422282 407264 422288
rect 407302 420336 407358 420345
rect 407302 420271 407358 420280
rect 407210 419656 407266 419665
rect 407316 419626 407344 420271
rect 407210 419591 407266 419600
rect 407304 419620 407356 419626
rect 407224 419558 407252 419591
rect 407304 419562 407356 419568
rect 407212 419552 407264 419558
rect 407212 419494 407264 419500
rect 407210 418976 407266 418985
rect 407210 418911 407266 418920
rect 407224 418266 407252 418911
rect 407212 418260 407264 418266
rect 407212 418202 407264 418208
rect 407580 416764 407632 416770
rect 407580 416706 407632 416712
rect 407592 416265 407620 416706
rect 407578 416256 407634 416265
rect 407578 416191 407634 416200
rect 407210 414896 407266 414905
rect 407210 414831 407266 414840
rect 407224 414050 407252 414831
rect 407212 414044 407264 414050
rect 407212 413986 407264 413992
rect 407302 412176 407358 412185
rect 407302 412111 407358 412120
rect 407210 411496 407266 411505
rect 407210 411431 407266 411440
rect 407224 411330 407252 411431
rect 407316 411398 407344 412111
rect 407304 411392 407356 411398
rect 407304 411334 407356 411340
rect 407212 411324 407264 411330
rect 407212 411266 407264 411272
rect 407210 410816 407266 410825
rect 407210 410751 407266 410760
rect 407224 409902 407252 410751
rect 407212 409896 407264 409902
rect 407212 409838 407264 409844
rect 407210 407416 407266 407425
rect 407210 407351 407266 407360
rect 407224 407182 407252 407351
rect 407212 407176 407264 407182
rect 407212 407118 407264 407124
rect 407210 406056 407266 406065
rect 407210 405991 407266 406000
rect 407224 405754 407252 405991
rect 407212 405748 407264 405754
rect 407212 405690 407264 405696
rect 407304 405680 407356 405686
rect 407304 405622 407356 405628
rect 407316 404705 407344 405622
rect 407302 404696 407358 404705
rect 407302 404631 407358 404640
rect 407210 401976 407266 401985
rect 407210 401911 407266 401920
rect 407224 401674 407252 401911
rect 407212 401668 407264 401674
rect 407212 401610 407264 401616
rect 407210 397896 407266 397905
rect 407210 397831 407266 397840
rect 407224 397594 407252 397831
rect 407212 397588 407264 397594
rect 407212 397530 407264 397536
rect 407210 395856 407266 395865
rect 407210 395791 407266 395800
rect 407224 394738 407252 395791
rect 407212 394732 407264 394738
rect 407212 394674 407264 394680
rect 407210 393816 407266 393825
rect 407210 393751 407266 393760
rect 407224 393378 407252 393751
rect 407212 393372 407264 393378
rect 407212 393314 407264 393320
rect 407302 391776 407358 391785
rect 407302 391711 407358 391720
rect 407210 391096 407266 391105
rect 407210 391031 407266 391040
rect 407224 390658 407252 391031
rect 407212 390652 407264 390658
rect 407212 390594 407264 390600
rect 407316 390590 407344 391711
rect 407304 390584 407356 390590
rect 407304 390526 407356 390532
rect 407212 386368 407264 386374
rect 407212 386310 407264 386316
rect 407224 385665 407252 386310
rect 407210 385656 407266 385665
rect 407210 385591 407266 385600
rect 407210 384976 407266 384985
rect 407210 384911 407266 384920
rect 407224 383722 407252 384911
rect 407212 383716 407264 383722
rect 407212 383658 407264 383664
rect 407210 381576 407266 381585
rect 407210 381511 407266 381520
rect 407224 381070 407252 381511
rect 407212 381064 407264 381070
rect 407212 381006 407264 381012
rect 407210 378856 407266 378865
rect 407210 378791 407266 378800
rect 407224 378214 407252 378791
rect 407212 378208 407264 378214
rect 407212 378150 407264 378156
rect 407210 374096 407266 374105
rect 407210 374031 407212 374040
rect 407264 374031 407266 374040
rect 407212 374002 407264 374008
rect 407210 373416 407266 373425
rect 407210 373351 407266 373360
rect 407224 372638 407252 373351
rect 407212 372632 407264 372638
rect 407212 372574 407264 372580
rect 407212 371204 407264 371210
rect 407212 371146 407264 371152
rect 407224 370705 407252 371146
rect 407210 370696 407266 370705
rect 407210 370631 407266 370640
rect 407210 369336 407266 369345
rect 407210 369271 407266 369280
rect 407224 368558 407252 369271
rect 407212 368552 407264 368558
rect 407212 368494 407264 368500
rect 407212 361548 407264 361554
rect 407212 361490 407264 361496
rect 407224 361185 407252 361490
rect 407210 361176 407266 361185
rect 407210 361111 407266 361120
rect 407210 360496 407266 360505
rect 407210 360431 407266 360440
rect 407224 360262 407252 360431
rect 407212 360256 407264 360262
rect 407212 360198 407264 360204
rect 407210 357776 407266 357785
rect 407210 357711 407266 357720
rect 407224 357474 407252 357711
rect 407212 357468 407264 357474
rect 407212 357410 407264 357416
rect 407210 357096 407266 357105
rect 407210 357031 407266 357040
rect 407224 356114 407252 357031
rect 407212 356108 407264 356114
rect 407212 356050 407264 356056
rect 407210 353696 407266 353705
rect 407210 353631 407266 353640
rect 407224 353326 407252 353631
rect 407212 353320 407264 353326
rect 407212 353262 407264 353268
rect 407302 353016 407358 353025
rect 407302 352951 407358 352960
rect 407210 352336 407266 352345
rect 407210 352271 407266 352280
rect 407224 352034 407252 352271
rect 407212 352028 407264 352034
rect 407212 351970 407264 351976
rect 407316 351966 407344 352951
rect 407304 351960 407356 351966
rect 407304 351902 407356 351908
rect 407210 351656 407266 351665
rect 407210 351591 407266 351600
rect 407224 350606 407252 351591
rect 407212 350600 407264 350606
rect 407212 350542 407264 350548
rect 407210 349344 407266 349353
rect 407210 349279 407266 349288
rect 407224 349246 407252 349279
rect 407212 349240 407264 349246
rect 407212 349182 407264 349188
rect 407212 346384 407264 346390
rect 407212 346326 407264 346332
rect 407224 345545 407252 346326
rect 407210 345536 407266 345545
rect 407210 345471 407266 345480
rect 407212 345024 407264 345030
rect 407212 344966 407264 344972
rect 407224 344865 407252 344966
rect 407210 344856 407266 344865
rect 407210 344791 407266 344800
rect 407210 343496 407266 343505
rect 407210 343431 407266 343440
rect 407224 342310 407252 343431
rect 407212 342304 407264 342310
rect 407212 342246 407264 342252
rect 407210 340776 407266 340785
rect 407210 340711 407266 340720
rect 407224 339522 407252 340711
rect 407212 339516 407264 339522
rect 407212 339458 407264 339464
rect 407212 336728 407264 336734
rect 407210 336696 407212 336705
rect 407264 336696 407266 336705
rect 407210 336631 407266 336640
rect 407302 332616 407358 332625
rect 407302 332551 407358 332560
rect 407212 331288 407264 331294
rect 407210 331256 407212 331265
rect 407264 331256 407266 331265
rect 407210 331191 407266 331200
rect 407210 330576 407266 330585
rect 407210 330511 407266 330520
rect 407224 329866 407252 330511
rect 407212 329860 407264 329866
rect 407212 329802 407264 329808
rect 407210 328536 407266 328545
rect 407210 328471 407212 328480
rect 407264 328471 407266 328480
rect 407212 328442 407264 328448
rect 407212 325644 407264 325650
rect 407212 325586 407264 325592
rect 407224 325145 407252 325586
rect 407210 325136 407266 325145
rect 407210 325071 407266 325080
rect 407210 323776 407266 323785
rect 407210 323711 407266 323720
rect 407120 323196 407172 323202
rect 407120 323138 407172 323144
rect 407118 323096 407174 323105
rect 407224 323066 407252 323711
rect 407118 323031 407174 323040
rect 407212 323060 407264 323066
rect 407132 322998 407160 323031
rect 407212 323002 407264 323008
rect 407120 322992 407172 322998
rect 407120 322934 407172 322940
rect 407212 322924 407264 322930
rect 407212 322866 407264 322872
rect 407120 322856 407172 322862
rect 407120 322798 407172 322804
rect 407132 322425 407160 322798
rect 407118 322416 407174 322425
rect 407118 322351 407174 322360
rect 407224 321745 407252 322866
rect 407210 321736 407266 321745
rect 407210 321671 407266 321680
rect 407118 321056 407174 321065
rect 407118 320991 407174 321000
rect 407132 320210 407160 320991
rect 407120 320204 407172 320210
rect 407120 320146 407172 320152
rect 407118 318336 407174 318345
rect 407118 318271 407174 318280
rect 407132 317490 407160 318271
rect 407120 317484 407172 317490
rect 407120 317426 407172 317432
rect 407118 312896 407174 312905
rect 407118 312831 407174 312840
rect 407132 311914 407160 312831
rect 407120 311908 407172 311914
rect 407120 311850 407172 311856
rect 407210 311128 407266 311137
rect 407210 311063 407266 311072
rect 407118 310856 407174 310865
rect 407118 310791 407174 310800
rect 407132 310622 407160 310791
rect 407120 310616 407172 310622
rect 407120 310558 407172 310564
rect 407224 310554 407252 311063
rect 407212 310548 407264 310554
rect 407212 310490 407264 310496
rect 407120 310480 407172 310486
rect 407120 310422 407172 310428
rect 407132 310185 407160 310422
rect 407118 310176 407174 310185
rect 407118 310111 407174 310120
rect 407118 308136 407174 308145
rect 407118 308071 407174 308080
rect 407132 307834 407160 308071
rect 407120 307828 407172 307834
rect 407120 307770 407172 307776
rect 407212 307760 407264 307766
rect 407212 307702 407264 307708
rect 407224 306785 407252 307702
rect 407210 306776 407266 306785
rect 407210 306711 407266 306720
rect 407118 305416 407174 305425
rect 407118 305351 407174 305360
rect 407132 305046 407160 305351
rect 407120 305040 407172 305046
rect 407120 304982 407172 304988
rect 407118 304056 407174 304065
rect 407118 303991 407174 304000
rect 407132 303686 407160 303991
rect 407120 303680 407172 303686
rect 407120 303622 407172 303628
rect 407210 302016 407266 302025
rect 407210 301951 407266 301960
rect 407118 301336 407174 301345
rect 407118 301271 407174 301280
rect 407132 300966 407160 301271
rect 407120 300960 407172 300966
rect 407120 300902 407172 300908
rect 407224 300898 407252 301951
rect 407212 300892 407264 300898
rect 407212 300834 407264 300840
rect 407118 299976 407174 299985
rect 407118 299911 407174 299920
rect 407132 299538 407160 299911
rect 407120 299532 407172 299538
rect 407120 299474 407172 299480
rect 407118 295896 407174 295905
rect 407118 295831 407174 295840
rect 407132 295390 407160 295831
rect 407120 295384 407172 295390
rect 407120 295326 407172 295332
rect 407210 293856 407266 293865
rect 407210 293791 407266 293800
rect 407118 293176 407174 293185
rect 407118 293111 407174 293120
rect 407132 292670 407160 293111
rect 407120 292664 407172 292670
rect 407120 292606 407172 292612
rect 407224 292602 407252 293791
rect 407212 292596 407264 292602
rect 407212 292538 407264 292544
rect 407120 292528 407172 292534
rect 407118 292496 407120 292505
rect 407172 292496 407174 292505
rect 407118 292431 407174 292440
rect 407212 292460 407264 292466
rect 407212 292402 407264 292408
rect 407224 291825 407252 292402
rect 407210 291816 407266 291825
rect 407210 291751 407266 291760
rect 407118 289096 407174 289105
rect 407118 289031 407174 289040
rect 407132 288522 407160 289031
rect 407120 288516 407172 288522
rect 407120 288458 407172 288464
rect 407118 288416 407174 288425
rect 407118 288351 407174 288360
rect 407132 287230 407160 288351
rect 407210 287736 407266 287745
rect 407210 287671 407266 287680
rect 407224 287434 407252 287671
rect 407212 287428 407264 287434
rect 407212 287370 407264 287376
rect 407120 287224 407172 287230
rect 407120 287166 407172 287172
rect 407118 287056 407174 287065
rect 407118 286991 407174 287000
rect 407132 285734 407160 286991
rect 407120 285728 407172 285734
rect 407120 285670 407172 285676
rect 407212 285660 407264 285666
rect 407212 285602 407264 285608
rect 407224 285025 407252 285602
rect 407210 285016 407266 285025
rect 407210 284951 407266 284960
rect 407120 284368 407172 284374
rect 407118 284336 407120 284345
rect 407172 284336 407174 284345
rect 407118 284271 407174 284280
rect 407212 284300 407264 284306
rect 407212 284242 407264 284248
rect 407224 283665 407252 284242
rect 407210 283656 407266 283665
rect 407210 283591 407266 283600
rect 407118 282976 407174 282985
rect 407118 282911 407120 282920
rect 407172 282911 407174 282920
rect 407120 282882 407172 282888
rect 407118 278896 407174 278905
rect 407118 278831 407174 278840
rect 407132 278798 407160 278831
rect 407120 278792 407172 278798
rect 407120 278734 407172 278740
rect 407120 277364 407172 277370
rect 407120 277306 407172 277312
rect 407132 276185 407160 277306
rect 407118 276176 407174 276185
rect 407118 276111 407174 276120
rect 407120 276004 407172 276010
rect 407120 275946 407172 275952
rect 407132 275505 407160 275946
rect 407118 275496 407174 275505
rect 407118 275431 407174 275440
rect 407118 272776 407174 272785
rect 407118 272711 407174 272720
rect 407132 271930 407160 272711
rect 407120 271924 407172 271930
rect 407120 271866 407172 271872
rect 407212 271856 407264 271862
rect 407212 271798 407264 271804
rect 407224 271425 407252 271798
rect 407210 271416 407266 271425
rect 407210 271351 407266 271360
rect 407118 270056 407174 270065
rect 407118 269991 407174 270000
rect 407132 269142 407160 269991
rect 407120 269136 407172 269142
rect 407120 269078 407172 269084
rect 407118 268016 407174 268025
rect 407118 267951 407174 267960
rect 407132 267782 407160 267951
rect 407120 267776 407172 267782
rect 407120 267718 407172 267724
rect 407118 263936 407174 263945
rect 407118 263871 407174 263880
rect 407132 263634 407160 263871
rect 407120 263628 407172 263634
rect 407120 263570 407172 263576
rect 407118 262576 407174 262585
rect 407118 262511 407174 262520
rect 407132 262274 407160 262511
rect 407120 262268 407172 262274
rect 407120 262210 407172 262216
rect 407118 261896 407174 261905
rect 407118 261831 407174 261840
rect 407132 260914 407160 261831
rect 407120 260908 407172 260914
rect 407120 260850 407172 260856
rect 407118 259856 407174 259865
rect 407118 259791 407174 259800
rect 407132 259486 407160 259791
rect 407120 259480 407172 259486
rect 407120 259422 407172 259428
rect 407210 257816 407266 257825
rect 407210 257751 407266 257760
rect 407118 257136 407174 257145
rect 407118 257071 407174 257080
rect 407132 256834 407160 257071
rect 407120 256828 407172 256834
rect 407120 256770 407172 256776
rect 407224 256766 407252 257751
rect 407212 256760 407264 256766
rect 407212 256702 407264 256708
rect 407118 255096 407174 255105
rect 407118 255031 407174 255040
rect 407132 253978 407160 255031
rect 407120 253972 407172 253978
rect 407120 253914 407172 253920
rect 407210 251696 407266 251705
rect 407210 251631 407266 251640
rect 407224 251258 407252 251631
rect 407212 251252 407264 251258
rect 407212 251194 407264 251200
rect 407120 251184 407172 251190
rect 407120 251126 407172 251132
rect 407132 250345 407160 251126
rect 407210 251016 407266 251025
rect 407210 250951 407266 250960
rect 407118 250336 407174 250345
rect 407118 250271 407174 250280
rect 407224 249898 407252 250951
rect 407212 249892 407264 249898
rect 407212 249834 407264 249840
rect 407210 246936 407266 246945
rect 407210 246871 407266 246880
rect 407118 246256 407174 246265
rect 407118 246191 407174 246200
rect 407132 245682 407160 246191
rect 407224 245750 407252 246871
rect 407212 245744 407264 245750
rect 407212 245686 407264 245692
rect 407120 245676 407172 245682
rect 407120 245618 407172 245624
rect 407210 245576 407266 245585
rect 407210 245511 407266 245520
rect 407224 244934 407252 245511
rect 407212 244928 407264 244934
rect 407118 244896 407174 244905
rect 407212 244870 407264 244876
rect 407118 244831 407174 244840
rect 407132 244322 407160 244831
rect 407120 244316 407172 244322
rect 407120 244258 407172 244264
rect 407120 242888 407172 242894
rect 407120 242830 407172 242836
rect 407132 242185 407160 242830
rect 407118 242176 407174 242185
rect 407118 242111 407174 242120
rect 407028 213308 407080 213314
rect 407028 213250 407080 213256
rect 407120 185768 407172 185774
rect 407120 185710 407172 185716
rect 406660 162172 406712 162178
rect 406660 162114 406712 162120
rect 406476 157888 406528 157894
rect 406476 157830 406528 157836
rect 406016 152720 406068 152726
rect 406016 152662 406068 152668
rect 405464 152652 405516 152658
rect 405464 152594 405516 152600
rect 403532 152516 403584 152522
rect 403532 152458 403584 152464
rect 402336 151904 402388 151910
rect 402336 151846 402388 151852
rect 403256 151904 403308 151910
rect 403256 151846 403308 151852
rect 403268 149940 403296 151846
rect 406488 149940 406516 157830
rect 407132 149940 407160 185710
rect 407212 183320 407264 183326
rect 407212 183262 407264 183268
rect 407224 149954 407252 183262
rect 407316 151026 407344 332551
rect 407396 323196 407448 323202
rect 407396 323138 407448 323144
rect 407408 319025 407436 323138
rect 407394 319016 407450 319025
rect 407394 318951 407450 318960
rect 407394 302696 407450 302705
rect 407394 302631 407450 302640
rect 407408 302258 407436 302631
rect 407396 302252 407448 302258
rect 407396 302194 407448 302200
rect 407670 298616 407726 298625
rect 407670 298551 407726 298560
rect 407488 272604 407540 272610
rect 407488 272546 407540 272552
rect 407500 262177 407528 272546
rect 407486 262168 407542 262177
rect 407486 262103 407542 262112
rect 407396 255264 407448 255270
rect 407396 255206 407448 255212
rect 407408 254425 407436 255206
rect 407394 254416 407450 254425
rect 407394 254351 407450 254360
rect 407684 242593 407712 298551
rect 407776 272610 407804 537911
rect 407854 483576 407910 483585
rect 407854 483511 407910 483520
rect 407868 483070 407896 483511
rect 407856 483064 407908 483070
rect 407856 483006 407908 483012
rect 407946 395176 408002 395185
rect 407946 395111 408002 395120
rect 407960 383654 407988 395111
rect 407868 383626 407988 383654
rect 407868 380186 407896 383626
rect 407946 383072 408002 383081
rect 407946 383007 408002 383016
rect 407856 380180 407908 380186
rect 407856 380122 407908 380128
rect 407856 320884 407908 320890
rect 407856 320826 407908 320832
rect 407764 272604 407816 272610
rect 407764 272546 407816 272552
rect 407762 267336 407818 267345
rect 407762 267271 407818 267280
rect 407776 266422 407804 267271
rect 407764 266416 407816 266422
rect 407764 266358 407816 266364
rect 407762 242992 407818 243001
rect 407762 242927 407818 242936
rect 407670 242584 407726 242593
rect 407670 242519 407726 242528
rect 407776 231674 407804 242927
rect 407764 231668 407816 231674
rect 407764 231610 407816 231616
rect 407868 183122 407896 320826
rect 407960 229770 407988 383007
rect 408052 362545 408080 558991
rect 408144 461145 408172 683606
rect 408316 683392 408368 683398
rect 408316 683334 408368 683340
rect 408224 681080 408276 681086
rect 408224 681022 408276 681028
rect 408236 650185 408264 681022
rect 408328 679425 408356 683334
rect 408960 680808 409012 680814
rect 408960 680750 409012 680756
rect 408408 679448 408460 679454
rect 408314 679416 408370 679425
rect 408408 679390 408460 679396
rect 408314 679351 408370 679360
rect 408316 678564 408368 678570
rect 408316 678506 408368 678512
rect 408222 650176 408278 650185
rect 408222 650111 408278 650120
rect 408328 635594 408356 678506
rect 408420 665145 408448 679390
rect 408406 665136 408462 665145
rect 408406 665071 408462 665080
rect 408406 646776 408462 646785
rect 408406 646711 408462 646720
rect 408316 635588 408368 635594
rect 408316 635530 408368 635536
rect 408316 635384 408368 635390
rect 408316 635326 408368 635332
rect 408224 628652 408276 628658
rect 408224 628594 408276 628600
rect 408236 476241 408264 628594
rect 408222 476232 408278 476241
rect 408222 476167 408278 476176
rect 408222 476096 408278 476105
rect 408222 476031 408278 476040
rect 408130 461136 408186 461145
rect 408130 461071 408186 461080
rect 408130 408776 408186 408785
rect 408130 408711 408186 408720
rect 408144 408542 408172 408711
rect 408132 408536 408184 408542
rect 408132 408478 408184 408484
rect 408130 382936 408186 382945
rect 408130 382871 408186 382880
rect 408038 362536 408094 362545
rect 408038 362471 408094 362480
rect 408038 346896 408094 346905
rect 408038 346831 408094 346840
rect 408052 278050 408080 346831
rect 408040 278044 408092 278050
rect 408040 277986 408092 277992
rect 408038 276856 408094 276865
rect 408038 276791 408094 276800
rect 407948 229764 408000 229770
rect 407948 229706 408000 229712
rect 408052 185638 408080 276791
rect 408040 185632 408092 185638
rect 408040 185574 408092 185580
rect 407856 183116 407908 183122
rect 407856 183058 407908 183064
rect 408144 164150 408172 382871
rect 408236 231742 408264 476031
rect 408328 457745 408356 635326
rect 408420 628658 408448 646711
rect 408408 628652 408460 628658
rect 408408 628594 408460 628600
rect 408406 594416 408462 594425
rect 408406 594351 408462 594360
rect 408420 586265 408448 594351
rect 408406 586256 408462 586265
rect 408406 586191 408462 586200
rect 408972 578105 409000 680750
rect 408958 578096 409014 578105
rect 408958 578031 409014 578040
rect 409064 510105 409092 685238
rect 409144 684888 409196 684894
rect 409144 684830 409196 684836
rect 409050 510096 409106 510105
rect 409050 510031 409106 510040
rect 409156 479505 409184 684830
rect 409328 684752 409380 684758
rect 409328 684694 409380 684700
rect 409236 684004 409288 684010
rect 409236 683946 409288 683952
rect 409142 479496 409198 479505
rect 409142 479431 409198 479440
rect 409248 476785 409276 683946
rect 409234 476776 409290 476785
rect 409234 476711 409290 476720
rect 409234 467256 409290 467265
rect 409234 467191 409290 467200
rect 408314 457736 408370 457745
rect 408314 457671 408370 457680
rect 408406 433936 408462 433945
rect 408406 433871 408462 433880
rect 408420 426426 408448 433871
rect 408408 426420 408460 426426
rect 408408 426362 408460 426368
rect 409144 426420 409196 426426
rect 409144 426362 409196 426368
rect 408314 421696 408370 421705
rect 408314 421631 408370 421640
rect 408224 231736 408276 231742
rect 408224 231678 408276 231684
rect 408132 164144 408184 164150
rect 408132 164086 408184 164092
rect 408328 155242 408356 421631
rect 408866 400344 408922 400353
rect 408866 400279 408922 400288
rect 408406 389736 408462 389745
rect 408406 389671 408462 389680
rect 408420 379522 408448 389671
rect 408420 379494 408540 379522
rect 408406 327856 408462 327865
rect 408406 327791 408462 327800
rect 408420 320890 408448 327791
rect 408408 320884 408460 320890
rect 408408 320826 408460 320832
rect 408406 259992 408462 260001
rect 408406 259927 408462 259936
rect 408420 239873 408448 259927
rect 408512 251122 408540 379494
rect 408500 251116 408552 251122
rect 408500 251058 408552 251064
rect 408406 239864 408462 239873
rect 408406 239799 408462 239808
rect 408880 232422 408908 400279
rect 409050 319696 409106 319705
rect 409050 319631 409106 319640
rect 408958 249656 409014 249665
rect 408958 249591 409014 249600
rect 408972 238542 409000 249591
rect 408960 238536 409012 238542
rect 408960 238478 409012 238484
rect 408868 232416 408920 232422
rect 408868 232358 408920 232364
rect 409064 229906 409092 319631
rect 409156 238270 409184 426362
rect 409248 281450 409276 467191
rect 409340 430545 409368 684694
rect 409420 683188 409472 683194
rect 409420 683130 409472 683136
rect 409326 430536 409382 430545
rect 409326 430471 409382 430480
rect 409432 428505 409460 683130
rect 409512 681896 409564 681902
rect 409512 681838 409564 681844
rect 409418 428496 409474 428505
rect 409418 428431 409474 428440
rect 409524 399265 409552 681838
rect 409604 680876 409656 680882
rect 409604 680818 409656 680824
rect 409510 399256 409566 399265
rect 409510 399191 409566 399200
rect 409326 393136 409382 393145
rect 409326 393071 409382 393080
rect 409340 300665 409368 393071
rect 409616 377505 409644 680818
rect 409602 377496 409658 377505
rect 409602 377431 409658 377440
rect 409708 364585 409736 685306
rect 411628 681828 411680 681834
rect 411628 681770 411680 681776
rect 409880 680740 409932 680746
rect 409880 680682 409932 680688
rect 409788 679516 409840 679522
rect 409788 679458 409840 679464
rect 409694 364576 409750 364585
rect 409694 364511 409750 364520
rect 409418 342816 409474 342825
rect 409418 342751 409474 342760
rect 409326 300656 409382 300665
rect 409326 300591 409382 300600
rect 409326 293992 409382 294001
rect 409326 293927 409382 293936
rect 409236 281444 409288 281450
rect 409236 281386 409288 281392
rect 409234 279576 409290 279585
rect 409234 279511 409290 279520
rect 409248 240582 409276 279511
rect 409236 240576 409288 240582
rect 409236 240518 409288 240524
rect 409144 238264 409196 238270
rect 409144 238206 409196 238212
rect 409340 236638 409368 293927
rect 409328 236632 409380 236638
rect 409328 236574 409380 236580
rect 409432 235210 409460 342751
rect 409694 339416 409750 339425
rect 409694 339351 409750 339360
rect 409602 289776 409658 289785
rect 409602 289711 409658 289720
rect 409510 241224 409566 241233
rect 409510 241159 409512 241168
rect 409564 241159 409566 241168
rect 409512 241130 409564 241136
rect 409510 240816 409566 240825
rect 409510 240751 409566 240760
rect 409524 240650 409552 240751
rect 409512 240644 409564 240650
rect 409512 240586 409564 240592
rect 409420 235204 409472 235210
rect 409420 235146 409472 235152
rect 409052 229900 409104 229906
rect 409052 229842 409104 229848
rect 409616 155718 409644 289711
rect 409604 155712 409656 155718
rect 409604 155654 409656 155660
rect 408316 155236 408368 155242
rect 408316 155178 408368 155184
rect 409708 154358 409736 339351
rect 409800 334665 409828 679458
rect 409892 678298 409920 680682
rect 411640 679946 411668 681770
rect 412916 681760 412968 681766
rect 412916 681702 412968 681708
rect 412928 679946 412956 681702
rect 413480 679946 413508 687210
rect 446404 686180 446456 686186
rect 446404 686122 446456 686128
rect 425794 684584 425850 684593
rect 425794 684519 425850 684528
rect 437572 684548 437624 684554
rect 424506 683496 424562 683505
rect 416688 683460 416740 683466
rect 424506 683431 424562 683440
rect 416688 683402 416740 683408
rect 416594 682952 416650 682961
rect 416594 682887 416650 682896
rect 416608 682174 416636 682887
rect 416596 682168 416648 682174
rect 416596 682110 416648 682116
rect 415490 682000 415546 682009
rect 415490 681935 415546 681944
rect 415504 679946 415532 681935
rect 416700 679946 416728 683402
rect 422392 682372 422444 682378
rect 422392 682314 422444 682320
rect 420000 681216 420052 681222
rect 420000 681158 420052 681164
rect 411640 679918 411976 679946
rect 412928 679918 413264 679946
rect 413480 679918 413908 679946
rect 415504 679918 415840 679946
rect 416484 679918 416728 679946
rect 420012 679946 420040 681158
rect 420012 679918 420348 679946
rect 422404 679810 422432 682314
rect 424520 679946 424548 683431
rect 424600 683188 424652 683194
rect 424600 683130 424652 683136
rect 424212 679918 424548 679946
rect 424612 679946 424640 683130
rect 425808 679946 425836 684519
rect 437572 684490 437624 684496
rect 436100 683868 436152 683874
rect 436100 683810 436152 683816
rect 429016 683800 429068 683806
rect 429016 683742 429068 683748
rect 427820 681216 427872 681222
rect 427820 681158 427872 681164
rect 427832 680785 427860 681158
rect 427912 681012 427964 681018
rect 427912 680954 427964 680960
rect 427818 680776 427874 680785
rect 427818 680711 427874 680720
rect 427084 680400 427136 680406
rect 427084 680342 427136 680348
rect 424612 679918 424856 679946
rect 425500 679918 425836 679946
rect 422280 679782 422432 679810
rect 427096 679658 427124 680342
rect 427924 679946 427952 680954
rect 429028 679946 429056 683742
rect 429660 683732 429712 683738
rect 429660 683674 429712 683680
rect 435456 683732 435508 683738
rect 435456 683674 435508 683680
rect 427924 679918 428076 679946
rect 428720 679918 429056 679946
rect 429672 679946 429700 683674
rect 432880 682168 432932 682174
rect 432880 682110 432932 682116
rect 432052 680944 432104 680950
rect 432052 680886 432104 680892
rect 429672 679918 430008 679946
rect 432064 679810 432092 680886
rect 432892 679946 432920 682110
rect 434628 680944 434680 680950
rect 434628 680886 434680 680892
rect 433844 680096 433900 680105
rect 433844 680031 433900 680040
rect 432584 679918 432920 679946
rect 433858 679932 433886 680031
rect 434640 679946 434668 680886
rect 435468 679946 435496 683674
rect 434516 679918 434668 679946
rect 435160 679918 435496 679946
rect 436112 679946 436140 683810
rect 437584 679946 437612 684490
rect 438676 683868 438728 683874
rect 438676 683810 438728 683816
rect 438688 679946 438716 683810
rect 445114 683768 445170 683777
rect 445114 683703 445170 683712
rect 442538 683224 442594 683233
rect 442538 683159 442594 683168
rect 442262 682816 442318 682825
rect 442262 682751 442318 682760
rect 440424 682440 440476 682446
rect 440424 682382 440476 682388
rect 440056 681760 440108 681766
rect 440056 681702 440108 681708
rect 439320 681080 439372 681086
rect 439320 681022 439372 681028
rect 439332 679946 439360 681022
rect 440068 681018 440096 681702
rect 440330 681184 440386 681193
rect 440330 681119 440386 681128
rect 440344 681086 440372 681119
rect 440332 681080 440384 681086
rect 440332 681022 440384 681028
rect 440056 681012 440108 681018
rect 440056 680954 440108 680960
rect 440148 680400 440200 680406
rect 440148 680342 440200 680348
rect 436112 679918 436448 679946
rect 437584 679918 437736 679946
rect 438380 679918 438716 679946
rect 439024 679918 439360 679946
rect 431940 679782 432092 679810
rect 440160 679658 440188 680342
rect 440436 679810 440464 682382
rect 441894 682272 441950 682281
rect 442276 682242 442304 682751
rect 441894 682207 441950 682216
rect 442264 682236 442316 682242
rect 441250 680776 441306 680785
rect 441250 680711 441306 680720
rect 441264 679946 441292 680711
rect 440956 679918 441292 679946
rect 441908 679946 441936 682207
rect 442264 682178 442316 682184
rect 442552 679946 442580 683159
rect 445128 679946 445156 683703
rect 446416 679946 446444 686122
rect 476578 686080 476634 686089
rect 476578 686015 476634 686024
rect 468392 685568 468444 685574
rect 468392 685510 468444 685516
rect 456800 685500 456852 685506
rect 456800 685442 456852 685448
rect 450268 685364 450320 685370
rect 450268 685306 450320 685312
rect 447690 682680 447746 682689
rect 447690 682615 447746 682624
rect 447704 679946 447732 682615
rect 450280 679946 450308 685306
rect 454224 685296 454276 685302
rect 454224 685238 454276 685244
rect 453856 684820 453908 684826
rect 453856 684762 453908 684768
rect 453868 680218 453896 684762
rect 453822 680190 453896 680218
rect 441908 679918 442244 679946
rect 442552 679918 442888 679946
rect 445128 679918 445464 679946
rect 446416 679918 446752 679946
rect 447704 679918 448040 679946
rect 450280 679918 450616 679946
rect 453822 679932 453850 680190
rect 454236 679946 454264 685238
rect 454774 684856 454830 684865
rect 454774 684791 454830 684800
rect 454788 679946 454816 684791
rect 456812 679946 456840 685442
rect 468300 685092 468352 685098
rect 468300 685034 468352 685040
rect 458638 682544 458694 682553
rect 458638 682479 458694 682488
rect 458180 682236 458232 682242
rect 458180 682178 458232 682184
rect 458192 681766 458220 682178
rect 458180 681760 458232 681766
rect 458180 681702 458232 681708
rect 457352 681284 457404 681290
rect 457352 681226 457404 681232
rect 457364 679946 457392 681226
rect 458192 679946 458220 681702
rect 458652 679946 458680 682479
rect 462502 682408 462558 682417
rect 462502 682343 462558 682352
rect 461216 680468 461268 680474
rect 461216 680410 461268 680416
rect 461228 679946 461256 680410
rect 462516 679946 462544 682343
rect 467010 681184 467066 681193
rect 463792 681148 463844 681154
rect 467010 681119 467066 681128
rect 463792 681090 463844 681096
rect 463804 679946 463832 681090
rect 467024 679946 467052 681119
rect 468312 679946 468340 685034
rect 454236 679918 454480 679946
rect 454788 679918 455124 679946
rect 456812 679918 457056 679946
rect 457364 679918 457700 679946
rect 458192 679918 458344 679946
rect 458652 679918 458988 679946
rect 461228 679918 461564 679946
rect 462516 679918 462852 679946
rect 463804 679918 464140 679946
rect 466716 679918 467052 679946
rect 468004 679918 468340 679946
rect 468404 679946 468432 685510
rect 470876 685228 470928 685234
rect 470876 685170 470928 685176
rect 470600 684956 470652 684962
rect 470600 684898 470652 684904
rect 470612 680218 470640 684898
rect 470566 680190 470640 680218
rect 468404 679918 468648 679946
rect 470566 679932 470594 680190
rect 470888 679946 470916 685170
rect 473544 685024 473596 685030
rect 473544 684966 473596 684972
rect 472162 681048 472218 681057
rect 472162 680983 472218 680992
rect 472176 679946 472204 680983
rect 473556 679946 473584 684966
rect 476488 684956 476540 684962
rect 476488 684898 476540 684904
rect 476500 679946 476528 684898
rect 470888 679918 471224 679946
rect 472176 679918 472512 679946
rect 473556 679918 473800 679946
rect 476376 679918 476528 679946
rect 476592 679946 476620 686015
rect 477512 682446 477540 702406
rect 484400 700732 484452 700738
rect 484400 700674 484452 700680
rect 484412 692774 484440 700674
rect 527192 700670 527220 703520
rect 543476 700738 543504 703520
rect 543464 700732 543516 700738
rect 543464 700674 543516 700680
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 551284 700596 551336 700602
rect 551284 700538 551336 700544
rect 498200 700460 498252 700466
rect 498200 700402 498252 700408
rect 484412 692746 484992 692774
rect 477500 682440 477552 682446
rect 477500 682382 477552 682388
rect 480352 682304 480404 682310
rect 480352 682246 480404 682252
rect 484860 682304 484912 682310
rect 484860 682246 484912 682252
rect 476592 679918 477020 679946
rect 480364 679810 480392 682246
rect 481178 681048 481234 681057
rect 481178 680983 481234 680992
rect 481192 679946 481220 680983
rect 484872 679946 484900 682246
rect 480884 679918 481220 679946
rect 484748 679918 484900 679946
rect 484964 679946 484992 692746
rect 487620 685024 487672 685030
rect 487620 684966 487672 684972
rect 487632 679946 487660 684966
rect 489552 684548 489604 684554
rect 489552 684490 489604 684496
rect 488722 680912 488778 680921
rect 488722 680847 488778 680856
rect 484964 679918 485392 679946
rect 487324 679918 487660 679946
rect 440312 679782 440464 679810
rect 480240 679782 480392 679810
rect 488736 679674 488764 680847
rect 489564 679946 489592 684490
rect 497280 684004 497332 684010
rect 497280 683946 497332 683952
rect 495164 682508 495216 682514
rect 495164 682450 495216 682456
rect 495176 679946 495204 682450
rect 496636 680468 496688 680474
rect 496636 680410 496688 680416
rect 496648 679946 496676 680410
rect 489256 679918 489592 679946
rect 495052 679918 495204 679946
rect 496340 679918 496676 679946
rect 497292 679946 497320 683946
rect 498212 680218 498240 700402
rect 550916 698964 550968 698970
rect 550916 698906 550968 698912
rect 550272 690668 550324 690674
rect 550272 690610 550324 690616
rect 538220 687948 538272 687954
rect 538220 687890 538272 687896
rect 528836 685976 528888 685982
rect 528836 685918 528888 685924
rect 514760 685432 514812 685438
rect 514760 685374 514812 685380
rect 509240 685160 509292 685166
rect 509240 685102 509292 685108
rect 502524 684072 502576 684078
rect 502524 684014 502576 684020
rect 499854 683632 499910 683641
rect 499854 683567 499910 683576
rect 499212 681148 499264 681154
rect 499212 681090 499264 681096
rect 498212 680190 498286 680218
rect 497292 679918 497628 679946
rect 498258 679932 498286 680190
rect 499224 679946 499252 681090
rect 498916 679918 499252 679946
rect 499868 679946 499896 683567
rect 502248 682372 502300 682378
rect 502248 682314 502300 682320
rect 501788 681284 501840 681290
rect 501788 681226 501840 681232
rect 500498 680640 500554 680649
rect 500498 680575 500554 680584
rect 500512 679946 500540 680575
rect 501800 679946 501828 681226
rect 502260 679946 502288 682314
rect 499868 679918 500204 679946
rect 500512 679918 500848 679946
rect 501492 679918 501828 679946
rect 502136 679918 502288 679946
rect 502536 679946 502564 684014
rect 507582 682680 507638 682689
rect 507582 682615 507638 682624
rect 505098 681864 505154 681873
rect 505098 681799 505154 681808
rect 504364 681216 504416 681222
rect 504364 681158 504416 681164
rect 504376 679946 504404 681158
rect 505112 679946 505140 681799
rect 507596 679946 507624 682615
rect 509252 680218 509280 685102
rect 509516 683256 509568 683262
rect 509516 683198 509568 683204
rect 502536 679918 502780 679946
rect 504376 679918 504712 679946
rect 505112 679918 505356 679946
rect 507288 679918 507624 679946
rect 509206 680190 509280 680218
rect 509206 679932 509234 680190
rect 509528 679946 509556 683198
rect 510528 683188 510580 683194
rect 510528 683130 510580 683136
rect 510540 680218 510568 683130
rect 512736 681828 512788 681834
rect 512736 681770 512788 681776
rect 510494 680190 510568 680218
rect 509528 679918 509864 679946
rect 510494 679932 510522 680190
rect 512748 679946 512776 681770
rect 512440 679918 512776 679946
rect 514772 679946 514800 685374
rect 523040 684888 523092 684894
rect 523040 684830 523092 684836
rect 521844 683936 521896 683942
rect 521844 683878 521896 683884
rect 517244 681216 517296 681222
rect 517244 681158 517296 681164
rect 517256 679946 517284 681158
rect 518990 680504 519046 680513
rect 518990 680439 519046 680448
rect 514772 679918 515016 679946
rect 516948 679918 517284 679946
rect 519004 679810 519032 680439
rect 521856 679946 521884 683878
rect 523052 679946 523080 684830
rect 528742 682408 528798 682417
rect 528742 682343 528798 682352
rect 524970 682136 525026 682145
rect 524970 682071 525026 682080
rect 526258 682136 526314 682145
rect 526258 682071 526314 682080
rect 524420 681080 524472 681086
rect 524420 681022 524472 681028
rect 524432 679946 524460 681022
rect 524984 679946 525012 682071
rect 526272 679946 526300 682071
rect 528756 679946 528784 682343
rect 521856 679918 522100 679946
rect 523052 679918 523388 679946
rect 524432 679918 524676 679946
rect 524984 679918 525320 679946
rect 525964 679918 526300 679946
rect 528540 679918 528784 679946
rect 528848 679946 528876 685918
rect 535460 684752 535512 684758
rect 535460 684694 535512 684700
rect 534078 682816 534134 682825
rect 534078 682751 534134 682760
rect 529664 682644 529716 682650
rect 529664 682586 529716 682592
rect 528848 679918 529184 679946
rect 518880 679782 519032 679810
rect 427084 679652 427136 679658
rect 427084 679594 427136 679600
rect 440148 679652 440200 679658
rect 488612 679646 488764 679674
rect 529676 679674 529704 682586
rect 532700 682576 532752 682582
rect 532700 682518 532752 682524
rect 531226 682272 531282 682281
rect 531226 682207 531282 682216
rect 530124 682032 530176 682038
rect 530124 681974 530176 681980
rect 530136 679946 530164 681974
rect 531240 679946 531268 682207
rect 530136 679918 530472 679946
rect 531116 679918 531268 679946
rect 532712 679946 532740 682518
rect 534092 679946 534120 682751
rect 535274 682544 535330 682553
rect 535274 682479 535330 682488
rect 535288 679946 535316 682479
rect 532712 679918 533048 679946
rect 534092 679918 534336 679946
rect 534980 679918 535316 679946
rect 535472 679946 535500 684694
rect 537852 682032 537904 682038
rect 537852 681974 537904 681980
rect 537864 679946 537892 681974
rect 538232 680218 538260 687890
rect 549996 686520 550048 686526
rect 549996 686462 550048 686468
rect 539140 684616 539192 684622
rect 539140 684558 539192 684564
rect 535472 679918 535624 679946
rect 537556 679918 537892 679946
rect 538186 680190 538260 680218
rect 538186 679932 538214 680190
rect 539152 679946 539180 684558
rect 545580 683596 545632 683602
rect 545580 683538 545632 683544
rect 545120 681964 545172 681970
rect 545120 681906 545172 681912
rect 541716 681760 541768 681766
rect 541716 681702 541768 681708
rect 541728 679946 541756 681702
rect 539152 679918 539488 679946
rect 541420 679918 541756 679946
rect 545132 679946 545160 681906
rect 545592 679946 545620 683538
rect 546958 682952 547014 682961
rect 546958 682887 547014 682896
rect 546866 682000 546922 682009
rect 546866 681935 546922 681944
rect 546880 679946 546908 681935
rect 545132 679918 545284 679946
rect 545592 679918 545928 679946
rect 546572 679918 546908 679946
rect 546972 679946 547000 682887
rect 547788 682100 547840 682106
rect 547788 682042 547840 682048
rect 549904 682100 549956 682106
rect 549904 682042 549956 682048
rect 547800 681086 547828 682042
rect 548800 681964 548852 681970
rect 548800 681906 548852 681912
rect 547788 681080 547840 681086
rect 547788 681022 547840 681028
rect 548812 679946 548840 681906
rect 549442 681864 549498 681873
rect 549442 681799 549498 681808
rect 549456 679946 549484 681799
rect 549916 679946 549944 682042
rect 546972 679918 547216 679946
rect 548504 679918 548840 679946
rect 549148 679918 549484 679946
rect 549792 679918 549944 679946
rect 550008 679810 550036 686462
rect 550178 680368 550234 680377
rect 550178 680303 550234 680312
rect 550008 679782 550128 679810
rect 529676 679646 529828 679674
rect 440148 679594 440200 679600
rect 489734 679552 489790 679561
rect 449820 679522 449972 679538
rect 449808 679516 449972 679522
rect 449860 679510 449972 679516
rect 489790 679510 489900 679538
rect 511152 679522 511488 679538
rect 511152 679516 511500 679522
rect 511152 679510 511448 679516
rect 489734 679487 489790 679496
rect 449808 679458 449860 679464
rect 511448 679458 511500 679464
rect 409880 678292 409932 678298
rect 409880 678234 409932 678240
rect 550100 378865 550128 679782
rect 550192 678745 550220 680303
rect 550178 678736 550234 678745
rect 550178 678671 550234 678680
rect 550180 674144 550232 674150
rect 550180 674086 550232 674092
rect 550192 576026 550220 674086
rect 550180 576020 550232 576026
rect 550180 575962 550232 575968
rect 550180 533384 550232 533390
rect 550180 533326 550232 533332
rect 550086 378856 550142 378865
rect 550086 378791 550142 378800
rect 409786 334656 409842 334665
rect 409786 334591 409842 334600
rect 409786 334520 409842 334529
rect 409786 334455 409842 334464
rect 409800 155854 409828 334455
rect 409878 315616 409934 315625
rect 409878 315551 409934 315560
rect 409892 222902 409920 315551
rect 550192 243982 550220 533326
rect 550284 507385 550312 690610
rect 550364 689308 550416 689314
rect 550364 689250 550416 689256
rect 550376 522345 550404 689250
rect 550640 683664 550692 683670
rect 550640 683606 550692 683612
rect 550456 682712 550508 682718
rect 550456 682654 550508 682660
rect 550468 674150 550496 682654
rect 550456 674144 550508 674150
rect 550456 674086 550508 674092
rect 550652 622985 550680 683606
rect 550732 680944 550784 680950
rect 550732 680886 550784 680892
rect 550638 622976 550694 622985
rect 550638 622911 550694 622920
rect 550456 576020 550508 576026
rect 550456 575962 550508 575968
rect 550468 564505 550496 575962
rect 550454 564496 550510 564505
rect 550454 564431 550510 564440
rect 550454 540016 550510 540025
rect 550454 539951 550510 539960
rect 550468 533390 550496 539951
rect 550456 533384 550508 533390
rect 550456 533326 550508 533332
rect 550362 522336 550418 522345
rect 550362 522271 550418 522280
rect 550270 507376 550326 507385
rect 550270 507311 550326 507320
rect 550638 282296 550694 282305
rect 550638 282231 550694 282240
rect 550270 266656 550326 266665
rect 550270 266591 550326 266600
rect 550180 243976 550232 243982
rect 550180 243918 550232 243924
rect 550178 242856 550234 242865
rect 550178 242791 550234 242800
rect 550086 240816 550142 240825
rect 550086 240751 550142 240760
rect 410156 240644 410208 240650
rect 410156 240586 410208 240592
rect 410248 240644 410300 240650
rect 410248 240586 410300 240592
rect 547328 240644 547380 240650
rect 547328 240586 547380 240592
rect 548708 240644 548760 240650
rect 548708 240586 548760 240592
rect 410030 239850 410058 240108
rect 410030 239822 410104 239850
rect 409972 233708 410024 233714
rect 409972 233650 410024 233656
rect 409880 222896 409932 222902
rect 409880 222838 409932 222844
rect 409984 190058 410012 233650
rect 410076 206310 410104 239822
rect 410064 206304 410116 206310
rect 410064 206246 410116 206252
rect 409972 190052 410024 190058
rect 409972 189994 410024 190000
rect 409788 155848 409840 155854
rect 409788 155790 409840 155796
rect 410168 155038 410196 240586
rect 410260 229094 410288 240586
rect 412272 240576 412324 240582
rect 412272 240518 412324 240524
rect 410800 240508 410852 240514
rect 410800 240450 410852 240456
rect 410352 240094 410688 240122
rect 410352 233714 410380 240094
rect 410340 233708 410392 233714
rect 410340 233650 410392 233656
rect 410812 231810 410840 240450
rect 411318 239850 411346 240108
rect 411318 239822 411392 239850
rect 410800 231804 410852 231810
rect 410800 231746 410852 231752
rect 410260 229066 410564 229094
rect 410156 155032 410208 155038
rect 410156 154974 410208 154980
rect 409696 154352 409748 154358
rect 409696 154294 409748 154300
rect 409050 152688 409106 152697
rect 409050 152623 409106 152632
rect 407304 151020 407356 151026
rect 407304 150962 407356 150968
rect 407224 149926 408434 149954
rect 409064 149940 409092 152623
rect 410340 152312 410392 152318
rect 410340 152254 410392 152260
rect 410352 149940 410380 152254
rect 410536 151337 410564 229066
rect 411364 202162 411392 239822
rect 412284 234297 412312 240518
rect 543996 240242 544332 240258
rect 543996 240236 544344 240242
rect 543996 240230 544292 240236
rect 544292 240178 544344 240184
rect 544752 240236 544804 240242
rect 544752 240178 544804 240184
rect 412620 240094 412864 240122
rect 412270 234288 412326 234297
rect 412270 234223 412326 234232
rect 412640 233708 412692 233714
rect 412640 233650 412692 233656
rect 411628 228948 411680 228954
rect 411628 228890 411680 228896
rect 411352 202156 411404 202162
rect 411352 202098 411404 202104
rect 410522 151328 410578 151337
rect 410522 151263 410578 151272
rect 411640 149940 411668 228890
rect 412652 151230 412680 233650
rect 412836 197130 412864 240094
rect 412928 240094 413264 240122
rect 414032 240094 414552 240122
rect 416484 240094 416728 240122
rect 412928 233714 412956 240094
rect 412916 233708 412968 233714
rect 412916 233650 412968 233656
rect 414032 231606 414060 240094
rect 416700 238134 416728 240094
rect 416976 240094 417128 240122
rect 420012 240094 420348 240122
rect 420992 240094 421328 240122
rect 416688 238128 416740 238134
rect 416688 238070 416740 238076
rect 416700 237998 416728 238070
rect 416688 237992 416740 237998
rect 416688 237934 416740 237940
rect 416780 232348 416832 232354
rect 416780 232290 416832 232296
rect 414020 231600 414072 231606
rect 414020 231542 414072 231548
rect 413560 222964 413612 222970
rect 413560 222906 413612 222912
rect 412824 197124 412876 197130
rect 412824 197066 412876 197072
rect 412824 181552 412876 181558
rect 412824 181494 412876 181500
rect 412640 151224 412692 151230
rect 412640 151166 412692 151172
rect 412836 149954 412864 181494
rect 412836 149926 412942 149954
rect 413572 149940 413600 222906
rect 414664 202904 414716 202910
rect 414664 202846 414716 202852
rect 414676 162858 414704 202846
rect 414664 162852 414716 162858
rect 414664 162794 414716 162800
rect 414848 153128 414900 153134
rect 414848 153070 414900 153076
rect 414860 149940 414888 153070
rect 416792 149940 416820 232290
rect 416976 211818 417004 240094
rect 417424 236700 417476 236706
rect 417424 236642 417476 236648
rect 416964 211812 417016 211818
rect 416964 211754 417016 211760
rect 417436 149940 417464 236642
rect 419356 236632 419408 236638
rect 419356 236574 419408 236580
rect 418804 233708 418856 233714
rect 418804 233650 418856 233656
rect 418068 227248 418120 227254
rect 418068 227190 418120 227196
rect 418080 149940 418108 227190
rect 418816 204270 418844 233650
rect 418804 204264 418856 204270
rect 418804 204206 418856 204212
rect 419368 149940 419396 236574
rect 420012 233714 420040 240094
rect 421300 238134 421328 240094
rect 422910 239850 422938 240108
rect 422864 239822 422938 239850
rect 423048 240094 423568 240122
rect 426452 240094 426788 240122
rect 426912 240094 427432 240122
rect 427832 240094 428076 240122
rect 428384 240094 428720 240122
rect 431940 240094 432092 240122
rect 421288 238128 421340 238134
rect 421288 238070 421340 238076
rect 422864 237930 422892 239822
rect 422852 237924 422904 237930
rect 422852 237866 422904 237872
rect 420000 233708 420052 233714
rect 420000 233650 420052 233656
rect 423048 219434 423076 240094
rect 422312 219406 423076 219434
rect 422312 197198 422340 219406
rect 422300 197192 422352 197198
rect 422300 197134 422352 197140
rect 420000 162852 420052 162858
rect 420000 162794 420052 162800
rect 420012 149940 420040 162794
rect 426452 160682 426480 240094
rect 426912 219434 426940 240094
rect 427832 238746 427860 240094
rect 427820 238740 427872 238746
rect 427820 238682 427872 238688
rect 428384 238610 428412 240094
rect 428372 238604 428424 238610
rect 428372 238546 428424 238552
rect 430304 236632 430356 236638
rect 430304 236574 430356 236580
rect 429200 224324 429252 224330
rect 429200 224266 429252 224272
rect 426544 219406 426940 219434
rect 426544 181490 426572 219406
rect 427082 188592 427138 188601
rect 427082 188527 427138 188536
rect 426532 181484 426584 181490
rect 426532 181426 426584 181432
rect 426440 160676 426492 160682
rect 426440 160618 426492 160624
rect 421932 152924 421984 152930
rect 421932 152866 421984 152872
rect 421944 149940 421972 152866
rect 425152 152448 425204 152454
rect 425152 152390 425204 152396
rect 425164 149940 425192 152390
rect 427096 149940 427124 188527
rect 429212 149954 429240 224266
rect 429212 149926 429686 149954
rect 430316 149940 430344 236574
rect 432064 178838 432092 240094
rect 432248 240094 432584 240122
rect 433352 240094 434516 240122
rect 436448 240094 436784 240122
rect 432248 238202 432276 240094
rect 432236 238196 432288 238202
rect 432236 238138 432288 238144
rect 433352 214606 433380 240094
rect 436756 238610 436784 240094
rect 438872 240094 439024 240122
rect 436744 238604 436796 238610
rect 436744 238546 436796 238552
rect 436744 224324 436796 224330
rect 436744 224266 436796 224272
rect 435456 220176 435508 220182
rect 435456 220118 435508 220124
rect 433340 214600 433392 214606
rect 433340 214542 433392 214548
rect 432052 178832 432104 178838
rect 432052 178774 432104 178780
rect 434168 152380 434220 152386
rect 434168 152322 434220 152328
rect 434180 149940 434208 152322
rect 435468 149940 435496 220118
rect 436756 149940 436784 224266
rect 438676 212016 438728 212022
rect 438676 211958 438728 211964
rect 438688 149940 438716 211958
rect 438872 185774 438900 240094
rect 440298 239850 440326 240108
rect 440252 239822 440326 239850
rect 442552 240094 442888 240122
rect 443656 240094 444176 240122
rect 444820 240094 445156 240122
rect 446752 240094 447088 240122
rect 440252 238678 440280 239822
rect 440240 238672 440292 238678
rect 440240 238614 440292 238620
rect 442552 238270 442580 240094
rect 442540 238264 442592 238270
rect 442540 238206 442592 238212
rect 443656 219434 443684 240094
rect 445128 238678 445156 240094
rect 447060 238882 447088 240094
rect 449912 240094 450616 240122
rect 451384 240094 451904 240122
rect 447048 238876 447100 238882
rect 447048 238818 447100 238824
rect 445116 238672 445168 238678
rect 445116 238614 445168 238620
rect 448336 229968 448388 229974
rect 448336 229910 448388 229916
rect 444472 224460 444524 224466
rect 444472 224402 444524 224408
rect 443012 219406 443684 219434
rect 441620 211948 441672 211954
rect 441620 211890 441672 211896
rect 438860 185768 438912 185774
rect 438860 185710 438912 185716
rect 439320 158704 439372 158710
rect 439320 158646 439372 158652
rect 439332 149940 439360 158646
rect 440606 156904 440662 156913
rect 440606 156839 440662 156848
rect 440620 149940 440648 156839
rect 441632 149954 441660 211890
rect 443012 204950 443040 219406
rect 443000 204944 443052 204950
rect 443000 204886 443052 204892
rect 443184 176044 443236 176050
rect 443184 175986 443236 175992
rect 441632 149926 441922 149954
rect 443196 149940 443224 175986
rect 444484 149940 444512 224402
rect 445760 217320 445812 217326
rect 445760 217262 445812 217268
rect 445772 149954 445800 217262
rect 447692 152992 447744 152998
rect 447692 152934 447744 152940
rect 445772 149926 446430 149954
rect 447704 149940 447732 152934
rect 448348 149940 448376 229910
rect 449912 194274 449940 240094
rect 451384 219434 451412 240094
rect 452534 239850 452562 240108
rect 452672 240094 453192 240122
rect 454144 240094 454480 240122
rect 454604 240094 455124 240122
rect 456412 240094 456748 240122
rect 457056 240094 457392 240122
rect 452534 239822 452608 239850
rect 452580 235686 452608 239822
rect 452568 235680 452620 235686
rect 452568 235622 452620 235628
rect 452672 231062 452700 240094
rect 454144 236570 454172 240094
rect 454132 236564 454184 236570
rect 454132 236506 454184 236512
rect 452660 231056 452712 231062
rect 452660 230998 452712 231004
rect 454604 219434 454632 240094
rect 456720 235550 456748 240094
rect 457364 238785 457392 240094
rect 458192 240094 458344 240122
rect 457350 238776 457406 238785
rect 457350 238711 457406 238720
rect 458192 238377 458220 240094
rect 459618 239850 459646 240108
rect 460906 239850 460934 240108
rect 461044 240094 461564 240122
rect 462424 240094 462852 240122
rect 463160 240094 463496 240122
rect 463712 240094 464140 240122
rect 465092 240094 465428 240122
rect 467852 240094 468004 240122
rect 468128 240094 468648 240122
rect 459618 239822 459692 239850
rect 460906 239822 460980 239850
rect 458178 238368 458234 238377
rect 458178 238303 458234 238312
rect 456708 235544 456760 235550
rect 456708 235486 456760 235492
rect 451292 219406 451412 219434
rect 454144 219406 454632 219434
rect 449900 194268 449952 194274
rect 449900 194210 449952 194216
rect 448980 153060 449032 153066
rect 448980 153002 449032 153008
rect 448992 149940 449020 153002
rect 451292 152930 451320 219406
rect 452844 195288 452896 195294
rect 452844 195230 452896 195236
rect 451280 152924 451332 152930
rect 451280 152866 451332 152872
rect 452856 149940 452884 195230
rect 453486 192672 453542 192681
rect 453486 192607 453542 192616
rect 453500 149940 453528 192607
rect 454144 159526 454172 219406
rect 459664 183054 459692 239822
rect 460952 235754 460980 239822
rect 460940 235748 460992 235754
rect 460940 235690 460992 235696
rect 459928 224392 459980 224398
rect 459928 224334 459980 224340
rect 459652 183048 459704 183054
rect 459652 182990 459704 182996
rect 458178 180160 458234 180169
rect 458178 180095 458234 180104
rect 454132 159520 454184 159526
rect 454132 159462 454184 159468
rect 458192 149954 458220 180095
rect 458192 149926 458666 149954
rect 459940 149940 459968 224334
rect 461044 219434 461072 240094
rect 461216 235884 461268 235890
rect 461216 235826 461268 235832
rect 460952 219406 461072 219434
rect 460952 178770 460980 219406
rect 460940 178764 460992 178770
rect 460940 178706 460992 178712
rect 460572 163532 460624 163538
rect 460572 163474 460624 163480
rect 460584 149940 460612 163474
rect 461228 149940 461256 235826
rect 462424 152998 462452 240094
rect 463160 238338 463188 240094
rect 463148 238332 463200 238338
rect 463148 238274 463200 238280
rect 463712 196382 463740 240094
rect 463700 196376 463752 196382
rect 463700 196318 463752 196324
rect 465092 195906 465120 240094
rect 465080 195900 465132 195906
rect 465080 195842 465132 195848
rect 467852 175030 467880 240094
rect 468128 219434 468156 240094
rect 469278 239850 469306 240108
rect 470566 239850 470594 240108
rect 470704 240094 471224 240122
rect 472512 240094 472664 240122
rect 469278 239822 469352 239850
rect 470566 239822 470640 239850
rect 467944 219406 468156 219434
rect 467944 198762 467972 219406
rect 467932 198756 467984 198762
rect 467932 198698 467984 198704
rect 469324 177818 469352 239822
rect 470612 238377 470640 239822
rect 470598 238368 470654 238377
rect 470598 238303 470654 238312
rect 470232 232416 470284 232422
rect 470232 232358 470284 232364
rect 469312 177812 469364 177818
rect 469312 177754 469364 177760
rect 467840 175024 467892 175030
rect 467840 174966 467892 174972
rect 468300 172032 468352 172038
rect 468300 171974 468352 171980
rect 463790 153096 463846 153105
rect 463790 153031 463846 153040
rect 462412 152992 462464 152998
rect 462412 152934 462464 152940
rect 463804 149940 463832 153031
rect 468312 149940 468340 171974
rect 470244 149940 470272 232358
rect 470704 219434 470732 240094
rect 472636 238338 472664 240094
rect 472728 240094 473156 240122
rect 474444 240094 474688 240122
rect 475088 240094 475424 240122
rect 472624 238332 472676 238338
rect 472624 238274 472676 238280
rect 471980 232484 472032 232490
rect 471980 232426 472032 232432
rect 470612 219406 470732 219434
rect 470612 166394 470640 219406
rect 470600 166388 470652 166394
rect 470600 166330 470652 166336
rect 471992 149954 472020 232426
rect 472728 219434 472756 240094
rect 474660 235822 474688 240094
rect 475396 238202 475424 240094
rect 476362 239850 476390 240108
rect 476500 240094 477020 240122
rect 476362 239822 476436 239850
rect 476408 238270 476436 239822
rect 476396 238264 476448 238270
rect 476396 238206 476448 238212
rect 475384 238196 475436 238202
rect 475384 238138 475436 238144
rect 474648 235816 474700 235822
rect 474648 235758 474700 235764
rect 472808 222896 472860 222902
rect 472808 222838 472860 222844
rect 472176 219406 472756 219434
rect 472176 191146 472204 219406
rect 472164 191140 472216 191146
rect 472164 191082 472216 191088
rect 471992 149926 472190 149954
rect 472820 149940 472848 222838
rect 476500 219434 476528 240094
rect 477650 239850 477678 240108
rect 478938 239850 478966 240108
rect 476224 219406 476528 219434
rect 477604 239822 477678 239850
rect 478892 239822 478966 239850
rect 480226 239850 480254 240108
rect 481514 239850 481542 240108
rect 483124 240094 483460 240122
rect 483768 240094 484104 240122
rect 484872 240094 485392 240122
rect 487448 240094 487968 240122
rect 480226 239822 480300 239850
rect 481514 239822 481588 239850
rect 476028 202156 476080 202162
rect 476028 202098 476080 202104
rect 476040 149940 476068 202098
rect 476224 194585 476252 219406
rect 476672 218748 476724 218754
rect 476672 218690 476724 218696
rect 476210 194576 476266 194585
rect 476210 194511 476266 194520
rect 476684 149940 476712 218690
rect 477604 212022 477632 239822
rect 478604 236564 478656 236570
rect 478604 236506 478656 236512
rect 477960 221468 478012 221474
rect 477960 221410 478012 221416
rect 477592 212016 477644 212022
rect 477592 211958 477644 211964
rect 477972 149940 478000 221410
rect 478616 149940 478644 236506
rect 478892 193186 478920 239822
rect 478880 193180 478932 193186
rect 478880 193122 478932 193128
rect 480272 159594 480300 239822
rect 481560 235958 481588 239822
rect 482928 237924 482980 237930
rect 482928 237866 482980 237872
rect 482940 237454 482968 237866
rect 482928 237448 482980 237454
rect 482928 237390 482980 237396
rect 481548 235952 481600 235958
rect 481548 235894 481600 235900
rect 481180 225616 481232 225622
rect 481180 225558 481232 225564
rect 480536 173188 480588 173194
rect 480536 173130 480588 173136
rect 480260 159588 480312 159594
rect 480260 159530 480312 159536
rect 480548 149940 480576 173130
rect 481192 149940 481220 225558
rect 481824 158160 481876 158166
rect 481824 158102 481876 158108
rect 481836 149940 481864 158102
rect 482940 153134 482968 237390
rect 483124 174690 483152 240094
rect 483768 237454 483796 240094
rect 483756 237448 483808 237454
rect 483756 237390 483808 237396
rect 484872 219434 484900 240094
rect 486976 233708 487028 233714
rect 486976 233650 487028 233656
rect 484412 219406 484900 219434
rect 483112 174684 483164 174690
rect 483112 174626 483164 174632
rect 484412 169590 484440 219406
rect 485044 213308 485096 213314
rect 485044 213250 485096 213256
rect 484400 169584 484452 169590
rect 484400 169526 484452 169532
rect 482928 153128 482980 153134
rect 482928 153070 482980 153076
rect 482466 152960 482522 152969
rect 482466 152895 482522 152904
rect 482480 149940 482508 152895
rect 485056 149940 485084 213250
rect 486988 149940 487016 233650
rect 487448 219434 487476 240094
rect 488598 239850 488626 240108
rect 487172 219406 487476 219434
rect 488552 239822 488626 239850
rect 488736 240094 489256 240122
rect 487172 197742 487200 219406
rect 487160 197736 487212 197742
rect 487160 197678 487212 197684
rect 488552 149938 488580 239822
rect 488736 219434 488764 240094
rect 490530 239850 490558 240108
rect 491174 239850 491202 240108
rect 492048 240094 492476 240122
rect 496832 240094 496984 240122
rect 497628 240094 497964 240122
rect 490530 239822 490604 239850
rect 491174 239822 491248 239850
rect 490576 237998 490604 239822
rect 490564 237992 490616 237998
rect 490564 237934 490616 237940
rect 491116 237992 491168 237998
rect 491116 237934 491168 237940
rect 491128 235142 491156 237934
rect 491116 235136 491168 235142
rect 491116 235078 491168 235084
rect 491220 235074 491248 239822
rect 491300 235204 491352 235210
rect 491300 235146 491352 235152
rect 491208 235068 491260 235074
rect 491208 235010 491260 235016
rect 488644 219406 488764 219434
rect 488644 178702 488672 219406
rect 490196 186992 490248 186998
rect 490196 186934 490248 186940
rect 488632 178696 488684 178702
rect 488632 178638 488684 178644
rect 488906 169008 488962 169017
rect 488906 168943 488962 168952
rect 488920 149940 488948 168943
rect 490208 149940 490236 186934
rect 491312 149954 491340 235146
rect 492048 219434 492076 240094
rect 496832 233714 496860 240094
rect 497936 238406 497964 240094
rect 498212 240094 498916 240122
rect 500328 240094 500848 240122
rect 501492 240094 501828 240122
rect 497924 238400 497976 238406
rect 497924 238342 497976 238348
rect 496820 233708 496872 233714
rect 496820 233650 496872 233656
rect 493416 232484 493468 232490
rect 493416 232426 493468 232432
rect 491404 219406 492076 219434
rect 491404 198422 491432 219406
rect 491392 198416 491444 198422
rect 491392 198358 491444 198364
rect 492770 185600 492826 185609
rect 492770 185535 492826 185544
rect 488540 149932 488592 149938
rect 387432 149874 387484 149880
rect 491312 149926 492154 149954
rect 492784 149940 492812 185535
rect 493428 149940 493456 232426
rect 497924 229832 497976 229838
rect 497924 229774 497976 229780
rect 494060 220108 494112 220114
rect 494060 220050 494112 220056
rect 494072 149940 494100 220050
rect 495438 195392 495494 195401
rect 495438 195327 495494 195336
rect 495452 149954 495480 195327
rect 497278 184240 497334 184249
rect 497278 184175 497334 184184
rect 495452 149926 496662 149954
rect 497292 149940 497320 184175
rect 497936 149940 497964 229774
rect 498212 152454 498240 240094
rect 500328 239442 500356 240094
rect 499684 239414 500356 239442
rect 499212 236496 499264 236502
rect 499212 236438 499264 236444
rect 498566 152824 498622 152833
rect 498566 152759 498622 152768
rect 498200 152448 498252 152454
rect 498200 152390 498252 152396
rect 498580 149940 498608 152759
rect 499224 149940 499252 236438
rect 499684 153066 499712 239414
rect 499856 238944 499908 238950
rect 499856 238886 499908 238892
rect 499672 153060 499724 153066
rect 499672 153002 499724 153008
rect 499868 149940 499896 238886
rect 501800 237998 501828 240094
rect 504376 240094 504712 240122
rect 505356 240094 505692 240122
rect 504376 238542 504404 240094
rect 505664 238950 505692 240094
rect 506630 239850 506658 240108
rect 506768 240094 507288 240122
rect 506630 239822 506704 239850
rect 505652 238944 505704 238950
rect 505652 238886 505704 238892
rect 506676 238542 506704 239822
rect 504364 238536 504416 238542
rect 504364 238478 504416 238484
rect 506664 238536 506716 238542
rect 506664 238478 506716 238484
rect 501788 237992 501840 237998
rect 501788 237934 501840 237940
rect 503720 229900 503772 229906
rect 503720 229842 503772 229848
rect 502430 167784 502486 167793
rect 502430 167719 502486 167728
rect 502444 149940 502472 167719
rect 503076 152380 503128 152386
rect 503076 152322 503128 152328
rect 503088 149940 503116 152322
rect 503732 149940 503760 229842
rect 506768 219434 506796 240094
rect 507918 239850 507946 240108
rect 509206 239850 509234 240108
rect 509344 240094 509864 240122
rect 514772 240094 515016 240122
rect 515324 240094 515660 240122
rect 507918 239822 507992 239850
rect 509206 239822 509280 239850
rect 506584 219406 506796 219434
rect 506584 192506 506612 219406
rect 507584 206304 507636 206310
rect 507584 206246 507636 206252
rect 506572 192500 506624 192506
rect 506572 192442 506624 192448
rect 506296 173324 506348 173330
rect 506296 173266 506348 173272
rect 505652 152312 505704 152318
rect 505652 152254 505704 152260
rect 505664 149940 505692 152254
rect 506308 149940 506336 173266
rect 506940 165096 506992 165102
rect 506940 165038 506992 165044
rect 506952 149940 506980 165038
rect 507596 149940 507624 206246
rect 507964 200802 507992 239822
rect 509252 238814 509280 239822
rect 509240 238808 509292 238814
rect 509240 238750 509292 238756
rect 509344 228954 509372 240094
rect 514772 238474 514800 240094
rect 514760 238468 514812 238474
rect 514760 238410 514812 238416
rect 515324 237862 515352 240094
rect 518866 239850 518894 240108
rect 519096 240094 519524 240122
rect 518866 239822 518940 239850
rect 515312 237856 515364 237862
rect 515312 237798 515364 237804
rect 511448 235612 511500 235618
rect 511448 235554 511500 235560
rect 509332 228948 509384 228954
rect 509332 228890 509384 228896
rect 508504 212560 508556 212566
rect 508504 212502 508556 212508
rect 508228 204944 508280 204950
rect 508228 204886 508280 204892
rect 507952 200796 508004 200802
rect 507952 200738 508004 200744
rect 508240 149940 508268 204886
rect 508516 166394 508544 212502
rect 508504 166388 508556 166394
rect 508504 166330 508556 166336
rect 510160 163464 510212 163470
rect 510160 163406 510212 163412
rect 510172 149940 510200 163406
rect 511460 149940 511488 235554
rect 518164 229900 518216 229906
rect 518164 229842 518216 229848
rect 512092 227180 512144 227186
rect 512092 227122 512144 227128
rect 512104 149940 512132 227122
rect 514024 166388 514076 166394
rect 514024 166330 514076 166336
rect 514036 149940 514064 166330
rect 518176 152318 518204 229842
rect 518164 152312 518216 152318
rect 518164 152254 518216 152260
rect 518912 151230 518940 239822
rect 519096 195974 519124 240094
rect 520154 239850 520182 240108
rect 524032 240094 524368 240122
rect 525320 240094 525656 240122
rect 527896 240094 528232 240122
rect 528540 240094 528784 240122
rect 520154 239822 520228 239850
rect 520200 238105 520228 239822
rect 524340 238241 524368 240094
rect 524326 238232 524382 238241
rect 524326 238167 524382 238176
rect 520186 238096 520242 238105
rect 520186 238031 520242 238040
rect 525628 232422 525656 240094
rect 528204 237930 528232 240094
rect 528756 237969 528784 240094
rect 528848 240094 529184 240122
rect 528848 238513 528876 240094
rect 529814 239850 529842 240108
rect 529952 240094 531116 240122
rect 531976 240094 532404 240122
rect 532712 240094 533048 240122
rect 534980 240094 535316 240122
rect 529814 239822 529888 239850
rect 528834 238504 528890 238513
rect 528834 238439 528890 238448
rect 528742 237960 528798 237969
rect 528192 237924 528244 237930
rect 528742 237895 528798 237904
rect 528192 237866 528244 237872
rect 529860 237862 529888 239822
rect 529848 237856 529900 237862
rect 529848 237798 529900 237804
rect 525616 232416 525668 232422
rect 525616 232358 525668 232364
rect 527548 227112 527600 227118
rect 527548 227054 527600 227060
rect 525800 227044 525852 227050
rect 525800 226986 525852 226992
rect 521660 224256 521712 224262
rect 521660 224198 521712 224204
rect 519176 203652 519228 203658
rect 519176 203594 519228 203600
rect 519084 195968 519136 195974
rect 519084 195910 519136 195916
rect 518900 151224 518952 151230
rect 518900 151166 518952 151172
rect 519188 149940 519216 203594
rect 519820 153944 519872 153950
rect 519820 153886 519872 153892
rect 519832 149940 519860 153886
rect 521672 149954 521700 224198
rect 524972 211880 525024 211886
rect 524972 211822 525024 211828
rect 523038 206272 523094 206281
rect 523038 206207 523094 206216
rect 521672 149926 521778 149954
rect 523052 149940 523080 206207
rect 523592 150068 523644 150074
rect 523592 150010 523644 150016
rect 523604 149938 523632 150010
rect 524984 149940 525012 211822
rect 525812 149954 525840 226986
rect 526444 175976 526496 175982
rect 526444 175918 526496 175924
rect 526456 151978 526484 175918
rect 526444 151972 526496 151978
rect 526444 151914 526496 151920
rect 523592 149932 523644 149938
rect 488540 149874 488592 149880
rect 525812 149926 526286 149954
rect 527560 149940 527588 227054
rect 529952 194342 529980 240094
rect 531976 219434 532004 240094
rect 532056 239352 532108 239358
rect 532056 239294 532108 239300
rect 531332 219406 532004 219434
rect 531332 195945 531360 219406
rect 531318 195936 531374 195945
rect 531318 195871 531374 195880
rect 529940 194336 529992 194342
rect 529940 194278 529992 194284
rect 529940 182912 529992 182918
rect 529940 182854 529992 182860
rect 529204 152856 529256 152862
rect 529204 152798 529256 152804
rect 529216 152318 529244 152798
rect 529204 152312 529256 152318
rect 529204 152254 529256 152260
rect 528836 151972 528888 151978
rect 528836 151914 528888 151920
rect 528848 149940 528876 151914
rect 529952 149954 529980 182854
rect 531412 152856 531464 152862
rect 531412 152798 531464 152804
rect 529952 149926 530150 149954
rect 531424 149940 531452 152798
rect 532068 149940 532096 239294
rect 532712 236774 532740 240094
rect 535288 238474 535316 240094
rect 536898 239850 536926 240108
rect 536852 239822 536926 239850
rect 542372 240094 543352 240122
rect 544212 240094 544640 240122
rect 535276 238468 535328 238474
rect 535276 238410 535328 238416
rect 532700 236768 532752 236774
rect 532700 236710 532752 236716
rect 536852 230994 536880 239822
rect 538862 239592 538918 239601
rect 538862 239527 538918 239536
rect 534724 230988 534776 230994
rect 534724 230930 534776 230936
rect 536840 230988 536892 230994
rect 536840 230930 536892 230936
rect 534736 152862 534764 230930
rect 535920 215960 535972 215966
rect 535920 215902 535972 215908
rect 534724 152856 534776 152862
rect 534724 152798 534776 152804
rect 534632 152312 534684 152318
rect 534632 152254 534684 152260
rect 534644 149940 534672 152254
rect 535932 149940 535960 215902
rect 536102 195256 536158 195265
rect 536102 195191 536158 195200
rect 536116 152862 536144 195191
rect 537484 157956 537536 157962
rect 537484 157898 537536 157904
rect 537116 155916 537168 155922
rect 537116 155858 537168 155864
rect 536104 152856 536156 152862
rect 536104 152798 536156 152804
rect 537128 150890 537156 155858
rect 537392 150952 537444 150958
rect 537392 150894 537444 150900
rect 537116 150884 537168 150890
rect 537116 150826 537168 150832
rect 537404 150006 537432 150894
rect 537496 150346 537524 157898
rect 537576 157820 537628 157826
rect 537576 157762 537628 157768
rect 537588 151745 537616 157762
rect 538876 152386 538904 239527
rect 540428 238060 540480 238066
rect 540428 238002 540480 238008
rect 540336 234388 540388 234394
rect 540336 234330 540388 234336
rect 540060 233164 540112 233170
rect 540060 233106 540112 233112
rect 538956 231804 539008 231810
rect 538956 231746 539008 231752
rect 538968 155922 538996 231746
rect 539048 208412 539100 208418
rect 539048 208354 539100 208360
rect 538956 155916 539008 155922
rect 538956 155858 539008 155864
rect 538956 155032 539008 155038
rect 538956 154974 539008 154980
rect 538864 152380 538916 152386
rect 538864 152322 538916 152328
rect 537574 151736 537630 151745
rect 537574 151671 537630 151680
rect 538864 150408 538916 150414
rect 538770 150376 538826 150385
rect 537484 150340 537536 150346
rect 538864 150350 538916 150356
rect 538770 150311 538826 150320
rect 537484 150282 537536 150288
rect 537392 150000 537444 150006
rect 537392 149942 537444 149948
rect 538784 149938 538812 150311
rect 538876 150249 538904 150350
rect 538862 150240 538918 150249
rect 538968 150210 538996 154974
rect 539060 150482 539088 208354
rect 539232 166456 539284 166462
rect 539232 166398 539284 166404
rect 539048 150476 539100 150482
rect 539048 150418 539100 150424
rect 538862 150175 538918 150184
rect 538956 150204 539008 150210
rect 538956 150146 539008 150152
rect 539046 149968 539102 149977
rect 538772 149932 538824 149938
rect 523592 149874 523644 149880
rect 539244 149954 539272 166398
rect 539968 159384 540020 159390
rect 539968 159326 540020 159332
rect 539324 158568 539376 158574
rect 539324 158510 539376 158516
rect 539336 150090 539364 158510
rect 539416 158228 539468 158234
rect 539416 158170 539468 158176
rect 539428 150278 539456 158170
rect 539508 155916 539560 155922
rect 539508 155858 539560 155864
rect 539520 150414 539548 155858
rect 539600 154420 539652 154426
rect 539600 154362 539652 154368
rect 539508 150408 539560 150414
rect 539508 150350 539560 150356
rect 539416 150272 539468 150278
rect 539416 150214 539468 150220
rect 539612 150142 539640 154362
rect 539784 152856 539836 152862
rect 539784 152798 539836 152804
rect 539600 150136 539652 150142
rect 539336 150062 539456 150090
rect 539600 150078 539652 150084
rect 539322 149968 539378 149977
rect 539244 149926 539322 149954
rect 539046 149903 539048 149912
rect 538772 149874 538824 149880
rect 539100 149903 539102 149912
rect 539428 149938 539456 150062
rect 539796 149940 539824 152798
rect 539876 150408 539928 150414
rect 539876 150350 539928 150356
rect 539888 150249 539916 150350
rect 539874 150240 539930 150249
rect 539874 150175 539930 150184
rect 539322 149903 539378 149912
rect 539416 149932 539468 149938
rect 539048 149874 539100 149880
rect 539416 149874 539468 149880
rect 60016 29889 60044 30124
rect 60002 29880 60058 29889
rect 60002 29815 60058 29824
rect 60738 29744 60794 29753
rect 60738 29679 60794 29688
rect 59912 17604 59964 17610
rect 59912 17546 59964 17552
rect 59820 17468 59872 17474
rect 59820 17410 59872 17416
rect 60752 16574 60780 29679
rect 61304 29617 61332 30124
rect 61290 29608 61346 29617
rect 61290 29543 61346 29552
rect 62592 28762 62620 30124
rect 63236 28830 63264 30124
rect 63500 29708 63552 29714
rect 63500 29650 63552 29656
rect 63224 28824 63276 28830
rect 63224 28766 63276 28772
rect 62580 28756 62632 28762
rect 62580 28698 62632 28704
rect 63512 28082 63540 29650
rect 63500 28076 63552 28082
rect 63500 28018 63552 28024
rect 65168 26234 65196 30124
rect 65812 28257 65840 30124
rect 65798 28248 65854 28257
rect 65798 28183 65854 28192
rect 66352 28144 66404 28150
rect 66352 28086 66404 28092
rect 64892 26206 65196 26234
rect 64892 23361 64920 26206
rect 64878 23352 64934 23361
rect 64878 23287 64934 23296
rect 66364 22642 66392 28086
rect 66456 27577 66484 30124
rect 67744 28898 67772 30124
rect 69048 29866 69076 30124
rect 69032 29838 69076 29866
rect 69032 29646 69060 29838
rect 69020 29640 69072 29646
rect 69020 29582 69072 29588
rect 69676 29510 69704 30124
rect 69664 29504 69716 29510
rect 69664 29446 69716 29452
rect 67732 28892 67784 28898
rect 67732 28834 67784 28840
rect 69940 28280 69992 28286
rect 69940 28222 69992 28228
rect 66442 27568 66498 27577
rect 66442 27503 66498 27512
rect 69662 27432 69718 27441
rect 69662 27367 69718 27376
rect 69676 26722 69704 27367
rect 69664 26716 69716 26722
rect 69664 26658 69716 26664
rect 67640 25492 67692 25498
rect 67640 25434 67692 25440
rect 66352 22636 66404 22642
rect 66352 22578 66404 22584
rect 60752 16546 60872 16574
rect 58808 16448 58860 16454
rect 58808 16390 58860 16396
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 53012 3392 53064 3398
rect 53012 3334 53064 3340
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 52932 462 53328 490
rect 57256 480 57284 3402
rect 60844 480 60872 16546
rect 64326 4856 64382 4865
rect 64326 4791 64382 4800
rect 64340 480 64368 4791
rect 53300 354 53328 462
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 25434
rect 69952 20670 69980 28222
rect 70320 27538 70348 30124
rect 70964 27606 70992 30124
rect 71608 28490 71636 30124
rect 72912 29866 72940 30124
rect 72896 29838 72940 29866
rect 71596 28484 71648 28490
rect 71596 28426 71648 28432
rect 72424 28484 72476 28490
rect 72424 28426 72476 28432
rect 72330 28248 72386 28257
rect 72330 28183 72386 28192
rect 70952 27600 71004 27606
rect 70952 27542 71004 27548
rect 70308 27532 70360 27538
rect 70308 27474 70360 27480
rect 70398 25392 70454 25401
rect 70398 25327 70454 25336
rect 69940 20664 69992 20670
rect 69940 20606 69992 20612
rect 70412 16574 70440 25327
rect 72344 22846 72372 28183
rect 72332 22840 72384 22846
rect 72332 22782 72384 22788
rect 72436 22574 72464 28426
rect 72896 28218 72924 29838
rect 73540 28558 73568 30124
rect 78048 28937 78076 30124
rect 78034 28928 78090 28937
rect 78034 28863 78090 28872
rect 82556 28694 82584 30124
rect 82544 28688 82596 28694
rect 82544 28630 82596 28636
rect 83464 28688 83516 28694
rect 83464 28630 83516 28636
rect 73528 28552 73580 28558
rect 73528 28494 73580 28500
rect 78772 28552 78824 28558
rect 78772 28494 78824 28500
rect 72884 28212 72936 28218
rect 72884 28154 72936 28160
rect 74540 28212 74592 28218
rect 74540 28154 74592 28160
rect 74552 24449 74580 28154
rect 77300 25628 77352 25634
rect 77300 25570 77352 25576
rect 74538 24440 74594 24449
rect 74538 24375 74594 24384
rect 72424 22568 72476 22574
rect 72424 22510 72476 22516
rect 77312 16574 77340 25570
rect 78784 22098 78812 28494
rect 81440 25560 81492 25566
rect 81440 25502 81492 25508
rect 78772 22092 78824 22098
rect 78772 22034 78824 22040
rect 81452 16574 81480 25502
rect 83476 18426 83504 28630
rect 84488 26234 84516 30124
rect 85792 29866 85820 30124
rect 85776 29838 85820 29866
rect 85776 29481 85804 29838
rect 85762 29472 85818 29481
rect 85762 29407 85818 29416
rect 87708 26858 87736 30124
rect 89656 29866 89684 30124
rect 89640 29838 89684 29866
rect 89640 27470 89668 29838
rect 91572 28393 91600 30124
rect 92216 28422 92244 30124
rect 92204 28416 92256 28422
rect 91558 28384 91614 28393
rect 92204 28358 92256 28364
rect 92478 28384 92534 28393
rect 91558 28319 91614 28328
rect 95436 28354 95464 30124
rect 92478 28319 92534 28328
rect 95424 28348 95476 28354
rect 89628 27464 89680 27470
rect 89628 27406 89680 27412
rect 92492 26926 92520 28319
rect 95424 28290 95476 28296
rect 96080 28257 96108 30124
rect 96804 28416 96856 28422
rect 96804 28358 96856 28364
rect 96066 28248 96122 28257
rect 96066 28183 96122 28192
rect 92572 27940 92624 27946
rect 92572 27882 92624 27888
rect 92480 26920 92532 26926
rect 92480 26862 92532 26868
rect 87696 26852 87748 26858
rect 87696 26794 87748 26800
rect 84212 26206 84516 26234
rect 83464 18420 83516 18426
rect 83464 18362 83516 18368
rect 84212 16969 84240 26206
rect 88338 25528 88394 25537
rect 88338 25463 88394 25472
rect 85580 24880 85632 24886
rect 85580 24822 85632 24828
rect 84198 16960 84254 16969
rect 84198 16895 84254 16904
rect 85592 16574 85620 24822
rect 88352 16574 88380 25463
rect 92584 21350 92612 27882
rect 92572 21344 92624 21350
rect 92572 21286 92624 21292
rect 96816 21282 96844 28358
rect 97354 28248 97410 28257
rect 97354 28183 97410 28192
rect 97368 21729 97396 28183
rect 98000 28076 98052 28082
rect 98000 28018 98052 28024
rect 97354 21720 97410 21729
rect 97354 21655 97410 21664
rect 96804 21276 96856 21282
rect 96804 21218 96856 21224
rect 98012 17950 98040 28018
rect 98656 26234 98684 30124
rect 99300 28082 99328 30124
rect 100588 28082 100616 30124
rect 99288 28076 99340 28082
rect 99288 28018 99340 28024
rect 99380 28076 99432 28082
rect 99380 28018 99432 28024
rect 100576 28076 100628 28082
rect 100576 28018 100628 28024
rect 98104 26206 98684 26234
rect 98104 23934 98132 26206
rect 99392 24002 99420 28018
rect 101232 26234 101260 30124
rect 103164 28014 103192 30124
rect 103808 28626 103836 30124
rect 103796 28620 103848 28626
rect 103796 28562 103848 28568
rect 103152 28008 103204 28014
rect 103152 27950 103204 27956
rect 104164 28008 104216 28014
rect 104164 27950 104216 27956
rect 103520 27668 103572 27674
rect 103520 27610 103572 27616
rect 100772 26206 101260 26234
rect 100772 24585 100800 26206
rect 100758 24576 100814 24585
rect 100758 24511 100814 24520
rect 99380 23996 99432 24002
rect 99380 23938 99432 23944
rect 98092 23928 98144 23934
rect 98092 23870 98144 23876
rect 103532 21418 103560 27610
rect 103520 21412 103572 21418
rect 103520 21354 103572 21360
rect 104176 18698 104204 27950
rect 105096 26234 105124 30124
rect 107028 26234 107056 30124
rect 104912 26206 105124 26234
rect 106384 26206 107056 26234
rect 104912 23458 104940 26206
rect 104900 23452 104952 23458
rect 104900 23394 104952 23400
rect 104164 18692 104216 18698
rect 104164 18634 104216 18640
rect 99380 18624 99432 18630
rect 99380 18566 99432 18572
rect 98000 17944 98052 17950
rect 98000 17886 98052 17892
rect 99392 16574 99420 18566
rect 106384 17882 106412 26206
rect 107672 21865 107700 30124
rect 108960 28082 108988 30124
rect 107752 28076 107804 28082
rect 107752 28018 107804 28024
rect 108948 28076 109000 28082
rect 108948 28018 109000 28024
rect 109040 28076 109092 28082
rect 109040 28018 109092 28024
rect 107764 22642 107792 28018
rect 109052 27674 109080 28018
rect 109040 27668 109092 27674
rect 109040 27610 109092 27616
rect 109604 26994 109632 30124
rect 116044 28234 116072 30124
rect 115952 28206 116072 28234
rect 109592 26988 109644 26994
rect 109592 26930 109644 26936
rect 110420 22772 110472 22778
rect 110420 22714 110472 22720
rect 107752 22636 107804 22642
rect 107752 22578 107804 22584
rect 107658 21856 107714 21865
rect 107658 21791 107714 21800
rect 106372 17876 106424 17882
rect 106372 17818 106424 17824
rect 106280 16652 106332 16658
rect 106280 16594 106332 16600
rect 70412 16546 71544 16574
rect 77312 16546 78168 16574
rect 81452 16546 81664 16574
rect 85592 16546 85712 16574
rect 88352 16546 89208 16574
rect 99392 16546 99880 16574
rect 71516 480 71544 16546
rect 74998 3496 75054 3505
rect 74998 3431 75054 3440
rect 75012 480 75040 3431
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 85684 480 85712 16546
rect 89180 480 89208 16546
rect 92756 3460 92808 3466
rect 92756 3402 92808 3408
rect 92768 480 92796 3402
rect 96252 3392 96304 3398
rect 96252 3334 96304 3340
rect 96264 480 96292 3334
rect 99852 480 99880 16546
rect 106292 6914 106320 16594
rect 110432 16574 110460 22714
rect 113180 18692 113232 18698
rect 113180 18634 113232 18640
rect 113192 16574 113220 18634
rect 115952 17338 115980 28206
rect 116688 26234 116716 30124
rect 117976 28121 118004 30124
rect 117962 28112 118018 28121
rect 117962 28047 118018 28056
rect 120552 26234 120580 30124
rect 123772 29442 123800 30124
rect 123760 29436 123812 29442
rect 123760 29378 123812 29384
rect 124416 26234 124444 30124
rect 125704 28234 125732 30124
rect 116044 26206 116716 26234
rect 120092 26206 120580 26234
rect 124232 26206 124444 26234
rect 125612 28206 125732 28234
rect 116044 17814 116072 26206
rect 120092 18358 120120 26206
rect 124232 24138 124260 26206
rect 124220 24132 124272 24138
rect 124220 24074 124272 24080
rect 124218 21312 124274 21321
rect 124218 21247 124274 21256
rect 120080 18352 120132 18358
rect 120080 18294 120132 18300
rect 116032 17808 116084 17814
rect 116032 17750 116084 17756
rect 115940 17332 115992 17338
rect 115940 17274 115992 17280
rect 120080 17264 120132 17270
rect 120080 17206 120132 17212
rect 120092 16574 120120 17206
rect 124232 16574 124260 21247
rect 125612 18766 125640 28206
rect 126348 26234 126376 30124
rect 127652 29866 127680 30124
rect 127636 29838 127680 29866
rect 127636 28937 127664 29838
rect 127622 28928 127678 28937
rect 127622 28863 127678 28872
rect 128924 27742 128952 30124
rect 128912 27736 128964 27742
rect 128912 27678 128964 27684
rect 129568 26234 129596 30124
rect 131516 29866 131544 30124
rect 131132 29838 131544 29866
rect 130200 28348 130252 28354
rect 130200 28290 130252 28296
rect 125704 26206 126376 26234
rect 128464 26206 129596 26234
rect 125704 23089 125732 26206
rect 128464 23322 128492 26206
rect 128452 23316 128504 23322
rect 128452 23258 128504 23264
rect 125690 23080 125746 23089
rect 125690 23015 125746 23024
rect 125690 21448 125746 21457
rect 125690 21383 125746 21392
rect 125600 18760 125652 18766
rect 125600 18702 125652 18708
rect 110432 16546 110552 16574
rect 113192 16546 114048 16574
rect 120092 16546 120672 16574
rect 124232 16546 124720 16574
rect 106292 6886 106504 6914
rect 103334 3360 103390 3369
rect 103334 3295 103390 3304
rect 103348 480 103376 3295
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 6886
rect 110524 480 110552 16546
rect 114020 480 114048 16546
rect 117596 4140 117648 4146
rect 117596 4082 117648 4088
rect 117608 480 117636 4082
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 124692 480 124720 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125704 354 125732 21383
rect 130212 19854 130240 28290
rect 131132 23390 131160 29838
rect 132144 26234 132172 30124
rect 138584 26234 138612 30124
rect 139888 29866 139916 30124
rect 131224 26206 132172 26234
rect 138032 26206 138612 26234
rect 139504 29838 139916 29866
rect 131224 24206 131252 26206
rect 131212 24200 131264 24206
rect 131212 24142 131264 24148
rect 131120 23384 131172 23390
rect 131120 23326 131172 23332
rect 138032 23089 138060 26206
rect 138018 23080 138074 23089
rect 138018 23015 138074 23024
rect 135258 21312 135314 21321
rect 135258 21247 135314 21256
rect 130200 19848 130252 19854
rect 130200 19790 130252 19796
rect 128358 18592 128414 18601
rect 128358 18527 128414 18536
rect 128372 16574 128400 18527
rect 128372 16546 128952 16574
rect 126978 3360 127034 3369
rect 126978 3295 127034 3304
rect 126992 480 127020 3295
rect 125846 354 125958 480
rect 125704 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130568 15972 130620 15978
rect 130568 15914 130620 15920
rect 130580 480 130608 15914
rect 132958 10296 133014 10305
rect 132958 10231 133014 10240
rect 132972 480 133000 10231
rect 135272 3534 135300 21247
rect 139400 19984 139452 19990
rect 139400 19926 139452 19932
rect 136640 18760 136692 18766
rect 136640 18702 136692 18708
rect 136652 16574 136680 18702
rect 139412 16574 139440 19926
rect 139504 18873 139532 29838
rect 141804 28490 141832 30124
rect 141792 28484 141844 28490
rect 141792 28426 141844 28432
rect 143092 28234 143120 30124
rect 143172 28620 143224 28626
rect 143172 28562 143224 28568
rect 142172 28206 143120 28234
rect 142172 24070 142200 28206
rect 143184 26234 143212 28562
rect 142816 26206 143212 26234
rect 142160 24064 142212 24070
rect 142160 24006 142212 24012
rect 139490 18864 139546 18873
rect 139490 18799 139546 18808
rect 142816 17406 142844 26206
rect 146312 18902 146340 30124
rect 148888 28490 148916 30124
rect 147680 28484 147732 28490
rect 147680 28426 147732 28432
rect 148876 28484 148928 28490
rect 148876 28426 148928 28432
rect 147692 21486 147720 28426
rect 149532 26234 149560 30124
rect 151464 26234 151492 30124
rect 154684 26234 154712 30124
rect 155972 27810 156000 30124
rect 157276 29918 157304 30124
rect 156052 29912 156104 29918
rect 156052 29854 156104 29860
rect 157264 29912 157316 29918
rect 157264 29854 157316 29860
rect 155960 27804 156012 27810
rect 155960 27746 156012 27752
rect 149072 26206 149560 26234
rect 150544 26206 151492 26234
rect 154592 26206 154712 26234
rect 147680 21480 147732 21486
rect 147680 21422 147732 21428
rect 146392 21412 146444 21418
rect 146392 21354 146444 21360
rect 146300 18896 146352 18902
rect 146300 18838 146352 18844
rect 142804 17400 142856 17406
rect 142804 17342 142856 17348
rect 146404 16574 146432 21354
rect 149072 18970 149100 26206
rect 150438 21448 150494 21457
rect 150438 21383 150494 21392
rect 149060 18964 149112 18970
rect 149060 18906 149112 18912
rect 147680 18556 147732 18562
rect 147680 18498 147732 18504
rect 147692 16574 147720 18498
rect 136652 16546 137232 16574
rect 139412 16546 139624 16574
rect 146404 16546 147168 16574
rect 147692 16546 147904 16574
rect 134156 3528 134208 3534
rect 134156 3470 134208 3476
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 136456 3528 136508 3534
rect 136456 3470 136508 3476
rect 134168 480 134196 3470
rect 136468 480 136496 3470
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 143538 16008 143594 16017
rect 143538 15943 143594 15952
rect 141240 10328 141292 10334
rect 141240 10270 141292 10276
rect 141252 480 141280 10270
rect 143552 3534 143580 15943
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144736 3528 144788 3534
rect 144736 3470 144788 3476
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 143540 2848 143592 2854
rect 143540 2790 143592 2796
rect 143552 480 143580 2790
rect 144748 480 144776 3470
rect 144840 2854 144868 3470
rect 144828 2848 144880 2854
rect 144828 2790 144880 2796
rect 147140 480 147168 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 150452 6914 150480 21383
rect 150544 16561 150572 26206
rect 151818 19952 151874 19961
rect 151818 19887 151874 19896
rect 153200 19916 153252 19922
rect 150530 16552 150586 16561
rect 150530 16487 150586 16496
rect 150452 6886 150664 6914
rect 150636 480 150664 6886
rect 151832 480 151860 19887
rect 153200 19858 153252 19864
rect 153212 16574 153240 19858
rect 154592 18494 154620 26206
rect 156064 21554 156092 29854
rect 157984 28484 158036 28490
rect 157984 28426 158036 28432
rect 157340 27532 157392 27538
rect 157340 27474 157392 27480
rect 156052 21548 156104 21554
rect 156052 21490 156104 21496
rect 154580 18488 154632 18494
rect 154580 18430 154632 18436
rect 157352 17814 157380 27474
rect 157340 17808 157392 17814
rect 157340 17750 157392 17756
rect 153212 16546 153792 16574
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 157996 16454 158024 28426
rect 158548 27538 158576 30124
rect 159836 29034 159864 30124
rect 161140 29866 161168 30124
rect 160112 29838 161168 29866
rect 159824 29028 159876 29034
rect 159824 28970 159876 28976
rect 158536 27532 158588 27538
rect 158536 27474 158588 27480
rect 160112 22574 160140 29838
rect 162412 26234 162440 30124
rect 161584 26206 162440 26234
rect 160100 22568 160152 22574
rect 160100 22510 160152 22516
rect 161478 21584 161534 21593
rect 161478 21519 161534 21528
rect 157984 16448 158036 16454
rect 157984 16390 158036 16396
rect 158904 15904 158956 15910
rect 157798 15872 157854 15881
rect 158904 15846 158956 15852
rect 157798 15807 157854 15816
rect 155406 7576 155462 7585
rect 155406 7511 155462 7520
rect 155420 480 155448 7511
rect 157812 480 157840 15807
rect 158916 480 158944 15846
rect 161492 6914 161520 21519
rect 161584 16522 161612 26206
rect 164238 24168 164294 24177
rect 164238 24103 164294 24112
rect 161572 16516 161624 16522
rect 161572 16458 161624 16464
rect 164252 6914 164280 24103
rect 164344 16590 164372 30124
rect 165648 29866 165676 30124
rect 165648 29838 165752 29866
rect 165724 25702 165752 29838
rect 166276 26234 166304 30124
rect 166920 27878 166948 30124
rect 168208 28150 168236 30124
rect 169512 29866 169540 30124
rect 169496 29838 169540 29866
rect 169496 28393 169524 29838
rect 169482 28384 169538 28393
rect 169482 28319 169538 28328
rect 170784 28234 170812 30124
rect 170864 28756 170916 28762
rect 170864 28698 170916 28704
rect 169772 28206 170812 28234
rect 168196 28144 168248 28150
rect 168196 28086 168248 28092
rect 166908 27872 166960 27878
rect 166908 27814 166960 27820
rect 165816 26206 166304 26234
rect 165712 25696 165764 25702
rect 165712 25638 165764 25644
rect 165816 24585 165844 26206
rect 165802 24576 165858 24585
rect 165802 24511 165858 24520
rect 168380 22772 168432 22778
rect 168380 22714 168432 22720
rect 165620 18828 165672 18834
rect 165620 18770 165672 18776
rect 164332 16584 164384 16590
rect 165632 16574 165660 18770
rect 165632 16546 166120 16574
rect 164332 16526 164384 16532
rect 161492 6886 162072 6914
rect 164252 6886 164464 6914
rect 161296 3800 161348 3806
rect 161296 3742 161348 3748
rect 161308 480 161336 3742
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 6886
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 6886
rect 166092 480 166120 16546
rect 168392 480 168420 22714
rect 169772 21622 169800 28206
rect 170876 27674 170904 28698
rect 170404 27668 170456 27674
rect 170404 27610 170456 27616
rect 170864 27668 170916 27674
rect 170864 27610 170916 27616
rect 169760 21616 169812 21622
rect 169760 21558 169812 21564
rect 170416 17202 170444 27610
rect 171428 26234 171456 30124
rect 174020 29866 174048 30124
rect 171152 26206 171456 26234
rect 173912 29838 174048 29866
rect 171152 22846 171180 26206
rect 171140 22840 171192 22846
rect 171140 22782 171192 22788
rect 173912 20097 173940 29838
rect 174648 27441 174676 30124
rect 175292 28529 175320 30124
rect 175278 28520 175334 28529
rect 175278 28455 175334 28464
rect 174634 27432 174690 27441
rect 174634 27367 174690 27376
rect 178512 26234 178540 30124
rect 179800 27946 179828 30124
rect 181088 28218 181116 30124
rect 182392 29866 182420 30124
rect 182376 29838 182420 29866
rect 182376 29034 182404 29838
rect 182364 29028 182416 29034
rect 182364 28970 182416 28976
rect 181076 28212 181128 28218
rect 181076 28154 181128 28160
rect 179788 27940 179840 27946
rect 179788 27882 179840 27888
rect 183020 26234 183048 30124
rect 183664 26234 183692 30124
rect 178052 26206 178540 26234
rect 182192 26206 183048 26234
rect 183572 26206 183692 26234
rect 176660 21480 176712 21486
rect 176660 21422 176712 21428
rect 173898 20088 173954 20097
rect 173898 20023 173954 20032
rect 170404 17196 170456 17202
rect 170404 17138 170456 17144
rect 171968 15904 172020 15910
rect 171968 15846 172020 15852
rect 169574 3496 169630 3505
rect 169574 3431 169630 3440
rect 169588 480 169616 3431
rect 171980 480 172008 15846
rect 175464 3800 175516 3806
rect 175464 3742 175516 3748
rect 173162 3632 173218 3641
rect 173162 3567 173218 3576
rect 173176 480 173204 3567
rect 175476 480 175504 3742
rect 176672 480 176700 21422
rect 178052 17785 178080 26206
rect 182192 24274 182220 26206
rect 182180 24268 182232 24274
rect 182180 24210 182232 24216
rect 179418 21720 179474 21729
rect 179418 21655 179474 21664
rect 178038 17776 178094 17785
rect 178038 17711 178094 17720
rect 179432 16574 179460 21655
rect 183572 19038 183600 26206
rect 184952 23390 184980 30124
rect 186256 29866 186284 30124
rect 186240 29838 186284 29866
rect 186240 28257 186268 29838
rect 186226 28248 186282 28257
rect 187528 28218 187556 30124
rect 188816 28558 188844 30124
rect 188804 28552 188856 28558
rect 188804 28494 188856 28500
rect 186226 28183 186282 28192
rect 186320 28212 186372 28218
rect 186320 28154 186372 28160
rect 187516 28212 187568 28218
rect 187516 28154 187568 28160
rect 186332 25770 186360 28154
rect 189460 26234 189488 30124
rect 190764 29866 190792 30124
rect 190748 29838 190792 29866
rect 190748 28694 190776 29838
rect 190736 28688 190788 28694
rect 190736 28630 190788 28636
rect 191392 26234 191420 30124
rect 191840 28212 191892 28218
rect 191840 28154 191892 28160
rect 189092 26206 189488 26234
rect 190564 26206 191420 26234
rect 186320 25764 186372 25770
rect 186320 25706 186372 25712
rect 184940 23384 184992 23390
rect 184940 23326 184992 23332
rect 184940 20052 184992 20058
rect 184940 19994 184992 20000
rect 183652 19984 183704 19990
rect 183652 19926 183704 19932
rect 183560 19032 183612 19038
rect 183560 18974 183612 18980
rect 183664 16574 183692 19926
rect 179432 16546 180288 16574
rect 183664 16546 183784 16574
rect 179050 6216 179106 6225
rect 179050 6151 179106 6160
rect 179064 480 179092 6151
rect 180260 480 180288 16546
rect 182548 4072 182600 4078
rect 182548 4014 182600 4020
rect 182560 480 182588 4014
rect 183756 480 183784 16546
rect 184952 3602 184980 19994
rect 189092 19718 189120 26206
rect 189080 19712 189132 19718
rect 189080 19654 189132 19660
rect 190564 12442 190592 26206
rect 190552 12436 190604 12442
rect 190552 12378 190604 12384
rect 191852 11014 191880 28154
rect 192036 26234 192064 30124
rect 192680 28218 192708 30124
rect 193324 29238 193352 30124
rect 195256 29306 195284 30124
rect 195244 29300 195296 29306
rect 195244 29242 195296 29248
rect 193312 29232 193364 29238
rect 193312 29174 193364 29180
rect 192668 28212 192720 28218
rect 192668 28154 192720 28160
rect 195900 28014 195928 30124
rect 195888 28008 195940 28014
rect 195888 27950 195940 27956
rect 197832 26234 197860 30124
rect 199764 29374 199792 30124
rect 199752 29368 199804 29374
rect 199752 29310 199804 29316
rect 201696 28082 201724 30124
rect 201684 28076 201736 28082
rect 201684 28018 201736 28024
rect 203628 26234 203656 30124
rect 204916 26234 204944 30124
rect 205560 29170 205588 30124
rect 205548 29164 205600 29170
rect 205548 29106 205600 29112
rect 206204 26234 206232 30124
rect 208136 26234 208164 30124
rect 210068 26234 210096 30124
rect 211372 29866 211400 30124
rect 211356 29838 211400 29866
rect 211356 28422 211384 29838
rect 211344 28416 211396 28422
rect 211344 28358 211396 28364
rect 212000 26234 212028 30124
rect 191944 26206 192064 26234
rect 197372 26206 197860 26234
rect 202892 26206 203656 26234
rect 204272 26206 204944 26234
rect 205652 26206 206232 26234
rect 207032 26206 208164 26234
rect 209792 26206 210096 26234
rect 211264 26206 212028 26234
rect 191944 24342 191972 26206
rect 191932 24336 191984 24342
rect 191932 24278 191984 24284
rect 197372 21690 197400 26206
rect 197360 21684 197412 21690
rect 197360 21626 197412 21632
rect 202892 19174 202920 26206
rect 204272 24410 204300 26206
rect 204260 24404 204312 24410
rect 204260 24346 204312 24352
rect 204258 19952 204314 19961
rect 204258 19887 204314 19896
rect 202880 19168 202932 19174
rect 202880 19110 202932 19116
rect 204272 16574 204300 19887
rect 205652 19106 205680 26206
rect 207032 25673 207060 26206
rect 207018 25664 207074 25673
rect 207018 25599 207074 25608
rect 207018 24304 207074 24313
rect 207018 24239 207074 24248
rect 205640 19100 205692 19106
rect 205640 19042 205692 19048
rect 204272 16546 205128 16574
rect 191840 11008 191892 11014
rect 191840 10950 191892 10956
rect 201498 10432 201554 10441
rect 201498 10367 201554 10376
rect 194416 7608 194468 7614
rect 194416 7550 194468 7556
rect 189724 4004 189776 4010
rect 189724 3946 189776 3952
rect 184848 3596 184900 3602
rect 184848 3538 184900 3544
rect 184940 3596 184992 3602
rect 184940 3538 184992 3544
rect 186136 3596 186188 3602
rect 186136 3538 186188 3544
rect 184860 3398 184888 3538
rect 184848 3392 184900 3398
rect 184848 3334 184900 3340
rect 186148 480 186176 3538
rect 187332 3392 187384 3398
rect 187332 3334 187384 3340
rect 187344 480 187372 3334
rect 189736 480 189764 3946
rect 193220 3936 193272 3942
rect 193220 3878 193272 3884
rect 190828 3596 190880 3602
rect 190828 3538 190880 3544
rect 190840 480 190868 3538
rect 193232 480 193260 3878
rect 194428 480 194456 7550
rect 196808 3868 196860 3874
rect 196808 3810 196860 3816
rect 196820 480 196848 3810
rect 197912 3732 197964 3738
rect 197912 3674 197964 3680
rect 197924 480 197952 3674
rect 200304 3188 200356 3194
rect 200304 3130 200356 3136
rect 200316 480 200344 3130
rect 201512 480 201540 10367
rect 203890 3632 203946 3641
rect 203890 3567 203946 3576
rect 203904 480 203932 3567
rect 205100 480 205128 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 24239
rect 209792 21894 209820 26206
rect 209872 24132 209924 24138
rect 209872 24074 209924 24080
rect 209780 21888 209832 21894
rect 209780 21830 209832 21836
rect 209884 16574 209912 24074
rect 211264 20126 211292 26206
rect 211252 20120 211304 20126
rect 211252 20062 211304 20068
rect 212644 17649 212672 30124
rect 213288 28286 213316 30124
rect 213932 28801 213960 30124
rect 213918 28792 213974 28801
rect 213918 28727 213974 28736
rect 213276 28280 213328 28286
rect 213276 28222 213328 28228
rect 216508 28218 216536 30124
rect 215300 28212 215352 28218
rect 215300 28154 215352 28160
rect 216496 28212 216548 28218
rect 216496 28154 216548 28160
rect 215312 22710 215340 28154
rect 217152 26234 217180 30124
rect 217796 29102 217824 30124
rect 219744 29866 219772 30124
rect 219452 29838 219772 29866
rect 217784 29096 217836 29102
rect 217784 29038 217836 29044
rect 216692 26206 217180 26234
rect 216692 25838 216720 26206
rect 216680 25832 216732 25838
rect 216680 25774 216732 25780
rect 215300 22704 215352 22710
rect 215300 22646 215352 22652
rect 219452 19310 219480 29838
rect 220372 26234 220400 30124
rect 221016 26234 221044 30124
rect 222948 26234 222976 30124
rect 224252 29866 224280 30124
rect 228116 29866 228144 30124
rect 219544 26206 220400 26234
rect 220924 26206 221044 26234
rect 222212 26206 222976 26234
rect 223592 29838 224280 29866
rect 227732 29838 228144 29866
rect 219544 20330 219572 26206
rect 220820 24200 220872 24206
rect 220820 24142 220872 24148
rect 219532 20324 219584 20330
rect 219532 20266 219584 20272
rect 219440 19304 219492 19310
rect 219440 19246 219492 19252
rect 212630 17640 212686 17649
rect 212630 17575 212686 17584
rect 218058 17232 218114 17241
rect 218058 17167 218114 17176
rect 209884 16546 211016 16574
rect 208584 8968 208636 8974
rect 208584 8910 208636 8916
rect 208596 480 208624 8910
rect 210988 480 211016 16546
rect 214470 16144 214526 16153
rect 214470 16079 214526 16088
rect 212172 3936 212224 3942
rect 212172 3878 212224 3884
rect 212184 480 212212 3878
rect 214484 480 214512 16079
rect 215668 3664 215720 3670
rect 215668 3606 215720 3612
rect 215680 480 215708 3606
rect 218072 3398 218100 17167
rect 220832 6914 220860 24142
rect 220924 15201 220952 26206
rect 222212 19009 222240 26206
rect 223592 21894 223620 29838
rect 224960 24268 225012 24274
rect 224960 24210 225012 24216
rect 223580 21888 223632 21894
rect 223580 21830 223632 21836
rect 222198 19000 222254 19009
rect 222198 18935 222254 18944
rect 224972 16574 225000 24210
rect 227732 20194 227760 29838
rect 230032 26234 230060 30124
rect 232624 29866 232652 30124
rect 229112 26206 230060 26234
rect 231964 29838 232652 29866
rect 229112 20398 229140 26206
rect 231860 24880 231912 24886
rect 231860 24822 231912 24828
rect 229100 20392 229152 20398
rect 229100 20334 229152 20340
rect 227720 20188 227772 20194
rect 227720 20130 227772 20136
rect 224972 16546 225184 16574
rect 220910 15192 220966 15201
rect 220910 15127 220966 15136
rect 220832 6886 221136 6914
rect 218152 3664 218204 3670
rect 218152 3606 218204 3612
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218164 1850 218192 3606
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 218072 1822 218192 1850
rect 218072 480 218100 1822
rect 219268 480 219296 3334
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 6886
rect 222752 4004 222804 4010
rect 222752 3946 222804 3952
rect 222764 480 222792 3946
rect 225156 480 225184 16546
rect 228272 16108 228324 16114
rect 228272 16050 228324 16056
rect 226340 16040 226392 16046
rect 226340 15982 226392 15988
rect 226352 480 226380 15982
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16050
rect 229376 15972 229428 15978
rect 229376 15914 229428 15920
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 15914
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 24822
rect 231964 20398 231992 29838
rect 231952 20392 232004 20398
rect 231952 20334 232004 20340
rect 233252 16590 233280 30124
rect 234540 28801 234568 30124
rect 234526 28792 234582 28801
rect 234526 28727 234582 28736
rect 235184 26234 235212 30124
rect 237116 26234 237144 30124
rect 238404 26234 238432 30124
rect 243556 26234 243584 30124
rect 244200 29345 244228 30124
rect 244186 29336 244242 29345
rect 244186 29271 244242 29280
rect 246776 26234 246804 30124
rect 247420 26234 247448 30124
rect 249996 28762 250024 30124
rect 249984 28756 250036 28762
rect 249984 28698 250036 28704
rect 251284 28626 251312 30124
rect 251272 28620 251324 28626
rect 251272 28562 251324 28568
rect 251928 26234 251956 30124
rect 252572 28354 252600 30124
rect 252560 28348 252612 28354
rect 252560 28290 252612 28296
rect 256436 26234 256464 30124
rect 257740 29866 257768 30124
rect 234632 26206 235212 26234
rect 236012 26206 237144 26234
rect 237392 26206 238432 26234
rect 242912 26206 243584 26234
rect 245764 26206 246804 26234
rect 247052 26206 247448 26234
rect 251284 26206 251956 26234
rect 255332 26206 256464 26234
rect 256712 29838 257768 29866
rect 234632 17474 234660 26206
rect 236012 21865 236040 26206
rect 235998 21856 236054 21865
rect 235998 21791 236054 21800
rect 237392 17542 237420 26206
rect 237380 17536 237432 17542
rect 237380 17478 237432 17484
rect 234620 17468 234672 17474
rect 234620 17410 234672 17416
rect 233240 16584 233292 16590
rect 233240 16526 233292 16532
rect 242912 15162 242940 26206
rect 245660 24336 245712 24342
rect 245660 24278 245712 24284
rect 245672 16574 245700 24278
rect 245764 17610 245792 26206
rect 247052 19310 247080 26206
rect 251284 20330 251312 26206
rect 255332 21758 255360 26206
rect 256712 24546 256740 29838
rect 259012 28558 259040 30124
rect 260944 29102 260972 30124
rect 266112 29866 266140 30124
rect 266096 29838 266140 29866
rect 260932 29096 260984 29102
rect 260932 29038 260984 29044
rect 259000 28552 259052 28558
rect 259000 28494 259052 28500
rect 266096 28286 266124 29838
rect 266084 28280 266136 28286
rect 266084 28222 266136 28228
rect 266740 27130 266768 30124
rect 268028 28354 268056 30124
rect 268016 28348 268068 28354
rect 268016 28290 268068 28296
rect 268672 27130 268700 30124
rect 270620 29866 270648 30124
rect 270512 29838 270648 29866
rect 266728 27124 266780 27130
rect 266728 27066 266780 27072
rect 268660 27124 268712 27130
rect 268660 27066 268712 27072
rect 256700 24540 256752 24546
rect 256700 24482 256752 24488
rect 270512 22914 270540 29838
rect 271248 28898 271276 30124
rect 271236 28892 271288 28898
rect 271236 28834 271288 28840
rect 272536 28490 272564 30124
rect 272524 28484 272576 28490
rect 272524 28426 272576 28432
rect 275112 26234 275140 30124
rect 275756 27878 275784 30124
rect 275744 27872 275796 27878
rect 275744 27814 275796 27820
rect 276400 26234 276428 30124
rect 280264 26234 280292 30124
rect 284128 29209 284156 30124
rect 284114 29200 284170 29209
rect 284114 29135 284170 29144
rect 286060 26234 286088 30124
rect 287364 29866 287392 30124
rect 287348 29838 287392 29866
rect 287348 29170 287376 29838
rect 287336 29164 287388 29170
rect 287336 29106 287388 29112
rect 289280 26234 289308 30124
rect 291228 29866 291256 30124
rect 274652 26206 275140 26234
rect 276032 26206 276428 26234
rect 280172 26206 280292 26234
rect 285692 26206 286088 26234
rect 288452 26206 289308 26234
rect 291212 29838 291256 29866
rect 274652 24449 274680 26206
rect 274638 24440 274694 24449
rect 274638 24375 274694 24384
rect 270500 22908 270552 22914
rect 270500 22850 270552 22856
rect 255320 21752 255372 21758
rect 255320 21694 255372 21700
rect 258080 21616 258132 21622
rect 258080 21558 258132 21564
rect 251272 20324 251324 20330
rect 251272 20266 251324 20272
rect 253940 20120 253992 20126
rect 253940 20062 253992 20068
rect 247040 19304 247092 19310
rect 247040 19246 247092 19252
rect 251180 18828 251232 18834
rect 251180 18770 251232 18776
rect 245752 17604 245804 17610
rect 245752 17546 245804 17552
rect 245672 16546 245976 16574
rect 242900 15156 242952 15162
rect 242900 15098 242952 15104
rect 236550 14512 236606 14521
rect 236550 14447 236606 14456
rect 234620 13184 234672 13190
rect 234620 13126 234672 13132
rect 234632 3398 234660 13126
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 235828 480 235856 3334
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 82 233506 480
rect 233394 66 233832 82
rect 233394 60 233844 66
rect 233394 54 233792 60
rect 233394 -960 233506 54
rect 233792 2 233844 8
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 14447
rect 242900 13116 242952 13122
rect 242900 13058 242952 13064
rect 239312 11756 239364 11762
rect 239312 11698 239364 11704
rect 239324 480 239352 11698
rect 240508 3868 240560 3874
rect 240508 3810 240560 3816
rect 240520 480 240548 3810
rect 242912 3398 242940 13058
rect 242990 3768 243046 3777
rect 242990 3703 243046 3712
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 243004 1850 243032 3703
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 242912 1822 243032 1850
rect 242912 480 242940 1822
rect 244108 480 244136 3334
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247592 14476 247644 14482
rect 247592 14418 247644 14424
rect 247604 480 247632 14418
rect 249984 9036 250036 9042
rect 249984 8978 250036 8984
rect 249996 480 250024 8978
rect 251192 480 251220 18770
rect 253952 16574 253980 20062
rect 258092 16574 258120 21558
rect 260840 21548 260892 21554
rect 260840 21490 260892 21496
rect 259460 17332 259512 17338
rect 259460 17274 259512 17280
rect 253952 16546 254256 16574
rect 258092 16546 258304 16574
rect 253480 16176 253532 16182
rect 253480 16118 253532 16124
rect 253492 480 253520 16118
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 256700 11824 256752 11830
rect 256700 11766 256752 11772
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 11766
rect 258276 480 258304 16546
rect 259472 3398 259500 17274
rect 260852 16574 260880 21490
rect 271880 18896 271932 18902
rect 267738 18864 267794 18873
rect 271880 18838 271932 18844
rect 267738 18799 267794 18808
rect 267752 16574 267780 18799
rect 271892 16574 271920 18838
rect 276032 16574 276060 26206
rect 280172 24546 280200 26206
rect 280160 24540 280212 24546
rect 280160 24482 280212 24488
rect 285692 23050 285720 26206
rect 285680 23044 285732 23050
rect 285680 22986 285732 22992
rect 282918 19000 282974 19009
rect 282918 18935 282974 18944
rect 278778 18728 278834 18737
rect 278778 18663 278834 18672
rect 278792 16574 278820 18663
rect 282932 16574 282960 18935
rect 260852 16546 261800 16574
rect 267752 16546 268424 16574
rect 271892 16546 272472 16574
rect 276032 16546 276152 16574
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 260668 480 260696 3334
rect 261772 480 261800 16546
rect 264980 16244 265032 16250
rect 264980 16186 265032 16192
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 16186
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 272444 480 272472 16546
rect 276018 7712 276074 7721
rect 276018 7647 276074 7656
rect 276032 480 276060 7647
rect 276124 1358 276152 16546
rect 276112 1352 276164 1358
rect 276112 1294 276164 1300
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 283116 480 283144 16546
rect 286600 13252 286652 13258
rect 286600 13194 286652 13200
rect 286612 480 286640 13194
rect 288452 5506 288480 26206
rect 291212 19145 291240 29838
rect 291856 28490 291884 30124
rect 291844 28484 291896 28490
rect 291844 28426 291896 28432
rect 293144 26234 293172 30124
rect 294432 26234 294460 30124
rect 295736 29866 295764 30124
rect 295720 29838 295764 29866
rect 295720 28830 295748 29838
rect 295708 28824 295760 28830
rect 295708 28766 295760 28772
rect 297008 27062 297036 30124
rect 299600 29866 299628 30124
rect 299492 29838 299628 29866
rect 296996 27056 297048 27062
rect 296996 26998 297048 27004
rect 292592 26206 293172 26234
rect 293972 26206 294460 26234
rect 292592 25906 292620 26206
rect 292580 25900 292632 25906
rect 292580 25842 292632 25848
rect 292580 20188 292632 20194
rect 292580 20130 292632 20136
rect 291198 19136 291254 19145
rect 291198 19071 291254 19080
rect 292592 16574 292620 20130
rect 293972 19242 294000 26206
rect 293960 19236 294012 19242
rect 293960 19178 294012 19184
rect 292592 16546 293264 16574
rect 289820 16312 289872 16318
rect 289820 16254 289872 16260
rect 288440 5500 288492 5506
rect 288440 5442 288492 5448
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 16254
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 297272 13320 297324 13326
rect 297272 13262 297324 13268
rect 297284 480 297312 13262
rect 299492 5438 299520 29838
rect 300872 28234 300900 30124
rect 300872 28206 300992 28234
rect 300860 28144 300912 28150
rect 300860 28086 300912 28092
rect 300872 19145 300900 28086
rect 300964 24041 300992 28206
rect 302160 28150 302188 30124
rect 304108 29866 304136 30124
rect 303632 29838 304136 29866
rect 302148 28144 302200 28150
rect 302148 28086 302200 28092
rect 300950 24032 301006 24041
rect 300950 23967 301006 23976
rect 303632 22982 303660 29838
rect 306024 26234 306052 30124
rect 306668 26234 306696 30124
rect 308600 26234 308628 30124
rect 311176 28626 311204 30124
rect 312480 29866 312508 30124
rect 311912 29838 312508 29866
rect 311164 28620 311216 28626
rect 311164 28562 311216 28568
rect 305012 26206 306052 26234
rect 306392 26206 306696 26234
rect 307772 26206 308628 26234
rect 303620 22976 303672 22982
rect 303620 22918 303672 22924
rect 305012 22545 305040 26206
rect 306392 25974 306420 26206
rect 307772 26042 307800 26206
rect 307760 26036 307812 26042
rect 307760 25978 307812 25984
rect 306380 25968 306432 25974
rect 306380 25910 306432 25916
rect 311912 24478 311940 29838
rect 313752 26234 313780 30124
rect 314396 29209 314424 30124
rect 314382 29200 314438 29209
rect 314382 29135 314438 29144
rect 315040 26234 315068 30124
rect 318904 26234 318932 30124
rect 319548 28665 319576 30124
rect 319534 28656 319590 28665
rect 319534 28591 319590 28600
rect 321480 28218 321508 30124
rect 320180 28212 320232 28218
rect 320180 28154 320232 28160
rect 321468 28212 321520 28218
rect 321468 28154 321520 28160
rect 321560 28212 321612 28218
rect 321560 28154 321612 28160
rect 313292 26206 313780 26234
rect 314764 26206 315068 26234
rect 318812 26206 318932 26234
rect 311900 24472 311952 24478
rect 311900 24414 311952 24420
rect 304998 22536 305054 22545
rect 304998 22471 305054 22480
rect 300858 19136 300914 19145
rect 300858 19071 300914 19080
rect 311440 13388 311492 13394
rect 311440 13330 311492 13336
rect 303896 10396 303948 10402
rect 303896 10338 303948 10344
rect 300768 6180 300820 6186
rect 300768 6122 300820 6128
rect 299480 5432 299532 5438
rect 299480 5374 299532 5380
rect 300780 480 300808 6122
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 10338
rect 307944 9104 307996 9110
rect 307944 9046 307996 9052
rect 307956 480 307984 9046
rect 311452 480 311480 13330
rect 313292 12374 313320 26206
rect 314660 24948 314712 24954
rect 314660 24890 314712 24896
rect 313280 12368 313332 12374
rect 313280 12310 313332 12316
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 24890
rect 314764 12306 314792 26206
rect 318812 26110 318840 26206
rect 318800 26104 318852 26110
rect 318800 26046 318852 26052
rect 317420 18964 317472 18970
rect 317420 18906 317472 18912
rect 317432 16574 317460 18906
rect 317432 16546 318104 16574
rect 314752 12300 314804 12306
rect 314752 12242 314804 12248
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 320192 13802 320220 28154
rect 321572 23118 321600 28154
rect 322124 26234 322152 30124
rect 322768 28218 322796 30124
rect 322756 28212 322808 28218
rect 322756 28154 322808 28160
rect 323412 26234 323440 30124
rect 324716 29866 324744 30124
rect 324424 29838 324744 29866
rect 324320 28212 324372 28218
rect 324320 28154 324372 28160
rect 321664 26206 322152 26234
rect 322952 26206 323440 26234
rect 321560 23112 321612 23118
rect 321560 23054 321612 23060
rect 320180 13796 320232 13802
rect 320180 13738 320232 13744
rect 321664 12238 321692 26206
rect 322952 26110 322980 26206
rect 322940 26104 322992 26110
rect 322940 26046 322992 26052
rect 321744 25560 321796 25566
rect 321744 25502 321796 25508
rect 321756 16574 321784 25502
rect 321756 16546 322152 16574
rect 321652 12232 321704 12238
rect 321652 12174 321704 12180
rect 322124 480 322152 16546
rect 324332 12170 324360 28154
rect 324424 22681 324452 29838
rect 325344 28218 325372 30124
rect 325988 28966 326016 30124
rect 325976 28960 326028 28966
rect 325976 28902 326028 28908
rect 325332 28212 325384 28218
rect 325332 28154 325384 28160
rect 326632 26234 326660 30124
rect 327276 28014 327304 30124
rect 329224 29866 329252 30124
rect 328472 29838 329252 29866
rect 327264 28008 327316 28014
rect 327264 27950 327316 27956
rect 325804 26206 326660 26234
rect 325804 26042 325832 26206
rect 325792 26036 325844 26042
rect 325792 25978 325844 25984
rect 324410 22672 324466 22681
rect 324410 22607 324466 22616
rect 324410 13016 324466 13025
rect 324410 12951 324466 12960
rect 324320 12164 324372 12170
rect 324320 12106 324372 12112
rect 324424 3398 324452 12951
rect 328472 12102 328500 29838
rect 331140 28218 331168 30124
rect 329840 28212 329892 28218
rect 329840 28154 329892 28160
rect 331128 28212 331180 28218
rect 331128 28154 331180 28160
rect 329852 17678 329880 28154
rect 333716 26234 333744 30124
rect 334360 26234 334388 30124
rect 336292 26234 336320 30124
rect 337596 29866 337624 30124
rect 332612 26206 333744 26234
rect 333992 26206 334388 26234
rect 335464 26206 336320 26234
rect 336752 29838 337624 29866
rect 332612 25673 332640 26206
rect 332598 25664 332654 25673
rect 332598 25599 332654 25608
rect 333992 24614 334020 26206
rect 333980 24608 334032 24614
rect 333980 24550 334032 24556
rect 332600 24404 332652 24410
rect 332600 24346 332652 24352
rect 329840 17672 329892 17678
rect 329840 17614 329892 17620
rect 332612 16574 332640 24346
rect 335358 17368 335414 17377
rect 335358 17303 335414 17312
rect 332612 16546 332732 16574
rect 328460 12096 328512 12102
rect 328460 12038 328512 12044
rect 328734 11792 328790 11801
rect 328734 11727 328790 11736
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 11727
rect 332704 480 332732 16546
rect 335372 6914 335400 17303
rect 335464 16454 335492 26206
rect 336752 19281 336780 29838
rect 338224 28762 338252 30124
rect 338212 28756 338264 28762
rect 338212 28698 338264 28704
rect 339512 26234 339540 30124
rect 342104 29918 342132 30124
rect 340880 29912 340932 29918
rect 340880 29854 340932 29860
rect 342092 29912 342144 29918
rect 342092 29854 342144 29860
rect 339512 26206 339632 26234
rect 339498 25528 339554 25537
rect 339498 25463 339554 25472
rect 336738 19272 336794 19281
rect 336738 19207 336794 19216
rect 335452 16448 335504 16454
rect 335452 16390 335504 16396
rect 335372 6886 336320 6914
rect 336292 480 336320 6886
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 25463
rect 339604 13705 339632 26206
rect 340892 17678 340920 29854
rect 343376 26234 343404 30124
rect 344020 27946 344048 30124
rect 344008 27940 344060 27946
rect 344008 27882 344060 27888
rect 347240 26234 347268 30124
rect 347780 28212 347832 28218
rect 347780 28154 347832 28160
rect 342272 26206 343404 26234
rect 346412 26206 347268 26234
rect 342272 23186 342300 26206
rect 342352 25628 342404 25634
rect 342352 25570 342404 25576
rect 342260 23180 342312 23186
rect 342260 23122 342312 23128
rect 340880 17672 340932 17678
rect 340880 17614 340932 17620
rect 342364 16574 342392 25570
rect 342364 16546 342944 16574
rect 339590 13696 339646 13705
rect 339590 13631 339646 13640
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 346412 11966 346440 26206
rect 347792 16386 347820 28154
rect 347884 24041 347912 30124
rect 348528 28218 348556 30124
rect 348516 28212 348568 28218
rect 348516 28154 348568 28160
rect 352392 26234 352420 30124
rect 354680 28212 354732 28218
rect 354680 28154 354732 28160
rect 351932 26206 352420 26234
rect 347870 24032 347926 24041
rect 347870 23967 347926 23976
rect 347780 16380 347832 16386
rect 347780 16322 347832 16328
rect 349160 13592 349212 13598
rect 349160 13534 349212 13540
rect 346952 13524 347004 13530
rect 346952 13466 347004 13472
rect 346400 11960 346452 11966
rect 346400 11902 346452 11908
rect 346964 480 346992 13466
rect 349172 3398 349200 13534
rect 351932 12034 351960 26206
rect 354692 23254 354720 28154
rect 354968 26234 354996 30124
rect 355612 28218 355640 30124
rect 355600 28212 355652 28218
rect 355600 28154 355652 28160
rect 356256 26234 356284 30124
rect 356900 29238 356928 30124
rect 356888 29232 356940 29238
rect 356888 29174 356940 29180
rect 357544 26234 357572 30124
rect 358848 29866 358876 30124
rect 358848 29838 358952 29866
rect 358820 28212 358872 28218
rect 358820 28154 358872 28160
rect 354784 26206 354996 26234
rect 356072 26206 356284 26234
rect 357452 26206 357572 26234
rect 354784 24682 354812 26206
rect 354772 24676 354824 24682
rect 354772 24618 354824 24624
rect 354680 23248 354732 23254
rect 354680 23190 354732 23196
rect 356072 22506 356100 26206
rect 356060 22500 356112 22506
rect 356060 22442 356112 22448
rect 353298 17504 353354 17513
rect 353298 17439 353354 17448
rect 353312 16574 353340 17439
rect 353312 16546 353616 16574
rect 351920 12028 351972 12034
rect 351920 11970 351972 11976
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 357452 11694 357480 26206
rect 358832 19242 358860 28154
rect 358924 26897 358952 29838
rect 359476 29345 359504 30124
rect 359462 29336 359518 29345
rect 359462 29271 359518 29280
rect 360120 28218 360148 30124
rect 362712 29918 362740 30124
rect 361580 29912 361632 29918
rect 361580 29854 361632 29860
rect 362700 29912 362752 29918
rect 362700 29854 362752 29860
rect 360108 28212 360160 28218
rect 360108 28154 360160 28160
rect 358910 26888 358966 26897
rect 358910 26823 358966 26832
rect 360200 19916 360252 19922
rect 360200 19858 360252 19864
rect 358820 19236 358872 19242
rect 358820 19178 358872 19184
rect 360212 16574 360240 19858
rect 360212 16546 361160 16574
rect 357532 13660 357584 13666
rect 357532 13602 357584 13608
rect 357440 11688 357492 11694
rect 357440 11630 357492 11636
rect 357544 480 357572 13602
rect 361132 480 361160 16546
rect 361592 16522 361620 29854
rect 363340 26234 363368 30124
rect 363984 27198 364012 30124
rect 364628 28234 364656 30124
rect 364352 28206 364656 28234
rect 363972 27192 364024 27198
rect 363972 27134 364024 27140
rect 363064 26206 363368 26234
rect 361580 16516 361632 16522
rect 361580 16458 361632 16464
rect 363064 11898 363092 26206
rect 364352 21826 364380 28206
rect 365272 26234 365300 30124
rect 365916 26234 365944 30124
rect 367220 29866 367248 30124
rect 367204 29838 367248 29866
rect 367100 28212 367152 28218
rect 367100 28154 367152 28160
rect 364444 26206 365300 26234
rect 365732 26206 365944 26234
rect 364444 25809 364472 26206
rect 364430 25800 364486 25809
rect 364430 25735 364486 25744
rect 365732 23186 365760 26206
rect 365720 23180 365772 23186
rect 365720 23122 365772 23128
rect 364340 21820 364392 21826
rect 364340 21762 364392 21768
rect 367112 20466 367140 28154
rect 367100 20460 367152 20466
rect 367100 20402 367152 20408
rect 367204 20262 367232 29838
rect 367848 28218 367876 30124
rect 367836 28212 367888 28218
rect 367836 28154 367888 28160
rect 368480 28212 368532 28218
rect 368480 28154 368532 28160
rect 368492 26178 368520 28154
rect 369136 27033 369164 30124
rect 369780 28218 369808 30124
rect 369768 28212 369820 28218
rect 369768 28154 369820 28160
rect 369122 27024 369178 27033
rect 369122 26959 369178 26968
rect 368480 26172 368532 26178
rect 368480 26114 368532 26120
rect 373000 22094 373028 30124
rect 373644 29073 373672 30124
rect 375592 29866 375620 30124
rect 375392 29838 375620 29866
rect 373630 29064 373686 29073
rect 373630 28999 373686 29008
rect 373998 25800 374054 25809
rect 373998 25735 374054 25744
rect 372632 22066 373028 22094
rect 371240 21684 371292 21690
rect 371240 21626 371292 21632
rect 367192 20256 367244 20262
rect 367192 20198 367244 20204
rect 367744 13456 367796 13462
rect 367744 13398 367796 13404
rect 364616 13048 364668 13054
rect 364616 12990 364668 12996
rect 363052 11892 363104 11898
rect 363052 11834 363104 11840
rect 364628 480 364656 12990
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 13398
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 21626
rect 372632 13734 372660 22066
rect 372620 13728 372672 13734
rect 372620 13670 372672 13676
rect 374012 3398 374040 25735
rect 375392 17746 375420 29838
rect 377508 28665 377536 30124
rect 378152 30002 378180 30124
rect 378060 29974 378180 30002
rect 378060 29578 378088 29974
rect 379456 29918 379484 30124
rect 378140 29912 378192 29918
rect 378140 29854 378192 29860
rect 379444 29912 379496 29918
rect 379444 29854 379496 29860
rect 378048 29572 378100 29578
rect 378048 29514 378100 29520
rect 377494 28656 377550 28665
rect 377494 28591 377550 28600
rect 378152 17746 378180 29854
rect 378232 29572 378284 29578
rect 378232 29514 378284 29520
rect 378244 27169 378272 29514
rect 381372 27198 381400 30124
rect 381360 27192 381412 27198
rect 378230 27160 378286 27169
rect 381360 27134 381412 27140
rect 378230 27095 378286 27104
rect 382016 26234 382044 30124
rect 382660 26761 382688 30124
rect 384592 29306 384620 30124
rect 384580 29300 384632 29306
rect 384580 29242 384632 29248
rect 385236 27266 385264 30124
rect 385224 27260 385276 27266
rect 385224 27202 385276 27208
rect 382646 26752 382702 26761
rect 382646 26687 382702 26696
rect 385880 26234 385908 30124
rect 386524 26234 386552 30124
rect 387828 29866 387856 30124
rect 380912 26206 382044 26234
rect 385144 26206 385908 26234
rect 386432 26206 386552 26234
rect 387812 29838 387856 29866
rect 375380 17740 375432 17746
rect 375380 17682 375432 17688
rect 378140 17740 378192 17746
rect 378140 17682 378192 17688
rect 380912 15094 380940 26206
rect 385040 22908 385092 22914
rect 385040 22850 385092 22856
rect 385052 16574 385080 22850
rect 385144 21826 385172 26206
rect 385132 21820 385184 21826
rect 385132 21762 385184 21768
rect 385052 16546 386000 16574
rect 380900 15088 380952 15094
rect 380900 15030 380952 15036
rect 382372 14612 382424 14618
rect 382372 14554 382424 14560
rect 378416 14544 378468 14550
rect 378416 14486 378468 14492
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 14486
rect 382384 480 382412 14554
rect 385972 480 386000 16546
rect 386432 15065 386460 26206
rect 387812 20534 387840 29838
rect 389100 28218 389128 30124
rect 389088 28212 389140 28218
rect 389088 28154 389140 28160
rect 389744 27305 389772 30124
rect 389730 27296 389786 27305
rect 389730 27231 389786 27240
rect 390388 26994 390416 30124
rect 390376 26988 390428 26994
rect 390376 26930 390428 26936
rect 391940 26240 391992 26246
rect 392964 26234 392992 30124
rect 394252 26234 394280 30124
rect 398116 26234 398144 30124
rect 398760 27266 398788 30124
rect 398748 27260 398800 27266
rect 398748 27202 398800 27208
rect 399404 26234 399432 30124
rect 401336 26234 401364 30124
rect 403268 26234 403296 30124
rect 404572 29866 404600 30124
rect 409080 29866 409108 30124
rect 391992 26206 392992 26234
rect 393332 26206 394280 26234
rect 397472 26206 398144 26234
rect 398852 26206 399432 26234
rect 400232 26206 401364 26234
rect 402992 26206 403296 26234
rect 404372 29838 404600 29866
rect 408512 29838 409108 29866
rect 391940 26182 391992 26188
rect 391938 22672 391994 22681
rect 391938 22607 391994 22616
rect 387800 20528 387852 20534
rect 387800 20470 387852 20476
rect 391952 16574 391980 22607
rect 391952 16546 392624 16574
rect 386418 15056 386474 15065
rect 386418 14991 386474 15000
rect 389456 6248 389508 6254
rect 389456 6190 389508 6196
rect 389468 480 389496 6190
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 393332 15026 393360 26206
rect 396080 25764 396132 25770
rect 396080 25706 396132 25712
rect 393320 15020 393372 15026
rect 393320 14962 393372 14968
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 25706
rect 397472 24750 397500 26206
rect 397460 24744 397512 24750
rect 397460 24686 397512 24692
rect 398852 15842 398880 26206
rect 400232 21962 400260 26206
rect 400220 21956 400272 21962
rect 400220 21898 400272 21904
rect 402992 17105 403020 26206
rect 402978 17096 403034 17105
rect 402978 17031 403034 17040
rect 398840 15836 398892 15842
rect 398840 15778 398892 15784
rect 404372 14958 404400 29838
rect 408512 25945 408540 29838
rect 409708 29374 409736 30124
rect 409696 29368 409748 29374
rect 409696 29310 409748 29316
rect 410352 27062 410380 30124
rect 410340 27056 410392 27062
rect 410340 26998 410392 27004
rect 410996 26234 411024 30124
rect 411640 26234 411668 30124
rect 416148 26234 416176 30124
rect 417452 29866 417480 30124
rect 417436 29838 417480 29866
rect 417436 28150 417464 29838
rect 417424 28144 417476 28150
rect 417424 28086 417476 28092
rect 420012 26234 420040 30124
rect 421316 29866 421344 30124
rect 409984 26206 411024 26234
rect 411272 26206 411668 26234
rect 415412 26206 416176 26234
rect 419552 26206 420040 26234
rect 421024 29838 421344 29866
rect 408498 25936 408554 25945
rect 408498 25871 408554 25880
rect 409878 25936 409934 25945
rect 409878 25871 409934 25880
rect 407118 21176 407174 21185
rect 407118 21111 407174 21120
rect 407132 16574 407160 21111
rect 409892 16574 409920 25871
rect 409984 23118 410012 26206
rect 409972 23112 410024 23118
rect 409972 23054 410024 23060
rect 411272 22030 411300 26206
rect 415412 22817 415440 26206
rect 416780 25696 416832 25702
rect 416780 25638 416832 25644
rect 416688 22840 416740 22846
rect 415398 22808 415454 22817
rect 415398 22743 415454 22752
rect 416686 22808 416688 22817
rect 416740 22808 416742 22817
rect 416686 22743 416742 22752
rect 411260 22024 411312 22030
rect 411260 21966 411312 21972
rect 414020 17400 414072 17406
rect 414020 17342 414072 17348
rect 414032 16574 414060 17342
rect 416792 16574 416820 25638
rect 419552 19174 419580 26206
rect 420920 21752 420972 21758
rect 420920 21694 420972 21700
rect 419540 19168 419592 19174
rect 419540 19110 419592 19116
rect 407132 16546 407252 16574
rect 409892 16546 410840 16574
rect 414032 16546 414336 16574
rect 416792 16546 417464 16574
rect 404360 14952 404412 14958
rect 404360 14894 404412 14900
rect 403624 14748 403676 14754
rect 403624 14690 403676 14696
rect 398840 14680 398892 14686
rect 398840 14622 398892 14628
rect 398852 3398 398880 14622
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 403636 480 403664 14690
rect 407224 480 407252 16546
rect 410812 480 410840 16546
rect 414308 480 414336 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 21694
rect 421024 20466 421052 29838
rect 421944 27305 421972 30124
rect 421930 27296 421986 27305
rect 421930 27231 421986 27240
rect 423876 26234 423904 30124
rect 426440 28076 426492 28082
rect 426440 28018 426492 28024
rect 423692 26206 423904 26234
rect 423692 20534 423720 26206
rect 423680 20528 423732 20534
rect 423680 20470 423732 20476
rect 421012 20460 421064 20466
rect 421012 20402 421064 20408
rect 426452 14822 426480 28018
rect 427096 26234 427124 30124
rect 427740 28082 427768 30124
rect 429028 28082 429056 30124
rect 427728 28076 427780 28082
rect 427728 28018 427780 28024
rect 427820 28076 427872 28082
rect 427820 28018 427872 28024
rect 429016 28076 429068 28082
rect 429016 28018 429068 28024
rect 426544 26206 427124 26234
rect 426544 22953 426572 26206
rect 426530 22944 426586 22953
rect 426530 22879 426586 22888
rect 427832 21214 427860 28018
rect 431604 26234 431632 30124
rect 432248 26234 432276 30124
rect 434196 29866 434224 30124
rect 430592 26206 431632 26234
rect 431972 26206 432276 26234
rect 433352 29838 434224 29866
rect 427820 21208 427872 21214
rect 427820 21150 427872 21156
rect 427820 17468 427872 17474
rect 427820 17410 427872 17416
rect 427832 16574 427860 17410
rect 427832 16546 428504 16574
rect 426440 14816 426492 14822
rect 426440 14758 426492 14764
rect 424968 6316 425020 6322
rect 424968 6258 425020 6264
rect 424980 480 425008 6258
rect 428476 480 428504 16546
rect 430592 14414 430620 26206
rect 431972 16561 432000 26206
rect 431958 16552 432014 16561
rect 431958 16487 432014 16496
rect 430580 14408 430632 14414
rect 430580 14350 430632 14356
rect 433352 14278 433380 29838
rect 435468 26234 435496 30124
rect 437400 28082 437428 30124
rect 436100 28076 436152 28082
rect 436100 28018 436152 28024
rect 437388 28076 437440 28082
rect 437388 28018 437440 28024
rect 434824 26206 435496 26234
rect 434720 20256 434772 20262
rect 434720 20198 434772 20204
rect 433340 14272 433392 14278
rect 433340 14214 433392 14220
rect 434732 6914 434760 20198
rect 434824 14346 434852 26206
rect 436112 24750 436140 28018
rect 439332 26234 439360 30124
rect 440620 26234 440648 30124
rect 441264 27334 441292 30124
rect 443196 28694 443224 30124
rect 443184 28688 443236 28694
rect 443184 28630 443236 28636
rect 444484 28234 444512 30124
rect 444392 28206 444512 28234
rect 441252 27328 441304 27334
rect 441252 27270 441304 27276
rect 438872 26206 439360 26234
rect 440344 26206 440648 26234
rect 436100 24744 436152 24750
rect 436100 24686 436152 24692
rect 438872 14929 438900 26206
rect 440344 16425 440372 26206
rect 440330 16416 440386 16425
rect 440330 16351 440386 16360
rect 438858 14920 438914 14929
rect 444392 14890 444420 28206
rect 445128 26234 445156 30124
rect 445772 28234 445800 30124
rect 447076 29866 447104 30124
rect 447060 29838 447104 29866
rect 445772 28206 445892 28234
rect 445760 28076 445812 28082
rect 445760 28018 445812 28024
rect 444484 26206 445156 26234
rect 444484 24818 444512 26206
rect 444472 24812 444524 24818
rect 444472 24754 444524 24760
rect 445772 22001 445800 28018
rect 445864 22953 445892 28206
rect 447060 28082 447088 29838
rect 448348 28082 448376 30124
rect 447048 28076 447100 28082
rect 447048 28018 447100 28024
rect 447140 28076 447192 28082
rect 447140 28018 447192 28024
rect 448336 28076 448388 28082
rect 448336 28018 448388 28024
rect 448520 28076 448572 28082
rect 448520 28018 448572 28024
rect 445850 22944 445906 22953
rect 445850 22879 445906 22888
rect 445758 21992 445814 22001
rect 445758 21927 445814 21936
rect 447152 15774 447180 28018
rect 448532 20233 448560 28018
rect 448992 26234 449020 30124
rect 449636 28082 449664 30124
rect 450940 29866 450968 30124
rect 449912 29838 450968 29866
rect 449624 28076 449676 28082
rect 449624 28018 449676 28024
rect 448624 26206 449020 26234
rect 448624 25401 448652 26206
rect 448610 25392 448666 25401
rect 448610 25327 448666 25336
rect 449912 22982 449940 29838
rect 451568 26234 451596 30124
rect 452856 28529 452884 30124
rect 459312 29918 459340 30124
rect 458180 29912 458232 29918
rect 458180 29854 458232 29860
rect 459300 29912 459352 29918
rect 459300 29854 459352 29860
rect 452842 28520 452898 28529
rect 452842 28455 452898 28464
rect 451924 28280 451976 28286
rect 451924 28222 451976 28228
rect 451292 26206 451596 26234
rect 451292 23050 451320 26206
rect 451280 23044 451332 23050
rect 451280 22986 451332 22992
rect 449900 22976 449952 22982
rect 449900 22918 449952 22924
rect 448518 20224 448574 20233
rect 448518 20159 448574 20168
rect 447140 15768 447192 15774
rect 447140 15710 447192 15716
rect 438858 14855 438914 14864
rect 444380 14884 444432 14890
rect 444380 14826 444432 14832
rect 434812 14340 434864 14346
rect 434812 14282 434864 14288
rect 451936 11626 451964 28222
rect 456800 22840 456852 22846
rect 456800 22782 456852 22788
rect 456812 16574 456840 22782
rect 458192 20602 458220 29854
rect 459940 26738 459968 30124
rect 459572 26710 459968 26738
rect 458180 20596 458232 20602
rect 458180 20538 458232 20544
rect 459572 19038 459600 26710
rect 460584 26234 460612 30124
rect 461228 28234 461256 30124
rect 459664 26206 460612 26234
rect 460952 28206 461256 28234
rect 459664 24721 459692 26206
rect 459650 24712 459706 24721
rect 459650 24647 459706 24656
rect 459560 19032 459612 19038
rect 459560 18974 459612 18980
rect 460952 17610 460980 28206
rect 461872 26234 461900 30124
rect 462516 26234 462544 30124
rect 463820 29866 463848 30124
rect 463804 29838 463848 29866
rect 463700 28280 463752 28286
rect 463700 28222 463752 28228
rect 461044 26206 461900 26234
rect 462332 26206 462544 26234
rect 461044 25362 461072 26206
rect 461032 25356 461084 25362
rect 461032 25298 461084 25304
rect 462332 19786 462360 26206
rect 462320 19780 462372 19786
rect 462320 19722 462372 19728
rect 463712 19106 463740 28222
rect 463804 20233 463832 29838
rect 464448 28286 464476 30124
rect 464436 28280 464488 28286
rect 464436 28222 464488 28228
rect 465092 28234 465120 30124
rect 465092 28206 465212 28234
rect 465080 28076 465132 28082
rect 465080 28018 465132 28024
rect 463790 20224 463846 20233
rect 463790 20159 463846 20168
rect 465092 19786 465120 28018
rect 465184 22001 465212 28206
rect 465736 26234 465764 30124
rect 466380 28082 466408 30124
rect 466368 28076 466420 28082
rect 466368 28018 466420 28024
rect 465276 26206 465764 26234
rect 465276 22710 465304 26206
rect 468956 23225 468984 30124
rect 468942 23216 468998 23225
rect 468942 23151 468998 23160
rect 465264 22704 465316 22710
rect 465264 22646 465316 22652
rect 469600 22094 469628 30124
rect 470888 27402 470916 30124
rect 470876 27396 470928 27402
rect 470876 27338 470928 27344
rect 473464 24857 473492 30124
rect 474004 28824 474056 28830
rect 474004 28766 474056 28772
rect 473450 24848 473506 24857
rect 473450 24783 473506 24792
rect 470600 24472 470652 24478
rect 470600 24414 470652 24420
rect 469232 22066 469628 22094
rect 465170 21992 465226 22001
rect 465170 21927 465226 21936
rect 465080 19780 465132 19786
rect 465080 19722 465132 19728
rect 463700 19100 463752 19106
rect 463700 19042 463752 19048
rect 466460 18556 466512 18562
rect 466460 18498 466512 18504
rect 460940 17604 460992 17610
rect 460940 17546 460992 17552
rect 466472 16574 466500 18498
rect 469232 18494 469260 22066
rect 469220 18488 469272 18494
rect 469220 18430 469272 18436
rect 456812 16546 456932 16574
rect 466472 16546 467512 16574
rect 453304 12980 453356 12986
rect 453304 12922 453356 12928
rect 451924 11620 451976 11626
rect 451924 11562 451976 11568
rect 434732 6886 435128 6914
rect 432052 6384 432104 6390
rect 432052 6326 432104 6332
rect 432064 480 432092 6326
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 6886
rect 446220 6792 446272 6798
rect 446220 6734 446272 6740
rect 439136 6724 439188 6730
rect 439136 6666 439188 6672
rect 439148 480 439176 6666
rect 442632 6452 442684 6458
rect 442632 6394 442684 6400
rect 442644 480 442672 6394
rect 446232 480 446260 6734
rect 449808 6520 449860 6526
rect 449808 6462 449860 6468
rect 449820 480 449848 6462
rect 453316 480 453344 12922
rect 456904 480 456932 16546
rect 463976 6860 464028 6866
rect 463976 6802 464028 6808
rect 460388 6588 460440 6594
rect 460388 6530 460440 6536
rect 460400 480 460428 6530
rect 463988 480 464016 6802
rect 467484 480 467512 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 24414
rect 474016 12918 474044 28766
rect 474752 28257 474780 30124
rect 476056 29866 476084 30124
rect 476040 29838 476084 29866
rect 474738 28248 474794 28257
rect 474738 28183 474794 28192
rect 476040 24682 476068 29838
rect 476684 29510 476712 30124
rect 476672 29504 476724 29510
rect 476672 29446 476724 29452
rect 477328 28286 477356 30124
rect 476120 28280 476172 28286
rect 476120 28222 476172 28228
rect 477316 28280 477368 28286
rect 477316 28222 477368 28228
rect 476132 24818 476160 28222
rect 478616 26234 478644 30124
rect 479260 26234 479288 30124
rect 480564 29866 480592 30124
rect 477512 26206 478644 26234
rect 478892 26206 479288 26234
rect 480272 29838 480592 29866
rect 476120 24812 476172 24818
rect 476120 24754 476172 24760
rect 476028 24676 476080 24682
rect 476028 24618 476080 24624
rect 477512 24614 477540 26206
rect 478892 26081 478920 26206
rect 478878 26072 478934 26081
rect 478878 26007 478934 26016
rect 479062 26072 479118 26081
rect 479062 26007 479118 26016
rect 479076 24954 479104 26007
rect 479064 24948 479116 24954
rect 479064 24890 479116 24896
rect 477500 24608 477552 24614
rect 477500 24550 477552 24556
rect 480272 20602 480300 29838
rect 481836 29442 481864 30124
rect 481824 29436 481876 29442
rect 481824 29378 481876 29384
rect 483124 26234 483152 30124
rect 484428 29866 484456 30124
rect 484428 29838 484624 29866
rect 484492 28280 484544 28286
rect 484492 28222 484544 28228
rect 484400 28076 484452 28082
rect 484400 28018 484452 28024
rect 483032 26206 483152 26234
rect 483032 22030 483060 26206
rect 483020 22024 483072 22030
rect 483020 21966 483072 21972
rect 480260 20596 480312 20602
rect 480260 20538 480312 20544
rect 474004 12912 474056 12918
rect 474004 12854 474056 12860
rect 484412 12345 484440 28018
rect 484504 24857 484532 28222
rect 484596 25265 484624 29838
rect 485056 28082 485084 30124
rect 485700 28286 485728 30124
rect 487632 28393 487660 30124
rect 487618 28384 487674 28393
rect 487618 28319 487674 28328
rect 485688 28280 485740 28286
rect 485688 28222 485740 28228
rect 485044 28076 485096 28082
rect 485044 28018 485096 28024
rect 489564 26234 489592 30124
rect 491496 27334 491524 30124
rect 492800 29866 492828 30124
rect 492692 29838 492828 29866
rect 491484 27328 491536 27334
rect 491484 27270 491536 27276
rect 485042 26208 485098 26217
rect 485042 26143 485098 26152
rect 488552 26206 489592 26234
rect 484582 25256 484638 25265
rect 484582 25191 484638 25200
rect 485056 24886 485084 26143
rect 485044 24880 485096 24886
rect 484490 24848 484546 24857
rect 485044 24822 485096 24828
rect 484490 24783 484546 24792
rect 488552 22098 488580 26206
rect 492692 26178 492720 29838
rect 493428 27538 493456 30124
rect 493416 27532 493468 27538
rect 493416 27474 493468 27480
rect 494072 26654 494100 30124
rect 494060 26648 494112 26654
rect 494060 26590 494112 26596
rect 499224 26234 499252 30124
rect 502444 28234 502472 30124
rect 502444 28206 502564 28234
rect 502432 28076 502484 28082
rect 502432 28018 502484 28024
rect 502340 27668 502392 27674
rect 502340 27610 502392 27616
rect 498212 26206 499252 26234
rect 492680 26172 492732 26178
rect 492680 26114 492732 26120
rect 498212 24070 498240 26206
rect 498200 24064 498252 24070
rect 498200 24006 498252 24012
rect 488540 22092 488592 22098
rect 488540 22034 488592 22040
rect 502352 16574 502380 27610
rect 502444 24002 502472 28018
rect 502536 25498 502564 28206
rect 503088 28082 503116 30124
rect 503076 28076 503128 28082
rect 503076 28018 503128 28024
rect 503168 28076 503220 28082
rect 503168 28018 503220 28024
rect 503180 27674 503208 28018
rect 503168 27668 503220 27674
rect 503168 27610 503220 27616
rect 504376 26234 504404 30124
rect 505680 29866 505708 30124
rect 505664 29838 505708 29866
rect 505664 28422 505692 29838
rect 505744 28552 505796 28558
rect 505744 28494 505796 28500
rect 505652 28416 505704 28422
rect 505652 28358 505704 28364
rect 505100 28280 505152 28286
rect 505100 28222 505152 28228
rect 503732 26206 504404 26234
rect 502524 25492 502576 25498
rect 502524 25434 502576 25440
rect 502432 23996 502484 24002
rect 502432 23938 502484 23944
rect 503732 20670 503760 26206
rect 503720 20664 503772 20670
rect 503720 20606 503772 20612
rect 504364 20664 504416 20670
rect 504364 20606 504416 20612
rect 504376 19854 504404 20606
rect 505112 20369 505140 28222
rect 505098 20360 505154 20369
rect 505098 20295 505154 20304
rect 504364 19848 504416 19854
rect 504364 19790 504416 19796
rect 502352 16546 503024 16574
rect 484398 12336 484454 12345
rect 484398 12271 484454 12280
rect 474556 6656 474608 6662
rect 474556 6598 474608 6604
rect 474568 480 474596 6598
rect 485226 6352 485282 6361
rect 485226 6287 485282 6296
rect 481732 6112 481784 6118
rect 481732 6054 481784 6060
rect 478144 4820 478196 4826
rect 478144 4762 478196 4768
rect 478156 480 478184 4762
rect 481744 480 481772 6054
rect 485240 480 485268 6287
rect 488816 6044 488868 6050
rect 488816 5986 488868 5992
rect 488828 480 488856 5986
rect 495900 4140 495952 4146
rect 495900 4082 495952 4088
rect 492312 4072 492364 4078
rect 492312 4014 492364 4020
rect 492324 480 492352 4014
rect 495912 480 495940 4082
rect 499396 3324 499448 3330
rect 499396 3266 499448 3272
rect 499408 480 499436 3266
rect 502996 480 503024 16546
rect 504376 10305 504404 19790
rect 505756 11558 505784 28494
rect 506308 28286 506336 30124
rect 506952 28558 506980 30124
rect 509544 29866 509572 30124
rect 509528 29838 509572 29866
rect 509528 29073 509556 29838
rect 509514 29064 509570 29073
rect 509514 28999 509570 29008
rect 506940 28552 506992 28558
rect 506940 28494 506992 28500
rect 506296 28280 506348 28286
rect 506296 28222 506348 28228
rect 510172 27402 510200 30124
rect 510712 27872 510764 27878
rect 510712 27814 510764 27820
rect 510160 27396 510212 27402
rect 510160 27338 510212 27344
rect 510724 21350 510752 27814
rect 510816 26761 510844 30124
rect 511460 27033 511488 30124
rect 512104 28830 512132 30124
rect 514052 29866 514080 30124
rect 514036 29838 514080 29866
rect 512092 28824 512144 28830
rect 512092 28766 512144 28772
rect 511446 27024 511502 27033
rect 511446 26959 511502 26968
rect 514036 26858 514064 29838
rect 515968 26926 515996 30124
rect 515956 26920 516008 26926
rect 515956 26862 516008 26868
rect 514024 26852 514076 26858
rect 514024 26794 514076 26800
rect 510802 26752 510858 26761
rect 510802 26687 510858 26696
rect 516612 26654 516640 30124
rect 517520 28348 517572 28354
rect 517520 28290 517572 28296
rect 516600 26648 516652 26654
rect 516600 26590 516652 26596
rect 513380 25900 513432 25906
rect 513380 25842 513432 25848
rect 510712 21344 510764 21350
rect 510712 21286 510764 21292
rect 505744 11552 505796 11558
rect 505744 11494 505796 11500
rect 504362 10296 504418 10305
rect 504362 10231 504418 10240
rect 506478 3904 506534 3913
rect 506478 3839 506534 3848
rect 506492 480 506520 3839
rect 510068 3392 510120 3398
rect 510068 3334 510120 3340
rect 510080 480 510108 3334
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 25842
rect 516140 25832 516192 25838
rect 516140 25774 516192 25780
rect 516152 16574 516180 25774
rect 517532 23458 517560 28290
rect 519188 28286 519216 30124
rect 519832 29481 519860 30124
rect 519818 29472 519874 29481
rect 519818 29407 519874 29416
rect 519176 28280 519228 28286
rect 519176 28222 519228 28228
rect 520476 26722 520504 30124
rect 521120 29782 521148 30124
rect 521108 29776 521160 29782
rect 521108 29718 521160 29724
rect 523052 29578 523080 30124
rect 523040 29572 523092 29578
rect 523040 29514 523092 29520
rect 523696 26790 523724 30124
rect 523684 26784 523736 26790
rect 523684 26726 523736 26732
rect 520464 26716 520516 26722
rect 520464 26658 520516 26664
rect 524340 26625 524368 30124
rect 524880 28756 524932 28762
rect 524880 28698 524932 28704
rect 524326 26616 524382 26625
rect 524326 26551 524382 26560
rect 520280 25968 520332 25974
rect 520280 25910 520332 25916
rect 517520 23452 517572 23458
rect 517520 23394 517572 23400
rect 516152 16546 517192 16574
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 25910
rect 524892 20670 524920 28698
rect 525628 27577 525656 30124
rect 526932 29918 526960 30124
rect 525800 29912 525852 29918
rect 525800 29854 525852 29860
rect 526920 29912 526972 29918
rect 526920 29854 526972 29860
rect 525614 27568 525670 27577
rect 525614 27503 525670 27512
rect 524880 20664 524932 20670
rect 524880 20606 524932 20612
rect 525812 20505 525840 29854
rect 528204 29510 528232 30124
rect 525892 29504 525944 29510
rect 525892 29446 525944 29452
rect 528192 29504 528244 29510
rect 528192 29446 528244 29452
rect 525904 28762 525932 29446
rect 527824 28892 527876 28898
rect 527824 28834 527876 28840
rect 525892 28756 525944 28762
rect 525892 28698 525944 28704
rect 525798 20496 525854 20505
rect 525798 20431 525854 20440
rect 526442 20360 526498 20369
rect 526442 20295 526498 20304
rect 522304 15700 522356 15706
rect 522304 15642 522356 15648
rect 522316 3806 522344 15642
rect 526456 4010 526484 20295
rect 527836 17542 527864 28834
rect 528848 26234 528876 30124
rect 529492 28354 529520 30124
rect 529940 28620 529992 28626
rect 529940 28562 529992 28568
rect 529480 28348 529532 28354
rect 529480 28290 529532 28296
rect 528572 26206 528876 26234
rect 528572 21962 528600 26206
rect 529952 23322 529980 28562
rect 531424 27606 531452 30124
rect 532068 28626 532096 30124
rect 536576 28966 536604 30124
rect 536564 28960 536616 28966
rect 536564 28902 536616 28908
rect 537220 28898 537248 30124
rect 537864 29617 537892 30124
rect 539168 29866 539196 30124
rect 538324 29838 539196 29866
rect 537850 29608 537906 29617
rect 537850 29543 537906 29552
rect 537208 28892 537260 28898
rect 537208 28834 537260 28840
rect 532056 28620 532108 28626
rect 532056 28562 532108 28568
rect 535460 28484 535512 28490
rect 535460 28426 535512 28432
rect 531412 27600 531464 27606
rect 531412 27542 531464 27548
rect 535472 27470 535500 28426
rect 536104 28212 536156 28218
rect 536104 28154 536156 28160
rect 535460 27464 535512 27470
rect 535460 27406 535512 27412
rect 536116 26246 536144 28154
rect 536104 26240 536156 26246
rect 536104 26182 536156 26188
rect 538220 25424 538272 25430
rect 538220 25366 538272 25372
rect 529940 23316 529992 23322
rect 529940 23258 529992 23264
rect 528560 21956 528612 21962
rect 528560 21898 528612 21904
rect 533344 18420 533396 18426
rect 533344 18362 533396 18368
rect 527824 17536 527876 17542
rect 527824 17478 527876 17484
rect 527824 5976 527876 5982
rect 527824 5918 527876 5924
rect 526444 4004 526496 4010
rect 526444 3946 526496 3952
rect 522304 3800 522356 3806
rect 522304 3742 522356 3748
rect 524236 3800 524288 3806
rect 524236 3742 524288 3748
rect 524248 480 524276 3742
rect 527836 480 527864 5918
rect 531318 4040 531374 4049
rect 531318 3975 531374 3984
rect 531332 480 531360 3975
rect 533356 3942 533384 18362
rect 533344 3936 533396 3942
rect 533344 3878 533396 3884
rect 534908 3936 534960 3942
rect 534908 3878 534960 3884
rect 534920 480 534948 3878
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 25366
rect 538324 20641 538352 29838
rect 539980 24614 540008 159326
rect 540072 147801 540100 233106
rect 540244 232688 540296 232694
rect 540244 232630 540296 232636
rect 540152 150476 540204 150482
rect 540152 150418 540204 150424
rect 540058 147792 540114 147801
rect 540058 147727 540114 147736
rect 540164 147674 540192 150418
rect 540072 147646 540192 147674
rect 540072 143449 540100 147646
rect 540150 147384 540206 147393
rect 540150 147319 540206 147328
rect 540058 143440 540114 143449
rect 540058 143375 540114 143384
rect 540164 142154 540192 147319
rect 540072 142126 540192 142154
rect 539968 24608 540020 24614
rect 539968 24550 540020 24556
rect 538310 20632 538366 20641
rect 538310 20567 538366 20576
rect 540072 15094 540100 142126
rect 540256 134094 540284 232630
rect 540244 134088 540296 134094
rect 540244 134030 540296 134036
rect 540244 129872 540296 129878
rect 540244 129814 540296 129820
rect 540060 15088 540112 15094
rect 540060 15030 540112 15036
rect 540256 11626 540284 129814
rect 540348 129062 540376 234330
rect 540440 152386 540468 238002
rect 542084 237516 542136 237522
rect 542084 237458 542136 237464
rect 541072 235272 541124 235278
rect 541072 235214 541124 235220
rect 540704 163600 540756 163606
rect 540704 163542 540756 163548
rect 540520 158636 540572 158642
rect 540520 158578 540572 158584
rect 540428 152380 540480 152386
rect 540428 152322 540480 152328
rect 540428 150340 540480 150346
rect 540428 150282 540480 150288
rect 540440 133210 540468 150282
rect 540428 133204 540480 133210
rect 540428 133146 540480 133152
rect 540336 129056 540388 129062
rect 540336 128998 540388 129004
rect 540336 125860 540388 125866
rect 540336 125802 540388 125808
rect 540348 13666 540376 125802
rect 540428 125316 540480 125322
rect 540428 125258 540480 125264
rect 540440 112062 540468 125258
rect 540532 116006 540560 158578
rect 540612 158432 540664 158438
rect 540612 158374 540664 158380
rect 540624 133958 540652 158374
rect 540716 150414 540744 163542
rect 540980 151700 541032 151706
rect 540980 151642 541032 151648
rect 540888 150884 540940 150890
rect 540888 150826 540940 150832
rect 540704 150408 540756 150414
rect 540704 150350 540756 150356
rect 540704 149864 540756 149870
rect 540704 149806 540756 149812
rect 540716 149705 540744 149806
rect 540702 149696 540758 149705
rect 540702 149631 540758 149640
rect 540900 149546 540928 150826
rect 540716 149518 540928 149546
rect 540716 147626 540744 149518
rect 540704 147620 540756 147626
rect 540704 147562 540756 147568
rect 540888 146940 540940 146946
rect 540888 146882 540940 146888
rect 540900 144914 540928 146882
rect 540992 145489 541020 151642
rect 540978 145480 541034 145489
rect 540978 145415 541034 145424
rect 540900 144886 541020 144914
rect 540612 133952 540664 133958
rect 540992 133906 541020 144886
rect 540612 133894 540664 133900
rect 540808 133878 541020 133906
rect 540808 126818 540836 133878
rect 541084 133521 541112 235214
rect 541624 233776 541676 233782
rect 541624 233718 541676 233724
rect 541256 163668 541308 163674
rect 541256 163610 541308 163616
rect 541164 156800 541216 156806
rect 541164 156742 541216 156748
rect 541070 133512 541126 133521
rect 541070 133447 541126 133456
rect 540886 133240 540942 133249
rect 540886 133175 540942 133184
rect 540980 133204 541032 133210
rect 540900 129742 540928 133175
rect 540980 133146 541032 133152
rect 540888 129736 540940 129742
rect 540992 129713 541020 133146
rect 541072 131096 541124 131102
rect 541072 131038 541124 131044
rect 540888 129678 540940 129684
rect 540978 129704 541034 129713
rect 540978 129639 541034 129648
rect 541084 128354 541112 131038
rect 540900 128326 541112 128354
rect 540796 126812 540848 126818
rect 540796 126754 540848 126760
rect 540796 126268 540848 126274
rect 540796 126210 540848 126216
rect 540704 121508 540756 121514
rect 540704 121450 540756 121456
rect 540520 116000 540572 116006
rect 540520 115942 540572 115948
rect 540610 115968 540666 115977
rect 540610 115903 540666 115912
rect 540428 112056 540480 112062
rect 540428 111998 540480 112004
rect 540428 110492 540480 110498
rect 540428 110434 540480 110440
rect 540440 26994 540468 110434
rect 540624 95198 540652 115903
rect 540716 108866 540744 121450
rect 540808 109614 540836 126210
rect 540900 125458 540928 128326
rect 540888 125452 540940 125458
rect 540888 125394 540940 125400
rect 541072 116000 541124 116006
rect 541072 115942 541124 115948
rect 540888 109948 540940 109954
rect 540888 109890 540940 109896
rect 540796 109608 540848 109614
rect 540796 109550 540848 109556
rect 540704 108860 540756 108866
rect 540704 108802 540756 108808
rect 540794 99512 540850 99521
rect 540900 99498 540928 109890
rect 540900 99470 541020 99498
rect 540794 99447 540850 99456
rect 540612 95192 540664 95198
rect 540612 95134 540664 95140
rect 540808 84194 540836 99447
rect 540992 96626 541020 99470
rect 540980 96620 541032 96626
rect 540980 96562 541032 96568
rect 541084 95169 541112 115942
rect 541176 101561 541204 156742
rect 541162 101552 541218 101561
rect 541162 101487 541218 101496
rect 541070 95160 541126 95169
rect 541070 95095 541126 95104
rect 540808 84166 541112 84194
rect 540612 82136 540664 82142
rect 540612 82078 540664 82084
rect 540520 75200 540572 75206
rect 540520 75142 540572 75148
rect 540428 26988 540480 26994
rect 540428 26930 540480 26936
rect 540336 13660 540388 13666
rect 540336 13602 540388 13608
rect 540532 12238 540560 75142
rect 540624 23458 540652 82078
rect 540704 31068 540756 31074
rect 540704 31010 540756 31016
rect 540716 25362 540744 31010
rect 540704 25356 540756 25362
rect 540704 25298 540756 25304
rect 540612 23452 540664 23458
rect 540612 23394 540664 23400
rect 540520 12232 540572 12238
rect 540520 12174 540572 12180
rect 540244 11620 540296 11626
rect 540244 11562 540296 11568
rect 541084 6730 541112 84166
rect 541268 43761 541296 163610
rect 541348 144900 541400 144906
rect 541348 144842 541400 144848
rect 541360 131170 541388 144842
rect 541530 141808 541586 141817
rect 541530 141743 541586 141752
rect 541440 133952 541492 133958
rect 541440 133894 541492 133900
rect 541348 131164 541400 131170
rect 541348 131106 541400 131112
rect 541348 130348 541400 130354
rect 541348 130290 541400 130296
rect 541360 125662 541388 130290
rect 541348 125656 541400 125662
rect 541348 125598 541400 125604
rect 541348 123956 541400 123962
rect 541348 123898 541400 123904
rect 541360 88330 541388 123898
rect 541452 109954 541480 133894
rect 541544 131102 541572 141743
rect 541636 136649 541664 233718
rect 541716 233028 541768 233034
rect 541716 232970 541768 232976
rect 541728 144430 541756 232970
rect 541900 232552 541952 232558
rect 541900 232494 541952 232500
rect 541808 228812 541860 228818
rect 541808 228754 541860 228760
rect 541716 144424 541768 144430
rect 541716 144366 541768 144372
rect 541820 140826 541848 228754
rect 541912 148306 541940 232494
rect 541992 207120 542044 207126
rect 541992 207062 542044 207068
rect 541900 148300 541952 148306
rect 541900 148242 541952 148248
rect 541898 147656 541954 147665
rect 541898 147591 541954 147600
rect 541808 140820 541860 140826
rect 541808 140762 541860 140768
rect 541622 136640 541678 136649
rect 541622 136575 541678 136584
rect 541716 134088 541768 134094
rect 541716 134030 541768 134036
rect 541624 134020 541676 134026
rect 541624 133962 541676 133968
rect 541532 131096 541584 131102
rect 541532 131038 541584 131044
rect 541636 125866 541664 133962
rect 541728 130898 541756 134030
rect 541806 133104 541862 133113
rect 541806 133039 541862 133048
rect 541716 130892 541768 130898
rect 541716 130834 541768 130840
rect 541716 130756 541768 130762
rect 541716 130698 541768 130704
rect 541624 125860 541676 125866
rect 541624 125802 541676 125808
rect 541728 125746 541756 130698
rect 541820 130422 541848 133039
rect 541912 132530 541940 147591
rect 542004 135182 542032 207062
rect 542096 198966 542124 237458
rect 542084 198960 542136 198966
rect 542084 198902 542136 198908
rect 542372 197305 542400 240094
rect 544212 238754 544240 240094
rect 543936 238726 544240 238754
rect 543094 236600 543150 236609
rect 543094 236535 543150 236544
rect 542452 232892 542504 232898
rect 542452 232834 542504 232840
rect 542358 197296 542414 197305
rect 542358 197231 542414 197240
rect 542464 157334 542492 232834
rect 543004 230512 543056 230518
rect 543004 230454 543056 230460
rect 542544 213240 542596 213246
rect 542544 213182 542596 213188
rect 542372 157306 542492 157334
rect 542176 150408 542228 150414
rect 542176 150350 542228 150356
rect 542188 147014 542216 150350
rect 542268 147620 542320 147626
rect 542268 147562 542320 147568
rect 542176 147008 542228 147014
rect 542176 146950 542228 146956
rect 542280 144786 542308 147562
rect 542372 144906 542400 157306
rect 542452 154284 542504 154290
rect 542452 154226 542504 154232
rect 542360 144900 542412 144906
rect 542360 144842 542412 144848
rect 542280 144758 542400 144786
rect 542268 144560 542320 144566
rect 542268 144502 542320 144508
rect 542280 138014 542308 144502
rect 542188 137986 542308 138014
rect 541992 135176 542044 135182
rect 541992 135118 542044 135124
rect 542084 132796 542136 132802
rect 542084 132738 542136 132744
rect 541992 132660 542044 132666
rect 541992 132602 542044 132608
rect 541900 132524 541952 132530
rect 541900 132466 541952 132472
rect 542004 130506 542032 132602
rect 541912 130478 542032 130506
rect 541808 130416 541860 130422
rect 541808 130358 541860 130364
rect 541808 129736 541860 129742
rect 541808 129678 541860 129684
rect 541820 127673 541848 129678
rect 541806 127664 541862 127673
rect 541912 127634 541940 130478
rect 541992 130416 542044 130422
rect 541992 130358 542044 130364
rect 541806 127599 541862 127608
rect 541900 127628 541952 127634
rect 541900 127570 541952 127576
rect 542004 127514 542032 130358
rect 541636 125718 541756 125746
rect 541820 127486 542032 127514
rect 541440 109948 541492 109954
rect 541440 109890 541492 109896
rect 541530 102232 541586 102241
rect 541530 102167 541586 102176
rect 541348 88324 541400 88330
rect 541348 88266 541400 88272
rect 541544 82929 541572 102167
rect 541530 82920 541586 82929
rect 541440 82884 541492 82890
rect 541530 82855 541586 82864
rect 541440 82826 541492 82832
rect 541254 43752 541310 43761
rect 541254 43687 541310 43696
rect 541452 16454 541480 82826
rect 541440 16448 541492 16454
rect 541440 16390 541492 16396
rect 541636 13530 541664 125718
rect 541716 125656 541768 125662
rect 541716 125598 541768 125604
rect 541728 115841 541756 125598
rect 541820 115977 541848 127486
rect 541992 127424 542044 127430
rect 541992 127366 542044 127372
rect 542004 126698 542032 127366
rect 542096 126868 542124 132738
rect 542188 131034 542216 137986
rect 542268 135312 542320 135318
rect 542268 135254 542320 135260
rect 542176 131028 542228 131034
rect 542176 130970 542228 130976
rect 542176 130892 542228 130898
rect 542176 130834 542228 130840
rect 542188 126970 542216 130834
rect 542280 129130 542308 135254
rect 542268 129124 542320 129130
rect 542268 129066 542320 129072
rect 542188 126942 542308 126970
rect 542096 126840 542216 126868
rect 542004 126670 542124 126698
rect 541992 124024 542044 124030
rect 541992 123966 542044 123972
rect 542004 121514 542032 123966
rect 541992 121508 542044 121514
rect 541992 121450 542044 121456
rect 541806 115968 541862 115977
rect 541806 115903 541862 115912
rect 541714 115832 541770 115841
rect 542096 115802 542124 126670
rect 541714 115767 541770 115776
rect 542084 115796 542136 115802
rect 542084 115738 542136 115744
rect 541808 111852 541860 111858
rect 541808 111794 541860 111800
rect 541716 110560 541768 110566
rect 541716 110502 541768 110508
rect 541624 13524 541676 13530
rect 541624 13466 541676 13472
rect 541728 12170 541756 110502
rect 541820 14278 541848 111794
rect 541900 106956 541952 106962
rect 541900 106898 541952 106904
rect 541912 17338 541940 106898
rect 542188 102678 542216 126840
rect 542280 113218 542308 126942
rect 542268 113212 542320 113218
rect 542268 113154 542320 113160
rect 542268 110356 542320 110362
rect 542268 110298 542320 110304
rect 542280 106214 542308 110298
rect 542268 106208 542320 106214
rect 542268 106150 542320 106156
rect 542176 102672 542228 102678
rect 542176 102614 542228 102620
rect 542084 100020 542136 100026
rect 542084 99962 542136 99968
rect 541992 92676 542044 92682
rect 541992 92618 542044 92624
rect 541900 17332 541952 17338
rect 541900 17274 541952 17280
rect 542004 14686 542032 92618
rect 542096 82618 542124 99962
rect 542176 95940 542228 95946
rect 542176 95882 542228 95888
rect 542188 84998 542216 95882
rect 542268 95192 542320 95198
rect 542268 95134 542320 95140
rect 542280 92546 542308 95134
rect 542268 92540 542320 92546
rect 542268 92482 542320 92488
rect 542268 88256 542320 88262
rect 542268 88198 542320 88204
rect 542176 84992 542228 84998
rect 542176 84934 542228 84940
rect 542280 84194 542308 88198
rect 542188 84166 542308 84194
rect 542084 82612 542136 82618
rect 542084 82554 542136 82560
rect 542188 21350 542216 84166
rect 542268 69284 542320 69290
rect 542268 69226 542320 69232
rect 542176 21344 542228 21350
rect 542176 21286 542228 21292
rect 542280 14754 542308 69226
rect 542268 14748 542320 14754
rect 542268 14690 542320 14696
rect 541992 14680 542044 14686
rect 541992 14622 542044 14628
rect 541808 14272 541860 14278
rect 541808 14214 541860 14220
rect 541716 12164 541768 12170
rect 541716 12106 541768 12112
rect 542372 11694 542400 144758
rect 542464 136678 542492 154226
rect 542556 145761 542584 213182
rect 542728 154556 542780 154562
rect 542728 154498 542780 154504
rect 542636 154488 542688 154494
rect 542636 154430 542688 154436
rect 542542 145752 542598 145761
rect 542542 145687 542598 145696
rect 542544 143472 542596 143478
rect 542544 143414 542596 143420
rect 542452 136672 542504 136678
rect 542452 136614 542504 136620
rect 542452 136536 542504 136542
rect 542452 136478 542504 136484
rect 542464 136241 542492 136478
rect 542450 136232 542506 136241
rect 542450 136167 542506 136176
rect 542452 135244 542504 135250
rect 542452 135186 542504 135192
rect 542464 134201 542492 135186
rect 542450 134192 542506 134201
rect 542450 134127 542506 134136
rect 542452 132456 542504 132462
rect 542452 132398 542504 132404
rect 542464 131481 542492 132398
rect 542450 131472 542506 131481
rect 542450 131407 542506 131416
rect 542452 131096 542504 131102
rect 542452 131038 542504 131044
rect 542464 130801 542492 131038
rect 542450 130792 542506 130801
rect 542450 130727 542506 130736
rect 542452 129736 542504 129742
rect 542452 129678 542504 129684
rect 542464 129441 542492 129678
rect 542450 129432 542506 129441
rect 542450 129367 542506 129376
rect 542556 125594 542584 143414
rect 542544 125588 542596 125594
rect 542544 125530 542596 125536
rect 542452 125384 542504 125390
rect 542450 125352 542452 125361
rect 542504 125352 542506 125361
rect 542450 125287 542506 125296
rect 542452 117292 542504 117298
rect 542452 117234 542504 117240
rect 542464 116521 542492 117234
rect 542450 116512 542506 116521
rect 542450 116447 542506 116456
rect 542450 113792 542506 113801
rect 542450 113727 542506 113736
rect 542464 113626 542492 113727
rect 542452 113620 542504 113626
rect 542452 113562 542504 113568
rect 542452 110424 542504 110430
rect 542452 110366 542504 110372
rect 542542 110392 542598 110401
rect 542464 109721 542492 110366
rect 542542 110327 542598 110336
rect 542450 109712 542506 109721
rect 542450 109647 542506 109656
rect 542452 109608 542504 109614
rect 542452 109550 542504 109556
rect 542464 92682 542492 109550
rect 542556 109478 542584 110327
rect 542544 109472 542596 109478
rect 542544 109414 542596 109420
rect 542648 109410 542676 154430
rect 542740 117162 542768 154498
rect 542912 147008 542964 147014
rect 542912 146950 542964 146956
rect 542820 146260 542872 146266
rect 542820 146202 542872 146208
rect 542832 140078 542860 146202
rect 542924 143410 542952 146950
rect 543016 144226 543044 230454
rect 543108 152862 543136 236535
rect 543554 231432 543610 231441
rect 543554 231367 543610 231376
rect 543188 228880 543240 228886
rect 543188 228822 543240 228828
rect 543200 171134 543228 228822
rect 543200 171106 543320 171134
rect 543096 152856 543148 152862
rect 543096 152798 543148 152804
rect 543188 150000 543240 150006
rect 543188 149942 543240 149948
rect 543004 144220 543056 144226
rect 543004 144162 543056 144168
rect 543096 144084 543148 144090
rect 543096 144026 543148 144032
rect 542912 143404 542964 143410
rect 542912 143346 542964 143352
rect 542912 141704 542964 141710
rect 542910 141672 542912 141681
rect 542964 141672 542966 141681
rect 542910 141607 542966 141616
rect 542820 140072 542872 140078
rect 542820 140014 542872 140020
rect 542912 136672 542964 136678
rect 542912 136614 542964 136620
rect 542820 136604 542872 136610
rect 542820 136546 542872 136552
rect 542832 135561 542860 136546
rect 542818 135552 542874 135561
rect 542818 135487 542874 135496
rect 542820 132524 542872 132530
rect 542820 132466 542872 132472
rect 542728 117156 542780 117162
rect 542728 117098 542780 117104
rect 542728 114844 542780 114850
rect 542728 114786 542780 114792
rect 542636 109404 542688 109410
rect 542636 109346 542688 109352
rect 542740 109154 542768 114786
rect 542556 109126 542768 109154
rect 542452 92676 542504 92682
rect 542452 92618 542504 92624
rect 542452 92540 542504 92546
rect 542452 92482 542504 92488
rect 542464 82890 542492 92482
rect 542452 82884 542504 82890
rect 542452 82826 542504 82832
rect 542556 30705 542584 109126
rect 542636 109064 542688 109070
rect 542636 109006 542688 109012
rect 542648 107681 542676 109006
rect 542634 107672 542690 107681
rect 542634 107607 542690 107616
rect 542832 92274 542860 132466
rect 542924 129577 542952 136614
rect 542910 129568 542966 129577
rect 542910 129503 542966 129512
rect 543108 126274 543136 144026
rect 543200 142154 543228 149942
rect 543292 146130 543320 171106
rect 543372 152380 543424 152386
rect 543372 152322 543424 152328
rect 543280 146124 543332 146130
rect 543280 146066 543332 146072
rect 543280 143540 543332 143546
rect 543280 143482 543332 143488
rect 543292 142361 543320 143482
rect 543384 142594 543412 152322
rect 543568 149734 543596 231367
rect 543936 229906 543964 238726
rect 544384 234116 544436 234122
rect 544384 234058 544436 234064
rect 544106 233880 544162 233889
rect 544106 233815 544162 233824
rect 544016 231736 544068 231742
rect 544016 231678 544068 231684
rect 543924 229900 543976 229906
rect 543924 229842 543976 229848
rect 543924 229764 543976 229770
rect 543924 229706 543976 229712
rect 543832 152788 543884 152794
rect 543832 152730 543884 152736
rect 543740 151632 543792 151638
rect 543740 151574 543792 151580
rect 543556 149728 543608 149734
rect 543556 149670 543608 149676
rect 543646 149696 543702 149705
rect 543646 149631 543702 149640
rect 543464 147620 543516 147626
rect 543464 147562 543516 147568
rect 543476 146441 543504 147562
rect 543462 146432 543518 146441
rect 543462 146367 543518 146376
rect 543372 142588 543424 142594
rect 543372 142530 543424 142536
rect 543464 142384 543516 142390
rect 543278 142352 543334 142361
rect 543464 142326 543516 142332
rect 543278 142287 543334 142296
rect 543200 142126 543320 142154
rect 543096 126268 543148 126274
rect 543096 126210 543148 126216
rect 543292 125594 543320 142126
rect 543372 139460 543424 139466
rect 543372 139402 543424 139408
rect 542924 125566 543320 125594
rect 542924 110362 542952 125566
rect 543004 120760 543056 120766
rect 543004 120702 543056 120708
rect 543016 115934 543044 120702
rect 543016 115906 543136 115934
rect 543108 115818 543136 115906
rect 543016 115790 543136 115818
rect 543280 115864 543332 115870
rect 543280 115806 543332 115812
rect 543016 110362 543044 115790
rect 543096 113824 543148 113830
rect 543096 113766 543148 113772
rect 542912 110356 542964 110362
rect 542912 110298 542964 110304
rect 543004 110356 543056 110362
rect 543004 110298 543056 110304
rect 543108 108338 543136 113766
rect 543292 112690 543320 115806
rect 543384 113898 543412 139402
rect 543476 138122 543504 142326
rect 543660 142154 543688 149631
rect 543752 143478 543780 151574
rect 543844 146266 543872 152730
rect 543832 146260 543884 146266
rect 543832 146202 543884 146208
rect 543740 143472 543792 143478
rect 543740 143414 543792 143420
rect 543660 142126 543780 142154
rect 543556 142112 543608 142118
rect 543556 142054 543608 142060
rect 543568 141001 543596 142054
rect 543554 140992 543610 141001
rect 543554 140927 543610 140936
rect 543556 139392 543608 139398
rect 543556 139334 543608 139340
rect 543568 138281 543596 139334
rect 543554 138272 543610 138281
rect 543554 138207 543610 138216
rect 543476 138094 543688 138122
rect 543660 134298 543688 138094
rect 543648 134292 543700 134298
rect 543648 134234 543700 134240
rect 543752 134178 543780 142126
rect 543660 134150 543780 134178
rect 543464 131028 543516 131034
rect 543464 130970 543516 130976
rect 543372 113892 543424 113898
rect 543372 113834 543424 113840
rect 543292 112662 543412 112690
rect 543188 111104 543240 111110
rect 543188 111046 543240 111052
rect 543016 108310 543136 108338
rect 542820 92268 542872 92274
rect 542820 92210 542872 92216
rect 542636 92200 542688 92206
rect 542636 92142 542688 92148
rect 542648 91361 542676 92142
rect 542634 91352 542690 91361
rect 542634 91287 542690 91296
rect 542820 91180 542872 91186
rect 542820 91122 542872 91128
rect 542728 89684 542780 89690
rect 542728 89626 542780 89632
rect 542740 88641 542768 89626
rect 542726 88632 542782 88641
rect 542726 88567 542782 88576
rect 542636 85128 542688 85134
rect 542636 85070 542688 85076
rect 542648 84561 542676 85070
rect 542634 84552 542690 84561
rect 542634 84487 542690 84496
rect 542832 82890 542860 91122
rect 542820 82884 542872 82890
rect 542820 82826 542872 82832
rect 542636 75744 542688 75750
rect 542634 75712 542636 75721
rect 542688 75712 542690 75721
rect 542634 75647 542690 75656
rect 542820 66224 542872 66230
rect 542820 66166 542872 66172
rect 542832 65521 542860 66166
rect 542818 65512 542874 65521
rect 542818 65447 542874 65456
rect 542728 53780 542780 53786
rect 542728 53722 542780 53728
rect 542740 52601 542768 53722
rect 542726 52592 542782 52601
rect 542726 52527 542782 52536
rect 542728 51060 542780 51066
rect 542728 51002 542780 51008
rect 542740 49881 542768 51002
rect 542726 49872 542782 49881
rect 542726 49807 542782 49816
rect 542728 49700 542780 49706
rect 542728 49642 542780 49648
rect 542740 48521 542768 49642
rect 542726 48512 542782 48521
rect 542726 48447 542782 48456
rect 542542 30696 542598 30705
rect 542542 30631 542598 30640
rect 543016 13598 543044 108310
rect 543200 107794 543228 111046
rect 543280 109064 543332 109070
rect 543280 109006 543332 109012
rect 543108 107766 543228 107794
rect 543004 13592 543056 13598
rect 543004 13534 543056 13540
rect 543108 12374 543136 107766
rect 543188 107636 543240 107642
rect 543188 107578 543240 107584
rect 543200 106321 543228 107578
rect 543186 106312 543242 106321
rect 543186 106247 543242 106256
rect 543188 105596 543240 105602
rect 543188 105538 543240 105544
rect 543200 14414 543228 105538
rect 543292 104802 543320 109006
rect 543384 104922 543412 112662
rect 543372 104916 543424 104922
rect 543372 104858 543424 104864
rect 543292 104774 543412 104802
rect 543280 103624 543332 103630
rect 543280 103566 543332 103572
rect 543292 18426 543320 103566
rect 543384 69290 543412 104774
rect 543476 102202 543504 130970
rect 543660 130762 543688 134150
rect 543740 131164 543792 131170
rect 543740 131106 543792 131112
rect 543648 130756 543700 130762
rect 543648 130698 543700 130704
rect 543556 128308 543608 128314
rect 543556 128250 543608 128256
rect 543568 128081 543596 128250
rect 543554 128072 543610 128081
rect 543554 128007 543610 128016
rect 543648 126948 543700 126954
rect 543648 126890 543700 126896
rect 543556 125520 543608 125526
rect 543556 125462 543608 125468
rect 543568 124681 543596 125462
rect 543554 124672 543610 124681
rect 543554 124607 543610 124616
rect 543660 124522 543688 126890
rect 543568 124494 543688 124522
rect 543568 121530 543596 124494
rect 543752 123962 543780 131106
rect 543832 127696 543884 127702
rect 543832 127638 543884 127644
rect 543844 125322 543872 127638
rect 543832 125316 543884 125322
rect 543832 125258 543884 125264
rect 543740 123956 543792 123962
rect 543740 123898 543792 123904
rect 543648 122800 543700 122806
rect 543648 122742 543700 122748
rect 543660 121961 543688 122742
rect 543646 121952 543702 121961
rect 543646 121887 543702 121896
rect 543568 121502 543688 121530
rect 543556 121440 543608 121446
rect 543556 121382 543608 121388
rect 543568 120601 543596 121382
rect 543554 120592 543610 120601
rect 543554 120527 543610 120536
rect 543660 118674 543688 121502
rect 543660 118646 543780 118674
rect 543554 118008 543610 118017
rect 543554 117943 543610 117952
rect 543568 110537 543596 117943
rect 543648 117360 543700 117366
rect 543648 117302 543700 117308
rect 543660 113150 543688 117302
rect 543648 113144 543700 113150
rect 543648 113086 543700 113092
rect 543752 111858 543780 118646
rect 543740 111852 543792 111858
rect 543740 111794 543792 111800
rect 543554 110528 543610 110537
rect 543554 110463 543610 110472
rect 543660 110486 543780 110514
rect 543660 110362 543688 110486
rect 543648 110356 543700 110362
rect 543648 110298 543700 110304
rect 543752 110294 543780 110486
rect 543740 110288 543792 110294
rect 543740 110230 543792 110236
rect 543648 108860 543700 108866
rect 543648 108802 543700 108808
rect 543660 107522 543688 108802
rect 543660 107494 543780 107522
rect 543752 104650 543780 107494
rect 543740 104644 543792 104650
rect 543740 104586 543792 104592
rect 543464 102196 543516 102202
rect 543464 102138 543516 102144
rect 543556 97980 543608 97986
rect 543556 97922 543608 97928
rect 543568 97481 543596 97922
rect 543554 97472 543610 97481
rect 543554 97407 543610 97416
rect 543464 96620 543516 96626
rect 543464 96562 543516 96568
rect 543648 96620 543700 96626
rect 543648 96562 543700 96568
rect 543476 89842 543504 96562
rect 543556 96552 543608 96558
rect 543556 96494 543608 96500
rect 543568 96121 543596 96494
rect 543554 96112 543610 96121
rect 543554 96047 543610 96056
rect 543660 95441 543688 96562
rect 543646 95432 543702 95441
rect 543646 95367 543702 95376
rect 543556 95192 543608 95198
rect 543556 95134 543608 95140
rect 543568 94081 543596 95134
rect 543554 94072 543610 94081
rect 543554 94007 543610 94016
rect 543556 93832 543608 93838
rect 543556 93774 543608 93780
rect 543568 92721 543596 93774
rect 543554 92712 543610 92721
rect 543554 92647 543610 92656
rect 543556 92472 543608 92478
rect 543556 92414 543608 92420
rect 543568 92041 543596 92414
rect 543554 92032 543610 92041
rect 543554 91967 543610 91976
rect 543476 89814 543780 89842
rect 543648 89752 543700 89758
rect 543648 89694 543700 89700
rect 543660 85542 543688 89694
rect 543648 85536 543700 85542
rect 543648 85478 543700 85484
rect 543464 83020 543516 83026
rect 543464 82962 543516 82968
rect 543372 69284 543424 69290
rect 543372 69226 543424 69232
rect 543280 18420 543332 18426
rect 543280 18362 543332 18368
rect 543188 14408 543240 14414
rect 543188 14350 543240 14356
rect 543096 12368 543148 12374
rect 543096 12310 543148 12316
rect 543476 12102 543504 82962
rect 543648 82952 543700 82958
rect 543648 82894 543700 82900
rect 543556 82816 543608 82822
rect 543556 82758 543608 82764
rect 543568 82521 543596 82758
rect 543554 82512 543610 82521
rect 543554 82447 543610 82456
rect 543556 78668 543608 78674
rect 543556 78610 543608 78616
rect 543568 77761 543596 78610
rect 543554 77752 543610 77761
rect 543554 77687 543610 77696
rect 543556 77240 543608 77246
rect 543556 77182 543608 77188
rect 543568 76401 543596 77182
rect 543554 76392 543610 76401
rect 543554 76327 543610 76336
rect 543556 75880 543608 75886
rect 543556 75822 543608 75828
rect 543568 75041 543596 75822
rect 543554 75032 543610 75041
rect 543554 74967 543610 74976
rect 543556 71732 543608 71738
rect 543556 71674 543608 71680
rect 543568 71641 543596 71674
rect 543554 71632 543610 71641
rect 543554 71567 543610 71576
rect 543556 70372 543608 70378
rect 543556 70314 543608 70320
rect 543568 70281 543596 70314
rect 543554 70272 543610 70281
rect 543554 70207 543610 70216
rect 543554 66192 543610 66201
rect 543554 66127 543556 66136
rect 543608 66127 543610 66136
rect 543556 66098 543608 66104
rect 543660 66094 543688 82894
rect 543648 66088 543700 66094
rect 543648 66030 543700 66036
rect 543554 64152 543610 64161
rect 543554 64087 543610 64096
rect 543568 63986 543596 64087
rect 543556 63980 543608 63986
rect 543556 63922 543608 63928
rect 543554 62112 543610 62121
rect 543554 62047 543556 62056
rect 543608 62047 543610 62056
rect 543556 62018 543608 62024
rect 543648 62008 543700 62014
rect 543648 61950 543700 61956
rect 543660 60761 543688 61950
rect 543646 60752 543702 60761
rect 543646 60687 543702 60696
rect 543556 57928 543608 57934
rect 543556 57870 543608 57876
rect 543568 56681 543596 57870
rect 543554 56672 543610 56681
rect 543554 56607 543610 56616
rect 543556 55888 543608 55894
rect 543556 55830 543608 55836
rect 543568 45121 543596 55830
rect 543648 48272 543700 48278
rect 543648 48214 543700 48220
rect 543660 47841 543688 48214
rect 543646 47832 543702 47841
rect 543646 47767 543702 47776
rect 543648 45552 543700 45558
rect 543648 45494 543700 45500
rect 543554 45112 543610 45121
rect 543554 45047 543610 45056
rect 543660 44441 543688 45494
rect 543646 44432 543702 44441
rect 543646 44367 543702 44376
rect 543648 42832 543700 42838
rect 543648 42774 543700 42780
rect 543556 41404 543608 41410
rect 543556 41346 543608 41352
rect 543568 41041 543596 41346
rect 543554 41032 543610 41041
rect 543554 40967 543610 40976
rect 543556 37256 543608 37262
rect 543556 37198 543608 37204
rect 543568 36281 543596 37198
rect 543554 36272 543610 36281
rect 543554 36207 543610 36216
rect 543660 36122 543688 42774
rect 543568 36094 543688 36122
rect 543464 12096 543516 12102
rect 543464 12038 543516 12044
rect 543568 11966 543596 36094
rect 543648 35896 543700 35902
rect 543648 35838 543700 35844
rect 543660 35601 543688 35838
rect 543646 35592 543702 35601
rect 543646 35527 543702 35536
rect 543646 31240 543702 31249
rect 543646 31175 543702 31184
rect 543660 30433 543688 31175
rect 543646 30424 543702 30433
rect 543646 30359 543702 30368
rect 543752 15026 543780 89814
rect 543832 82612 543884 82618
rect 543832 82554 543884 82560
rect 543740 15020 543792 15026
rect 543740 14962 543792 14968
rect 543556 11960 543608 11966
rect 543556 11902 543608 11908
rect 542360 11688 542412 11694
rect 542360 11630 542412 11636
rect 543844 11558 543872 82554
rect 543936 78441 543964 229706
rect 544028 125746 544056 231678
rect 544120 144809 544148 233815
rect 544200 154012 544252 154018
rect 544200 153954 544252 153960
rect 544106 144800 544162 144809
rect 544106 144735 544162 144744
rect 544108 140072 544160 140078
rect 544108 140014 544160 140020
rect 544120 127702 544148 140014
rect 544108 127696 544160 127702
rect 544108 127638 544160 127644
rect 544028 125718 544148 125746
rect 544016 125588 544068 125594
rect 544016 125530 544068 125536
rect 543922 78432 543978 78441
rect 543922 78367 543978 78376
rect 544028 14822 544056 125530
rect 544120 125390 544148 125718
rect 544108 125384 544160 125390
rect 544108 125326 544160 125332
rect 544108 112056 544160 112062
rect 544108 111998 544160 112004
rect 544120 15842 544148 111998
rect 544212 85134 544240 153954
rect 544396 144906 544424 234058
rect 544474 146568 544530 146577
rect 544474 146503 544530 146512
rect 544384 144900 544436 144906
rect 544384 144842 544436 144848
rect 544384 136468 544436 136474
rect 544384 136410 544436 136416
rect 544292 128376 544344 128382
rect 544292 128318 544344 128324
rect 544304 118046 544332 128318
rect 544396 124234 544424 136410
rect 544488 126886 544516 146503
rect 544658 146296 544714 146305
rect 544658 146231 544714 146240
rect 544568 144288 544620 144294
rect 544568 144230 544620 144236
rect 544580 139466 544608 144230
rect 544672 139505 544700 146231
rect 544658 139496 544714 139505
rect 544568 139460 544620 139466
rect 544658 139431 544714 139440
rect 544568 139402 544620 139408
rect 544660 139256 544712 139262
rect 544660 139198 544712 139204
rect 544566 136640 544622 136649
rect 544566 136575 544622 136584
rect 544580 131209 544608 136575
rect 544672 135318 544700 139198
rect 544660 135312 544712 135318
rect 544660 135254 544712 135260
rect 544566 131200 544622 131209
rect 544566 131135 544622 131144
rect 544476 126880 544528 126886
rect 544476 126822 544528 126828
rect 544476 125452 544528 125458
rect 544476 125394 544528 125400
rect 544384 124228 544436 124234
rect 544384 124170 544436 124176
rect 544384 123480 544436 123486
rect 544384 123422 544436 123428
rect 544292 118040 544344 118046
rect 544292 117982 544344 117988
rect 544290 114472 544346 114481
rect 544290 114407 544346 114416
rect 544304 92206 544332 114407
rect 544292 92200 544344 92206
rect 544292 92142 544344 92148
rect 544292 88324 544344 88330
rect 544292 88266 544344 88272
rect 544200 85128 544252 85134
rect 544200 85070 544252 85076
rect 544304 17542 544332 88266
rect 544396 22030 544424 123422
rect 544488 115938 544516 125394
rect 544566 124128 544622 124137
rect 544566 124063 544622 124072
rect 544580 117337 544608 124063
rect 544566 117328 544622 117337
rect 544566 117263 544622 117272
rect 544568 117224 544620 117230
rect 544568 117166 544620 117172
rect 544476 115932 544528 115938
rect 544476 115874 544528 115880
rect 544580 106962 544608 117166
rect 544568 106956 544620 106962
rect 544568 106898 544620 106904
rect 544476 102196 544528 102202
rect 544476 102138 544528 102144
rect 544488 89078 544516 102138
rect 544476 89072 544528 89078
rect 544476 89014 544528 89020
rect 544476 82884 544528 82890
rect 544476 82826 544528 82832
rect 544384 22024 544436 22030
rect 544384 21966 544436 21972
rect 544292 17536 544344 17542
rect 544292 17478 544344 17484
rect 544488 16386 544516 82826
rect 544568 67380 544620 67386
rect 544568 67322 544620 67328
rect 544476 16380 544528 16386
rect 544476 16322 544528 16328
rect 544108 15836 544160 15842
rect 544108 15778 544160 15784
rect 544016 14816 544068 14822
rect 544016 14758 544068 14764
rect 544580 12306 544608 67322
rect 544764 29238 544792 240178
rect 545592 240094 545928 240122
rect 544844 237924 544896 237930
rect 544844 237866 544896 237872
rect 544752 29232 544804 29238
rect 544752 29174 544804 29180
rect 544856 28150 544884 237866
rect 545592 236842 545620 240094
rect 547234 239456 547290 239465
rect 547234 239391 547290 239400
rect 545856 237924 545908 237930
rect 545856 237866 545908 237872
rect 545672 237856 545724 237862
rect 545672 237798 545724 237804
rect 545580 236836 545632 236842
rect 545580 236778 545632 236784
rect 545304 203584 545356 203590
rect 545304 203526 545356 203532
rect 545316 157334 545344 203526
rect 545396 161356 545448 161362
rect 545396 161298 545448 161304
rect 545132 157306 545344 157334
rect 545132 150362 545160 157306
rect 545040 150334 545160 150362
rect 545304 150408 545356 150414
rect 545304 150350 545356 150356
rect 545040 146946 545068 150334
rect 545028 146940 545080 146946
rect 545028 146882 545080 146888
rect 545028 144152 545080 144158
rect 545028 144094 545080 144100
rect 544936 139460 544988 139466
rect 544936 139402 544988 139408
rect 544948 136406 544976 139402
rect 545040 138038 545068 144094
rect 545120 143404 545172 143410
rect 545120 143346 545172 143352
rect 545028 138032 545080 138038
rect 545028 137974 545080 137980
rect 544936 136400 544988 136406
rect 544936 136342 544988 136348
rect 545028 134564 545080 134570
rect 545028 134506 545080 134512
rect 545040 128228 545068 134506
rect 545132 128382 545160 143346
rect 545210 138136 545266 138145
rect 545210 138071 545266 138080
rect 545224 128489 545252 138071
rect 545210 128480 545266 128489
rect 545210 128415 545266 128424
rect 545120 128376 545172 128382
rect 545120 128318 545172 128324
rect 545040 128200 545252 128228
rect 545118 127120 545174 127129
rect 545118 127055 545174 127064
rect 545028 127016 545080 127022
rect 545028 126958 545080 126964
rect 544936 126812 544988 126818
rect 544936 126754 544988 126760
rect 544948 110498 544976 126754
rect 545040 122834 545068 126958
rect 545132 124001 545160 127055
rect 545224 125594 545252 128200
rect 545212 125588 545264 125594
rect 545212 125530 545264 125536
rect 545118 123992 545174 124001
rect 545118 123927 545174 123936
rect 545040 122806 545160 122834
rect 545132 117230 545160 122806
rect 545120 117224 545172 117230
rect 545120 117166 545172 117172
rect 545212 113144 545264 113150
rect 545212 113086 545264 113092
rect 544936 110492 544988 110498
rect 544936 110434 544988 110440
rect 545028 106276 545080 106282
rect 545028 106218 545080 106224
rect 545040 89486 545068 106218
rect 545028 89480 545080 89486
rect 545028 89422 545080 89428
rect 544936 85536 544988 85542
rect 544936 85478 544988 85484
rect 544948 82210 544976 85478
rect 544936 82204 544988 82210
rect 544936 82146 544988 82152
rect 544844 28144 544896 28150
rect 544844 28086 544896 28092
rect 544568 12300 544620 12306
rect 544568 12242 544620 12248
rect 543832 11552 543884 11558
rect 543832 11494 543884 11500
rect 541072 6724 541124 6730
rect 541072 6666 541124 6672
rect 541990 3224 542046 3233
rect 541990 3159 542046 3168
rect 542004 480 542032 3159
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545224 66 545252 113086
rect 545316 18494 545344 150350
rect 545408 141710 545436 161298
rect 545580 150204 545632 150210
rect 545580 150146 545632 150152
rect 545488 148300 545540 148306
rect 545488 148242 545540 148248
rect 545396 141704 545448 141710
rect 545396 141646 545448 141652
rect 545396 138032 545448 138038
rect 545396 137974 545448 137980
rect 545408 110362 545436 137974
rect 545500 129878 545528 148242
rect 545592 139466 545620 150146
rect 545580 139460 545632 139466
rect 545580 139402 545632 139408
rect 545488 129872 545540 129878
rect 545488 129814 545540 129820
rect 545580 115932 545632 115938
rect 545580 115874 545632 115880
rect 545488 115796 545540 115802
rect 545488 115738 545540 115744
rect 545396 110356 545448 110362
rect 545396 110298 545448 110304
rect 545304 18488 545356 18494
rect 545304 18430 545356 18436
rect 545500 6798 545528 115738
rect 545592 89758 545620 115874
rect 545580 89752 545632 89758
rect 545580 89694 545632 89700
rect 545684 25770 545712 237798
rect 545764 237448 545816 237454
rect 545764 237390 545816 237396
rect 545672 25764 545724 25770
rect 545672 25706 545724 25712
rect 545488 6792 545540 6798
rect 545488 6734 545540 6740
rect 545776 6186 545804 237390
rect 545868 75750 545896 237866
rect 545948 234524 546000 234530
rect 545948 234466 546000 234472
rect 545960 140486 545988 234466
rect 547052 233844 547104 233850
rect 547052 233786 547104 233792
rect 546040 231668 546092 231674
rect 546040 231610 546092 231616
rect 546052 149870 546080 231610
rect 546776 228472 546828 228478
rect 546776 228414 546828 228420
rect 546224 159656 546276 159662
rect 546224 159598 546276 159604
rect 546130 155544 546186 155553
rect 546130 155479 546186 155488
rect 546040 149864 546092 149870
rect 546040 149806 546092 149812
rect 546144 149054 546172 155479
rect 546132 149048 546184 149054
rect 546132 148990 546184 148996
rect 545948 140480 546000 140486
rect 545948 140422 546000 140428
rect 546038 139496 546094 139505
rect 546038 139431 546094 139440
rect 546052 126993 546080 139431
rect 546038 126984 546094 126993
rect 546038 126919 546094 126928
rect 545948 124908 546000 124914
rect 545948 124850 546000 124856
rect 545856 75744 545908 75750
rect 545856 75686 545908 75692
rect 545960 13054 545988 124850
rect 546040 124296 546092 124302
rect 546040 124238 546092 124244
rect 546052 115870 546080 124238
rect 546132 117224 546184 117230
rect 546132 117166 546184 117172
rect 546040 115864 546092 115870
rect 546040 115806 546092 115812
rect 546144 111790 546172 117166
rect 546132 111784 546184 111790
rect 546132 111726 546184 111732
rect 546040 90364 546092 90370
rect 546040 90306 546092 90312
rect 546052 14958 546080 90306
rect 546132 89752 546184 89758
rect 546132 89694 546184 89700
rect 546144 82958 546172 89694
rect 546132 82952 546184 82958
rect 546132 82894 546184 82900
rect 546236 25498 546264 159598
rect 546500 146192 546552 146198
rect 546500 146134 546552 146140
rect 546512 144090 546540 146134
rect 546788 144566 546816 228414
rect 546868 163736 546920 163742
rect 546868 163678 546920 163684
rect 546776 144560 546828 144566
rect 546776 144502 546828 144508
rect 546776 144424 546828 144430
rect 546776 144366 546828 144372
rect 546500 144084 546552 144090
rect 546500 144026 546552 144032
rect 546592 140956 546644 140962
rect 546592 140898 546644 140904
rect 546604 134026 546632 140898
rect 546684 135176 546736 135182
rect 546684 135118 546736 135124
rect 546592 134020 546644 134026
rect 546592 133962 546644 133968
rect 546500 129668 546552 129674
rect 546500 129610 546552 129616
rect 546408 129192 546460 129198
rect 546408 129134 546460 129140
rect 546420 91798 546448 129134
rect 546512 127022 546540 129610
rect 546500 127016 546552 127022
rect 546500 126958 546552 126964
rect 546592 118040 546644 118046
rect 546592 117982 546644 117988
rect 546500 110356 546552 110362
rect 546500 110298 546552 110304
rect 546512 106282 546540 110298
rect 546500 106276 546552 106282
rect 546500 106218 546552 106224
rect 546604 105602 546632 117982
rect 546592 105596 546644 105602
rect 546592 105538 546644 105544
rect 546408 91792 546460 91798
rect 546408 91734 546460 91740
rect 546500 71460 546552 71466
rect 546500 71402 546552 71408
rect 546512 67386 546540 71402
rect 546500 67380 546552 67386
rect 546500 67322 546552 67328
rect 546224 25492 546276 25498
rect 546224 25434 546276 25440
rect 546696 20466 546724 135118
rect 546788 120766 546816 144366
rect 546880 126954 546908 163678
rect 546958 146840 547014 146849
rect 546958 146775 547014 146784
rect 546972 145926 547000 146775
rect 546960 145920 547012 145926
rect 546960 145862 547012 145868
rect 546960 144900 547012 144906
rect 546960 144842 547012 144848
rect 546972 132802 547000 144842
rect 547064 140962 547092 233786
rect 547144 233096 547196 233102
rect 547144 233038 547196 233044
rect 547156 152538 547184 233038
rect 547248 152794 547276 239391
rect 547236 152788 547288 152794
rect 547236 152730 547288 152736
rect 547156 152510 547276 152538
rect 547144 147688 547196 147694
rect 547144 147630 547196 147636
rect 547052 140956 547104 140962
rect 547052 140898 547104 140904
rect 547052 140820 547104 140826
rect 547052 140762 547104 140768
rect 546960 132796 547012 132802
rect 546960 132738 547012 132744
rect 546868 126948 546920 126954
rect 546868 126890 546920 126896
rect 546868 125588 546920 125594
rect 546868 125530 546920 125536
rect 546776 120760 546828 120766
rect 546776 120702 546828 120708
rect 546776 117156 546828 117162
rect 546776 117098 546828 117104
rect 546684 20460 546736 20466
rect 546684 20402 546736 20408
rect 546040 14952 546092 14958
rect 546040 14894 546092 14900
rect 546788 14346 546816 117098
rect 546880 109070 546908 125530
rect 547064 122834 547092 140762
rect 547156 122874 547184 147630
rect 547248 146062 547276 152510
rect 547236 146056 547288 146062
rect 547236 145998 547288 146004
rect 547236 145920 547288 145926
rect 547236 145862 547288 145868
rect 547248 140894 547276 145862
rect 547236 140888 547288 140894
rect 547236 140830 547288 140836
rect 546972 122806 547092 122834
rect 547144 122868 547196 122874
rect 547144 122810 547196 122816
rect 546972 110566 547000 122806
rect 547340 114850 547368 240586
rect 547860 240094 548104 240122
rect 547512 238128 547564 238134
rect 547512 238070 547564 238076
rect 547420 141432 547472 141438
rect 547420 141374 547472 141380
rect 547432 138145 547460 141374
rect 547418 138136 547474 138145
rect 547418 138071 547474 138080
rect 547418 126984 547474 126993
rect 547418 126919 547474 126928
rect 547432 117366 547460 126919
rect 547420 117360 547472 117366
rect 547420 117302 547472 117308
rect 547328 114844 547380 114850
rect 547328 114786 547380 114792
rect 547144 114572 547196 114578
rect 547144 114514 547196 114520
rect 547052 111920 547104 111926
rect 547052 111862 547104 111868
rect 546960 110560 547012 110566
rect 546960 110502 547012 110508
rect 546868 109064 546920 109070
rect 546868 109006 546920 109012
rect 546960 106208 547012 106214
rect 546960 106150 547012 106156
rect 546868 102672 546920 102678
rect 546868 102614 546920 102620
rect 546776 14340 546828 14346
rect 546776 14282 546828 14288
rect 545948 13048 546000 13054
rect 545948 12990 546000 12996
rect 545764 6180 545816 6186
rect 545764 6122 545816 6128
rect 546880 5506 546908 102614
rect 546972 17746 547000 106150
rect 547064 89758 547092 111862
rect 547052 89752 547104 89758
rect 547052 89694 547104 89700
rect 547052 66088 547104 66094
rect 547052 66030 547104 66036
rect 547064 42838 547092 66030
rect 547052 42832 547104 42838
rect 547052 42774 547104 42780
rect 546960 17740 547012 17746
rect 546960 17682 547012 17688
rect 546868 5500 546920 5506
rect 546868 5442 546920 5448
rect 547156 5438 547184 114514
rect 547236 111852 547288 111858
rect 547236 111794 547288 111800
rect 547248 88398 547276 111794
rect 547328 89480 547380 89486
rect 547328 89422 547380 89428
rect 547236 88392 547288 88398
rect 547236 88334 547288 88340
rect 547236 84244 547288 84250
rect 547236 84186 547288 84192
rect 547248 14618 547276 84186
rect 547340 71670 547368 89422
rect 547420 89072 547472 89078
rect 547420 89014 547472 89020
rect 547432 82890 547460 89014
rect 547420 82884 547472 82890
rect 547420 82826 547472 82832
rect 547328 71664 547380 71670
rect 547328 71606 547380 71612
rect 547524 26246 547552 238070
rect 548076 238066 548104 240094
rect 548168 240094 548504 240122
rect 548168 238649 548196 240094
rect 548720 239630 548748 240586
rect 549996 240372 550048 240378
rect 549996 240314 550048 240320
rect 549536 240168 549588 240174
rect 548812 240094 549148 240122
rect 549536 240110 549588 240116
rect 548708 239624 548760 239630
rect 548708 239566 548760 239572
rect 548154 238640 548210 238649
rect 548154 238575 548210 238584
rect 548064 238060 548116 238066
rect 548064 238002 548116 238008
rect 547604 237992 547656 237998
rect 547604 237934 547656 237940
rect 547512 26240 547564 26246
rect 547512 26182 547564 26188
rect 547616 19922 547644 237934
rect 548812 237454 548840 240094
rect 548982 238232 549038 238241
rect 548982 238167 549038 238176
rect 548800 237448 548852 237454
rect 548800 237390 548852 237396
rect 548064 234320 548116 234326
rect 548064 234262 548116 234268
rect 547972 232824 548024 232830
rect 547972 232766 548024 232772
rect 547788 155304 547840 155310
rect 547788 155246 547840 155252
rect 547800 148374 547828 155246
rect 547788 148368 547840 148374
rect 547788 148310 547840 148316
rect 547984 147694 548012 232766
rect 547972 147688 548024 147694
rect 547972 147630 548024 147636
rect 548076 146282 548104 234262
rect 548156 232620 548208 232626
rect 548156 232562 548208 232568
rect 547800 146254 548104 146282
rect 547800 144158 547828 146254
rect 547972 146124 548024 146130
rect 547972 146066 548024 146072
rect 547788 144152 547840 144158
rect 547788 144094 547840 144100
rect 547880 140888 547932 140894
rect 547880 140830 547932 140836
rect 547788 140820 547840 140826
rect 547788 140762 547840 140768
rect 547696 128240 547748 128246
rect 547696 128182 547748 128188
rect 547708 117230 547736 128182
rect 547800 117230 547828 140762
rect 547892 136474 547920 140830
rect 547984 139262 548012 146066
rect 548168 142390 548196 232562
rect 548248 231464 548300 231470
rect 548248 231406 548300 231412
rect 548260 146198 548288 231406
rect 548340 164212 548392 164218
rect 548340 164154 548392 164160
rect 548248 146192 548300 146198
rect 548248 146134 548300 146140
rect 548248 146056 548300 146062
rect 548248 145998 548300 146004
rect 548156 142384 548208 142390
rect 548156 142326 548208 142332
rect 548156 140480 548208 140486
rect 548156 140422 548208 140428
rect 547972 139256 548024 139262
rect 547972 139198 548024 139204
rect 547880 136468 547932 136474
rect 547880 136410 547932 136416
rect 547880 134292 547932 134298
rect 547880 134234 547932 134240
rect 547892 132494 547920 134234
rect 547892 132466 548012 132494
rect 547878 130520 547934 130529
rect 547878 130455 547934 130464
rect 547892 128246 547920 130455
rect 547880 128240 547932 128246
rect 547880 128182 547932 128188
rect 547984 124302 548012 132466
rect 548064 129804 548116 129810
rect 548064 129746 548116 129752
rect 547972 124296 548024 124302
rect 547972 124238 548024 124244
rect 547880 122868 547932 122874
rect 547880 122810 547932 122816
rect 547696 117224 547748 117230
rect 547696 117166 547748 117172
rect 547788 117224 547840 117230
rect 547788 117166 547840 117172
rect 547892 111858 547920 122810
rect 547880 111852 547932 111858
rect 547880 111794 547932 111800
rect 547880 110288 547932 110294
rect 547880 110230 547932 110236
rect 547788 103556 547840 103562
rect 547788 103498 547840 103504
rect 547800 85649 547828 103498
rect 547892 91186 547920 110230
rect 547972 92268 548024 92274
rect 547972 92210 548024 92216
rect 547880 91180 547932 91186
rect 547880 91122 547932 91128
rect 547786 85640 547842 85649
rect 547786 85575 547842 85584
rect 547984 83026 548012 92210
rect 547972 83020 548024 83026
rect 547972 82962 548024 82968
rect 547880 82204 547932 82210
rect 547880 82146 547932 82152
rect 547892 75206 547920 82146
rect 547880 75200 547932 75206
rect 547880 75142 547932 75148
rect 547604 19916 547656 19922
rect 547604 19858 547656 19864
rect 547236 14612 547288 14618
rect 547236 14554 547288 14560
rect 548076 11898 548104 129746
rect 548168 129674 548196 140422
rect 548156 129668 548208 129674
rect 548156 129610 548208 129616
rect 548156 126880 548208 126886
rect 548156 126822 548208 126828
rect 548168 20126 548196 126822
rect 548260 111110 548288 145998
rect 548352 113626 548380 164154
rect 548524 160608 548576 160614
rect 548524 160550 548576 160556
rect 548432 153876 548484 153882
rect 548432 153818 548484 153824
rect 548340 113620 548392 113626
rect 548340 113562 548392 113568
rect 548248 111104 548300 111110
rect 548248 111046 548300 111052
rect 548444 109478 548472 153818
rect 548536 130354 548564 160550
rect 548708 149048 548760 149054
rect 548708 148990 548760 148996
rect 548616 142588 548668 142594
rect 548616 142530 548668 142536
rect 548628 135182 548656 142530
rect 548720 140826 548748 148990
rect 548708 140820 548760 140826
rect 548708 140762 548760 140768
rect 548616 135176 548668 135182
rect 548616 135118 548668 135124
rect 548524 130348 548576 130354
rect 548524 130290 548576 130296
rect 548616 128376 548668 128382
rect 548616 128318 548668 128324
rect 548432 109472 548484 109478
rect 548432 109414 548484 109420
rect 548248 104848 548300 104854
rect 548248 104790 548300 104796
rect 548260 82142 548288 104790
rect 548248 82136 548300 82142
rect 548248 82078 548300 82084
rect 548628 21894 548656 128318
rect 548708 112532 548760 112538
rect 548708 112474 548760 112480
rect 548616 21888 548668 21894
rect 548616 21830 548668 21836
rect 548156 20120 548208 20126
rect 548156 20062 548208 20068
rect 548720 14550 548748 112474
rect 548892 111852 548944 111858
rect 548892 111794 548944 111800
rect 548800 111784 548852 111790
rect 548800 111726 548852 111732
rect 548812 98734 548840 111726
rect 548904 103630 548932 111794
rect 548892 103624 548944 103630
rect 548892 103566 548944 103572
rect 548800 98728 548852 98734
rect 548800 98670 548852 98676
rect 548800 83496 548852 83502
rect 548800 83438 548852 83444
rect 548812 16590 548840 83438
rect 548892 82884 548944 82890
rect 548892 82826 548944 82832
rect 548904 63374 548932 82826
rect 548892 63368 548944 63374
rect 548892 63310 548944 63316
rect 548996 22574 549024 238167
rect 549442 238096 549498 238105
rect 549442 238031 549498 238040
rect 549076 159724 549128 159730
rect 549076 159666 549128 159672
rect 549088 26926 549116 159666
rect 549168 151768 549220 151774
rect 549168 151710 549220 151716
rect 549076 26920 549128 26926
rect 549076 26862 549128 26868
rect 549180 26858 549208 151710
rect 549352 151496 549404 151502
rect 549352 151438 549404 151444
rect 549364 138009 549392 151438
rect 549350 138000 549406 138009
rect 549350 137935 549406 137944
rect 549260 136400 549312 136406
rect 549260 136342 549312 136348
rect 549272 132666 549300 136342
rect 549352 135176 549404 135182
rect 549352 135118 549404 135124
rect 549260 132660 549312 132666
rect 549260 132602 549312 132608
rect 549364 129810 549392 135118
rect 549352 129804 549404 129810
rect 549352 129746 549404 129752
rect 549352 129056 549404 129062
rect 549352 128998 549404 129004
rect 549364 114578 549392 128998
rect 549352 114572 549404 114578
rect 549352 114514 549404 114520
rect 549352 114436 549404 114442
rect 549352 114378 549404 114384
rect 549260 113212 549312 113218
rect 549260 113154 549312 113160
rect 549272 100026 549300 113154
rect 549364 111926 549392 114378
rect 549352 111920 549404 111926
rect 549352 111862 549404 111868
rect 549260 100020 549312 100026
rect 549260 99962 549312 99968
rect 549260 98728 549312 98734
rect 549260 98670 549312 98676
rect 549272 71466 549300 98670
rect 549260 71460 549312 71466
rect 549260 71402 549312 71408
rect 549168 26852 549220 26858
rect 549168 26794 549220 26800
rect 548984 22568 549036 22574
rect 548984 22510 549036 22516
rect 549456 18698 549484 238031
rect 549548 195770 549576 240110
rect 549640 240094 549792 240122
rect 549640 237522 549668 240094
rect 549904 239556 549956 239562
rect 549904 239498 549956 239504
rect 549628 237516 549680 237522
rect 549628 237458 549680 237464
rect 549720 228744 549772 228750
rect 549720 228686 549772 228692
rect 549536 195764 549588 195770
rect 549536 195706 549588 195712
rect 549536 166796 549588 166802
rect 549536 166738 549588 166744
rect 549548 26654 549576 166738
rect 549628 161424 549680 161430
rect 549628 161366 549680 161372
rect 549640 63986 549668 161366
rect 549732 139330 549760 228686
rect 549812 149796 549864 149802
rect 549812 149738 549864 149744
rect 549720 139324 549772 139330
rect 549720 139266 549772 139272
rect 549720 129124 549772 129130
rect 549720 129066 549772 129072
rect 549732 114442 549760 129066
rect 549824 128382 549852 149738
rect 549812 128376 549864 128382
rect 549812 128318 549864 128324
rect 549812 117224 549864 117230
rect 549812 117166 549864 117172
rect 549720 114436 549772 114442
rect 549720 114378 549772 114384
rect 549718 113248 549774 113257
rect 549718 113183 549774 113192
rect 549732 111790 549760 113183
rect 549720 111784 549772 111790
rect 549720 111726 549772 111732
rect 549720 104644 549772 104650
rect 549720 104586 549772 104592
rect 549628 63980 549680 63986
rect 549628 63922 549680 63928
rect 549628 63368 549680 63374
rect 549628 63310 549680 63316
rect 549536 26648 549588 26654
rect 549536 26590 549588 26596
rect 549444 18692 549496 18698
rect 549444 18634 549496 18640
rect 548800 16584 548852 16590
rect 548800 16526 548852 16532
rect 548708 14544 548760 14550
rect 548708 14486 548760 14492
rect 548064 11892 548116 11898
rect 548064 11834 548116 11840
rect 547144 5432 547196 5438
rect 547144 5374 547196 5380
rect 549076 4004 549128 4010
rect 549076 3946 549128 3952
rect 545488 3256 545540 3262
rect 545488 3198 545540 3204
rect 545500 480 545528 3198
rect 549088 480 549116 3946
rect 549640 1358 549668 63310
rect 549732 12918 549760 104586
rect 549824 103562 549852 117166
rect 549812 103556 549864 103562
rect 549812 103498 549864 103504
rect 549812 84992 549864 84998
rect 549812 84934 549864 84940
rect 549824 15774 549852 84934
rect 549812 15768 549864 15774
rect 549812 15710 549864 15716
rect 549720 12912 549772 12918
rect 549720 12854 549772 12860
rect 549916 3466 549944 239498
rect 550008 239426 550036 240314
rect 550100 240174 550128 240751
rect 550088 240168 550140 240174
rect 550088 240110 550140 240116
rect 549996 239420 550048 239426
rect 549996 239362 550048 239368
rect 550192 239290 550220 242791
rect 550180 239284 550232 239290
rect 550180 239226 550232 239232
rect 549996 231532 550048 231538
rect 549996 231474 550048 231480
rect 550008 134638 550036 231474
rect 549996 134632 550048 134638
rect 549996 134574 550048 134580
rect 549996 129804 550048 129810
rect 549996 129746 550048 129752
rect 550008 24682 550036 129746
rect 550086 126304 550142 126313
rect 550086 126239 550142 126248
rect 550100 121514 550128 126239
rect 550088 121508 550140 121514
rect 550088 121450 550140 121456
rect 550088 112464 550140 112470
rect 550088 112406 550140 112412
rect 550100 84250 550128 112406
rect 550088 84244 550140 84250
rect 550088 84186 550140 84192
rect 550088 71664 550140 71670
rect 550088 71606 550140 71612
rect 549996 24676 550048 24682
rect 549996 24618 550048 24624
rect 550100 14482 550128 71606
rect 550284 29306 550312 266591
rect 550362 262576 550418 262585
rect 550362 262511 550418 262520
rect 550272 29300 550324 29306
rect 550272 29242 550324 29248
rect 550376 29034 550404 262511
rect 550548 243976 550600 243982
rect 550548 243918 550600 243924
rect 550560 235890 550588 243918
rect 550652 238474 550680 282231
rect 550744 271425 550772 680886
rect 550824 674144 550876 674150
rect 550824 674086 550876 674092
rect 550836 363905 550864 674086
rect 550928 431905 550956 698906
rect 551100 688016 551152 688022
rect 551100 687958 551152 687964
rect 551008 681012 551060 681018
rect 551008 680954 551060 680960
rect 551020 468625 551048 680954
rect 551112 524385 551140 687958
rect 551192 679312 551244 679318
rect 551192 679254 551244 679260
rect 551098 524376 551154 524385
rect 551098 524311 551154 524320
rect 551204 520985 551232 679254
rect 551190 520976 551246 520985
rect 551190 520911 551246 520920
rect 551296 484362 551324 700538
rect 559668 700534 559696 703520
rect 559656 700528 559708 700534
rect 559656 700470 559708 700476
rect 564716 700392 564768 700398
rect 564716 700334 564768 700340
rect 552940 694816 552992 694822
rect 552940 694758 552992 694764
rect 551374 684720 551430 684729
rect 551374 684655 551430 684664
rect 552480 684684 552532 684690
rect 551388 674150 551416 684655
rect 552480 684626 552532 684632
rect 551468 682644 551520 682650
rect 551468 682586 551520 682592
rect 551376 674144 551428 674150
rect 551376 674086 551428 674092
rect 551376 572756 551428 572762
rect 551376 572698 551428 572704
rect 551284 484356 551336 484362
rect 551284 484298 551336 484304
rect 551006 468616 551062 468625
rect 551006 468551 551062 468560
rect 551284 458380 551336 458386
rect 551284 458322 551336 458328
rect 550914 431896 550970 431905
rect 550914 431831 550970 431840
rect 551006 422376 551062 422385
rect 551006 422311 551062 422320
rect 550914 407416 550970 407425
rect 550914 407351 550970 407360
rect 550822 363896 550878 363905
rect 550822 363831 550878 363840
rect 550822 287736 550878 287745
rect 550822 287671 550878 287680
rect 550730 271416 550786 271425
rect 550730 271351 550786 271360
rect 550640 238468 550692 238474
rect 550640 238410 550692 238416
rect 550548 235884 550600 235890
rect 550548 235826 550600 235832
rect 550730 234152 550786 234161
rect 550730 234087 550786 234096
rect 550640 149932 550692 149938
rect 550640 149874 550692 149880
rect 550652 129810 550680 149874
rect 550744 141438 550772 234087
rect 550732 141432 550784 141438
rect 550732 141374 550784 141380
rect 550640 129804 550692 129810
rect 550640 129746 550692 129752
rect 550640 121508 550692 121514
rect 550640 121450 550692 121456
rect 550652 111858 550680 121450
rect 550640 111852 550692 111858
rect 550640 111794 550692 111800
rect 550364 29028 550416 29034
rect 550364 28970 550416 28976
rect 550088 14476 550140 14482
rect 550088 14418 550140 14424
rect 550836 9110 550864 287671
rect 550928 236910 550956 407351
rect 551020 371385 551048 422311
rect 551006 371376 551062 371385
rect 551006 371311 551062 371320
rect 551098 365256 551154 365265
rect 551098 365191 551154 365200
rect 551006 333976 551062 333985
rect 551006 333911 551062 333920
rect 550916 236904 550968 236910
rect 550916 236846 550968 236852
rect 551020 198354 551048 333911
rect 551112 239494 551140 365191
rect 551190 327856 551246 327865
rect 551190 327791 551246 327800
rect 551100 239488 551152 239494
rect 551100 239430 551152 239436
rect 551204 238882 551232 327791
rect 551192 238876 551244 238882
rect 551192 238818 551244 238824
rect 551008 198348 551060 198354
rect 551008 198290 551060 198296
rect 550916 163872 550968 163878
rect 550916 163814 550968 163820
rect 550928 28898 550956 163814
rect 551100 163804 551152 163810
rect 551100 163746 551152 163752
rect 551008 158092 551060 158098
rect 551008 158034 551060 158040
rect 551020 51066 551048 158034
rect 551112 62014 551140 163746
rect 551192 150136 551244 150142
rect 551192 150078 551244 150084
rect 551204 95946 551232 150078
rect 551192 95940 551244 95946
rect 551192 95882 551244 95888
rect 551192 91792 551244 91798
rect 551192 91734 551244 91740
rect 551100 62008 551152 62014
rect 551100 61950 551152 61956
rect 551008 51060 551060 51066
rect 551008 51002 551060 51008
rect 550916 28892 550968 28898
rect 550916 28834 550968 28840
rect 551204 12034 551232 91734
rect 551296 78674 551324 458322
rect 551388 238338 551416 572698
rect 551480 545358 551508 682586
rect 551560 682508 551612 682514
rect 551560 682450 551612 682456
rect 551572 676598 551600 682450
rect 552112 681352 552164 681358
rect 552112 681294 552164 681300
rect 552018 679416 552074 679425
rect 551928 679380 551980 679386
rect 552018 679351 552074 679360
rect 551928 679322 551980 679328
rect 551940 678994 551968 679322
rect 552032 679114 552060 679351
rect 552020 679108 552072 679114
rect 552020 679050 552072 679056
rect 551940 678966 552060 678994
rect 552032 678162 552060 678966
rect 552020 678156 552072 678162
rect 552020 678098 552072 678104
rect 552018 678056 552074 678065
rect 552018 677991 552074 678000
rect 552032 677618 552060 677991
rect 552020 677612 552072 677618
rect 552020 677554 552072 677560
rect 551560 676592 551612 676598
rect 551560 676534 551612 676540
rect 552018 676016 552074 676025
rect 552018 675951 552074 675960
rect 552032 674898 552060 675951
rect 552020 674892 552072 674898
rect 552020 674834 552072 674840
rect 552124 674098 552152 681294
rect 552388 680876 552440 680882
rect 552388 680818 552440 680824
rect 552204 680808 552256 680814
rect 552204 680750 552256 680756
rect 552216 674218 552244 680750
rect 552296 678156 552348 678162
rect 552296 678098 552348 678104
rect 552308 674665 552336 678098
rect 552294 674656 552350 674665
rect 552294 674591 552350 674600
rect 552204 674212 552256 674218
rect 552204 674154 552256 674160
rect 552124 674070 552336 674098
rect 552204 674008 552256 674014
rect 552204 673950 552256 673956
rect 552018 672480 552074 672489
rect 552018 672415 552074 672424
rect 552032 672110 552060 672415
rect 552020 672104 552072 672110
rect 552020 672046 552072 672052
rect 552216 661745 552244 673950
rect 552202 661736 552258 661745
rect 552202 661671 552258 661680
rect 552110 653576 552166 653585
rect 552110 653511 552166 653520
rect 552124 653274 552152 653511
rect 552112 653268 552164 653274
rect 552112 653210 552164 653216
rect 551558 650176 551614 650185
rect 551558 650111 551614 650120
rect 551468 545352 551520 545358
rect 551468 545294 551520 545300
rect 551468 239420 551520 239426
rect 551468 239362 551520 239368
rect 551376 238332 551428 238338
rect 551376 238274 551428 238280
rect 551376 235476 551428 235482
rect 551376 235418 551428 235424
rect 551388 149802 551416 235418
rect 551480 196450 551508 239362
rect 551572 238785 551600 650111
rect 552110 645416 552166 645425
rect 552110 645351 552166 645360
rect 552124 644502 552152 645351
rect 552112 644496 552164 644502
rect 552112 644438 552164 644444
rect 552020 642592 552072 642598
rect 552020 642534 552072 642540
rect 552032 642025 552060 642534
rect 552018 642016 552074 642025
rect 552018 641951 552074 641960
rect 552110 638344 552166 638353
rect 552110 638279 552166 638288
rect 552018 637936 552074 637945
rect 552124 637906 552152 638279
rect 552018 637871 552074 637880
rect 552112 637900 552164 637906
rect 552032 637634 552060 637871
rect 552112 637842 552164 637848
rect 552020 637628 552072 637634
rect 552020 637570 552072 637576
rect 552018 631816 552074 631825
rect 552018 631751 552074 631760
rect 552032 631242 552060 631751
rect 552020 631236 552072 631242
rect 552020 631178 552072 631184
rect 552018 625424 552074 625433
rect 552018 625359 552020 625368
rect 552072 625359 552074 625368
rect 552020 625330 552072 625336
rect 552018 624336 552074 624345
rect 552018 624271 552074 624280
rect 552032 623830 552060 624271
rect 552020 623824 552072 623830
rect 552020 623766 552072 623772
rect 552202 607336 552258 607345
rect 552202 607271 552204 607280
rect 552256 607271 552258 607280
rect 552204 607242 552256 607248
rect 552020 603968 552072 603974
rect 552018 603936 552020 603945
rect 552072 603936 552074 603945
rect 552018 603871 552074 603880
rect 552032 598505 552060 603871
rect 552308 600545 552336 674070
rect 552400 634545 552428 680818
rect 552492 642705 552520 684626
rect 552846 679824 552902 679833
rect 552846 679759 552902 679768
rect 552572 679244 552624 679250
rect 552572 679186 552624 679192
rect 552584 654265 552612 679186
rect 552756 676592 552808 676598
rect 552756 676534 552808 676540
rect 552570 654256 552626 654265
rect 552570 654191 552626 654200
rect 552570 646776 552626 646785
rect 552570 646711 552626 646720
rect 552584 645930 552612 646711
rect 552572 645924 552624 645930
rect 552572 645866 552624 645872
rect 552478 642696 552534 642705
rect 552478 642631 552534 642640
rect 552386 634536 552442 634545
rect 552386 634471 552442 634480
rect 552570 620256 552626 620265
rect 552570 620191 552626 620200
rect 552584 619682 552612 620191
rect 552572 619676 552624 619682
rect 552572 619618 552624 619624
rect 552478 608696 552534 608705
rect 552478 608631 552480 608640
rect 552532 608631 552534 608640
rect 552480 608602 552532 608608
rect 552294 600536 552350 600545
rect 552294 600471 552350 600480
rect 552018 598496 552074 598505
rect 552018 598431 552074 598440
rect 552294 597544 552350 597553
rect 552294 597479 552350 597488
rect 552018 596456 552074 596465
rect 552018 596391 552074 596400
rect 552032 572762 552060 596391
rect 552112 589008 552164 589014
rect 552110 588976 552112 588985
rect 552164 588976 552166 588985
rect 552110 588911 552166 588920
rect 552112 574048 552164 574054
rect 552110 574016 552112 574025
rect 552164 574016 552166 574025
rect 552110 573951 552166 573960
rect 552020 572756 552072 572762
rect 552020 572698 552072 572704
rect 552018 562456 552074 562465
rect 552018 562391 552020 562400
rect 552072 562391 552074 562400
rect 552020 562362 552072 562368
rect 552018 557016 552074 557025
rect 552018 556951 552074 556960
rect 552032 556578 552060 556951
rect 552020 556572 552072 556578
rect 552020 556514 552072 556520
rect 552308 555665 552336 597479
rect 552570 586256 552626 586265
rect 552570 586191 552626 586200
rect 552584 585206 552612 586191
rect 552572 585200 552624 585206
rect 552572 585142 552624 585148
rect 552570 569936 552626 569945
rect 552570 569871 552626 569880
rect 552584 568614 552612 569871
rect 552572 568608 552624 568614
rect 552478 568576 552534 568585
rect 552572 568550 552624 568556
rect 552478 568511 552534 568520
rect 552492 567254 552520 568511
rect 552480 567248 552532 567254
rect 552480 567190 552532 567196
rect 552294 555656 552350 555665
rect 552294 555591 552350 555600
rect 552020 553852 552072 553858
rect 552020 553794 552072 553800
rect 552032 553625 552060 553794
rect 552018 553616 552074 553625
rect 552018 553551 552074 553560
rect 552386 552936 552442 552945
rect 552386 552871 552442 552880
rect 552400 552090 552428 552871
rect 552388 552084 552440 552090
rect 552388 552026 552440 552032
rect 552110 545456 552166 545465
rect 552110 545391 552166 545400
rect 552020 545352 552072 545358
rect 552020 545294 552072 545300
rect 552032 536625 552060 545294
rect 552018 536616 552074 536625
rect 552018 536551 552074 536560
rect 552020 532568 552072 532574
rect 552018 532536 552020 532545
rect 552072 532536 552074 532545
rect 552018 532471 552074 532480
rect 552020 530936 552072 530942
rect 552020 530878 552072 530884
rect 552032 530505 552060 530878
rect 552018 530496 552074 530505
rect 552018 530431 552074 530440
rect 552018 526416 552074 526425
rect 552018 526351 552074 526360
rect 552032 526114 552060 526351
rect 552020 526108 552072 526114
rect 552020 526050 552072 526056
rect 552020 525768 552072 525774
rect 552018 525736 552020 525745
rect 552072 525736 552074 525745
rect 552018 525671 552074 525680
rect 552018 521656 552074 521665
rect 552018 521591 552074 521600
rect 552032 520334 552060 521591
rect 552020 520328 552072 520334
rect 552020 520270 552072 520276
rect 552018 519480 552074 519489
rect 552018 519415 552074 519424
rect 552032 519314 552060 519415
rect 552020 519308 552072 519314
rect 552020 519250 552072 519256
rect 552020 518968 552072 518974
rect 552018 518936 552020 518945
rect 552072 518936 552074 518945
rect 552018 518871 552074 518880
rect 552018 516896 552074 516905
rect 552018 516831 552074 516840
rect 552032 516186 552060 516831
rect 552020 516180 552072 516186
rect 552020 516122 552072 516128
rect 552018 514856 552074 514865
rect 552018 514791 552020 514800
rect 552072 514791 552074 514800
rect 552020 514762 552072 514768
rect 552020 484356 552072 484362
rect 552020 484298 552072 484304
rect 552032 480185 552060 484298
rect 552018 480176 552074 480185
rect 552018 480111 552074 480120
rect 552018 465896 552074 465905
rect 552018 465831 552074 465840
rect 552032 465118 552060 465831
rect 552020 465112 552072 465118
rect 552020 465054 552072 465060
rect 552018 464400 552074 464409
rect 552018 464335 552074 464344
rect 552032 463962 552060 464335
rect 552020 463956 552072 463962
rect 552020 463898 552072 463904
rect 552018 463176 552074 463185
rect 552018 463111 552074 463120
rect 552032 462398 552060 463111
rect 552020 462392 552072 462398
rect 552020 462334 552072 462340
rect 552018 459776 552074 459785
rect 552018 459711 552074 459720
rect 552032 459610 552060 459711
rect 552020 459604 552072 459610
rect 552020 459546 552072 459552
rect 552018 459096 552074 459105
rect 552018 459031 552020 459040
rect 552072 459031 552074 459040
rect 552020 459002 552072 459008
rect 552018 457736 552074 457745
rect 552018 457671 552074 457680
rect 552032 456822 552060 457671
rect 552020 456816 552072 456822
rect 552020 456758 552072 456764
rect 552018 456376 552074 456385
rect 552018 456311 552020 456320
rect 552072 456311 552074 456320
rect 552020 456282 552072 456288
rect 552018 416256 552074 416265
rect 552018 416191 552074 416200
rect 552032 416090 552060 416191
rect 552020 416084 552072 416090
rect 552020 416026 552072 416032
rect 552018 415576 552074 415585
rect 552018 415511 552074 415520
rect 552032 415478 552060 415511
rect 552020 415472 552072 415478
rect 552020 415414 552072 415420
rect 552018 412856 552074 412865
rect 552018 412791 552020 412800
rect 552072 412791 552074 412800
rect 552020 412762 552072 412768
rect 552018 393816 552074 393825
rect 552018 393751 552074 393760
rect 552032 393514 552060 393751
rect 552020 393508 552072 393514
rect 552020 393450 552072 393456
rect 552020 368144 552072 368150
rect 552020 368086 552072 368092
rect 552032 367985 552060 368086
rect 552018 367976 552074 367985
rect 552018 367911 552074 367920
rect 552018 350976 552074 350985
rect 552018 350911 552020 350920
rect 552072 350911 552074 350920
rect 552020 350882 552072 350888
rect 552020 342848 552072 342854
rect 552018 342816 552020 342825
rect 552072 342816 552074 342825
rect 552018 342751 552074 342760
rect 552018 322416 552074 322425
rect 552018 322351 552074 322360
rect 552032 321842 552060 322351
rect 552020 321836 552072 321842
rect 552020 321778 552072 321784
rect 552020 307488 552072 307494
rect 552018 307456 552020 307465
rect 552072 307456 552074 307465
rect 552018 307391 552074 307400
rect 552018 293176 552074 293185
rect 552018 293111 552020 293120
rect 552072 293111 552074 293120
rect 552020 293082 552072 293088
rect 552018 290456 552074 290465
rect 552018 290391 552074 290400
rect 552032 290154 552060 290391
rect 552020 290148 552072 290154
rect 552020 290090 552072 290096
rect 551928 270088 551980 270094
rect 551928 270030 551980 270036
rect 551558 238776 551614 238785
rect 551558 238711 551614 238720
rect 551468 196444 551520 196450
rect 551468 196386 551520 196392
rect 551940 195294 551968 270030
rect 552018 263256 552074 263265
rect 552018 263191 552074 263200
rect 552032 262410 552060 263191
rect 552020 262404 552072 262410
rect 552020 262346 552072 262352
rect 552018 243400 552074 243409
rect 552018 243335 552074 243344
rect 552032 237386 552060 243335
rect 552124 237930 552152 545391
rect 552570 540696 552626 540705
rect 552570 540631 552626 540640
rect 552584 539646 552612 540631
rect 552572 539640 552624 539646
rect 552572 539582 552624 539588
rect 552570 539336 552626 539345
rect 552570 539271 552626 539280
rect 552584 538286 552612 539271
rect 552572 538280 552624 538286
rect 552572 538222 552624 538228
rect 552386 534576 552442 534585
rect 552386 534511 552442 534520
rect 552400 534206 552428 534511
rect 552388 534200 552440 534206
rect 552388 534142 552440 534148
rect 552478 533896 552534 533905
rect 552478 533831 552534 533840
rect 552294 515536 552350 515545
rect 552294 515471 552350 515480
rect 552204 496596 552256 496602
rect 552204 496538 552256 496544
rect 552216 496505 552244 496538
rect 552202 496496 552258 496505
rect 552202 496431 552258 496440
rect 552202 460456 552258 460465
rect 552202 460391 552258 460400
rect 552216 459678 552244 460391
rect 552204 459672 552256 459678
rect 552204 459614 552256 459620
rect 552202 451480 552258 451489
rect 552202 451415 552258 451424
rect 552216 432585 552244 451415
rect 552202 432576 552258 432585
rect 552202 432511 552258 432520
rect 552308 421705 552336 515471
rect 552386 500576 552442 500585
rect 552386 500511 552442 500520
rect 552400 454345 552428 500511
rect 552492 492425 552520 533831
rect 552662 531176 552718 531185
rect 552662 531111 552718 531120
rect 552676 529990 552704 531111
rect 552664 529984 552716 529990
rect 552664 529926 552716 529932
rect 552570 493776 552626 493785
rect 552570 493711 552626 493720
rect 552584 492726 552612 493711
rect 552572 492720 552624 492726
rect 552572 492662 552624 492668
rect 552478 492416 552534 492425
rect 552478 492351 552534 492360
rect 552570 484256 552626 484265
rect 552570 484191 552626 484200
rect 552584 483070 552612 484191
rect 552572 483064 552624 483070
rect 552572 483006 552624 483012
rect 552570 478816 552626 478825
rect 552570 478751 552626 478760
rect 552584 477562 552612 478751
rect 552572 477556 552624 477562
rect 552572 477498 552624 477504
rect 552478 455016 552534 455025
rect 552478 454951 552534 454960
rect 552386 454336 552442 454345
rect 552386 454271 552442 454280
rect 552492 454102 552520 454951
rect 552480 454096 552532 454102
rect 552480 454038 552532 454044
rect 552570 453656 552626 453665
rect 552570 453591 552626 453600
rect 552584 452674 552612 453591
rect 552572 452668 552624 452674
rect 552572 452610 552624 452616
rect 552386 446856 552442 446865
rect 552386 446791 552442 446800
rect 552294 421696 552350 421705
rect 552294 421631 552350 421640
rect 552296 421048 552348 421054
rect 552294 421016 552296 421025
rect 552348 421016 552350 421025
rect 552294 420951 552350 420960
rect 552202 413400 552258 413409
rect 552202 413335 552258 413344
rect 552216 412690 552244 413335
rect 552204 412684 552256 412690
rect 552204 412626 552256 412632
rect 552294 390416 552350 390425
rect 552294 390351 552350 390360
rect 552308 389230 552336 390351
rect 552296 389224 552348 389230
rect 552296 389166 552348 389172
rect 552202 360496 552258 360505
rect 552202 360431 552204 360440
rect 552256 360431 552258 360440
rect 552204 360402 552256 360408
rect 552294 351656 552350 351665
rect 552294 351591 552350 351600
rect 552308 350606 552336 351591
rect 552296 350600 552348 350606
rect 552296 350542 552348 350548
rect 552294 306096 552350 306105
rect 552294 306031 552350 306040
rect 552308 305386 552336 306031
rect 552296 305380 552348 305386
rect 552296 305322 552348 305328
rect 552202 291816 552258 291825
rect 552202 291751 552204 291760
rect 552256 291751 552258 291760
rect 552204 291722 552256 291728
rect 552294 274816 552350 274825
rect 552294 274751 552296 274760
rect 552348 274751 552350 274760
rect 552296 274722 552348 274728
rect 552400 240378 552428 446791
rect 552570 445496 552626 445505
rect 552570 445431 552626 445440
rect 552584 444446 552612 445431
rect 552572 444440 552624 444446
rect 552572 444382 552624 444388
rect 552662 437336 552718 437345
rect 552662 437271 552718 437280
rect 552676 436150 552704 437271
rect 552664 436144 552716 436150
rect 552664 436086 552716 436092
rect 552662 435976 552718 435985
rect 552662 435911 552718 435920
rect 552676 434790 552704 435911
rect 552664 434784 552716 434790
rect 552664 434726 552716 434732
rect 552662 358456 552718 358465
rect 552662 358391 552718 358400
rect 552676 357678 552704 358391
rect 552664 357672 552716 357678
rect 552664 357614 552716 357620
rect 552662 347576 552718 347585
rect 552662 347511 552718 347520
rect 552676 346458 552704 347511
rect 552664 346452 552716 346458
rect 552664 346394 552716 346400
rect 552478 331256 552534 331265
rect 552478 331191 552534 331200
rect 552388 240372 552440 240378
rect 552388 240314 552440 240320
rect 552112 237924 552164 237930
rect 552112 237866 552164 237872
rect 552020 237380 552072 237386
rect 552020 237322 552072 237328
rect 551928 195288 551980 195294
rect 551928 195230 551980 195236
rect 552492 183258 552520 331191
rect 552570 314936 552626 314945
rect 552570 314871 552626 314880
rect 552480 183252 552532 183258
rect 552480 183194 552532 183200
rect 552584 180334 552612 314871
rect 552662 301336 552718 301345
rect 552662 301271 552718 301280
rect 552572 180328 552624 180334
rect 552572 180270 552624 180276
rect 552676 174622 552704 301271
rect 552768 235385 552796 676534
rect 552860 665825 552888 679759
rect 552846 665816 552902 665825
rect 552846 665751 552902 665760
rect 552952 597825 552980 694758
rect 554136 687540 554188 687546
rect 554136 687482 554188 687488
rect 553952 687472 554004 687478
rect 553952 687414 554004 687420
rect 553768 686112 553820 686118
rect 553768 686054 553820 686060
rect 553492 680740 553544 680746
rect 553492 680682 553544 680688
rect 553400 680672 553452 680678
rect 553400 680614 553452 680620
rect 553124 679448 553176 679454
rect 553124 679390 553176 679396
rect 553030 670576 553086 670585
rect 553030 670511 553086 670520
rect 552938 597816 552994 597825
rect 552938 597751 552994 597760
rect 552938 584896 552994 584905
rect 552938 584831 552994 584840
rect 552952 583778 552980 584831
rect 552940 583772 552992 583778
rect 552940 583714 552992 583720
rect 552938 561096 552994 561105
rect 552938 561031 552994 561040
rect 552952 560386 552980 561031
rect 552940 560380 552992 560386
rect 552940 560322 552992 560328
rect 552938 558376 552994 558385
rect 552938 558311 552994 558320
rect 552952 557666 552980 558311
rect 552940 557660 552992 557666
rect 552940 557602 552992 557608
rect 552846 484936 552902 484945
rect 552846 484871 552902 484880
rect 552860 484634 552888 484871
rect 552848 484628 552900 484634
rect 552848 484570 552900 484576
rect 552938 476096 552994 476105
rect 552938 476031 552994 476040
rect 552952 474774 552980 476031
rect 552940 474768 552992 474774
rect 552940 474710 552992 474716
rect 553044 458386 553072 670511
rect 553136 547505 553164 679390
rect 553306 667856 553362 667865
rect 553306 667791 553362 667800
rect 553320 666602 553348 667791
rect 553308 666596 553360 666602
rect 553308 666538 553360 666544
rect 553306 656976 553362 656985
rect 553306 656911 553308 656920
rect 553360 656911 553362 656920
rect 553308 656882 553360 656888
rect 553306 648816 553362 648825
rect 553306 648751 553362 648760
rect 553320 648650 553348 648751
rect 553308 648644 553360 648650
rect 553308 648586 553360 648592
rect 553214 644736 553270 644745
rect 553214 644671 553216 644680
rect 553268 644671 553270 644680
rect 553216 644642 553268 644648
rect 553306 641336 553362 641345
rect 553306 641271 553362 641280
rect 553320 640354 553348 641271
rect 553308 640348 553360 640354
rect 553308 640290 553360 640296
rect 553306 617536 553362 617545
rect 553306 617471 553362 617480
rect 553320 616894 553348 617471
rect 553308 616888 553360 616894
rect 553308 616830 553360 616836
rect 553214 613456 553270 613465
rect 553214 613391 553270 613400
rect 553228 612814 553256 613391
rect 553308 612876 553360 612882
rect 553308 612818 553360 612824
rect 553216 612808 553268 612814
rect 553320 612785 553348 612818
rect 553216 612750 553268 612756
rect 553306 612776 553362 612785
rect 553306 612711 553362 612720
rect 553306 611416 553362 611425
rect 553306 611351 553308 611360
rect 553360 611351 553362 611360
rect 553308 611322 553360 611328
rect 553306 610736 553362 610745
rect 553306 610671 553362 610680
rect 553320 610026 553348 610671
rect 553308 610020 553360 610026
rect 553308 609962 553360 609968
rect 553306 605976 553362 605985
rect 553412 605962 553440 680614
rect 553362 605934 553440 605962
rect 553306 605911 553362 605920
rect 553306 603256 553362 603265
rect 553306 603191 553362 603200
rect 553320 603158 553348 603191
rect 553308 603152 553360 603158
rect 553308 603094 553360 603100
rect 553306 599856 553362 599865
rect 553306 599791 553362 599800
rect 553320 599010 553348 599791
rect 553308 599004 553360 599010
rect 553308 598946 553360 598952
rect 553306 586936 553362 586945
rect 553306 586871 553362 586880
rect 553320 586566 553348 586871
rect 553308 586560 553360 586566
rect 553308 586502 553360 586508
rect 553214 585576 553270 585585
rect 553214 585511 553270 585520
rect 553122 547496 553178 547505
rect 553122 547431 553178 547440
rect 553124 506456 553176 506462
rect 553124 506398 553176 506404
rect 553136 505345 553164 506398
rect 553122 505336 553178 505345
rect 553122 505271 553178 505280
rect 553122 501936 553178 501945
rect 553122 501871 553178 501880
rect 553136 501090 553164 501871
rect 553124 501084 553176 501090
rect 553124 501026 553176 501032
rect 553122 493096 553178 493105
rect 553122 493031 553178 493040
rect 553032 458380 553084 458386
rect 553032 458322 553084 458328
rect 553030 449576 553086 449585
rect 553030 449511 553086 449520
rect 553044 448594 553072 449511
rect 553032 448588 553084 448594
rect 553032 448530 553084 448536
rect 552846 428496 552902 428505
rect 552846 428431 552902 428440
rect 552860 418154 552888 428431
rect 553032 426488 553084 426494
rect 553030 426456 553032 426465
rect 553084 426456 553086 426465
rect 553030 426391 553086 426400
rect 553032 425128 553084 425134
rect 553030 425096 553032 425105
rect 553084 425096 553086 425105
rect 553030 425031 553086 425040
rect 552938 424416 552994 424425
rect 552938 424351 552994 424360
rect 552952 423774 552980 424351
rect 552940 423768 552992 423774
rect 552940 423710 552992 423716
rect 553030 423736 553086 423745
rect 553030 423671 553032 423680
rect 553084 423671 553086 423680
rect 553032 423642 553084 423648
rect 553030 420336 553086 420345
rect 553030 420271 553086 420280
rect 553044 419898 553072 420271
rect 553032 419892 553084 419898
rect 553032 419834 553084 419840
rect 552860 418126 553072 418154
rect 552940 405680 552992 405686
rect 552940 405622 552992 405628
rect 552952 405385 552980 405622
rect 552938 405376 552994 405385
rect 552938 405311 552994 405320
rect 552846 404016 552902 404025
rect 552846 403951 552902 403960
rect 552860 403034 552888 403951
rect 552938 403336 552994 403345
rect 552938 403271 552994 403280
rect 552952 403102 552980 403271
rect 552940 403096 552992 403102
rect 552940 403038 552992 403044
rect 552848 403028 552900 403034
rect 552848 402970 552900 402976
rect 552938 395176 552994 395185
rect 552938 395111 552994 395120
rect 552952 394738 552980 395111
rect 552940 394732 552992 394738
rect 552940 394674 552992 394680
rect 552846 391776 552902 391785
rect 552846 391711 552902 391720
rect 552860 390658 552888 391711
rect 552938 391096 552994 391105
rect 552938 391031 552994 391040
rect 552848 390652 552900 390658
rect 552848 390594 552900 390600
rect 552952 390590 552980 391031
rect 552940 390584 552992 390590
rect 552940 390526 552992 390532
rect 552938 388376 552994 388385
rect 552938 388311 552994 388320
rect 552952 387870 552980 388311
rect 552940 387864 552992 387870
rect 552940 387806 552992 387812
rect 552938 387696 552994 387705
rect 552938 387631 552994 387640
rect 552952 386442 552980 387631
rect 552940 386436 552992 386442
rect 552940 386378 552992 386384
rect 552938 385656 552994 385665
rect 552938 385591 552994 385600
rect 552952 385082 552980 385591
rect 552940 385076 552992 385082
rect 552940 385018 552992 385024
rect 552938 381576 552994 381585
rect 552938 381511 552994 381520
rect 552952 381138 552980 381511
rect 552940 381132 552992 381138
rect 552940 381074 552992 381080
rect 552938 377496 552994 377505
rect 552938 377431 552994 377440
rect 552952 376786 552980 377431
rect 552940 376780 552992 376786
rect 552940 376722 552992 376728
rect 552938 372736 552994 372745
rect 552938 372671 552940 372680
rect 552992 372671 552994 372680
rect 552940 372642 552992 372648
rect 552938 370696 552994 370705
rect 552938 370631 552994 370640
rect 552952 369918 552980 370631
rect 552940 369912 552992 369918
rect 552940 369854 552992 369860
rect 552846 369336 552902 369345
rect 552846 369271 552902 369280
rect 552860 368558 552888 369271
rect 552938 368656 552994 368665
rect 552938 368591 552940 368600
rect 552992 368591 552994 368600
rect 552940 368562 552992 368568
rect 552848 368552 552900 368558
rect 552848 368494 552900 368500
rect 552846 366480 552902 366489
rect 552846 366415 552902 366424
rect 552860 365770 552888 366415
rect 552938 365936 552994 365945
rect 552938 365871 552994 365880
rect 552952 365838 552980 365871
rect 552940 365832 552992 365838
rect 552940 365774 552992 365780
rect 552848 365764 552900 365770
rect 552848 365706 552900 365712
rect 552848 362976 552900 362982
rect 552848 362918 552900 362924
rect 552860 270094 552888 362918
rect 552938 361176 552994 361185
rect 552938 361111 552994 361120
rect 552952 360262 552980 361111
rect 552940 360256 552992 360262
rect 552940 360198 552992 360204
rect 552940 358760 552992 358766
rect 552940 358702 552992 358708
rect 552952 357785 552980 358702
rect 552938 357776 552994 357785
rect 552938 357711 552994 357720
rect 552938 355736 552994 355745
rect 552938 355671 552994 355680
rect 552952 354754 552980 355671
rect 552940 354748 552992 354754
rect 552940 354690 552992 354696
rect 552940 354476 552992 354482
rect 552940 354418 552992 354424
rect 552952 340105 552980 354418
rect 552938 340096 552994 340105
rect 552938 340031 552994 340040
rect 552938 336016 552994 336025
rect 552938 335951 552994 335960
rect 552952 335374 552980 335951
rect 552940 335368 552992 335374
rect 552940 335310 552992 335316
rect 552938 326496 552994 326505
rect 552938 326431 552994 326440
rect 552952 325718 552980 326431
rect 552940 325712 552992 325718
rect 552940 325654 552992 325660
rect 552938 323776 552994 323785
rect 552938 323711 552994 323720
rect 552952 323338 552980 323711
rect 552940 323332 552992 323338
rect 552940 323274 552992 323280
rect 552938 318336 552994 318345
rect 552938 318271 552994 318280
rect 552952 317490 552980 318271
rect 552940 317484 552992 317490
rect 552940 317426 552992 317432
rect 552938 314256 552994 314265
rect 552938 314191 552994 314200
rect 552952 313342 552980 314191
rect 552940 313336 552992 313342
rect 552940 313278 552992 313284
rect 552938 311400 552994 311409
rect 552938 311335 552994 311344
rect 552952 310622 552980 311335
rect 552940 310616 552992 310622
rect 552940 310558 552992 310564
rect 552938 289776 552994 289785
rect 552938 289711 552994 289720
rect 552952 288522 552980 289711
rect 552940 288516 552992 288522
rect 552940 288458 552992 288464
rect 552940 280152 552992 280158
rect 552940 280094 552992 280100
rect 552952 279585 552980 280094
rect 552938 279576 552994 279585
rect 552938 279511 552994 279520
rect 552848 270088 552900 270094
rect 552848 270030 552900 270036
rect 552938 264616 552994 264625
rect 552938 264551 552994 264560
rect 552952 263634 552980 264551
rect 552940 263628 552992 263634
rect 552940 263570 552992 263576
rect 552938 260400 552994 260409
rect 552938 260335 552994 260344
rect 552952 259554 552980 260335
rect 552940 259548 552992 259554
rect 552940 259490 552992 259496
rect 552938 255096 552994 255105
rect 552938 255031 552994 255040
rect 552952 254046 552980 255031
rect 552940 254040 552992 254046
rect 552940 253982 552992 253988
rect 552938 250336 552994 250345
rect 552938 250271 552994 250280
rect 552952 249830 552980 250271
rect 552940 249824 552992 249830
rect 552940 249766 552992 249772
rect 552754 235376 552810 235385
rect 552754 235311 552810 235320
rect 552756 235068 552808 235074
rect 552756 235010 552808 235016
rect 552664 174616 552716 174622
rect 552664 174558 552716 174564
rect 552572 169040 552624 169046
rect 552572 168982 552624 168988
rect 552112 163940 552164 163946
rect 552112 163882 552164 163888
rect 551468 162172 551520 162178
rect 551468 162114 551520 162120
rect 551376 149796 551428 149802
rect 551376 149738 551428 149744
rect 551376 111784 551428 111790
rect 551376 111726 551428 111732
rect 551388 92546 551416 111726
rect 551376 92540 551428 92546
rect 551376 92482 551428 92488
rect 551376 91792 551428 91798
rect 551376 91734 551428 91740
rect 551284 78668 551336 78674
rect 551284 78610 551336 78616
rect 551284 76288 551336 76294
rect 551284 76230 551336 76236
rect 551296 20670 551324 76230
rect 551284 20664 551336 20670
rect 551284 20606 551336 20612
rect 551388 19242 551416 91734
rect 551480 24002 551508 162114
rect 552020 158296 552072 158302
rect 552020 158238 552072 158244
rect 551560 157072 551612 157078
rect 551560 157014 551612 157020
rect 551468 23996 551520 24002
rect 551468 23938 551520 23944
rect 551572 22098 551600 157014
rect 551928 139460 551980 139466
rect 551928 139402 551980 139408
rect 551940 122834 551968 139402
rect 552032 129198 552060 158238
rect 552020 129192 552072 129198
rect 552020 129134 552072 129140
rect 551940 122806 552060 122834
rect 552032 114510 552060 122806
rect 552020 114504 552072 114510
rect 552020 114446 552072 114452
rect 552020 92540 552072 92546
rect 552020 92482 552072 92488
rect 552032 81569 552060 92482
rect 552018 81560 552074 81569
rect 552018 81495 552074 81504
rect 552124 28966 552152 163882
rect 552202 163568 552258 163577
rect 552202 163503 552258 163512
rect 552216 29646 552244 163503
rect 552480 161288 552532 161294
rect 552480 161230 552532 161236
rect 552294 151464 552350 151473
rect 552294 151399 552350 151408
rect 552204 29640 552256 29646
rect 552204 29582 552256 29588
rect 552112 28960 552164 28966
rect 552112 28902 552164 28908
rect 552308 24818 552336 151399
rect 552388 151156 552440 151162
rect 552388 151098 552440 151104
rect 552400 29510 552428 151098
rect 552492 49706 552520 161230
rect 552584 93838 552612 168982
rect 552662 146976 552718 146985
rect 552662 146911 552718 146920
rect 552676 133113 552704 146911
rect 552662 133104 552718 133113
rect 552662 133039 552718 133048
rect 552768 123486 552796 235010
rect 552848 231328 552900 231334
rect 552848 231270 552900 231276
rect 552860 147558 552888 231270
rect 553044 159458 553072 418126
rect 553136 354482 553164 493031
rect 553124 354476 553176 354482
rect 553124 354418 553176 354424
rect 553122 354376 553178 354385
rect 553122 354311 553178 354320
rect 553136 353802 553164 354311
rect 553124 353796 553176 353802
rect 553124 353738 553176 353744
rect 553122 353696 553178 353705
rect 553122 353631 553178 353640
rect 553136 353326 553164 353631
rect 553124 353320 553176 353326
rect 553124 353262 553176 353268
rect 553122 349480 553178 349489
rect 553122 349415 553178 349424
rect 553136 349178 553164 349415
rect 553124 349172 553176 349178
rect 553124 349114 553176 349120
rect 553122 346896 553178 346905
rect 553122 346831 553178 346840
rect 553136 346526 553164 346831
rect 553124 346520 553176 346526
rect 553124 346462 553176 346468
rect 553122 343496 553178 343505
rect 553122 343431 553178 343440
rect 553136 342310 553164 343431
rect 553124 342304 553176 342310
rect 553124 342246 553176 342252
rect 553122 338736 553178 338745
rect 553122 338671 553178 338680
rect 553136 338162 553164 338671
rect 553124 338156 553176 338162
rect 553124 338098 553176 338104
rect 553122 335336 553178 335345
rect 553122 335271 553124 335280
rect 553176 335271 553178 335280
rect 553124 335242 553176 335248
rect 553122 334656 553178 334665
rect 553122 334591 553178 334600
rect 553136 334014 553164 334591
rect 553124 334008 553176 334014
rect 553124 333950 553176 333956
rect 553122 327176 553178 327185
rect 553122 327111 553124 327120
rect 553176 327111 553178 327120
rect 553124 327082 553176 327088
rect 553122 325816 553178 325825
rect 553122 325751 553124 325760
rect 553176 325751 553178 325760
rect 553124 325722 553176 325728
rect 553122 317656 553178 317665
rect 553122 317591 553178 317600
rect 553136 317558 553164 317591
rect 553124 317552 553176 317558
rect 553124 317494 553176 317500
rect 553122 316296 553178 316305
rect 553122 316231 553178 316240
rect 553136 316062 553164 316231
rect 553124 316056 553176 316062
rect 553124 315998 553176 316004
rect 553124 313268 553176 313274
rect 553124 313210 553176 313216
rect 553136 312905 553164 313210
rect 553122 312896 553178 312905
rect 553122 312831 553178 312840
rect 553122 310856 553178 310865
rect 553122 310791 553178 310800
rect 553136 310554 553164 310791
rect 553124 310548 553176 310554
rect 553124 310490 553176 310496
rect 553122 310176 553178 310185
rect 553122 310111 553178 310120
rect 553136 309194 553164 310111
rect 553124 309188 553176 309194
rect 553124 309130 553176 309136
rect 553122 308816 553178 308825
rect 553122 308751 553178 308760
rect 553136 307834 553164 308751
rect 553124 307828 553176 307834
rect 553124 307770 553176 307776
rect 553122 305416 553178 305425
rect 553122 305351 553178 305360
rect 553136 305046 553164 305351
rect 553124 305040 553176 305046
rect 553124 304982 553176 304988
rect 553122 302016 553178 302025
rect 553122 301951 553178 301960
rect 553136 300898 553164 301951
rect 553124 300892 553176 300898
rect 553124 300834 553176 300840
rect 553122 300656 553178 300665
rect 553122 300591 553178 300600
rect 553136 299538 553164 300591
rect 553124 299532 553176 299538
rect 553124 299474 553176 299480
rect 553122 297936 553178 297945
rect 553122 297871 553124 297880
rect 553176 297871 553178 297880
rect 553124 297842 553176 297848
rect 553122 297256 553178 297265
rect 553122 297191 553178 297200
rect 553136 296750 553164 297191
rect 553124 296744 553176 296750
rect 553124 296686 553176 296692
rect 553122 292496 553178 292505
rect 553122 292431 553178 292440
rect 553136 291242 553164 292431
rect 553124 291236 553176 291242
rect 553124 291178 553176 291184
rect 553122 289096 553178 289105
rect 553122 289031 553178 289040
rect 553136 288454 553164 289031
rect 553124 288448 553176 288454
rect 553124 288390 553176 288396
rect 553122 286376 553178 286385
rect 553122 286311 553178 286320
rect 553136 285734 553164 286311
rect 553124 285728 553176 285734
rect 553124 285670 553176 285676
rect 553122 283656 553178 283665
rect 553122 283591 553124 283600
rect 553176 283591 553178 283600
rect 553124 283562 553176 283568
rect 553124 282872 553176 282878
rect 553124 282814 553176 282820
rect 553136 281625 553164 282814
rect 553122 281616 553178 281625
rect 553122 281551 553178 281560
rect 553122 280936 553178 280945
rect 553122 280871 553124 280880
rect 553176 280871 553178 280880
rect 553124 280842 553176 280848
rect 553122 280256 553178 280265
rect 553122 280191 553124 280200
rect 553176 280191 553178 280200
rect 553124 280162 553176 280168
rect 553122 278896 553178 278905
rect 553122 278831 553178 278840
rect 553136 278798 553164 278831
rect 553124 278792 553176 278798
rect 553124 278734 553176 278740
rect 553122 277536 553178 277545
rect 553122 277471 553178 277480
rect 553136 277438 553164 277471
rect 553124 277432 553176 277438
rect 553124 277374 553176 277380
rect 553122 276176 553178 276185
rect 553122 276111 553178 276120
rect 553136 276078 553164 276111
rect 553124 276072 553176 276078
rect 553124 276014 553176 276020
rect 553122 273456 553178 273465
rect 553122 273391 553178 273400
rect 553136 273290 553164 273391
rect 553124 273284 553176 273290
rect 553124 273226 553176 273232
rect 553122 270736 553178 270745
rect 553122 270671 553178 270680
rect 553136 270570 553164 270671
rect 553124 270564 553176 270570
rect 553124 270506 553176 270512
rect 553122 268696 553178 268705
rect 553122 268631 553124 268640
rect 553176 268631 553178 268640
rect 553124 268602 553176 268608
rect 553122 265296 553178 265305
rect 553122 265231 553178 265240
rect 553136 264994 553164 265231
rect 553124 264988 553176 264994
rect 553124 264930 553176 264936
rect 553122 263936 553178 263945
rect 553122 263871 553178 263880
rect 553136 263702 553164 263871
rect 553124 263696 553176 263702
rect 553124 263638 553176 263644
rect 553122 261896 553178 261905
rect 553122 261831 553178 261840
rect 553136 260914 553164 261831
rect 553124 260908 553176 260914
rect 553124 260850 553176 260856
rect 553122 259856 553178 259865
rect 553122 259791 553178 259800
rect 553136 259486 553164 259791
rect 553124 259480 553176 259486
rect 553124 259422 553176 259428
rect 553122 259176 553178 259185
rect 553122 259111 553178 259120
rect 553136 258126 553164 259111
rect 553124 258120 553176 258126
rect 553124 258062 553176 258068
rect 553122 257816 553178 257825
rect 553122 257751 553178 257760
rect 553136 256766 553164 257751
rect 553124 256760 553176 256766
rect 553124 256702 553176 256708
rect 553122 254416 553178 254425
rect 553122 254351 553178 254360
rect 553136 253978 553164 254351
rect 553124 253972 553176 253978
rect 553124 253914 553176 253920
rect 553122 253736 553178 253745
rect 553122 253671 553178 253680
rect 553136 252618 553164 253671
rect 553124 252612 553176 252618
rect 553124 252554 553176 252560
rect 553122 252376 553178 252385
rect 553122 252311 553178 252320
rect 553136 251258 553164 252311
rect 553124 251252 553176 251258
rect 553124 251194 553176 251200
rect 553124 249756 553176 249762
rect 553124 249698 553176 249704
rect 553136 249665 553164 249698
rect 553122 249656 553178 249665
rect 553122 249591 553178 249600
rect 553122 248296 553178 248305
rect 553122 248231 553178 248240
rect 553136 247178 553164 248231
rect 553124 247172 553176 247178
rect 553124 247114 553176 247120
rect 553122 246256 553178 246265
rect 553122 246191 553178 246200
rect 553136 245682 553164 246191
rect 553124 245676 553176 245682
rect 553124 245618 553176 245624
rect 553122 244896 553178 244905
rect 553122 244831 553178 244840
rect 553136 244322 553164 244831
rect 553124 244316 553176 244322
rect 553124 244258 553176 244264
rect 553228 174593 553256 585511
rect 553306 578096 553362 578105
rect 553306 578031 553362 578040
rect 553320 577250 553348 578031
rect 553308 577244 553360 577250
rect 553308 577186 553360 577192
rect 553306 576056 553362 576065
rect 553306 575991 553362 576000
rect 553320 575550 553348 575991
rect 553308 575544 553360 575550
rect 553308 575486 553360 575492
rect 553306 567896 553362 567905
rect 553306 567831 553362 567840
rect 553320 567322 553348 567831
rect 553308 567316 553360 567322
rect 553308 567258 553360 567264
rect 553306 560416 553362 560425
rect 553306 560351 553362 560360
rect 553320 560318 553348 560351
rect 553308 560312 553360 560318
rect 553308 560254 553360 560260
rect 553306 557696 553362 557705
rect 553306 557631 553362 557640
rect 553320 557598 553348 557631
rect 553308 557592 553360 557598
rect 553308 557534 553360 557540
rect 553306 550896 553362 550905
rect 553306 550831 553308 550840
rect 553360 550831 553362 550840
rect 553308 550802 553360 550808
rect 553306 549536 553362 549545
rect 553306 549471 553362 549480
rect 553320 549302 553348 549471
rect 553308 549296 553360 549302
rect 553308 549238 553360 549244
rect 553306 546816 553362 546825
rect 553306 546751 553362 546760
rect 553320 546514 553348 546751
rect 553308 546508 553360 546514
rect 553308 546450 553360 546456
rect 553306 544096 553362 544105
rect 553306 544031 553362 544040
rect 553320 543794 553348 544031
rect 553308 543788 553360 543794
rect 553308 543730 553360 543736
rect 553306 535936 553362 535945
rect 553306 535871 553308 535880
rect 553360 535871 553362 535880
rect 553308 535842 553360 535848
rect 553306 535256 553362 535265
rect 553306 535191 553362 535200
rect 553320 534138 553348 535191
rect 553308 534132 553360 534138
rect 553308 534074 553360 534080
rect 553306 528456 553362 528465
rect 553306 528391 553362 528400
rect 553320 527202 553348 528391
rect 553308 527196 553360 527202
rect 553308 527138 553360 527144
rect 553306 510096 553362 510105
rect 553306 510031 553362 510040
rect 553320 509930 553348 510031
rect 553308 509924 553360 509930
rect 553308 509866 553360 509872
rect 553306 506016 553362 506025
rect 553306 505951 553362 505960
rect 553320 505170 553348 505951
rect 553308 505164 553360 505170
rect 553308 505106 553360 505112
rect 553306 504656 553362 504665
rect 553306 504591 553362 504600
rect 553320 503742 553348 504591
rect 553308 503736 553360 503742
rect 553308 503678 553360 503684
rect 553306 502480 553362 502489
rect 553306 502415 553308 502424
rect 553360 502415 553362 502424
rect 553308 502386 553360 502392
rect 553306 501256 553362 501265
rect 553306 501191 553362 501200
rect 553320 501022 553348 501191
rect 553308 501016 553360 501022
rect 553308 500958 553360 500964
rect 553306 499896 553362 499905
rect 553306 499831 553308 499840
rect 553360 499831 553362 499840
rect 553308 499802 553360 499808
rect 553306 498536 553362 498545
rect 553306 498471 553362 498480
rect 553320 498234 553348 498471
rect 553308 498228 553360 498234
rect 553308 498170 553360 498176
rect 553306 495816 553362 495825
rect 553306 495751 553362 495760
rect 553320 495514 553348 495751
rect 553308 495508 553360 495514
rect 553308 495450 553360 495456
rect 553306 489016 553362 489025
rect 553306 488951 553362 488960
rect 553320 488850 553348 488951
rect 553308 488844 553360 488850
rect 553308 488786 553360 488792
rect 553306 488336 553362 488345
rect 553306 488271 553362 488280
rect 553320 487218 553348 488271
rect 553308 487212 553360 487218
rect 553308 487154 553360 487160
rect 553306 479496 553362 479505
rect 553306 479431 553362 479440
rect 553320 478922 553348 479431
rect 553308 478916 553360 478922
rect 553308 478858 553360 478864
rect 553306 475416 553362 475425
rect 553306 475351 553362 475360
rect 553320 474842 553348 475351
rect 553308 474836 553360 474842
rect 553308 474778 553360 474784
rect 553306 470656 553362 470665
rect 553306 470591 553308 470600
rect 553360 470591 553362 470600
rect 553308 470562 553360 470568
rect 553306 469976 553362 469985
rect 553306 469911 553362 469920
rect 553320 469266 553348 469911
rect 553308 469260 553360 469266
rect 553308 469202 553360 469208
rect 553306 466576 553362 466585
rect 553306 466511 553362 466520
rect 553320 466478 553348 466511
rect 553308 466472 553360 466478
rect 553308 466414 553360 466420
rect 553306 448896 553362 448905
rect 553306 448831 553362 448840
rect 553320 448662 553348 448831
rect 553308 448656 553360 448662
rect 553308 448598 553360 448604
rect 553306 443456 553362 443465
rect 553306 443391 553362 443400
rect 553320 443018 553348 443391
rect 553308 443012 553360 443018
rect 553308 442954 553360 442960
rect 553306 438696 553362 438705
rect 553306 438631 553362 438640
rect 553320 438122 553348 438631
rect 553308 438116 553360 438122
rect 553308 438058 553360 438064
rect 553306 438016 553362 438025
rect 553306 437951 553362 437960
rect 553320 437510 553348 437951
rect 553308 437504 553360 437510
rect 553308 437446 553360 437452
rect 553306 436656 553362 436665
rect 553306 436591 553362 436600
rect 553214 174584 553270 174593
rect 553214 174519 553270 174528
rect 553320 160750 553348 436591
rect 553504 429865 553532 680682
rect 553582 679688 553638 679697
rect 553582 679623 553638 679632
rect 553490 429856 553546 429865
rect 553490 429791 553546 429800
rect 553596 378185 553624 679623
rect 553676 679584 553728 679590
rect 553676 679526 553728 679532
rect 553688 525774 553716 679526
rect 553780 532574 553808 686054
rect 553860 679176 553912 679182
rect 553860 679118 553912 679124
rect 553768 532568 553820 532574
rect 553768 532510 553820 532516
rect 553872 530942 553900 679118
rect 553964 553858 553992 687414
rect 554044 686044 554096 686050
rect 554044 685986 554096 685992
rect 554056 574054 554084 685986
rect 554148 589014 554176 687482
rect 554228 687404 554280 687410
rect 554228 687346 554280 687352
rect 554240 642598 554268 687346
rect 563704 683800 563756 683806
rect 563704 683742 563756 683748
rect 555240 683528 555292 683534
rect 555240 683470 555292 683476
rect 554872 682236 554924 682242
rect 554872 682178 554924 682184
rect 554228 642592 554280 642598
rect 554228 642534 554280 642540
rect 554228 631236 554280 631242
rect 554228 631178 554280 631184
rect 554136 589008 554188 589014
rect 554136 588950 554188 588956
rect 554044 574048 554096 574054
rect 554044 573990 554096 573996
rect 553952 553852 554004 553858
rect 553952 553794 554004 553800
rect 553860 530936 553912 530942
rect 553860 530878 553912 530884
rect 553768 526108 553820 526114
rect 553768 526050 553820 526056
rect 553676 525768 553728 525774
rect 553676 525710 553728 525716
rect 553676 519308 553728 519314
rect 553676 519250 553728 519256
rect 553582 378176 553638 378185
rect 553582 378111 553638 378120
rect 553688 342854 553716 519250
rect 553780 368150 553808 526050
rect 553952 459060 554004 459066
rect 553952 459002 554004 459008
rect 553860 456340 553912 456346
rect 553860 456282 553912 456288
rect 553768 368144 553820 368150
rect 553768 368086 553820 368092
rect 553676 342848 553728 342854
rect 553676 342790 553728 342796
rect 553582 340776 553638 340785
rect 553582 340711 553638 340720
rect 553398 258496 553454 258505
rect 553398 258431 553454 258440
rect 553308 160744 553360 160750
rect 553308 160686 553360 160692
rect 553032 159452 553084 159458
rect 553032 159394 553084 159400
rect 552848 147552 552900 147558
rect 552848 147494 552900 147500
rect 552846 138680 552902 138689
rect 552846 138615 552902 138624
rect 552756 123480 552808 123486
rect 552756 123422 552808 123428
rect 552664 101448 552716 101454
rect 552664 101390 552716 101396
rect 552572 93832 552624 93838
rect 552572 93774 552624 93780
rect 552480 49700 552532 49706
rect 552480 49642 552532 49648
rect 552388 29504 552440 29510
rect 552388 29446 552440 29452
rect 552296 24812 552348 24818
rect 552296 24754 552348 24760
rect 551560 22092 551612 22098
rect 551560 22034 551612 22040
rect 552676 21826 552704 101390
rect 552756 80096 552808 80102
rect 552756 80038 552808 80044
rect 552664 21820 552716 21826
rect 552664 21762 552716 21768
rect 551376 19236 551428 19242
rect 551376 19178 551428 19184
rect 552768 15162 552796 80038
rect 552756 15156 552808 15162
rect 552756 15098 552808 15104
rect 551192 12028 551244 12034
rect 551192 11970 551244 11976
rect 550824 9104 550876 9110
rect 550824 9046 550876 9052
rect 552664 3732 552716 3738
rect 552664 3674 552716 3680
rect 549904 3460 549956 3466
rect 549904 3402 549956 3408
rect 549628 1352 549680 1358
rect 549628 1294 549680 1300
rect 552676 480 552704 3674
rect 552860 3194 552888 138615
rect 553308 113892 553360 113898
rect 553308 113834 553360 113840
rect 553320 111042 553348 113834
rect 553308 111036 553360 111042
rect 553308 110978 553360 110984
rect 553412 9042 553440 258431
rect 553490 247616 553546 247625
rect 553490 247551 553546 247560
rect 553504 236706 553532 247551
rect 553492 236700 553544 236706
rect 553492 236642 553544 236648
rect 553490 89040 553546 89049
rect 553490 88975 553546 88984
rect 553504 27334 553532 88975
rect 553492 27328 553544 27334
rect 553492 27270 553544 27276
rect 553596 20058 553624 340711
rect 553676 321836 553728 321842
rect 553676 321778 553728 321784
rect 553688 21690 553716 321778
rect 553872 307494 553900 456282
rect 553860 307488 553912 307494
rect 553860 307430 553912 307436
rect 553768 293140 553820 293146
rect 553768 293082 553820 293088
rect 553676 21684 553728 21690
rect 553676 21626 553728 21632
rect 553584 20052 553636 20058
rect 553584 19994 553636 20000
rect 553780 13190 553808 293082
rect 553860 290148 553912 290154
rect 553860 290090 553912 290096
rect 553872 22778 553900 290090
rect 553964 198558 553992 459002
rect 554044 350940 554096 350946
rect 554044 350882 554096 350888
rect 554056 239358 554084 350882
rect 554044 239352 554096 239358
rect 554044 239294 554096 239300
rect 554044 238128 554096 238134
rect 554044 238070 554096 238076
rect 553952 198552 554004 198558
rect 553952 198494 554004 198500
rect 553952 155100 554004 155106
rect 553952 155042 554004 155048
rect 553860 22772 553912 22778
rect 553860 22714 553912 22720
rect 553768 13184 553820 13190
rect 553768 13126 553820 13132
rect 553400 9036 553452 9042
rect 553400 8978 553452 8984
rect 553964 4078 553992 155042
rect 554056 22710 554084 238070
rect 554240 235414 554268 631178
rect 554884 603974 554912 682178
rect 555146 681184 555202 681193
rect 555146 681119 555202 681128
rect 554964 653268 555016 653274
rect 554964 653210 555016 653216
rect 554872 603968 554924 603974
rect 554872 603910 554924 603916
rect 554872 556572 554924 556578
rect 554872 556514 554924 556520
rect 554320 393508 554372 393514
rect 554320 393450 554372 393456
rect 554228 235408 554280 235414
rect 554228 235350 554280 235356
rect 554136 155644 554188 155650
rect 554136 155586 554188 155592
rect 554148 29374 554176 155586
rect 554226 151056 554282 151065
rect 554226 150991 554282 151000
rect 554240 89185 554268 150991
rect 554226 89176 554282 89185
rect 554226 89111 554282 89120
rect 554136 29368 554188 29374
rect 554136 29310 554188 29316
rect 554044 22704 554096 22710
rect 554044 22646 554096 22652
rect 554332 20194 554360 393450
rect 554780 262404 554832 262410
rect 554780 262346 554832 262352
rect 554792 238270 554820 262346
rect 554780 238264 554832 238270
rect 554780 238206 554832 238212
rect 554884 25945 554912 556514
rect 554976 239873 555004 653210
rect 555056 607300 555108 607306
rect 555056 607242 555108 607248
rect 554962 239864 555018 239873
rect 554962 239799 555018 239808
rect 554964 232416 555016 232422
rect 554964 232358 555016 232364
rect 554870 25936 554926 25945
rect 554870 25871 554926 25880
rect 554976 22642 555004 232358
rect 555068 196625 555096 607242
rect 555160 362982 555188 681119
rect 555252 421054 555280 683470
rect 561036 682372 561088 682378
rect 561036 682314 561088 682320
rect 555332 681080 555384 681086
rect 555332 681022 555384 681028
rect 555344 496602 555372 681022
rect 558920 656940 558972 656946
rect 558920 656882 558972 656888
rect 556436 645924 556488 645930
rect 556436 645866 556488 645872
rect 555700 608660 555752 608666
rect 555700 608602 555752 608608
rect 555332 496596 555384 496602
rect 555332 496538 555384 496544
rect 555240 421048 555292 421054
rect 555240 420990 555292 420996
rect 555332 412820 555384 412826
rect 555332 412762 555384 412768
rect 555148 362976 555200 362982
rect 555148 362918 555200 362924
rect 555148 360460 555200 360466
rect 555148 360402 555200 360408
rect 555054 196616 555110 196625
rect 555054 196551 555110 196560
rect 555056 155576 555108 155582
rect 555056 155518 555108 155524
rect 554964 22636 555016 22642
rect 554964 22578 555016 22584
rect 554320 20188 554372 20194
rect 554320 20130 554372 20136
rect 553952 4072 554004 4078
rect 553952 4014 554004 4020
rect 555068 3330 555096 155518
rect 555160 10334 555188 360402
rect 555240 274780 555292 274786
rect 555240 274722 555292 274728
rect 555252 19990 555280 274722
rect 555344 238542 555372 412762
rect 555424 305380 555476 305386
rect 555424 305322 555476 305328
rect 555332 238536 555384 238542
rect 555332 238478 555384 238484
rect 555436 188329 555464 305322
rect 555516 291780 555568 291786
rect 555516 291722 555568 291728
rect 555528 233986 555556 291722
rect 555608 234456 555660 234462
rect 555608 234398 555660 234404
rect 555516 233980 555568 233986
rect 555516 233922 555568 233928
rect 555514 231568 555570 231577
rect 555514 231503 555570 231512
rect 555422 188320 555478 188329
rect 555422 188255 555478 188264
rect 555424 153128 555476 153134
rect 555424 153070 555476 153076
rect 555332 152720 555384 152726
rect 555332 152662 555384 152668
rect 555344 23118 555372 152662
rect 555332 23112 555384 23118
rect 555332 23054 555384 23060
rect 555436 22982 555464 153070
rect 555528 139466 555556 231503
rect 555620 146946 555648 234398
rect 555608 146940 555660 146946
rect 555608 146882 555660 146888
rect 555516 139460 555568 139466
rect 555516 139402 555568 139408
rect 555516 139324 555568 139330
rect 555516 139266 555568 139272
rect 555528 115938 555556 139266
rect 555516 115932 555568 115938
rect 555516 115874 555568 115880
rect 555516 114504 555568 114510
rect 555516 114446 555568 114452
rect 555528 80102 555556 114446
rect 555516 80096 555568 80102
rect 555516 80038 555568 80044
rect 555712 25430 555740 608602
rect 556252 484628 556304 484634
rect 556252 484570 556304 484576
rect 556158 150240 556214 150249
rect 556158 150175 556214 150184
rect 556172 134570 556200 150175
rect 556160 134564 556212 134570
rect 556160 134506 556212 134512
rect 556160 111036 556212 111042
rect 556160 110978 556212 110984
rect 556172 90370 556200 110978
rect 556160 90364 556212 90370
rect 556160 90306 556212 90312
rect 555700 25424 555752 25430
rect 555700 25366 555752 25372
rect 555424 22976 555476 22982
rect 555424 22918 555476 22924
rect 555240 19984 555292 19990
rect 555240 19926 555292 19932
rect 555148 10328 555200 10334
rect 555148 10270 555200 10276
rect 556264 7614 556292 484570
rect 556344 463956 556396 463962
rect 556344 463898 556396 463904
rect 556356 24410 556384 463898
rect 556448 238377 556476 645866
rect 556804 644700 556856 644706
rect 556804 644642 556856 644648
rect 556816 632058 556844 644642
rect 557816 637900 557868 637906
rect 557816 637842 557868 637848
rect 556804 632052 556856 632058
rect 556804 631994 556856 632000
rect 557080 625388 557132 625394
rect 557080 625330 557132 625336
rect 556620 562420 556672 562426
rect 556620 562362 556672 562368
rect 556528 372700 556580 372706
rect 556528 372642 556580 372648
rect 556434 238368 556490 238377
rect 556434 238303 556490 238312
rect 556434 234696 556490 234705
rect 556434 234631 556490 234640
rect 556448 189854 556476 234631
rect 556436 189848 556488 189854
rect 556436 189790 556488 189796
rect 556436 155168 556488 155174
rect 556436 155110 556488 155116
rect 556344 24404 556396 24410
rect 556344 24346 556396 24352
rect 556252 7608 556304 7614
rect 556252 7550 556304 7556
rect 556448 4146 556476 155110
rect 556540 8974 556568 372642
rect 556632 236570 556660 562362
rect 556804 357672 556856 357678
rect 556804 357614 556856 357620
rect 556712 323332 556764 323338
rect 556712 323274 556764 323280
rect 556620 236564 556672 236570
rect 556620 236506 556672 236512
rect 556620 157004 556672 157010
rect 556620 156946 556672 156952
rect 556632 20602 556660 156946
rect 556724 22846 556752 323274
rect 556816 236638 556844 357614
rect 556896 297900 556948 297906
rect 556896 297842 556948 297848
rect 556804 236632 556856 236638
rect 556804 236574 556856 236580
rect 556804 195288 556856 195294
rect 556804 195230 556856 195236
rect 556816 110945 556844 195230
rect 556908 189922 556936 297842
rect 556988 268660 557040 268666
rect 556988 268602 557040 268608
rect 557000 196654 557028 268602
rect 556988 196648 557040 196654
rect 556988 196590 557040 196596
rect 556896 189916 556948 189922
rect 556896 189858 556948 189864
rect 556896 151224 556948 151230
rect 556896 151166 556948 151172
rect 556908 117298 556936 151166
rect 556896 117292 556948 117298
rect 556896 117234 556948 117240
rect 556896 115932 556948 115938
rect 556896 115874 556948 115880
rect 556802 110936 556858 110945
rect 556802 110871 556858 110880
rect 556908 76294 556936 115874
rect 556896 76288 556948 76294
rect 556896 76230 556948 76236
rect 556712 22840 556764 22846
rect 556712 22782 556764 22788
rect 556620 20596 556672 20602
rect 556620 20538 556672 20544
rect 557092 16318 557120 625330
rect 557632 577244 557684 577250
rect 557632 577186 557684 577192
rect 557540 152448 557592 152454
rect 557540 152390 557592 152396
rect 557552 136542 557580 152390
rect 557540 136536 557592 136542
rect 557540 136478 557592 136484
rect 557644 24478 557672 577186
rect 557724 499860 557776 499866
rect 557724 499802 557776 499808
rect 557632 24472 557684 24478
rect 557632 24414 557684 24420
rect 557080 16312 557132 16318
rect 557080 16254 557132 16260
rect 557736 10402 557764 499802
rect 557828 197985 557856 637842
rect 558552 612876 558604 612882
rect 558552 612818 558604 612824
rect 558000 438116 558052 438122
rect 558000 438058 558052 438064
rect 557908 368620 557960 368626
rect 557908 368562 557960 368568
rect 557814 197976 557870 197985
rect 557814 197911 557870 197920
rect 557816 155780 557868 155786
rect 557816 155722 557868 155728
rect 557828 41410 557856 155722
rect 557816 41404 557868 41410
rect 557816 41346 557868 41352
rect 557724 10396 557776 10402
rect 557724 10338 557776 10344
rect 556528 8968 556580 8974
rect 556528 8910 556580 8916
rect 557920 4826 557948 368562
rect 558012 238406 558040 438058
rect 558092 419892 558144 419898
rect 558092 419834 558144 419840
rect 558000 238400 558052 238406
rect 558000 238342 558052 238348
rect 558000 238060 558052 238066
rect 558000 238002 558052 238008
rect 558012 18970 558040 238002
rect 558104 235346 558132 419834
rect 558184 353796 558236 353802
rect 558184 353738 558236 353744
rect 558092 235340 558144 235346
rect 558092 235282 558144 235288
rect 558196 182986 558224 353738
rect 558276 280900 558328 280906
rect 558276 280842 558328 280848
rect 558288 198490 558316 280842
rect 558368 231600 558420 231606
rect 558368 231542 558420 231548
rect 558276 198484 558328 198490
rect 558276 198426 558328 198432
rect 558184 182980 558236 182986
rect 558184 182922 558236 182928
rect 558092 156732 558144 156738
rect 558092 156674 558144 156680
rect 558104 121446 558132 156674
rect 558276 140888 558328 140894
rect 558276 140830 558328 140836
rect 558184 134020 558236 134026
rect 558184 133962 558236 133968
rect 558092 121440 558144 121446
rect 558092 121382 558144 121388
rect 558000 18964 558052 18970
rect 558000 18906 558052 18912
rect 558196 13326 558224 133962
rect 558288 20369 558316 140830
rect 558380 140826 558408 231542
rect 558458 148608 558514 148617
rect 558458 148543 558514 148552
rect 558368 140820 558420 140826
rect 558368 140762 558420 140768
rect 558472 135114 558500 148543
rect 558460 135108 558512 135114
rect 558460 135050 558512 135056
rect 558564 22914 558592 612818
rect 558932 143546 558960 656882
rect 560484 599004 560536 599010
rect 560484 598946 560536 598952
rect 560392 583772 560444 583778
rect 560392 583714 560444 583720
rect 559472 550860 559524 550866
rect 559472 550802 559524 550808
rect 559380 535900 559432 535906
rect 559380 535842 559432 535848
rect 559104 509924 559156 509930
rect 559104 509866 559156 509872
rect 559012 502444 559064 502450
rect 559012 502386 559064 502392
rect 558920 143540 558972 143546
rect 558920 143482 558972 143488
rect 558920 140820 558972 140826
rect 558920 140762 558972 140768
rect 558552 22908 558604 22914
rect 558552 22850 558604 22856
rect 558274 20360 558330 20369
rect 558274 20295 558330 20304
rect 558932 16114 558960 140762
rect 558920 16108 558972 16114
rect 558920 16050 558972 16056
rect 558184 13320 558236 13326
rect 558184 13262 558236 13268
rect 559024 12986 559052 502386
rect 559116 21758 559144 509866
rect 559196 488844 559248 488850
rect 559196 488786 559248 488792
rect 559104 21752 559156 21758
rect 559104 21694 559156 21700
rect 559208 20262 559236 488786
rect 559288 452668 559340 452674
rect 559288 452610 559340 452616
rect 559196 20256 559248 20262
rect 559196 20198 559248 20204
rect 559012 12980 559064 12986
rect 559012 12922 559064 12928
rect 559300 6254 559328 452610
rect 559392 198898 559420 535842
rect 559484 234054 559512 550802
rect 559564 538280 559616 538286
rect 559564 538222 559616 538228
rect 559576 238610 559604 538222
rect 559656 416084 559708 416090
rect 559656 416026 559708 416032
rect 559564 238604 559616 238610
rect 559564 238546 559616 238552
rect 559472 234048 559524 234054
rect 559472 233990 559524 233996
rect 559564 228608 559616 228614
rect 559564 228550 559616 228556
rect 559380 198892 559432 198898
rect 559380 198834 559432 198840
rect 559472 158500 559524 158506
rect 559472 158442 559524 158448
rect 559380 158024 559432 158030
rect 559380 157966 559432 157972
rect 559392 139398 559420 157966
rect 559380 139392 559432 139398
rect 559380 139334 559432 139340
rect 559484 122806 559512 158442
rect 559576 140962 559604 228550
rect 559668 198830 559696 416026
rect 559748 381132 559800 381138
rect 559748 381074 559800 381080
rect 559656 198824 559708 198830
rect 559656 198766 559708 198772
rect 559760 187610 559788 381074
rect 560300 258120 560352 258126
rect 560300 258062 560352 258068
rect 560312 239426 560340 258062
rect 560300 239420 560352 239426
rect 560300 239362 560352 239368
rect 560298 231296 560354 231305
rect 560298 231231 560354 231240
rect 559748 187604 559800 187610
rect 559748 187546 559800 187552
rect 559840 151292 559892 151298
rect 559840 151234 559892 151240
rect 559748 147552 559800 147558
rect 559748 147494 559800 147500
rect 559564 140956 559616 140962
rect 559564 140898 559616 140904
rect 559760 137766 559788 147494
rect 559748 137760 559800 137766
rect 559748 137702 559800 137708
rect 559564 137352 559616 137358
rect 559564 137294 559616 137300
rect 559654 137320 559710 137329
rect 559472 122800 559524 122806
rect 559472 122742 559524 122748
rect 559576 13258 559604 137294
rect 559654 137255 559710 137264
rect 559668 86193 559696 137255
rect 559654 86184 559710 86193
rect 559654 86119 559710 86128
rect 559852 24070 559880 151234
rect 560312 140894 560340 231231
rect 560404 164898 560432 583714
rect 560496 197169 560524 598946
rect 560668 575544 560720 575550
rect 560668 575486 560720 575492
rect 560576 567316 560628 567322
rect 560576 567258 560628 567264
rect 560482 197160 560538 197169
rect 560482 197095 560538 197104
rect 560588 184346 560616 567258
rect 560680 197033 560708 575486
rect 560760 546508 560812 546514
rect 560760 546450 560812 546456
rect 560772 198801 560800 546450
rect 560852 390652 560904 390658
rect 560852 390594 560904 390600
rect 560758 198792 560814 198801
rect 560758 198727 560814 198736
rect 560666 197024 560722 197033
rect 560666 196959 560722 196968
rect 560864 189990 560892 390594
rect 560944 386436 560996 386442
rect 560944 386378 560996 386384
rect 560956 199170 560984 386378
rect 561048 238134 561076 682314
rect 562600 637628 562652 637634
rect 562600 637570 562652 637576
rect 561864 557660 561916 557666
rect 561864 557602 561916 557608
rect 561772 448656 561824 448662
rect 561772 448598 561824 448604
rect 561036 238128 561088 238134
rect 561036 238070 561088 238076
rect 561036 234184 561088 234190
rect 561036 234126 561088 234132
rect 560944 199164 560996 199170
rect 560944 199106 560996 199112
rect 560852 189984 560904 189990
rect 560852 189926 560904 189932
rect 560576 184340 560628 184346
rect 560576 184282 560628 184288
rect 560484 166592 560536 166598
rect 560484 166534 560536 166540
rect 560392 164892 560444 164898
rect 560392 164834 560444 164840
rect 560392 149864 560444 149870
rect 560392 149806 560444 149812
rect 560404 144294 560432 149806
rect 560392 144288 560444 144294
rect 560392 144230 560444 144236
rect 560300 140888 560352 140894
rect 560300 140830 560352 140836
rect 560300 134632 560352 134638
rect 560300 134574 560352 134580
rect 560312 112538 560340 134574
rect 560300 112532 560352 112538
rect 560300 112474 560352 112480
rect 560496 27606 560524 166534
rect 560576 164144 560628 164150
rect 560576 164086 560628 164092
rect 560588 35902 560616 164086
rect 560944 164008 560996 164014
rect 560944 163950 560996 163956
rect 560668 161084 560720 161090
rect 560668 161026 560720 161032
rect 560680 37262 560708 161026
rect 560760 152652 560812 152658
rect 560760 152594 560812 152600
rect 560668 37256 560720 37262
rect 560668 37198 560720 37204
rect 560576 35896 560628 35902
rect 560576 35838 560628 35844
rect 560772 31113 560800 152594
rect 560852 144220 560904 144226
rect 560852 144162 560904 144168
rect 560758 31104 560814 31113
rect 560758 31039 560814 31048
rect 560484 27600 560536 27606
rect 560484 27542 560536 27548
rect 560864 26178 560892 144162
rect 560956 62082 560984 163950
rect 561048 135182 561076 234126
rect 561220 166728 561272 166734
rect 561220 166670 561272 166676
rect 561128 140956 561180 140962
rect 561128 140898 561180 140904
rect 561036 135176 561088 135182
rect 561036 135118 561088 135124
rect 561140 83502 561168 140898
rect 561128 83496 561180 83502
rect 561128 83438 561180 83444
rect 560944 62076 560996 62082
rect 560944 62018 560996 62024
rect 560852 26172 560904 26178
rect 560852 26114 560904 26120
rect 559840 24064 559892 24070
rect 559840 24006 559892 24012
rect 560298 17640 560354 17649
rect 560298 17575 560354 17584
rect 560312 16658 560340 17575
rect 560300 16652 560352 16658
rect 560300 16594 560352 16600
rect 559564 13252 559616 13258
rect 559564 13194 559616 13200
rect 561232 6866 561260 166670
rect 561680 152856 561732 152862
rect 561680 152798 561732 152804
rect 561312 152584 561364 152590
rect 561312 152526 561364 152532
rect 561220 6860 561272 6866
rect 561220 6802 561272 6808
rect 559288 6248 559340 6254
rect 559288 6190 559340 6196
rect 561324 6050 561352 152526
rect 561692 129742 561720 152798
rect 561680 129736 561732 129742
rect 561680 129678 561732 129684
rect 561784 27198 561812 448598
rect 561876 185706 561904 557602
rect 561956 543788 562008 543794
rect 561956 543730 562008 543736
rect 561864 185700 561916 185706
rect 561864 185642 561916 185648
rect 561968 182034 561996 543730
rect 562232 437504 562284 437510
rect 562232 437446 562284 437452
rect 562048 403096 562100 403102
rect 562048 403038 562100 403044
rect 561956 182028 562008 182034
rect 561956 181970 562008 181976
rect 561864 152924 561916 152930
rect 561864 152866 561916 152872
rect 561772 27192 561824 27198
rect 561772 27134 561824 27140
rect 561312 6044 561364 6050
rect 561312 5986 561364 5992
rect 557908 4820 557960 4826
rect 557908 4762 557960 4768
rect 556436 4140 556488 4146
rect 556436 4082 556488 4088
rect 556160 4072 556212 4078
rect 556160 4014 556212 4020
rect 555056 3324 555108 3330
rect 555056 3266 555108 3272
rect 552848 3188 552900 3194
rect 552848 3130 552900 3136
rect 556172 480 556200 4014
rect 561876 3738 561904 152866
rect 561954 149288 562010 149297
rect 561954 149223 562010 149232
rect 561968 18834 561996 149223
rect 562060 55894 562088 403038
rect 562140 369912 562192 369918
rect 562140 369854 562192 369860
rect 562048 55888 562100 55894
rect 562048 55830 562100 55836
rect 562152 28014 562180 369854
rect 562244 193866 562272 437446
rect 562324 291236 562376 291242
rect 562324 291178 562376 291184
rect 562336 240854 562364 291178
rect 562416 247172 562468 247178
rect 562416 247114 562468 247120
rect 562324 240848 562376 240854
rect 562324 240790 562376 240796
rect 562324 235136 562376 235142
rect 562324 235078 562376 235084
rect 562232 193860 562284 193866
rect 562232 193802 562284 193808
rect 562232 155508 562284 155514
rect 562232 155450 562284 155456
rect 562244 107642 562272 155450
rect 562232 107636 562284 107642
rect 562232 107578 562284 107584
rect 562140 28008 562192 28014
rect 562140 27950 562192 27956
rect 562336 23322 562364 235078
rect 562428 199889 562456 247114
rect 562508 231396 562560 231402
rect 562508 231338 562560 231344
rect 562414 199880 562470 199889
rect 562414 199815 562470 199824
rect 562416 127628 562468 127634
rect 562416 127570 562468 127576
rect 562324 23316 562376 23322
rect 562324 23258 562376 23264
rect 561956 18828 562008 18834
rect 561956 18770 562008 18776
rect 562428 13394 562456 127570
rect 562520 126954 562548 231338
rect 562508 126948 562560 126954
rect 562508 126890 562560 126896
rect 562612 28286 562640 637570
rect 563336 567248 563388 567254
rect 563336 567190 563388 567196
rect 563152 474836 563204 474842
rect 563152 474778 563204 474784
rect 563060 135108 563112 135114
rect 563060 135050 563112 135056
rect 563072 112470 563100 135050
rect 563060 112464 563112 112470
rect 563060 112406 563112 112412
rect 563164 28694 563192 474778
rect 563244 385076 563296 385082
rect 563244 385018 563296 385024
rect 563152 28688 563204 28694
rect 563152 28630 563204 28636
rect 562600 28280 562652 28286
rect 562600 28222 562652 28228
rect 563256 27946 563284 385018
rect 563348 224330 563376 567190
rect 563428 529984 563480 529990
rect 563428 529926 563480 529932
rect 563440 232490 563468 529926
rect 563612 495508 563664 495514
rect 563612 495450 563664 495456
rect 563520 436144 563572 436150
rect 563520 436086 563572 436092
rect 563428 232484 563480 232490
rect 563428 232426 563480 232432
rect 563428 228540 563480 228546
rect 563428 228482 563480 228488
rect 563336 224324 563388 224330
rect 563336 224266 563388 224272
rect 563336 152992 563388 152998
rect 563336 152934 563388 152940
rect 563244 27940 563296 27946
rect 563244 27882 563296 27888
rect 562416 13388 562468 13394
rect 562416 13330 562468 13336
rect 563348 4078 563376 152934
rect 563440 13802 563468 228482
rect 563532 169114 563560 436086
rect 563624 237114 563652 495450
rect 563716 247722 563744 683742
rect 564532 648644 564584 648650
rect 564532 648586 564584 648592
rect 563980 477556 564032 477562
rect 563980 477498 564032 477504
rect 563888 288516 563940 288522
rect 563888 288458 563940 288464
rect 563796 277432 563848 277438
rect 563796 277374 563848 277380
rect 563704 247716 563756 247722
rect 563704 247658 563756 247664
rect 563704 245676 563756 245682
rect 563704 245618 563756 245624
rect 563612 237108 563664 237114
rect 563612 237050 563664 237056
rect 563612 235680 563664 235686
rect 563612 235622 563664 235628
rect 563520 169108 563572 169114
rect 563520 169050 563572 169056
rect 563520 166660 563572 166666
rect 563520 166602 563572 166608
rect 563532 19038 563560 166602
rect 563624 27470 563652 235622
rect 563612 27464 563664 27470
rect 563612 27406 563664 27412
rect 563716 24342 563744 245618
rect 563808 25566 563836 277374
rect 563900 241262 563928 288458
rect 563888 241256 563940 241262
rect 563888 241198 563940 241204
rect 563888 231260 563940 231266
rect 563888 231202 563940 231208
rect 563900 134026 563928 231202
rect 563888 134020 563940 134026
rect 563888 133962 563940 133968
rect 563796 25560 563848 25566
rect 563796 25502 563848 25508
rect 563704 24336 563756 24342
rect 563704 24278 563756 24284
rect 563520 19032 563572 19038
rect 563520 18974 563572 18980
rect 563428 13796 563480 13802
rect 563428 13738 563480 13744
rect 563992 6914 564020 477498
rect 564440 256760 564492 256766
rect 564440 256702 564492 256708
rect 564452 239562 564480 256702
rect 564440 239556 564492 239562
rect 564440 239498 564492 239504
rect 564544 147626 564572 648586
rect 564624 518968 564676 518974
rect 564624 518910 564676 518916
rect 564532 147620 564584 147626
rect 564532 147562 564584 147568
rect 564532 146940 564584 146946
rect 564532 146882 564584 146888
rect 564440 135176 564492 135182
rect 564440 135118 564492 135124
rect 564452 113830 564480 135118
rect 564544 127634 564572 146882
rect 564636 136610 564664 518910
rect 564728 335306 564756 700334
rect 567200 700324 567252 700330
rect 567200 700266 567252 700272
rect 565912 682032 565964 682038
rect 565912 681974 565964 681980
rect 565268 644496 565320 644502
rect 565268 644438 565320 644444
rect 564808 527196 564860 527202
rect 564808 527138 564860 527144
rect 564716 335300 564768 335306
rect 564716 335242 564768 335248
rect 564716 317552 564768 317558
rect 564716 317494 564768 317500
rect 564728 283626 564756 317494
rect 564716 283620 564768 283626
rect 564716 283562 564768 283568
rect 564728 277394 564756 283562
rect 564820 280158 564848 527138
rect 564992 280220 565044 280226
rect 564992 280162 565044 280168
rect 564808 280152 564860 280158
rect 564808 280094 564860 280100
rect 564728 277366 564940 277394
rect 564808 260908 564860 260914
rect 564808 260850 564860 260856
rect 564716 254040 564768 254046
rect 564716 253982 564768 253988
rect 564624 136604 564676 136610
rect 564624 136546 564676 136552
rect 564532 127628 564584 127634
rect 564532 127570 564584 127576
rect 564440 113824 564492 113830
rect 564440 113766 564492 113772
rect 564622 99512 564678 99521
rect 564622 99447 564678 99456
rect 564636 20398 564664 99447
rect 564728 24138 564756 253982
rect 564820 239902 564848 260850
rect 564808 239896 564860 239902
rect 564808 239838 564860 239844
rect 564912 239698 564940 277366
rect 564900 239692 564952 239698
rect 564900 239634 564952 239640
rect 564900 235952 564952 235958
rect 564900 235894 564952 235900
rect 564808 235748 564860 235754
rect 564808 235690 564860 235696
rect 564716 24132 564768 24138
rect 564716 24074 564768 24080
rect 564624 20392 564676 20398
rect 564624 20334 564676 20340
rect 564820 15910 564848 235690
rect 564912 16250 564940 235894
rect 565004 193905 565032 280162
rect 565174 231160 565230 231169
rect 565174 231095 565230 231104
rect 564990 193896 565046 193905
rect 564990 193831 565046 193840
rect 565084 155848 565136 155854
rect 565084 155790 565136 155796
rect 564992 151564 565044 151570
rect 564992 151506 565044 151512
rect 564900 16244 564952 16250
rect 564900 16186 564952 16192
rect 564808 15904 564860 15910
rect 564808 15846 564860 15852
rect 563440 6886 564020 6914
rect 563336 4072 563388 4078
rect 563336 4014 563388 4020
rect 561864 3732 561916 3738
rect 561864 3674 561916 3680
rect 559748 3460 559800 3466
rect 559748 3402 559800 3408
rect 559760 480 559788 3402
rect 563440 3244 563468 6886
rect 565004 6322 565032 151506
rect 565096 19174 565124 155790
rect 565188 149161 565216 231095
rect 565174 149152 565230 149161
rect 565174 149087 565230 149096
rect 565176 111852 565228 111858
rect 565176 111794 565228 111800
rect 565188 91798 565216 111794
rect 565176 91792 565228 91798
rect 565176 91734 565228 91740
rect 565280 29442 565308 644438
rect 565924 239601 565952 681974
rect 566740 666596 566792 666602
rect 566740 666538 566792 666544
rect 566280 503736 566332 503742
rect 566280 503678 566332 503684
rect 566188 501084 566240 501090
rect 566188 501026 566240 501032
rect 566004 454096 566056 454102
rect 566004 454038 566056 454044
rect 565910 239592 565966 239601
rect 565910 239527 565966 239536
rect 565912 167680 565964 167686
rect 565912 167622 565964 167628
rect 565360 155440 565412 155446
rect 565360 155382 565412 155388
rect 565268 29436 565320 29442
rect 565268 29378 565320 29384
rect 565084 19168 565136 19174
rect 565084 19110 565136 19116
rect 564992 6316 565044 6322
rect 564992 6258 565044 6264
rect 565372 3942 565400 155382
rect 565452 149796 565504 149802
rect 565452 149738 565504 149744
rect 565464 101454 565492 149738
rect 565820 149728 565872 149734
rect 565820 149670 565872 149676
rect 565832 136649 565860 149670
rect 565818 136640 565874 136649
rect 565818 136575 565874 136584
rect 565820 126948 565872 126954
rect 565820 126890 565872 126896
rect 565832 111858 565860 126890
rect 565820 111852 565872 111858
rect 565820 111794 565872 111800
rect 565452 101448 565504 101454
rect 565452 101390 565504 101396
rect 565924 16574 565952 167622
rect 566016 28558 566044 454038
rect 566096 415472 566148 415478
rect 566096 415414 566148 415420
rect 566108 29578 566136 415414
rect 566200 160818 566228 501026
rect 566292 236978 566320 503678
rect 566372 365832 566424 365838
rect 566372 365774 566424 365780
rect 566280 236972 566332 236978
rect 566280 236914 566332 236920
rect 566384 194410 566412 365774
rect 566464 335368 566516 335374
rect 566464 335310 566516 335316
rect 566476 194478 566504 335310
rect 566648 234252 566700 234258
rect 566648 234194 566700 234200
rect 566556 207052 566608 207058
rect 566556 206994 566608 207000
rect 566464 194472 566516 194478
rect 566464 194414 566516 194420
rect 566372 194404 566424 194410
rect 566372 194346 566424 194352
rect 566280 166524 566332 166530
rect 566280 166466 566332 166472
rect 566188 160812 566240 160818
rect 566188 160754 566240 160760
rect 566186 152688 566242 152697
rect 566186 152623 566242 152632
rect 566096 29572 566148 29578
rect 566096 29514 566148 29520
rect 566004 28552 566056 28558
rect 566004 28494 566056 28500
rect 565924 16546 566136 16574
rect 565360 3936 565412 3942
rect 565360 3878 565412 3884
rect 565820 3732 565872 3738
rect 565820 3674 565872 3680
rect 565832 3398 565860 3674
rect 566108 3482 566136 16546
rect 566200 5982 566228 152623
rect 566188 5976 566240 5982
rect 566188 5918 566240 5924
rect 566292 3738 566320 166466
rect 566372 152788 566424 152794
rect 566372 152730 566424 152736
rect 566384 6526 566412 152730
rect 566464 137760 566516 137766
rect 566464 137702 566516 137708
rect 566476 124914 566504 137702
rect 566464 124908 566516 124914
rect 566464 124850 566516 124856
rect 566568 70378 566596 206994
rect 566660 137358 566688 234194
rect 566648 137352 566700 137358
rect 566648 137294 566700 137300
rect 566556 70372 566608 70378
rect 566556 70314 566608 70320
rect 566752 28393 566780 666538
rect 567212 249762 567240 700266
rect 579066 697232 579122 697241
rect 579066 697167 579122 697176
rect 569960 687336 570012 687342
rect 569960 687278 570012 687284
rect 568764 686588 568816 686594
rect 568764 686530 568816 686536
rect 567936 683868 567988 683874
rect 567936 683810 567988 683816
rect 567292 682440 567344 682446
rect 567292 682382 567344 682388
rect 567304 313274 567332 682382
rect 567384 539640 567436 539646
rect 567384 539582 567436 539588
rect 567292 313268 567344 313274
rect 567292 313210 567344 313216
rect 567292 259548 567344 259554
rect 567292 259490 567344 259496
rect 567200 249756 567252 249762
rect 567200 249698 567252 249704
rect 567200 151020 567252 151026
rect 567200 150962 567252 150968
rect 567212 128246 567240 150962
rect 567200 128240 567252 128246
rect 567200 128182 567252 128188
rect 566738 28384 566794 28393
rect 566738 28319 566794 28328
rect 567304 25906 567332 259490
rect 567396 189786 567424 539582
rect 567568 514820 567620 514826
rect 567568 514762 567620 514768
rect 567476 342304 567528 342310
rect 567476 342246 567528 342252
rect 567384 189780 567436 189786
rect 567384 189722 567436 189728
rect 567384 155712 567436 155718
rect 567384 155654 567436 155660
rect 567292 25900 567344 25906
rect 567292 25842 567344 25848
rect 566372 6520 566424 6526
rect 566372 6462 566424 6468
rect 566280 3732 566332 3738
rect 566280 3674 566332 3680
rect 566108 3454 566872 3482
rect 565820 3392 565872 3398
rect 565820 3334 565872 3340
rect 563256 3216 563468 3244
rect 563256 480 563284 3216
rect 566844 480 566872 3454
rect 567396 3262 567424 155654
rect 567488 18902 567516 342246
rect 567580 237726 567608 514762
rect 567844 470620 567896 470626
rect 567844 470562 567896 470568
rect 567660 466472 567712 466478
rect 567660 466414 567712 466420
rect 567672 239766 567700 466414
rect 567752 263696 567804 263702
rect 567752 263638 567804 263644
rect 567764 240038 567792 263638
rect 567752 240032 567804 240038
rect 567752 239974 567804 239980
rect 567660 239760 567712 239766
rect 567660 239702 567712 239708
rect 567658 237960 567714 237969
rect 567658 237895 567714 237904
rect 567568 237720 567620 237726
rect 567568 237662 567620 237668
rect 567672 237538 567700 237895
rect 567580 237510 567700 237538
rect 567476 18896 567528 18902
rect 567476 18838 567528 18844
rect 567580 15706 567608 237510
rect 567660 235340 567712 235346
rect 567660 235282 567712 235288
rect 567672 235249 567700 235282
rect 567658 235240 567714 235249
rect 567658 235175 567714 235184
rect 567672 19854 567700 235175
rect 567752 166320 567804 166326
rect 567752 166262 567804 166268
rect 567764 82822 567792 166262
rect 567752 82816 567804 82822
rect 567752 82758 567804 82764
rect 567660 19848 567712 19854
rect 567660 19790 567712 19796
rect 567568 15700 567620 15706
rect 567568 15642 567620 15648
rect 567856 7614 567884 470562
rect 567948 139398 567976 683810
rect 568672 557592 568724 557598
rect 568672 557534 568724 557540
rect 568580 263628 568632 263634
rect 568580 263570 568632 263576
rect 568028 249824 568080 249830
rect 568028 249766 568080 249772
rect 567936 139392 567988 139398
rect 567936 139334 567988 139340
rect 567844 7608 567896 7614
rect 567844 7550 567896 7556
rect 568040 3534 568068 249766
rect 568592 240145 568620 263570
rect 568578 240136 568634 240145
rect 568578 240071 568634 240080
rect 568580 148368 568632 148374
rect 568580 148310 568632 148316
rect 568592 131102 568620 148310
rect 568580 131096 568632 131102
rect 568580 131038 568632 131044
rect 568684 24206 568712 557534
rect 568776 282878 568804 686530
rect 569408 611380 569460 611386
rect 569408 611322 569460 611328
rect 569224 560380 569276 560386
rect 569224 560322 569276 560328
rect 568948 425128 569000 425134
rect 568948 425070 569000 425076
rect 568856 390584 568908 390590
rect 568856 390526 568908 390532
rect 568764 282872 568816 282878
rect 568764 282814 568816 282820
rect 568764 235816 568816 235822
rect 568764 235758 568816 235764
rect 568672 24200 568724 24206
rect 568672 24142 568724 24148
rect 568776 18562 568804 235758
rect 568868 21622 568896 390526
rect 568960 150385 568988 425070
rect 569040 423768 569092 423774
rect 569040 423710 569092 423716
rect 569052 235346 569080 423710
rect 569132 325780 569184 325786
rect 569132 325722 569184 325728
rect 569040 235340 569092 235346
rect 569040 235282 569092 235288
rect 568946 150376 569002 150385
rect 568946 150311 569002 150320
rect 569144 142118 569172 325722
rect 569236 238270 569264 560322
rect 569316 252612 569368 252618
rect 569316 252554 569368 252560
rect 569224 238264 569276 238270
rect 569224 238206 569276 238212
rect 569328 195838 569356 252554
rect 569316 195832 569368 195838
rect 569316 195774 569368 195780
rect 569316 154352 569368 154358
rect 569316 154294 569368 154300
rect 569224 151428 569276 151434
rect 569224 151370 569276 151376
rect 569132 142112 569184 142118
rect 569132 142054 569184 142060
rect 569236 24750 569264 151370
rect 569328 89690 569356 154294
rect 569316 89684 569368 89690
rect 569316 89626 569368 89632
rect 569420 28082 569448 611322
rect 569592 285728 569644 285734
rect 569592 285670 569644 285676
rect 569498 157176 569554 157185
rect 569498 157111 569554 157120
rect 569408 28076 569460 28082
rect 569408 28018 569460 28024
rect 569224 24744 569276 24750
rect 569224 24686 569276 24692
rect 568856 21616 568908 21622
rect 568856 21558 568908 21564
rect 568764 18556 568816 18562
rect 568764 18498 568816 18504
rect 569512 6594 569540 157111
rect 569604 21418 569632 285670
rect 569592 21412 569644 21418
rect 569592 21354 569644 21360
rect 569500 6588 569552 6594
rect 569500 6530 569552 6536
rect 569972 6118 570000 687278
rect 571340 685092 571392 685098
rect 571340 685034 571392 685040
rect 570050 684584 570106 684593
rect 570050 684519 570106 684528
rect 570064 16046 570092 684519
rect 570604 682168 570656 682174
rect 570604 682110 570656 682116
rect 570144 534200 570196 534206
rect 570144 534142 570196 534148
rect 570156 18766 570184 534142
rect 570236 448588 570288 448594
rect 570236 448530 570288 448536
rect 570144 18760 570196 18766
rect 570144 18702 570196 18708
rect 570052 16040 570104 16046
rect 570052 15982 570104 15988
rect 569960 6112 570012 6118
rect 569960 6054 570012 6060
rect 570248 3806 570276 448530
rect 570512 300892 570564 300898
rect 570512 300834 570564 300840
rect 570328 264988 570380 264994
rect 570328 264930 570380 264936
rect 570340 238678 570368 264930
rect 570420 253972 570472 253978
rect 570420 253914 570472 253920
rect 570328 238672 570380 238678
rect 570328 238614 570380 238620
rect 570328 238264 570380 238270
rect 570328 238206 570380 238212
rect 570236 3800 570288 3806
rect 570236 3742 570288 3748
rect 568028 3528 568080 3534
rect 568028 3470 568080 3476
rect 567384 3256 567436 3262
rect 567384 3198 567436 3204
rect 570340 480 570368 238206
rect 570432 27538 570460 253914
rect 570524 173233 570552 300834
rect 570616 259418 570644 682110
rect 570696 643136 570748 643142
rect 570696 643078 570748 643084
rect 570708 506462 570736 643078
rect 570880 516180 570932 516186
rect 570880 516122 570932 516128
rect 570696 506456 570748 506462
rect 570696 506398 570748 506404
rect 570788 470620 570840 470626
rect 570788 470562 570840 470568
rect 570696 423700 570748 423706
rect 570696 423642 570748 423648
rect 570604 259412 570656 259418
rect 570604 259354 570656 259360
rect 570510 173224 570566 173233
rect 570510 173159 570566 173168
rect 570604 164076 570656 164082
rect 570604 164018 570656 164024
rect 570512 155236 570564 155242
rect 570512 155178 570564 155184
rect 570420 27532 570472 27538
rect 570420 27474 570472 27480
rect 570524 6390 570552 155178
rect 570616 21962 570644 164018
rect 570708 33114 570736 423642
rect 570800 238950 570828 470562
rect 570892 420238 570920 516122
rect 570880 420232 570932 420238
rect 570880 420174 570932 420180
rect 570880 278792 570932 278798
rect 570880 278734 570932 278740
rect 570788 238944 570840 238950
rect 570788 238886 570840 238892
rect 570892 198626 570920 278734
rect 570880 198620 570932 198626
rect 570880 198562 570932 198568
rect 570786 158128 570842 158137
rect 570786 158063 570842 158072
rect 570800 125526 570828 158063
rect 570788 125520 570840 125526
rect 570788 125462 570840 125468
rect 570696 33108 570748 33114
rect 570696 33050 570748 33056
rect 570604 21956 570656 21962
rect 570604 21898 570656 21904
rect 571352 17406 571380 685034
rect 576860 684820 576912 684826
rect 576860 684762 576912 684768
rect 572812 683732 572864 683738
rect 572812 683674 572864 683680
rect 571616 672104 571668 672110
rect 571616 672046 571668 672052
rect 571432 585200 571484 585206
rect 571432 585142 571484 585148
rect 571444 24274 571472 585142
rect 571524 520328 571576 520334
rect 571524 520270 571576 520276
rect 571536 25974 571564 520270
rect 571628 241194 571656 672046
rect 571984 610020 572036 610026
rect 571984 609962 572036 609968
rect 571996 525774 572024 609962
rect 571984 525768 572036 525774
rect 571984 525710 572036 525716
rect 572076 501016 572128 501022
rect 572076 500958 572128 500964
rect 571800 368552 571852 368558
rect 571800 368494 571852 368500
rect 571708 354748 571760 354754
rect 571708 354690 571760 354696
rect 571616 241188 571668 241194
rect 571616 241130 571668 241136
rect 571616 238196 571668 238202
rect 571616 238138 571668 238144
rect 571524 25968 571576 25974
rect 571524 25910 571576 25916
rect 571432 24268 571484 24274
rect 571432 24210 571484 24216
rect 571628 17474 571656 238138
rect 571720 25838 571748 354690
rect 571812 236502 571840 368494
rect 571984 360256 572036 360262
rect 571984 360198 572036 360204
rect 571892 299532 571944 299538
rect 571892 299474 571944 299480
rect 571800 236496 571852 236502
rect 571800 236438 571852 236444
rect 571904 177546 571932 299474
rect 571892 177540 571944 177546
rect 571892 177482 571944 177488
rect 571800 158364 571852 158370
rect 571800 158306 571852 158312
rect 571708 25832 571760 25838
rect 571708 25774 571760 25780
rect 571812 19786 571840 158306
rect 571892 156936 571944 156942
rect 571892 156878 571944 156884
rect 571904 75886 571932 156878
rect 571892 75880 571944 75886
rect 571892 75822 571944 75828
rect 571996 60722 572024 360198
rect 572088 325650 572116 500958
rect 572076 325644 572128 325650
rect 572076 325586 572128 325592
rect 572076 307828 572128 307834
rect 572076 307770 572128 307776
rect 572088 273222 572116 307770
rect 572168 296744 572220 296750
rect 572168 296686 572220 296692
rect 572076 273216 572128 273222
rect 572076 273158 572128 273164
rect 572076 228948 572128 228954
rect 572076 228890 572128 228896
rect 571984 60716 572036 60722
rect 571984 60658 572036 60664
rect 571800 19780 571852 19786
rect 571800 19722 571852 19728
rect 571616 17468 571668 17474
rect 571616 17410 571668 17416
rect 571340 17400 571392 17406
rect 571340 17342 571392 17348
rect 570512 6384 570564 6390
rect 570512 6326 570564 6332
rect 572088 3058 572116 228890
rect 572180 194546 572208 296686
rect 572168 194540 572220 194546
rect 572168 194482 572220 194488
rect 572168 154148 572220 154154
rect 572168 154090 572220 154096
rect 572180 110430 572208 154090
rect 572720 151088 572772 151094
rect 572720 151030 572772 151036
rect 572732 135250 572760 151030
rect 572720 135244 572772 135250
rect 572720 135186 572772 135192
rect 572168 110424 572220 110430
rect 572168 110366 572220 110372
rect 572824 16182 572852 683674
rect 573640 683460 573692 683466
rect 573640 683402 573692 683408
rect 572904 681216 572956 681222
rect 572904 681158 572956 681164
rect 572916 57934 572944 681158
rect 572996 505164 573048 505170
rect 572996 505106 573048 505112
rect 572904 57928 572956 57934
rect 572904 57870 572956 57876
rect 573008 21554 573036 505106
rect 573088 487212 573140 487218
rect 573088 487154 573140 487160
rect 572996 21548 573048 21554
rect 572996 21490 573048 21496
rect 573100 21486 573128 487154
rect 573272 459672 573324 459678
rect 573272 459614 573324 459620
rect 573180 346520 573232 346526
rect 573180 346462 573232 346468
rect 573192 25634 573220 346462
rect 573284 195634 573312 459614
rect 573364 443012 573416 443018
rect 573364 442954 573416 442960
rect 573376 239834 573404 442954
rect 573456 338156 573508 338162
rect 573456 338098 573508 338104
rect 573364 239828 573416 239834
rect 573364 239770 573416 239776
rect 573468 237046 573496 338098
rect 573548 251252 573600 251258
rect 573548 251194 573600 251200
rect 573456 237040 573508 237046
rect 573456 236982 573508 236988
rect 573364 235544 573416 235550
rect 573364 235486 573416 235492
rect 573272 195628 573324 195634
rect 573272 195570 573324 195576
rect 573272 151360 573324 151366
rect 573272 151302 573324 151308
rect 573180 25628 573232 25634
rect 573180 25570 573232 25576
rect 573088 21480 573140 21486
rect 573088 21422 573140 21428
rect 573284 17610 573312 151302
rect 573376 19310 573404 235486
rect 573560 182850 573588 251194
rect 573548 182844 573600 182850
rect 573548 182786 573600 182792
rect 573456 154216 573508 154222
rect 573456 154158 573508 154164
rect 573468 27402 573496 154158
rect 573456 27396 573508 27402
rect 573456 27338 573508 27344
rect 573364 19304 573416 19310
rect 573364 19246 573416 19252
rect 573272 17604 573324 17610
rect 573272 17546 573324 17552
rect 572812 16176 572864 16182
rect 572812 16118 572864 16124
rect 573652 4010 573680 683402
rect 575480 682304 575532 682310
rect 575480 682246 575532 682252
rect 574100 682100 574152 682106
rect 574100 682042 574152 682048
rect 574112 105505 574140 682042
rect 574744 681284 574796 681290
rect 574744 681226 574796 681232
rect 574284 640348 574336 640354
rect 574284 640290 574336 640296
rect 574192 568608 574244 568614
rect 574192 568550 574244 568556
rect 574098 105496 574154 105505
rect 574098 105431 574154 105440
rect 573640 4004 573692 4010
rect 573640 3946 573692 3952
rect 574204 3874 574232 568550
rect 574296 174554 574324 640290
rect 574468 465112 574520 465118
rect 574468 465054 574520 465060
rect 574376 353320 574428 353326
rect 574376 353262 574428 353268
rect 574284 174548 574336 174554
rect 574284 174490 574336 174496
rect 574284 156868 574336 156874
rect 574284 156810 574336 156816
rect 574296 19106 574324 156810
rect 574388 24546 574416 353262
rect 574480 191826 574508 465054
rect 574652 462392 574704 462398
rect 574652 462334 574704 462340
rect 574560 310616 574612 310622
rect 574560 310558 574612 310564
rect 574572 237250 574600 310558
rect 574664 240786 574692 462334
rect 574652 240780 574704 240786
rect 574652 240722 574704 240728
rect 574560 237244 574612 237250
rect 574560 237186 574612 237192
rect 574652 231056 574704 231062
rect 574652 230998 574704 231004
rect 574468 191820 574520 191826
rect 574468 191762 574520 191768
rect 574468 156664 574520 156670
rect 574468 156606 574520 156612
rect 574480 28422 574508 156606
rect 574468 28416 574520 28422
rect 574468 28358 574520 28364
rect 574376 24540 574428 24546
rect 574376 24482 574428 24488
rect 574284 19100 574336 19106
rect 574284 19042 574336 19048
rect 574192 3868 574244 3874
rect 574192 3810 574244 3816
rect 574664 3670 574692 230998
rect 574756 73166 574784 681226
rect 574836 426488 574888 426494
rect 574836 426430 574888 426436
rect 574744 73160 574796 73166
rect 574744 73102 574796 73108
rect 574848 4282 574876 426430
rect 574928 378208 574980 378214
rect 574928 378150 574980 378156
rect 574940 358766 574968 378150
rect 574928 358760 574980 358766
rect 574928 358702 574980 358708
rect 575020 247716 575072 247722
rect 575020 247658 575072 247664
rect 574926 157992 574982 158001
rect 574926 157927 574982 157936
rect 574940 92478 574968 157927
rect 574928 92472 574980 92478
rect 574928 92414 574980 92420
rect 575032 6458 575060 247658
rect 575492 97986 575520 682246
rect 575664 674892 575716 674898
rect 575664 674834 575716 674840
rect 575572 549296 575624 549302
rect 575572 549238 575624 549244
rect 575480 97980 575532 97986
rect 575480 97922 575532 97928
rect 575478 29200 575534 29209
rect 575478 29135 575480 29144
rect 575532 29135 575534 29144
rect 575480 29106 575532 29112
rect 575584 25537 575612 549238
rect 575676 193118 575704 674834
rect 576124 619676 576176 619682
rect 576124 619618 576176 619624
rect 575756 483064 575808 483070
rect 575756 483006 575808 483012
rect 575664 193112 575716 193118
rect 575664 193054 575716 193060
rect 575662 157040 575718 157049
rect 575662 156975 575718 156984
rect 575570 25528 575626 25537
rect 575570 25463 575626 25472
rect 575020 6452 575072 6458
rect 575020 6394 575072 6400
rect 574836 4276 574888 4282
rect 574836 4218 574888 4224
rect 574652 3664 574704 3670
rect 574652 3606 574704 3612
rect 575676 3466 575704 156975
rect 575768 15978 575796 483006
rect 575848 403028 575900 403034
rect 575848 402970 575900 402976
rect 575860 25702 575888 402970
rect 575940 309188 575992 309194
rect 575940 309130 575992 309136
rect 575952 28354 575980 309130
rect 576032 276072 576084 276078
rect 576032 276014 576084 276020
rect 575940 28348 575992 28354
rect 575940 28290 575992 28296
rect 576044 27062 576072 276014
rect 576136 181490 576164 619618
rect 576308 616888 576360 616894
rect 576308 616830 576360 616836
rect 576216 456816 576268 456822
rect 576216 456758 576268 456764
rect 576124 181484 576176 181490
rect 576124 181426 576176 181432
rect 576124 155372 576176 155378
rect 576124 155314 576176 155320
rect 576032 27056 576084 27062
rect 576032 26998 576084 27004
rect 575848 25696 575900 25702
rect 575848 25638 575900 25644
rect 575756 15972 575808 15978
rect 575756 15914 575808 15920
rect 576136 14890 576164 155314
rect 576228 113150 576256 456758
rect 576320 431934 576348 616830
rect 576308 431928 576360 431934
rect 576308 431870 576360 431876
rect 576308 316056 576360 316062
rect 576308 315998 576360 316004
rect 576320 240553 576348 315998
rect 576306 240544 576362 240553
rect 576306 240479 576362 240488
rect 576308 228676 576360 228682
rect 576308 228618 576360 228624
rect 576216 113144 576268 113150
rect 576216 113086 576268 113092
rect 576124 14884 576176 14890
rect 576124 14826 576176 14832
rect 576320 11762 576348 228618
rect 576308 11756 576360 11762
rect 576308 11698 576360 11704
rect 576872 3602 576900 684762
rect 576952 681964 577004 681970
rect 576952 681906 577004 681912
rect 576964 26081 576992 681906
rect 577228 681828 577280 681834
rect 577228 681770 577280 681776
rect 577136 680468 577188 680474
rect 577136 680410 577188 680416
rect 577044 679516 577096 679522
rect 577044 679458 577096 679464
rect 577056 28665 577084 679458
rect 577148 48278 577176 680410
rect 577240 96558 577268 681770
rect 577504 681760 577556 681766
rect 577504 681702 577556 681708
rect 577320 498228 577372 498234
rect 577320 498170 577372 498176
rect 577228 96552 577280 96558
rect 577228 96494 577280 96500
rect 577136 48272 577188 48278
rect 577136 48214 577188 48220
rect 577042 28656 577098 28665
rect 577042 28591 577098 28600
rect 576950 26072 577006 26081
rect 576950 26007 577006 26016
rect 577332 25809 577360 498170
rect 577412 478916 577464 478922
rect 577412 478858 577464 478864
rect 577318 25800 577374 25809
rect 577318 25735 577374 25744
rect 577424 18630 577452 478858
rect 577516 315382 577544 681702
rect 578884 612808 578936 612814
rect 578884 612750 578936 612756
rect 578332 469260 578384 469266
rect 578332 469202 578384 469208
rect 577596 327140 577648 327146
rect 577596 327082 577648 327088
rect 577504 315376 577556 315382
rect 577504 315318 577556 315324
rect 577504 270564 577556 270570
rect 577504 270506 577556 270512
rect 577516 27130 577544 270506
rect 577608 240106 577636 327082
rect 577688 310548 577740 310554
rect 577688 310490 577740 310496
rect 577596 240100 577648 240106
rect 577596 240042 577648 240048
rect 577700 237289 577728 310490
rect 577686 237280 577742 237289
rect 577686 237215 577742 237224
rect 577688 232756 577740 232762
rect 577688 232698 577740 232704
rect 577596 228404 577648 228410
rect 577596 228346 577648 228352
rect 577504 27124 577556 27130
rect 577504 27066 577556 27072
rect 577412 18624 577464 18630
rect 577412 18566 577464 18572
rect 577608 11830 577636 228346
rect 577700 17678 577728 232698
rect 578240 161016 578292 161022
rect 578240 160958 578292 160964
rect 578252 132462 578280 160958
rect 578240 132456 578292 132462
rect 578240 132398 578292 132404
rect 578344 66162 578372 469202
rect 578608 412684 578660 412690
rect 578608 412626 578660 412632
rect 578424 365764 578476 365770
rect 578424 365706 578476 365712
rect 578332 66156 578384 66162
rect 578332 66098 578384 66104
rect 578436 26042 578464 365706
rect 578516 288448 578568 288454
rect 578516 288390 578568 288396
rect 578528 26110 578556 288390
rect 578620 177682 578648 412626
rect 578792 389224 578844 389230
rect 578792 389166 578844 389172
rect 578700 346452 578752 346458
rect 578700 346394 578752 346400
rect 578712 237318 578740 346394
rect 578700 237312 578752 237318
rect 578700 237254 578752 237260
rect 578700 232960 578752 232966
rect 578700 232902 578752 232908
rect 578608 177676 578660 177682
rect 578608 177618 578660 177624
rect 578608 161152 578660 161158
rect 578608 161094 578660 161100
rect 578620 31074 578648 161094
rect 578608 31068 578660 31074
rect 578608 31010 578660 31016
rect 578516 26104 578568 26110
rect 578516 26046 578568 26052
rect 578424 26036 578476 26042
rect 578424 25978 578476 25984
rect 577688 17672 577740 17678
rect 577688 17614 577740 17620
rect 578712 13122 578740 232902
rect 578804 190466 578832 389166
rect 578792 190460 578844 190466
rect 578792 190402 578844 190408
rect 578792 160948 578844 160954
rect 578792 160890 578844 160896
rect 578804 96626 578832 160890
rect 578792 96620 578844 96626
rect 578792 96562 578844 96568
rect 578896 19825 578924 612750
rect 578976 586560 579028 586566
rect 578976 586502 579028 586508
rect 578882 19816 578938 19825
rect 578882 19751 578938 19760
rect 578700 13116 578752 13122
rect 578700 13058 578752 13064
rect 577596 11824 577648 11830
rect 577596 11766 577648 11772
rect 577412 4276 577464 4282
rect 577412 4218 577464 4224
rect 576860 3596 576912 3602
rect 576860 3538 576912 3544
rect 575664 3460 575716 3466
rect 575664 3402 575716 3408
rect 572076 3052 572128 3058
rect 572076 2994 572128 3000
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 577424 480 577452 4218
rect 578988 3330 579016 586502
rect 579080 405686 579108 697167
rect 582380 687268 582432 687274
rect 582380 687210 582432 687216
rect 580908 685908 580960 685914
rect 580908 685850 580960 685856
rect 580356 683324 580408 683330
rect 580356 683266 580408 683272
rect 579160 683188 579212 683194
rect 579160 683130 579212 683136
rect 579068 405680 579120 405686
rect 579068 405622 579120 405628
rect 579172 13462 579200 683130
rect 580264 681148 580316 681154
rect 580264 681090 580316 681096
rect 579620 677612 579672 677618
rect 579620 677554 579672 677560
rect 579632 23254 579660 677554
rect 579986 644056 580042 644065
rect 579986 643991 580042 644000
rect 580000 643142 580028 643991
rect 579988 643136 580040 643142
rect 579988 643078 580040 643084
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 579712 552084 579764 552090
rect 579712 552026 579764 552032
rect 579620 23248 579672 23254
rect 579620 23190 579672 23196
rect 579724 20097 579752 552026
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 579804 387864 579856 387870
rect 579804 387806 579856 387812
rect 579816 23186 579844 387806
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580080 334008 580132 334014
rect 580080 333950 580132 333956
rect 579896 317484 579948 317490
rect 579896 317426 579948 317432
rect 579908 28937 579936 317426
rect 579988 273284 580040 273290
rect 579988 273226 580040 273232
rect 579894 28928 579950 28937
rect 579894 28863 579950 28872
rect 579804 23180 579856 23186
rect 579804 23122 579856 23128
rect 579710 20088 579766 20097
rect 579710 20023 579766 20032
rect 580000 17270 580028 273226
rect 580092 237182 580120 333950
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580080 237176 580132 237182
rect 580080 237118 580132 237124
rect 580080 233912 580132 233918
rect 580080 233854 580132 233860
rect 580092 20534 580120 233854
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 681090
rect 580368 484673 580396 683266
rect 580448 681896 580500 681902
rect 580448 681838 580500 681844
rect 580460 537849 580488 681838
rect 580632 680604 580684 680610
rect 580632 680546 580684 680552
rect 580540 679652 580592 679658
rect 580540 679594 580592 679600
rect 580552 564369 580580 679594
rect 580644 577697 580672 680546
rect 580724 680536 580776 680542
rect 580724 680478 580776 680484
rect 580736 591025 580764 680478
rect 580816 679040 580868 679046
rect 580816 678982 580868 678988
rect 580828 617545 580856 678982
rect 580920 670721 580948 685850
rect 581092 684956 581144 684962
rect 581092 684898 581144 684904
rect 581000 684548 581052 684554
rect 581000 684490 581052 684496
rect 580906 670712 580962 670721
rect 580906 670647 580962 670656
rect 580814 617536 580870 617545
rect 580814 617471 580870 617480
rect 580722 591016 580778 591025
rect 580722 590951 580778 590960
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580538 564360 580594 564369
rect 580538 564295 580594 564304
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580354 484664 580410 484673
rect 580354 484599 580410 484608
rect 580448 420232 580500 420238
rect 580448 420174 580500 420180
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580368 234598 580396 418231
rect 580460 365129 580488 420174
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580448 315376 580500 315382
rect 580448 315318 580500 315324
rect 580356 234592 580408 234598
rect 580356 234534 580408 234540
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 580460 192545 580488 315318
rect 580538 312080 580594 312089
rect 580538 312015 580594 312024
rect 580552 239970 580580 312015
rect 580540 239964 580592 239970
rect 580540 239906 580592 239912
rect 580446 192536 580502 192545
rect 580446 192471 580502 192480
rect 580724 181484 580776 181490
rect 580724 181426 580776 181432
rect 580736 179217 580764 181426
rect 580722 179208 580778 179217
rect 580722 179143 580778 179152
rect 580264 161220 580316 161226
rect 580264 161162 580316 161168
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580170 152416 580226 152425
rect 580170 152351 580226 152360
rect 580080 20528 580132 20534
rect 580080 20470 580132 20476
rect 579988 17264 580040 17270
rect 579988 17206 580040 17212
rect 579160 13456 579212 13462
rect 579160 13398 579212 13404
rect 580184 12345 580212 152351
rect 580276 53786 580304 161162
rect 580356 153060 580408 153066
rect 580356 153002 580408 153008
rect 580368 77246 580396 153002
rect 580448 152516 580500 152522
rect 580448 152458 580500 152464
rect 580460 99521 580488 152458
rect 580540 139392 580592 139398
rect 580538 139360 580540 139369
rect 580592 139360 580594 139369
rect 580538 139295 580594 139304
rect 580540 113144 580592 113150
rect 580540 113086 580592 113092
rect 580552 112849 580580 113086
rect 580538 112840 580594 112849
rect 580538 112775 580594 112784
rect 580446 99512 580502 99521
rect 580446 99447 580502 99456
rect 580356 77240 580408 77246
rect 580356 77182 580408 77188
rect 580356 73160 580408 73166
rect 580356 73102 580408 73108
rect 580368 73001 580396 73102
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580356 60716 580408 60722
rect 580356 60658 580408 60664
rect 580368 59673 580396 60658
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580264 53780 580316 53786
rect 580264 53722 580316 53728
rect 580262 33144 580318 33153
rect 580262 33079 580264 33088
rect 580316 33079 580318 33088
rect 580264 33050 580316 33056
rect 581012 16153 581040 684490
rect 581104 28762 581132 684898
rect 581184 683392 581236 683398
rect 581184 683334 581236 683340
rect 581092 28756 581144 28762
rect 581092 28698 581144 28704
rect 581196 28626 581224 683334
rect 581552 534132 581604 534138
rect 581552 534074 581604 534080
rect 581460 492720 581512 492726
rect 581460 492662 581512 492668
rect 581276 459604 581328 459610
rect 581276 459546 581328 459552
rect 581184 28620 581236 28626
rect 581184 28562 581236 28568
rect 581288 23361 581316 459546
rect 581368 434784 581420 434790
rect 581368 434726 581420 434732
rect 581274 23352 581330 23361
rect 581274 23287 581330 23296
rect 581380 17882 581408 434726
rect 581472 154086 581500 492662
rect 581564 241330 581592 534074
rect 581828 394732 581880 394738
rect 581828 394674 581880 394680
rect 581644 325712 581696 325718
rect 581644 325654 581696 325660
rect 581552 241324 581604 241330
rect 581552 241266 581604 241272
rect 581552 214600 581604 214606
rect 581552 214542 581604 214548
rect 581460 154080 581512 154086
rect 581460 154022 581512 154028
rect 581368 17876 581420 17882
rect 581368 17818 581420 17824
rect 580998 16144 581054 16153
rect 580998 16079 581054 16088
rect 580170 12336 580226 12345
rect 580170 12271 580226 12280
rect 579804 7608 579856 7614
rect 579804 7550 579856 7556
rect 578976 3324 579028 3330
rect 578976 3266 579028 3272
rect 579816 480 579844 7550
rect 581564 6914 581592 214542
rect 581656 23390 581684 325654
rect 581736 231124 581788 231130
rect 581736 231066 581788 231072
rect 581644 23384 581696 23390
rect 581644 23326 581696 23332
rect 581748 16522 581776 231066
rect 581840 200977 581868 394674
rect 581826 200968 581882 200977
rect 581826 200903 581882 200912
rect 581828 160880 581880 160886
rect 581828 160822 581880 160828
rect 581840 95198 581868 160822
rect 581828 95192 581880 95198
rect 581828 95134 581880 95140
rect 581736 16516 581788 16522
rect 581736 16458 581788 16464
rect 581472 6886 581592 6914
rect 545212 60 545264 66
rect 545212 2 545264 8
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 354 581082 480
rect 581472 354 581500 6886
rect 582392 6662 582420 687210
rect 582472 685024 582524 685030
rect 582472 684966 582524 684972
rect 582484 15881 582512 684966
rect 582840 679108 582892 679114
rect 582840 679050 582892 679056
rect 582656 623824 582708 623830
rect 582656 623766 582708 623772
rect 582564 603152 582616 603158
rect 582564 603094 582616 603100
rect 582576 45558 582604 603094
rect 582668 71738 582696 623766
rect 582748 560312 582800 560318
rect 582748 560254 582800 560260
rect 582656 71732 582708 71738
rect 582656 71674 582708 71680
rect 582760 66230 582788 560254
rect 582852 189038 582880 679050
rect 582932 474768 582984 474774
rect 582932 474710 582984 474716
rect 582840 189032 582892 189038
rect 582840 188974 582892 188980
rect 582748 66224 582800 66230
rect 582748 66166 582800 66172
rect 582564 45552 582616 45558
rect 582564 45494 582616 45500
rect 582944 23050 582972 474710
rect 583024 444440 583076 444446
rect 583024 444382 583076 444388
rect 583036 29102 583064 444382
rect 583116 376780 583168 376786
rect 583116 376722 583168 376728
rect 583024 29096 583076 29102
rect 583024 29038 583076 29044
rect 583128 27266 583156 376722
rect 583208 350600 583260 350606
rect 583208 350542 583260 350548
rect 583116 27260 583168 27266
rect 583116 27202 583168 27208
rect 582932 23044 582984 23050
rect 582932 22986 582984 22992
rect 583220 20330 583248 350542
rect 583300 349172 583352 349178
rect 583300 349114 583352 349120
rect 583312 240009 583340 349114
rect 583392 313336 583444 313342
rect 583392 313278 583444 313284
rect 583298 240000 583354 240009
rect 583298 239935 583354 239944
rect 583300 211812 583352 211818
rect 583300 211754 583352 211760
rect 583208 20324 583260 20330
rect 583208 20266 583260 20272
rect 583312 16574 583340 211754
rect 583404 17950 583432 313278
rect 583484 305040 583536 305046
rect 583484 304982 583536 304988
rect 583496 28830 583524 304982
rect 583576 259480 583628 259486
rect 583576 259422 583628 259428
rect 583484 28824 583536 28830
rect 583484 28766 583536 28772
rect 583392 17944 583444 17950
rect 583392 17886 583444 17892
rect 583588 17814 583616 259422
rect 583668 244316 583720 244322
rect 583668 244258 583720 244264
rect 583576 17808 583628 17814
rect 583576 17750 583628 17756
rect 583312 16546 583432 16574
rect 582470 15872 582526 15881
rect 582470 15807 582526 15816
rect 582380 6656 582432 6662
rect 582380 6598 582432 6604
rect 582196 3324 582248 3330
rect 582196 3266 582248 3272
rect 582208 480 582236 3266
rect 583404 480 583432 16546
rect 583680 12442 583708 244258
rect 583760 231192 583812 231198
rect 583760 231134 583812 231140
rect 583772 13734 583800 231134
rect 583760 13728 583812 13734
rect 583760 13670 583812 13676
rect 583668 12436 583720 12442
rect 583668 12378 583720 12384
rect 580970 326 581500 354
rect 580970 -960 581082 326
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3330 658180 3332 658200
rect 3332 658180 3384 658200
rect 3384 658180 3386 658200
rect 3330 658144 3386 658180
rect 3238 566888 3294 566944
rect 3514 671200 3570 671256
rect 3606 619112 3662 619168
rect 3698 606056 3754 606112
rect 3698 588512 3754 588568
rect 3422 553832 3478 553888
rect 3422 501744 3478 501800
rect 3146 449520 3202 449576
rect 2962 410488 3018 410544
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3514 462576 3570 462632
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 4066 201864 4122 201920
rect 3422 197240 3478 197296
rect 4066 194384 4122 194440
rect 1398 192480 1454 192536
rect 2778 190984 2834 191040
rect 3422 188808 3478 188864
rect 3330 149776 3386 149832
rect 2870 97552 2926 97608
rect 3514 136720 3570 136776
rect 3514 84632 3570 84688
rect 3422 58520 3478 58576
rect 9678 680040 9734 680096
rect 3422 6432 3478 6488
rect 17866 584296 17922 584352
rect 19062 156576 19118 156632
rect 19154 152632 19210 152688
rect 19982 198600 20038 198656
rect 21270 198464 21326 198520
rect 25778 587424 25834 587480
rect 21914 23160 21970 23216
rect 20534 20304 20590 20360
rect 24674 565800 24730 565856
rect 24214 153720 24270 153776
rect 25870 587288 25926 587344
rect 25870 198192 25926 198248
rect 26054 561992 26110 562048
rect 30102 562128 30158 562184
rect 26882 158072 26938 158128
rect 27250 560904 27306 560960
rect 27250 194248 27306 194304
rect 27066 157936 27122 157992
rect 28814 561720 28870 561776
rect 27618 192752 27674 192808
rect 27526 29144 27582 29200
rect 24490 22888 24546 22944
rect 23294 22752 23350 22808
rect 22742 20440 22798 20496
rect 28630 152496 28686 152552
rect 28814 160656 28870 160712
rect 30286 560224 30342 560280
rect 30194 27376 30250 27432
rect 35254 679496 35310 679552
rect 34242 625912 34298 625968
rect 34150 622784 34206 622840
rect 34426 623736 34482 623792
rect 34334 598304 34390 598360
rect 34242 598032 34298 598088
rect 30286 24656 30342 24712
rect 31666 560632 31722 560688
rect 31758 171808 31814 171864
rect 31482 29280 31538 29336
rect 31298 29008 31354 29064
rect 33874 558728 33930 558784
rect 34150 561040 34206 561096
rect 33966 203496 34022 203552
rect 24214 3440 24270 3496
rect 34886 619928 34942 619984
rect 34426 570560 34482 570616
rect 34426 560768 34482 560824
rect 34334 196832 34390 196888
rect 89166 700304 89222 700360
rect 166906 676132 166908 676152
rect 166908 676132 166960 676152
rect 166960 676132 166962 676152
rect 166906 676096 166962 676132
rect 154486 674892 154542 674928
rect 154486 674872 154488 674892
rect 154488 674872 154540 674892
rect 154540 674872 154542 674892
rect 172610 668616 172666 668672
rect 35622 626864 35678 626920
rect 35438 621016 35494 621072
rect 35530 618160 35586 618216
rect 35714 599936 35770 599992
rect 35622 587152 35678 587208
rect 35806 220088 35862 220144
rect 35714 199008 35770 199064
rect 35622 198328 35678 198384
rect 84382 589464 84438 589520
rect 36542 198056 36598 198112
rect 36450 184456 36506 184512
rect 35990 3440 36046 3496
rect 38014 559952 38070 560008
rect 37186 199688 37242 199744
rect 37738 220768 37794 220824
rect 37738 205672 37794 205728
rect 38106 218048 38162 218104
rect 38290 198872 38346 198928
rect 38566 28600 38622 28656
rect 39210 199824 39266 199880
rect 39578 560088 39634 560144
rect 40774 510448 40830 510504
rect 40774 275984 40830 276040
rect 40682 204856 40738 204912
rect 40498 100000 40554 100056
rect 41234 189896 41290 189952
rect 41050 180240 41106 180296
rect 41878 199960 41934 200016
rect 41786 24792 41842 24848
rect 42982 205672 43038 205728
rect 43442 317328 43498 317384
rect 43994 563080 44050 563136
rect 44178 264832 44234 264888
rect 44178 220768 44234 220824
rect 44914 561312 44970 561368
rect 45006 359352 45062 359408
rect 44914 310256 44970 310312
rect 44822 283192 44878 283248
rect 44638 177656 44694 177712
rect 45190 339496 45246 339552
rect 45098 264696 45154 264752
rect 45098 244296 45154 244352
rect 45098 200504 45154 200560
rect 45098 155352 45154 155408
rect 45282 257896 45338 257952
rect 45650 525136 45706 525192
rect 46110 556144 46166 556200
rect 46110 546508 46166 546544
rect 46110 546488 46112 546508
rect 46112 546488 46164 546508
rect 46164 546488 46166 546508
rect 46018 545672 46074 545728
rect 46110 544312 46166 544368
rect 45926 544176 45982 544232
rect 46110 541048 46166 541104
rect 46110 538056 46166 538112
rect 46018 532208 46074 532264
rect 46110 529932 46112 529952
rect 46112 529932 46164 529952
rect 46164 529932 46166 529952
rect 46110 529896 46166 529932
rect 45834 528944 45890 529000
rect 46294 556552 46350 556608
rect 46294 551384 46350 551440
rect 46294 550860 46350 550896
rect 46294 550840 46296 550860
rect 46296 550840 46348 550860
rect 46348 550840 46350 550860
rect 46294 549752 46350 549808
rect 46202 526496 46258 526552
rect 46202 520376 46258 520432
rect 46018 516568 46074 516624
rect 45926 513848 45982 513904
rect 45742 510856 45798 510912
rect 46110 509496 46166 509552
rect 45650 500656 45706 500712
rect 45926 494536 45982 494592
rect 45834 484472 45890 484528
rect 45926 445032 45982 445088
rect 45926 439592 45982 439648
rect 45926 403552 45982 403608
rect 45926 345344 45982 345400
rect 45834 328752 45890 328808
rect 45834 264560 45890 264616
rect 45926 256672 45982 256728
rect 45834 242956 45890 242992
rect 45834 242936 45836 242956
rect 45836 242936 45888 242956
rect 45888 242936 45890 242956
rect 45650 234660 45706 234696
rect 45650 234640 45652 234660
rect 45652 234640 45704 234660
rect 45704 234640 45706 234660
rect 46110 506912 46166 506968
rect 46110 505164 46166 505200
rect 46110 505144 46112 505164
rect 46112 505144 46164 505164
rect 46164 505144 46166 505164
rect 46110 501336 46166 501392
rect 46110 496032 46166 496088
rect 46110 400288 46166 400344
rect 46110 373088 46166 373144
rect 45650 203632 45706 203688
rect 45558 202836 45614 202872
rect 45558 202816 45560 202836
rect 45560 202816 45612 202836
rect 45612 202816 45614 202836
rect 45742 201456 45798 201512
rect 46018 217232 46074 217288
rect 45926 195336 45982 195392
rect 45374 181464 45430 181520
rect 46294 489776 46350 489832
rect 46478 497256 46534 497312
rect 46478 495896 46534 495952
rect 46478 495216 46534 495272
rect 46478 493176 46534 493232
rect 46478 489932 46534 489968
rect 46478 489912 46480 489932
rect 46480 489912 46532 489932
rect 46532 489912 46534 489932
rect 46478 482296 46534 482352
rect 46386 480256 46442 480312
rect 46754 485852 46810 485888
rect 46754 485832 46756 485852
rect 46756 485832 46808 485852
rect 46808 485832 46810 485852
rect 46754 485152 46810 485208
rect 46754 480528 46810 480584
rect 46662 475496 46718 475552
rect 46570 474136 46626 474192
rect 46754 473456 46810 473512
rect 46754 469648 46810 469704
rect 46662 468288 46718 468344
rect 46754 468016 46810 468072
rect 46754 464208 46810 464264
rect 46754 463800 46810 463856
rect 46662 463256 46718 463312
rect 46754 460964 46810 461000
rect 46754 460944 46756 460964
rect 46756 460944 46808 460964
rect 46808 460944 46810 460964
rect 46478 445984 46534 446040
rect 46662 459856 46718 459912
rect 46754 456456 46810 456512
rect 46662 455776 46718 455832
rect 46754 450336 46810 450392
rect 46754 443264 46810 443320
rect 46570 442856 46626 442912
rect 46294 438776 46350 438832
rect 46754 436464 46810 436520
rect 46754 434732 46756 434752
rect 46756 434732 46808 434752
rect 46808 434732 46810 434752
rect 46754 434696 46810 434732
rect 46754 433608 46810 433664
rect 46386 431996 46442 432032
rect 46386 431976 46388 431996
rect 46388 431976 46440 431996
rect 46440 431976 46442 431996
rect 46386 429936 46442 429992
rect 46754 429256 46810 429312
rect 46754 427896 46810 427952
rect 46570 425312 46626 425368
rect 46478 421232 46534 421288
rect 46754 425176 46810 425232
rect 46662 424496 46718 424552
rect 46754 423700 46810 423736
rect 46754 423680 46756 423700
rect 46756 423680 46808 423700
rect 46808 423680 46810 423700
rect 46754 420980 46810 421016
rect 46754 420960 46756 420980
rect 46756 420960 46808 420980
rect 46808 420960 46810 420980
rect 46662 420008 46718 420064
rect 46754 419600 46810 419656
rect 46662 418648 46718 418704
rect 46754 418240 46810 418296
rect 46662 415928 46718 415984
rect 46754 415540 46810 415576
rect 46754 415520 46756 415540
rect 46756 415520 46808 415540
rect 46808 415520 46810 415540
rect 46754 414044 46810 414080
rect 46754 414024 46756 414044
rect 46756 414024 46808 414044
rect 46808 414024 46810 414044
rect 46570 411324 46626 411360
rect 46570 411304 46572 411324
rect 46572 411304 46624 411324
rect 46624 411304 46626 411324
rect 46570 407632 46626 407688
rect 46570 399472 46626 399528
rect 46478 396616 46534 396672
rect 46570 394984 46626 395040
rect 46570 393624 46626 393680
rect 46478 392672 46534 392728
rect 46570 392128 46626 392184
rect 46478 390904 46534 390960
rect 46570 390516 46626 390552
rect 46570 390496 46572 390516
rect 46572 390496 46624 390516
rect 46624 390496 46626 390516
rect 46570 389544 46626 389600
rect 46570 386436 46626 386472
rect 46570 386416 46572 386436
rect 46572 386416 46624 386436
rect 46624 386416 46626 386436
rect 46478 385736 46534 385792
rect 46570 385076 46626 385112
rect 46570 385056 46572 385076
rect 46572 385056 46624 385076
rect 46624 385056 46626 385076
rect 46570 382336 46626 382392
rect 46478 380976 46534 381032
rect 46570 379888 46626 379944
rect 46570 378256 46626 378312
rect 46478 374060 46534 374096
rect 46478 374040 46480 374060
rect 46480 374040 46532 374060
rect 46532 374040 46534 374060
rect 46478 372680 46534 372736
rect 46478 371456 46534 371512
rect 46478 369008 46534 369064
rect 46386 367648 46442 367704
rect 46478 366016 46534 366072
rect 46478 363432 46534 363488
rect 46478 357856 46534 357912
rect 46478 354748 46534 354784
rect 46478 354728 46480 354748
rect 46480 354728 46532 354748
rect 46532 354728 46534 354748
rect 46478 353096 46534 353152
rect 46478 349424 46534 349480
rect 46478 347112 46534 347168
rect 46478 336796 46534 336832
rect 46478 336776 46480 336796
rect 46480 336776 46532 336796
rect 46532 336776 46534 336796
rect 46386 329840 46442 329896
rect 46478 302912 46534 302968
rect 46478 292576 46534 292632
rect 46478 284280 46534 284336
rect 46386 252456 46442 252512
rect 46202 204312 46258 204368
rect 46202 201592 46258 201648
rect 46386 245384 46442 245440
rect 46386 222128 46442 222184
rect 46386 188808 46442 188864
rect 46570 254224 46626 254280
rect 46846 330656 46902 330712
rect 46846 327936 46902 327992
rect 46846 325216 46902 325272
rect 46846 323040 46902 323096
rect 46846 321680 46902 321736
rect 46846 320204 46902 320240
rect 46846 320184 46848 320204
rect 46848 320184 46900 320204
rect 46900 320184 46902 320204
rect 46846 318980 46902 319016
rect 46846 318960 46848 318980
rect 46848 318960 46900 318980
rect 46900 318960 46902 318980
rect 46846 318416 46902 318472
rect 46846 314744 46902 314800
rect 46846 310936 46902 310992
rect 46846 309188 46902 309224
rect 46846 309168 46848 309188
rect 46848 309168 46900 309188
rect 46900 309168 46902 309188
rect 46846 303728 46902 303784
rect 46846 302132 46848 302152
rect 46848 302132 46900 302152
rect 46900 302132 46902 302152
rect 46846 302096 46902 302132
rect 46846 300892 46902 300928
rect 46846 300872 46848 300892
rect 46848 300872 46900 300892
rect 46900 300872 46902 300892
rect 46846 298172 46902 298208
rect 46846 298152 46848 298172
rect 46848 298152 46900 298172
rect 46900 298152 46902 298172
rect 46846 296792 46902 296848
rect 46846 292848 46902 292904
rect 46846 291488 46902 291544
rect 46846 288496 46902 288552
rect 46846 285776 46902 285832
rect 46938 285232 46994 285288
rect 46846 281580 46902 281616
rect 46846 281560 46848 281580
rect 46848 281560 46900 281580
rect 46900 281560 46902 281580
rect 46846 277752 46902 277808
rect 46846 268232 46902 268288
rect 46754 247560 46810 247616
rect 46754 247424 46810 247480
rect 46754 245792 46810 245848
rect 46662 244296 46718 244352
rect 46570 226616 46626 226672
rect 46662 221312 46718 221368
rect 46570 218592 46626 218648
rect 46846 238176 46902 238232
rect 46846 237496 46902 237552
rect 46846 236000 46902 236056
rect 46846 232328 46902 232384
rect 46846 230560 46902 230616
rect 46846 227840 46902 227896
rect 47214 376216 47270 376272
rect 47214 335416 47270 335472
rect 47122 270136 47178 270192
rect 47030 233416 47086 233472
rect 47030 230832 47086 230888
rect 46846 224032 46902 224088
rect 46846 222400 46902 222456
rect 46846 221040 46902 221096
rect 46846 218068 46902 218104
rect 46846 218048 46848 218068
rect 46848 218048 46900 218068
rect 46900 218048 46902 218068
rect 46846 215348 46902 215384
rect 46846 215328 46848 215348
rect 46848 215328 46900 215348
rect 46900 215328 46902 215348
rect 46846 213988 46902 214024
rect 46846 213968 46848 213988
rect 46848 213968 46900 213988
rect 46900 213968 46902 213988
rect 46846 211248 46902 211304
rect 46846 207576 46902 207632
rect 46846 206932 46848 206952
rect 46848 206932 46900 206952
rect 46900 206932 46902 206952
rect 46846 206896 46902 206932
rect 46846 205692 46902 205728
rect 46846 205672 46848 205692
rect 46848 205672 46900 205692
rect 46900 205672 46902 205692
rect 46662 178744 46718 178800
rect 46478 156712 46534 156768
rect 46386 155896 46442 155952
rect 46662 11600 46718 11656
rect 43074 3440 43130 3496
rect 47490 521736 47546 521792
rect 47398 504056 47454 504112
rect 47306 298016 47362 298072
rect 47398 281832 47454 281888
rect 47306 273264 47362 273320
rect 47490 259528 47546 259584
rect 47490 241440 47546 241496
rect 47490 216688 47546 216744
rect 52458 587832 52514 587888
rect 53838 587832 53894 587888
rect 56598 587832 56654 587888
rect 57886 587832 57942 587888
rect 58070 587832 58126 587888
rect 59358 587832 59414 587888
rect 62118 587832 62174 587888
rect 63498 587832 63554 587888
rect 63682 587832 63738 587888
rect 64970 587832 65026 587888
rect 66350 587832 66406 587888
rect 67638 587832 67694 587888
rect 69018 587832 69074 587888
rect 70398 587832 70454 587888
rect 71778 587832 71834 587888
rect 72422 587832 72478 587888
rect 74630 587832 74686 587888
rect 77298 587832 77354 587888
rect 78678 587832 78734 587888
rect 48962 561720 49018 561776
rect 49606 560244 49662 560280
rect 49606 560224 49608 560244
rect 49608 560224 49660 560244
rect 49660 560224 49662 560244
rect 51078 559952 51134 560008
rect 56506 587696 56562 587752
rect 56506 578856 56562 578912
rect 51630 560088 51686 560144
rect 57426 562128 57482 562184
rect 57978 561992 58034 562048
rect 59174 562128 59230 562184
rect 58070 560904 58126 560960
rect 59266 561992 59322 562048
rect 62026 587696 62082 587752
rect 59818 564440 59874 564496
rect 59266 561176 59322 561232
rect 59910 561856 59966 561912
rect 63590 587696 63646 587752
rect 63222 560496 63278 560552
rect 67546 586336 67602 586392
rect 64970 561040 65026 561096
rect 70306 587696 70362 587752
rect 70306 571920 70362 571976
rect 73066 587696 73122 587752
rect 74538 587696 74594 587752
rect 72422 581576 72478 581632
rect 74446 587560 74502 587616
rect 77206 587696 77262 587752
rect 77114 586336 77170 586392
rect 78770 587696 78826 587752
rect 77758 568656 77814 568712
rect 79782 587832 79838 587888
rect 81162 587832 81218 587888
rect 81806 587832 81862 587888
rect 82910 587832 82966 587888
rect 81898 587696 81954 587752
rect 85486 586336 85542 586392
rect 87142 587832 87198 587888
rect 88338 587832 88394 587888
rect 91098 587832 91154 587888
rect 93122 587832 93178 587888
rect 93858 587832 93914 587888
rect 95146 587832 95202 587888
rect 99470 587832 99526 587888
rect 101954 587832 102010 587888
rect 106922 587832 106978 587888
rect 109038 587832 109094 587888
rect 111798 587832 111854 587888
rect 115202 587832 115258 587888
rect 118698 587832 118754 587888
rect 124402 587832 124458 587888
rect 128358 587832 128414 587888
rect 131762 587832 131818 587888
rect 133970 587832 134026 587888
rect 136638 587832 136694 587888
rect 139398 587832 139454 587888
rect 86958 587696 87014 587752
rect 86866 586336 86922 586392
rect 85486 567160 85542 567216
rect 83094 563216 83150 563272
rect 86314 562400 86370 562456
rect 87050 586336 87106 586392
rect 89626 586336 89682 586392
rect 91006 586336 91062 586392
rect 92386 586336 92442 586392
rect 93122 582936 93178 582992
rect 92386 576000 92442 576056
rect 95238 587696 95294 587752
rect 97906 586336 97962 586392
rect 104806 586336 104862 586392
rect 89718 562264 89774 562320
rect 117226 586336 117282 586392
rect 106094 567296 106150 567352
rect 109590 565936 109646 565992
rect 128266 587696 128322 587752
rect 122746 586336 122802 586392
rect 141974 587832 142030 587888
rect 159086 587832 159142 587888
rect 125690 562128 125746 562184
rect 160006 586336 160062 586392
rect 153842 563624 153898 563680
rect 157798 566072 157854 566128
rect 164330 562536 164386 562592
rect 170770 561992 170826 562048
rect 328550 674908 328552 674928
rect 328552 674908 328604 674928
rect 328604 674908 328606 674928
rect 328550 674872 328606 674908
rect 329746 674892 329802 674928
rect 329746 674872 329748 674892
rect 329748 674872 329800 674892
rect 329800 674872 329802 674892
rect 340878 674872 340934 674928
rect 208306 626592 208362 626648
rect 207662 625368 207718 625424
rect 175278 608776 175334 608832
rect 176566 607280 176622 607336
rect 176566 605920 176622 605976
rect 175370 604424 175426 604480
rect 175462 603064 175518 603120
rect 190366 566208 190422 566264
rect 174542 561856 174598 561912
rect 188710 563352 188766 563408
rect 189446 561992 189502 562048
rect 195886 564576 195942 564632
rect 192574 562128 192630 562184
rect 207018 599392 207074 599448
rect 207754 623736 207810 623792
rect 208214 622376 208270 622432
rect 208122 621016 208178 621072
rect 208030 617616 208086 617672
rect 207938 597624 207994 597680
rect 209686 619928 209742 619984
rect 209134 598304 209190 598360
rect 224958 587832 225014 587888
rect 207478 560904 207534 560960
rect 227810 587832 227866 587888
rect 231674 587832 231730 587888
rect 234526 587832 234582 587888
rect 235998 587832 236054 587888
rect 237378 587832 237434 587888
rect 238666 587832 238722 587888
rect 238850 587832 238906 587888
rect 231766 586336 231822 586392
rect 233146 586336 233202 586392
rect 234618 587696 234674 587752
rect 238758 586764 238814 586800
rect 238758 586744 238760 586764
rect 238760 586744 238812 586764
rect 238812 586744 238814 586764
rect 257342 588920 257398 588976
rect 240506 587832 240562 587888
rect 242438 587832 242494 587888
rect 243542 587832 243598 587888
rect 245566 587832 245622 587888
rect 245842 587832 245898 587888
rect 247038 587832 247094 587888
rect 248142 587832 248198 587888
rect 248418 587832 248474 587888
rect 249706 587832 249762 587888
rect 252650 587832 252706 587888
rect 253938 587832 253994 587888
rect 255318 587832 255374 587888
rect 256606 587832 256662 587888
rect 240782 587696 240838 587752
rect 246946 587696 247002 587752
rect 244186 586336 244242 586392
rect 241426 566344 241482 566400
rect 240046 562264 240102 562320
rect 249798 587696 249854 587752
rect 252558 587696 252614 587752
rect 252466 586336 252522 586392
rect 257986 587832 258042 587888
rect 260654 587832 260710 587888
rect 261022 587832 261078 587888
rect 262034 587832 262090 587888
rect 262218 587832 262274 587888
rect 264886 587832 264942 587888
rect 266266 587832 266322 587888
rect 268934 587832 268990 587888
rect 269762 587832 269818 587888
rect 270498 587832 270554 587888
rect 273534 587832 273590 587888
rect 274638 587832 274694 587888
rect 281078 587832 281134 587888
rect 282918 587832 282974 587888
rect 286322 587832 286378 587888
rect 288438 587832 288494 587888
rect 291014 587832 291070 587888
rect 252650 569200 252706 569256
rect 258170 586744 258226 586800
rect 258078 586336 258134 586392
rect 264426 587696 264482 587752
rect 263506 586336 263562 586392
rect 260746 563488 260802 563544
rect 264978 587696 265034 587752
rect 267646 586336 267702 586392
rect 269026 586336 269082 586392
rect 277490 586472 277546 586528
rect 270498 577496 270554 577552
rect 268014 560768 268070 560824
rect 288438 583072 288494 583128
rect 298098 587832 298154 587888
rect 300858 587832 300914 587888
rect 302238 587832 302294 587888
rect 305090 587832 305146 587888
rect 308494 587832 308550 587888
rect 310518 587832 310574 587888
rect 313278 587832 313334 587888
rect 316038 587832 316094 587888
rect 293866 586336 293922 586392
rect 296626 586336 296682 586392
rect 277490 570696 277546 570752
rect 274454 562536 274510 562592
rect 289174 568792 289230 568848
rect 294326 562672 294382 562728
rect 297638 564712 297694 564768
rect 305090 574640 305146 574696
rect 308034 562400 308090 562456
rect 333886 587832 333942 587888
rect 333794 586336 333850 586392
rect 313278 567840 313334 567896
rect 315578 559952 315634 560008
rect 322110 564848 322166 564904
rect 328366 563624 328422 563680
rect 330482 560632 330538 560688
rect 335358 567432 335414 567488
rect 336370 561040 336426 561096
rect 339406 560360 339462 560416
rect 341982 561720 342038 561776
rect 349158 669160 349214 669216
rect 347870 522824 347926 522880
rect 347778 477944 347834 478000
rect 347778 474952 347834 475008
rect 47766 229336 47822 229392
rect 47766 226344 47822 226400
rect 47766 220224 47822 220280
rect 347686 200912 347742 200968
rect 347686 200232 347742 200288
rect 47858 199552 47914 199608
rect 48686 187040 48742 187096
rect 48686 149096 48742 149152
rect 53838 198192 53894 198248
rect 50434 177520 50490 177576
rect 50342 124072 50398 124128
rect 51722 155488 51778 155544
rect 51722 147736 51778 147792
rect 51814 147600 51870 147656
rect 51538 142024 51594 142080
rect 51538 124072 51594 124128
rect 52182 142160 52238 142216
rect 52366 146512 52422 146568
rect 50158 3440 50214 3496
rect 53746 135904 53802 135960
rect 53746 124752 53802 124808
rect 53654 25472 53710 25528
rect 56138 195472 56194 195528
rect 54666 122032 54722 122088
rect 55034 29688 55090 29744
rect 55770 151136 55826 151192
rect 55862 98096 55918 98152
rect 55954 77016 56010 77072
rect 56322 184320 56378 184376
rect 56230 148960 56286 149016
rect 56138 70216 56194 70272
rect 56046 41656 56102 41712
rect 56322 54576 56378 54632
rect 56690 141616 56746 141672
rect 56690 140256 56746 140312
rect 56690 125296 56746 125352
rect 56598 107616 56654 107672
rect 56874 159568 56930 159624
rect 57794 159296 57850 159352
rect 56966 158480 57022 158536
rect 57518 153992 57574 154048
rect 57242 139576 57298 139632
rect 56966 119856 57022 119912
rect 56966 117952 57022 118008
rect 57058 117136 57114 117192
rect 56874 113056 56930 113112
rect 56874 104216 56930 104272
rect 57426 120536 57482 120592
rect 57426 119176 57482 119232
rect 57426 115096 57482 115152
rect 57426 114452 57428 114472
rect 57428 114452 57480 114472
rect 57480 114452 57482 114472
rect 57426 114416 57482 114452
rect 57150 90616 57206 90672
rect 57150 68176 57206 68232
rect 56782 55936 56838 55992
rect 57150 47096 57206 47152
rect 57058 46416 57114 46472
rect 57150 45056 57206 45112
rect 56690 40976 56746 41032
rect 56414 32136 56470 32192
rect 57610 143520 57666 143576
rect 57610 137536 57666 137592
rect 57610 134816 57666 134872
rect 57610 132776 57666 132832
rect 57610 131416 57666 131472
rect 57610 130736 57666 130792
rect 57610 129376 57666 129432
rect 57610 128016 57666 128072
rect 57610 126656 57666 126712
rect 57610 123256 57666 123312
rect 57242 19216 57298 19272
rect 57518 110336 57574 110392
rect 57518 108296 57574 108352
rect 57518 103536 57574 103592
rect 57518 102856 57574 102912
rect 57518 101496 57574 101552
rect 57518 99456 57574 99512
rect 57518 94016 57574 94072
rect 57518 92656 57574 92712
rect 57610 89256 57666 89312
rect 57610 86536 57666 86592
rect 57886 145696 57942 145752
rect 57794 142976 57850 143032
rect 58070 124072 58126 124128
rect 57886 102176 57942 102232
rect 57610 82456 57666 82512
rect 57518 81776 57574 81832
rect 57610 75656 57666 75712
rect 57518 21664 57574 21720
rect 57886 81096 57942 81152
rect 57886 68856 57942 68912
rect 57886 67532 57888 67552
rect 57888 67532 57940 67552
rect 57940 67532 57942 67552
rect 57886 67496 57942 67532
rect 57886 64096 57942 64152
rect 57886 63452 57888 63472
rect 57888 63452 57940 63472
rect 57940 63452 57942 63472
rect 57886 63416 57942 63452
rect 57886 62076 57942 62112
rect 57886 62056 57888 62076
rect 57888 62056 57940 62076
rect 57940 62056 57942 62076
rect 57886 58656 57942 58712
rect 57886 57296 57942 57352
rect 57886 55256 57942 55312
rect 57886 40296 57942 40352
rect 57886 39616 57942 39672
rect 57886 33496 57942 33552
rect 57886 32816 57942 32872
rect 58254 115776 58310 115832
rect 58162 45736 58218 45792
rect 58990 197104 59046 197160
rect 60278 195744 60334 195800
rect 59082 144880 59138 144936
rect 59450 151680 59506 151736
rect 59634 151680 59690 151736
rect 59542 150048 59598 150104
rect 59726 151408 59782 151464
rect 59726 151272 59782 151328
rect 59726 148960 59782 149016
rect 59634 147600 59690 147656
rect 58898 143520 58954 143576
rect 59266 139168 59322 139224
rect 58898 136584 58954 136640
rect 58898 111832 58954 111888
rect 59082 137264 59138 137320
rect 59266 125432 59322 125488
rect 59266 120128 59322 120184
rect 60002 151408 60058 151464
rect 61934 153040 61990 153096
rect 60002 150048 60058 150104
rect 59910 149912 59966 149968
rect 68006 186904 68062 186960
rect 73342 177248 73398 177304
rect 72882 152360 72938 152416
rect 77390 179968 77446 180024
rect 77390 167592 77446 167648
rect 83462 198736 83518 198792
rect 82818 198328 82874 198384
rect 94410 198328 94466 198384
rect 93122 197920 93178 197976
rect 108302 180648 108358 180704
rect 110418 160792 110474 160848
rect 111890 153856 111946 153912
rect 120170 196968 120226 197024
rect 122746 198192 122802 198248
rect 117318 151272 117374 151328
rect 133050 194112 133106 194168
rect 139398 192888 139454 192944
rect 146298 192888 146354 192944
rect 147678 181600 147734 181656
rect 153658 198056 153714 198112
rect 158166 191664 158222 191720
rect 153382 152632 153438 152688
rect 157890 170312 157946 170368
rect 170402 198056 170458 198112
rect 174910 199008 174966 199064
rect 172058 179832 172114 179888
rect 168378 153040 168434 153096
rect 170126 152768 170182 152824
rect 179142 152768 179198 152824
rect 187790 196696 187846 196752
rect 196806 193976 196862 194032
rect 195242 172352 195298 172408
rect 200026 199008 200082 199064
rect 208122 197920 208178 197976
rect 199106 152632 199162 152688
rect 204902 152904 204958 152960
rect 211986 190304 212042 190360
rect 235170 196560 235226 196616
rect 240966 152496 241022 152552
rect 251270 162016 251326 162072
rect 257894 198872 257950 198928
rect 270590 196560 270646 196616
rect 271234 163376 271290 163432
rect 278594 191528 278650 191584
rect 317602 155760 317658 155816
rect 59082 96736 59138 96792
rect 58990 53216 59046 53272
rect 321466 163648 321522 163704
rect 330758 194248 330814 194304
rect 329194 180512 329250 180568
rect 325054 152496 325110 152552
rect 334070 158616 334126 158672
rect 346122 199280 346178 199336
rect 342350 196832 342406 196888
rect 341798 152904 341854 152960
rect 347594 199552 347650 199608
rect 347686 198464 347742 198520
rect 348330 523504 348386 523560
rect 348238 456456 348294 456512
rect 348146 433336 348202 433392
rect 348146 396616 348202 396672
rect 348054 390632 348110 390688
rect 347962 377032 348018 377088
rect 347962 368464 348018 368520
rect 347870 275984 347926 276040
rect 348330 295976 348386 296032
rect 350446 609320 350502 609376
rect 349250 607688 349306 607744
rect 350446 606328 350502 606384
rect 350446 604832 350502 604888
rect 349342 603608 349398 603664
rect 349158 541456 349214 541512
rect 348882 433200 348938 433256
rect 349158 489776 349214 489832
rect 348698 200232 348754 200288
rect 349434 554376 349490 554432
rect 349434 532072 349490 532128
rect 349342 451696 349398 451752
rect 349250 346976 349306 347032
rect 349158 299376 349214 299432
rect 349618 499976 349674 500032
rect 349526 409536 349582 409592
rect 349434 296656 349490 296712
rect 349342 279656 349398 279712
rect 349710 470736 349766 470792
rect 349710 456864 349766 456920
rect 349618 336096 349674 336152
rect 349618 280472 349674 280528
rect 349434 262792 349490 262848
rect 349250 262656 349306 262712
rect 349158 233824 349214 233880
rect 348698 198872 348754 198928
rect 349526 258712 349582 258768
rect 349526 210024 349582 210080
rect 349342 202272 349398 202328
rect 350170 547032 350226 547088
rect 350170 533432 350226 533488
rect 349894 521736 349950 521792
rect 350078 516568 350134 516624
rect 350078 513460 350134 513496
rect 350078 513440 350080 513460
rect 350080 513440 350132 513460
rect 350132 513440 350134 513460
rect 349986 506912 350042 506968
rect 350078 505552 350134 505608
rect 349986 485152 350042 485208
rect 350078 480664 350134 480720
rect 350078 476448 350134 476504
rect 350078 465976 350134 466032
rect 350078 462848 350134 462904
rect 350078 461352 350134 461408
rect 349802 455776 349858 455832
rect 350078 445848 350134 445904
rect 350078 437824 350134 437880
rect 350078 430888 350134 430944
rect 350078 421232 350134 421288
rect 350078 404912 350134 404968
rect 350078 395392 350134 395448
rect 349802 394848 349858 394904
rect 350078 391312 350134 391368
rect 349986 356632 350042 356688
rect 350170 343984 350226 344040
rect 349894 331200 349950 331256
rect 350170 319096 350226 319152
rect 350170 315152 350226 315208
rect 349894 302912 349950 302968
rect 349710 257896 349766 257952
rect 349710 200504 349766 200560
rect 350078 288496 350134 288552
rect 350446 551112 350502 551168
rect 350446 546508 350502 546544
rect 350446 546488 350448 546508
rect 350448 546488 350500 546508
rect 350500 546488 350502 546508
rect 350446 542952 350502 543008
rect 350446 538328 350502 538384
rect 350446 536852 350502 536888
rect 350446 536832 350448 536852
rect 350448 536832 350500 536852
rect 350500 536832 350502 536852
rect 350446 534656 350502 534712
rect 350446 532772 350502 532808
rect 350446 532752 350448 532772
rect 350448 532752 350500 532772
rect 350500 532752 350502 532772
rect 350446 530712 350502 530768
rect 350446 527196 350502 527232
rect 350446 527176 350448 527196
rect 350448 527176 350500 527196
rect 350500 527176 350502 527196
rect 350446 525972 350502 526008
rect 350446 525952 350448 525972
rect 350448 525952 350500 525972
rect 350500 525952 350502 525972
rect 350446 523232 350502 523288
rect 350538 522960 350594 523016
rect 350446 517540 350502 517576
rect 350446 517520 350448 517540
rect 350448 517520 350500 517540
rect 350500 517520 350502 517540
rect 350446 516316 350502 516352
rect 350446 516296 350448 516316
rect 350448 516296 350500 516316
rect 350500 516296 350502 516316
rect 350446 513712 350502 513768
rect 350446 511536 350502 511592
rect 350446 508816 350502 508872
rect 350446 505416 350502 505472
rect 350446 503784 350502 503840
rect 350446 500112 350502 500168
rect 350446 498228 350502 498264
rect 350446 498208 350448 498228
rect 350448 498208 350500 498228
rect 350500 498208 350502 498228
rect 350446 495508 350502 495544
rect 350446 495488 350448 495508
rect 350448 495488 350500 495508
rect 350500 495488 350502 495508
rect 350446 494556 350502 494592
rect 350446 494536 350448 494556
rect 350448 494536 350500 494556
rect 350500 494536 350502 494556
rect 350354 493856 350410 493912
rect 350354 491952 350410 492008
rect 350446 491408 350502 491464
rect 350446 490048 350502 490104
rect 350446 487736 350502 487792
rect 350446 483112 350502 483168
rect 350446 481652 350448 481672
rect 350448 481652 350500 481672
rect 350500 481652 350502 481672
rect 350446 481616 350502 481652
rect 350446 480276 350502 480312
rect 350446 480256 350448 480276
rect 350448 480256 350500 480276
rect 350500 480256 350502 480276
rect 350446 476176 350502 476232
rect 350446 473456 350502 473512
rect 350446 466520 350502 466576
rect 350446 465160 350502 465216
rect 350446 462440 350502 462496
rect 350446 461080 350502 461136
rect 350446 459604 350502 459640
rect 350446 459584 350448 459604
rect 350448 459584 350500 459604
rect 350500 459584 350502 459604
rect 350446 457292 350502 457328
rect 350446 457272 350448 457292
rect 350448 457272 350500 457292
rect 350500 457272 350502 457292
rect 350446 454164 350502 454200
rect 350446 454144 350448 454164
rect 350448 454144 350500 454164
rect 350500 454144 350502 454164
rect 350446 451832 350502 451888
rect 350446 451016 350502 451072
rect 350446 449948 350502 449984
rect 350446 449928 350448 449948
rect 350448 449928 350500 449948
rect 350500 449928 350502 449948
rect 350446 447752 350502 447808
rect 350446 446392 350502 446448
rect 350446 445576 350502 445632
rect 350446 441652 350502 441688
rect 350446 441632 350448 441652
rect 350448 441632 350500 441652
rect 350500 441632 350502 441652
rect 350446 440292 350502 440328
rect 350446 440272 350448 440292
rect 350448 440272 350500 440292
rect 350500 440272 350502 440292
rect 350446 436736 350502 436792
rect 350446 434732 350448 434752
rect 350448 434732 350500 434752
rect 350500 434732 350502 434752
rect 350446 434696 350502 434732
rect 350446 430652 350448 430672
rect 350448 430652 350500 430672
rect 350500 430652 350502 430672
rect 350446 430616 350502 430652
rect 350446 427896 350502 427952
rect 350446 426536 350502 426592
rect 350446 425312 350502 425368
rect 350446 422340 350502 422376
rect 350446 422320 350448 422340
rect 350448 422320 350500 422340
rect 350500 422320 350502 422340
rect 350446 420980 350502 421016
rect 350446 420960 350448 420980
rect 350448 420960 350500 420980
rect 350500 420960 350502 420980
rect 350446 419600 350502 419656
rect 350446 418376 350502 418432
rect 350446 416880 350502 416936
rect 350446 414452 350502 414488
rect 350446 414432 350448 414452
rect 350448 414432 350500 414452
rect 350500 414432 350502 414452
rect 350446 414044 350502 414080
rect 350446 414024 350448 414044
rect 350448 414024 350500 414044
rect 350500 414024 350502 414044
rect 350446 411324 350502 411360
rect 350446 411304 350448 411324
rect 350448 411304 350500 411324
rect 350500 411304 350502 411324
rect 350446 407244 350502 407280
rect 350446 407224 350448 407244
rect 350448 407224 350500 407244
rect 350500 407224 350502 407244
rect 350446 404504 350502 404560
rect 350446 400288 350502 400344
rect 350446 399472 350502 399528
rect 350446 397568 350502 397624
rect 350446 396752 350502 396808
rect 350446 394612 350448 394632
rect 350448 394612 350500 394632
rect 350500 394612 350502 394632
rect 350446 394576 350502 394612
rect 350446 392012 350502 392048
rect 350446 391992 350448 392012
rect 350448 391992 350500 392012
rect 350500 391992 350502 392012
rect 350354 389952 350410 390008
rect 350446 389816 350502 389872
rect 350446 387812 350448 387832
rect 350448 387812 350500 387832
rect 350500 387812 350502 387832
rect 350446 387776 350502 387812
rect 350354 387096 350410 387152
rect 350446 382336 350502 382392
rect 350354 381384 350410 381440
rect 350446 380976 350502 381032
rect 350446 377168 350502 377224
rect 350354 375808 350410 375864
rect 350446 374856 350502 374912
rect 350446 372816 350502 372872
rect 350446 371320 350502 371376
rect 350446 365336 350502 365392
rect 350446 364404 350502 364440
rect 350446 364384 350448 364404
rect 350448 364384 350500 364404
rect 350500 364384 350502 364404
rect 350446 358012 350502 358048
rect 350446 357992 350448 358012
rect 350448 357992 350500 358012
rect 350500 357992 350502 358012
rect 350446 355816 350502 355872
rect 350446 354748 350502 354784
rect 350446 354728 350448 354748
rect 350448 354728 350500 354748
rect 350500 354728 350502 354748
rect 350446 350648 350502 350704
rect 350354 349832 350410 349888
rect 350446 349288 350502 349344
rect 350354 345752 350410 345808
rect 350354 344392 350410 344448
rect 350354 342216 350410 342272
rect 350354 338156 350410 338192
rect 350354 338136 350356 338156
rect 350356 338136 350408 338156
rect 350408 338136 350410 338156
rect 350354 334056 350410 334112
rect 350354 332696 350410 332752
rect 350354 329860 350410 329896
rect 350354 329840 350356 329860
rect 350356 329840 350408 329860
rect 350408 329840 350410 329860
rect 350354 328888 350410 328944
rect 350354 325760 350410 325816
rect 350354 321680 350410 321736
rect 350354 320592 350410 320648
rect 350354 319232 350410 319288
rect 350354 317736 350410 317792
rect 350354 315016 350410 315072
rect 350354 312296 350410 312352
rect 350354 311072 350410 311128
rect 350354 308352 350410 308408
rect 350354 304272 350410 304328
rect 350354 302368 350410 302424
rect 350354 300892 350410 300928
rect 350354 300872 350356 300892
rect 350356 300872 350408 300892
rect 350408 300872 350410 300892
rect 350354 300192 350410 300248
rect 350354 298832 350410 298888
rect 350262 295332 350264 295352
rect 350264 295332 350316 295352
rect 350316 295332 350318 295352
rect 350262 295296 350318 295332
rect 350262 293972 350264 293992
rect 350264 293972 350316 293992
rect 350316 293972 350318 293992
rect 350262 293936 350318 293972
rect 350262 288632 350318 288688
rect 350262 287156 350318 287192
rect 350262 287136 350264 287156
rect 350264 287136 350316 287156
rect 350316 287136 350318 287156
rect 350262 286456 350318 286512
rect 350262 285096 350318 285152
rect 350262 277480 350318 277536
rect 350262 275576 350318 275632
rect 350170 273808 350226 273864
rect 350262 273420 350318 273456
rect 350262 273400 350264 273420
rect 350264 273400 350316 273420
rect 350316 273400 350318 273420
rect 350262 272176 350318 272232
rect 350262 270136 350318 270192
rect 350262 268776 350318 268832
rect 350262 266736 350318 266792
rect 350262 263880 350318 263936
rect 350262 261296 350318 261352
rect 349986 255992 350042 256048
rect 350078 247696 350134 247752
rect 350078 244296 350134 244352
rect 350170 242936 350226 242992
rect 350722 330656 350778 330712
rect 350906 385056 350962 385112
rect 351090 383696 351146 383752
rect 351090 379752 351146 379808
rect 350998 370096 351054 370152
rect 350998 363296 351054 363352
rect 350814 324536 350870 324592
rect 350630 284280 350686 284336
rect 350446 255332 350502 255368
rect 350446 255312 350448 255332
rect 350448 255312 350500 255332
rect 350500 255312 350502 255332
rect 350446 253972 350502 254008
rect 350446 253952 350448 253972
rect 350448 253952 350500 253972
rect 350500 253952 350502 253972
rect 350446 249872 350502 249928
rect 350446 248512 350502 248568
rect 350354 246064 350410 246120
rect 350446 245792 350502 245848
rect 350446 245692 350448 245712
rect 350448 245692 350500 245712
rect 350500 245692 350502 245712
rect 350446 245656 350502 245692
rect 350538 244432 350594 244488
rect 350446 243208 350502 243264
rect 350354 239264 350410 239320
rect 350446 238876 350502 238912
rect 350446 238856 350448 238876
rect 350448 238856 350500 238876
rect 350500 238856 350502 238876
rect 350446 236136 350502 236192
rect 350446 234932 350502 234968
rect 350446 234912 350448 234932
rect 350448 234912 350500 234932
rect 350500 234912 350502 234932
rect 350446 232192 350502 232248
rect 350446 230560 350502 230616
rect 350446 229200 350502 229256
rect 350446 225004 350502 225040
rect 350446 224984 350448 225004
rect 350448 224984 350500 225004
rect 350500 224984 350502 225004
rect 350446 222536 350502 222592
rect 350446 221196 350502 221232
rect 350446 221176 350448 221196
rect 350448 221176 350500 221196
rect 350500 221176 350502 221196
rect 350354 219952 350410 220008
rect 350262 217096 350318 217152
rect 350262 207712 350318 207768
rect 350262 204992 350318 205048
rect 350446 218068 350502 218104
rect 350446 218048 350448 218068
rect 350448 218048 350500 218068
rect 350500 218048 350502 218068
rect 350446 217504 350502 217560
rect 350446 215348 350502 215384
rect 350446 215328 350448 215348
rect 350448 215328 350500 215348
rect 350500 215328 350502 215348
rect 350446 213152 350502 213208
rect 350446 209072 350502 209128
rect 350446 207168 350502 207224
rect 350446 206932 350448 206952
rect 350448 206932 350500 206952
rect 350500 206932 350502 206952
rect 350446 206896 350502 206932
rect 350446 204212 350448 204232
rect 350448 204212 350500 204232
rect 350500 204212 350502 204232
rect 350446 204176 350502 204212
rect 350446 203088 350502 203144
rect 350446 201728 350502 201784
rect 352654 304952 352710 305008
rect 353298 201048 353354 201104
rect 355414 456728 355470 456784
rect 355506 285796 355562 285832
rect 355506 285776 355508 285796
rect 355508 285776 355560 285796
rect 355560 285776 355562 285796
rect 359554 159432 359610 159488
rect 362406 199688 362462 199744
rect 362958 177792 363014 177848
rect 363234 187584 363290 187640
rect 363694 680856 363750 680912
rect 369858 680448 369914 680504
rect 363694 199008 363750 199064
rect 365902 190168 365958 190224
rect 365718 155624 365774 155680
rect 366546 240080 366602 240136
rect 366638 232464 366694 232520
rect 367098 187448 367154 187504
rect 368478 194112 368534 194168
rect 368938 563624 368994 563680
rect 368662 187312 368718 187368
rect 368938 341400 368994 341456
rect 370962 191256 371018 191312
rect 371974 562400 372030 562456
rect 371238 173304 371294 173360
rect 372158 561992 372214 562048
rect 372158 210296 372214 210352
rect 372618 174936 372674 174992
rect 373354 564576 373410 564632
rect 373354 158480 373410 158536
rect 373538 185680 373594 185736
rect 373906 302232 373962 302288
rect 373722 190032 373778 190088
rect 374918 187176 374974 187232
rect 374734 163376 374790 163432
rect 373998 158344 374054 158400
rect 376022 174800 376078 174856
rect 375286 155352 375342 155408
rect 376206 561040 376262 561096
rect 376206 251776 376262 251832
rect 376390 178608 376446 178664
rect 377218 236544 377274 236600
rect 376114 152360 376170 152416
rect 377402 152768 377458 152824
rect 380438 235320 380494 235376
rect 384302 684800 384358 684856
rect 381726 154128 381782 154184
rect 382922 199280 382978 199336
rect 383566 231376 383622 231432
rect 383934 166232 383990 166288
rect 384210 155488 384266 155544
rect 384578 562536 384634 562592
rect 384578 166504 384634 166560
rect 384578 156984 384634 157040
rect 384670 155624 384726 155680
rect 387154 564712 387210 564768
rect 387062 562264 387118 562320
rect 385958 237224 386014 237280
rect 386326 149912 386382 149968
rect 387154 161064 387210 161120
rect 389086 311888 389142 311944
rect 388994 233824 389050 233880
rect 390006 563216 390062 563272
rect 394238 680312 394294 680368
rect 393042 239400 393098 239456
rect 394054 564440 394110 564496
rect 393962 166368 394018 166424
rect 393226 159432 393282 159488
rect 396446 239944 396502 240000
rect 396538 198600 396594 198656
rect 395986 166232 396042 166288
rect 397366 243480 397422 243536
rect 398194 559952 398250 560008
rect 398286 238448 398342 238504
rect 398102 152632 398158 152688
rect 399574 238584 399630 238640
rect 400678 231648 400734 231704
rect 399942 150048 399998 150104
rect 401138 159568 401194 159624
rect 402150 558184 402206 558240
rect 402426 161200 402482 161256
rect 404266 166368 404322 166424
rect 404818 588784 404874 588840
rect 405370 679632 405426 679688
rect 406382 642096 406438 642152
rect 406566 531800 406622 531856
rect 406474 459720 406530 459776
rect 406474 429800 406530 429856
rect 406750 667800 406806 667856
rect 406750 556280 406806 556336
rect 406658 372000 406714 372056
rect 406658 356360 406714 356416
rect 406566 262928 406622 262984
rect 407118 678000 407174 678056
rect 407118 670520 407174 670576
rect 407118 669160 407174 669216
rect 407210 667120 407266 667176
rect 407118 666440 407174 666496
rect 407026 644000 407082 644056
rect 406934 631760 406990 631816
rect 406842 467880 406898 467936
rect 407026 625368 407082 625424
rect 407210 663740 407266 663776
rect 407210 663720 407212 663740
rect 407212 663720 407264 663740
rect 407264 663720 407266 663740
rect 407394 662360 407450 662416
rect 407210 661680 407266 661736
rect 407302 661000 407358 661056
rect 407302 658960 407358 659016
rect 407210 654880 407266 654936
rect 407210 654220 407266 654256
rect 407210 654200 407212 654220
rect 407212 654200 407264 654220
rect 407264 654200 407266 654220
rect 407210 652840 407266 652896
rect 407210 650120 407266 650176
rect 407210 649440 407266 649496
rect 407486 648760 407542 648816
rect 407210 644680 407266 644736
rect 407210 641960 407266 642016
rect 407210 641280 407266 641336
rect 407302 638016 407358 638072
rect 407210 637880 407266 637936
rect 407210 637200 407266 637256
rect 407210 633800 407266 633856
rect 407210 632440 407266 632496
rect 407210 629040 407266 629096
rect 407302 619520 407358 619576
rect 407210 618840 407266 618896
rect 407302 616800 407358 616856
rect 407302 614896 407358 614952
rect 407210 612756 407212 612776
rect 407212 612756 407264 612776
rect 407264 612756 407266 612776
rect 407210 612720 407266 612756
rect 407210 608660 407266 608696
rect 407210 608640 407212 608660
rect 407212 608640 407264 608660
rect 407264 608640 407266 608660
rect 407302 602520 407358 602576
rect 407302 601840 407358 601896
rect 407302 599120 407358 599176
rect 407302 597080 407358 597136
rect 407302 595040 407358 595096
rect 407302 593000 407358 593056
rect 407394 591096 407450 591152
rect 407302 590960 407358 591016
rect 407302 588920 407358 588976
rect 407670 614760 407726 614816
rect 407486 588648 407542 588704
rect 407302 586880 407358 586936
rect 407946 605920 408002 605976
rect 407670 585520 407726 585576
rect 407302 584840 407358 584896
rect 407302 580080 407358 580136
rect 407302 577360 407358 577416
rect 407302 576680 407358 576736
rect 407302 573996 407304 574016
rect 407304 573996 407356 574016
rect 407356 573996 407358 574016
rect 407302 573960 407358 573996
rect 407302 573280 407358 573336
rect 407302 572600 407358 572656
rect 407946 570560 408002 570616
rect 407302 569880 407358 569936
rect 407302 567840 407358 567896
rect 408038 565120 408094 565176
rect 407394 564460 407450 564496
rect 407394 564440 407396 564460
rect 407396 564440 407448 564460
rect 407448 564440 407450 564460
rect 407854 561312 407910 561368
rect 407302 561040 407358 561096
rect 407578 555600 407634 555656
rect 407302 552880 407358 552936
rect 407394 551520 407450 551576
rect 407302 550840 407358 550896
rect 407302 550160 407358 550216
rect 407302 547440 407358 547496
rect 408038 559000 408094 559056
rect 407946 556960 408002 557016
rect 407854 548800 407910 548856
rect 407762 546080 407818 546136
rect 407302 544720 407358 544776
rect 407394 544040 407450 544096
rect 407302 542000 407358 542056
rect 407762 537920 407818 537976
rect 407302 535200 407358 535256
rect 407302 529080 407358 529136
rect 407394 525680 407450 525736
rect 407302 525036 407304 525056
rect 407304 525036 407356 525056
rect 407356 525036 407358 525056
rect 407302 525000 407358 525036
rect 407302 523640 407358 523696
rect 407394 522960 407450 523016
rect 407302 522280 407358 522336
rect 407302 521600 407358 521656
rect 407394 518200 407450 518256
rect 407302 517556 407304 517576
rect 407304 517556 407356 517576
rect 407356 517556 407358 517576
rect 407302 517520 407358 517556
rect 407394 516840 407450 516896
rect 407302 516196 407304 516216
rect 407304 516196 407356 516216
rect 407356 516196 407358 516216
rect 407302 516160 407358 516196
rect 407670 514800 407726 514856
rect 407302 512760 407358 512816
rect 407302 512080 407358 512136
rect 407302 509360 407358 509416
rect 407302 508000 407358 508056
rect 407302 506640 407358 506696
rect 407302 501200 407358 501256
rect 407394 500520 407450 500576
rect 407302 495760 407358 495816
rect 407302 493040 407358 493096
rect 407302 491000 407358 491056
rect 407302 489640 407358 489696
rect 407302 487600 407358 487656
rect 407302 486920 407358 486976
rect 407486 485560 407542 485616
rect 407302 484880 407358 484936
rect 407302 484200 407358 484256
rect 407302 482160 407358 482216
rect 407302 478080 407358 478136
rect 407302 475360 407358 475416
rect 407394 474680 407450 474736
rect 407302 474000 407358 474056
rect 407302 471996 407304 472016
rect 407304 471996 407356 472016
rect 407356 471996 407358 472016
rect 407302 471960 407358 471996
rect 407302 469920 407358 469976
rect 407302 468152 407358 468208
rect 407302 465840 407358 465896
rect 407302 463800 407358 463856
rect 407394 463120 407450 463176
rect 407302 462440 407358 462496
rect 407302 459040 407358 459096
rect 407302 457000 407358 457056
rect 407394 455640 407450 455696
rect 407302 454960 407358 455016
rect 407394 454280 407450 454336
rect 407670 452920 407726 452976
rect 407302 451560 407358 451616
rect 407302 449520 407358 449576
rect 407302 447208 407358 447264
rect 407394 446120 407450 446176
rect 407302 444760 407358 444816
rect 407302 442040 407358 442096
rect 407394 441360 407450 441416
rect 407210 440000 407266 440056
rect 407210 437960 407266 438016
rect 407210 437280 407266 437336
rect 407210 435920 407266 435976
rect 407486 438640 407542 438696
rect 407302 434560 407358 434616
rect 407210 433200 407266 433256
rect 407210 429120 407266 429176
rect 407302 427760 407358 427816
rect 407210 427080 407266 427136
rect 407210 425720 407266 425776
rect 407210 423700 407266 423736
rect 407210 423680 407212 423700
rect 407212 423680 407264 423700
rect 407264 423680 407266 423700
rect 407210 423000 407266 423056
rect 407302 420280 407358 420336
rect 407210 419600 407266 419656
rect 407210 418920 407266 418976
rect 407578 416200 407634 416256
rect 407210 414840 407266 414896
rect 407302 412120 407358 412176
rect 407210 411440 407266 411496
rect 407210 410760 407266 410816
rect 407210 407360 407266 407416
rect 407210 406000 407266 406056
rect 407302 404640 407358 404696
rect 407210 401920 407266 401976
rect 407210 397840 407266 397896
rect 407210 395800 407266 395856
rect 407210 393760 407266 393816
rect 407302 391720 407358 391776
rect 407210 391040 407266 391096
rect 407210 385600 407266 385656
rect 407210 384920 407266 384976
rect 407210 381520 407266 381576
rect 407210 378800 407266 378856
rect 407210 374060 407266 374096
rect 407210 374040 407212 374060
rect 407212 374040 407264 374060
rect 407264 374040 407266 374060
rect 407210 373360 407266 373416
rect 407210 370640 407266 370696
rect 407210 369280 407266 369336
rect 407210 361120 407266 361176
rect 407210 360440 407266 360496
rect 407210 357720 407266 357776
rect 407210 357040 407266 357096
rect 407210 353640 407266 353696
rect 407302 352960 407358 353016
rect 407210 352280 407266 352336
rect 407210 351600 407266 351656
rect 407210 349288 407266 349344
rect 407210 345480 407266 345536
rect 407210 344800 407266 344856
rect 407210 343440 407266 343496
rect 407210 340720 407266 340776
rect 407210 336676 407212 336696
rect 407212 336676 407264 336696
rect 407264 336676 407266 336696
rect 407210 336640 407266 336676
rect 407302 332560 407358 332616
rect 407210 331236 407212 331256
rect 407212 331236 407264 331256
rect 407264 331236 407266 331256
rect 407210 331200 407266 331236
rect 407210 330520 407266 330576
rect 407210 328500 407266 328536
rect 407210 328480 407212 328500
rect 407212 328480 407264 328500
rect 407264 328480 407266 328500
rect 407210 325080 407266 325136
rect 407210 323720 407266 323776
rect 407118 323040 407174 323096
rect 407118 322360 407174 322416
rect 407210 321680 407266 321736
rect 407118 321000 407174 321056
rect 407118 318280 407174 318336
rect 407118 312840 407174 312896
rect 407210 311072 407266 311128
rect 407118 310800 407174 310856
rect 407118 310120 407174 310176
rect 407118 308080 407174 308136
rect 407210 306720 407266 306776
rect 407118 305360 407174 305416
rect 407118 304000 407174 304056
rect 407210 301960 407266 302016
rect 407118 301280 407174 301336
rect 407118 299920 407174 299976
rect 407118 295840 407174 295896
rect 407210 293800 407266 293856
rect 407118 293120 407174 293176
rect 407118 292476 407120 292496
rect 407120 292476 407172 292496
rect 407172 292476 407174 292496
rect 407118 292440 407174 292476
rect 407210 291760 407266 291816
rect 407118 289040 407174 289096
rect 407118 288360 407174 288416
rect 407210 287680 407266 287736
rect 407118 287000 407174 287056
rect 407210 284960 407266 285016
rect 407118 284316 407120 284336
rect 407120 284316 407172 284336
rect 407172 284316 407174 284336
rect 407118 284280 407174 284316
rect 407210 283600 407266 283656
rect 407118 282940 407174 282976
rect 407118 282920 407120 282940
rect 407120 282920 407172 282940
rect 407172 282920 407174 282940
rect 407118 278840 407174 278896
rect 407118 276120 407174 276176
rect 407118 275440 407174 275496
rect 407118 272720 407174 272776
rect 407210 271360 407266 271416
rect 407118 270000 407174 270056
rect 407118 267960 407174 268016
rect 407118 263880 407174 263936
rect 407118 262520 407174 262576
rect 407118 261840 407174 261896
rect 407118 259800 407174 259856
rect 407210 257760 407266 257816
rect 407118 257080 407174 257136
rect 407118 255040 407174 255096
rect 407210 251640 407266 251696
rect 407210 250960 407266 251016
rect 407118 250280 407174 250336
rect 407210 246880 407266 246936
rect 407118 246200 407174 246256
rect 407210 245520 407266 245576
rect 407118 244840 407174 244896
rect 407118 242120 407174 242176
rect 407394 318960 407450 319016
rect 407394 302640 407450 302696
rect 407670 298560 407726 298616
rect 407486 262112 407542 262168
rect 407394 254360 407450 254416
rect 407854 483520 407910 483576
rect 407946 395120 408002 395176
rect 407946 383016 408002 383072
rect 407762 267280 407818 267336
rect 407762 242936 407818 242992
rect 407670 242528 407726 242584
rect 408314 679360 408370 679416
rect 408222 650120 408278 650176
rect 408406 665080 408462 665136
rect 408406 646720 408462 646776
rect 408222 476176 408278 476232
rect 408222 476040 408278 476096
rect 408130 461080 408186 461136
rect 408130 408720 408186 408776
rect 408130 382880 408186 382936
rect 408038 362480 408094 362536
rect 408038 346840 408094 346896
rect 408038 276800 408094 276856
rect 408406 594360 408462 594416
rect 408406 586200 408462 586256
rect 408958 578040 409014 578096
rect 409050 510040 409106 510096
rect 409142 479440 409198 479496
rect 409234 476720 409290 476776
rect 409234 467200 409290 467256
rect 408314 457680 408370 457736
rect 408406 433880 408462 433936
rect 408314 421640 408370 421696
rect 408866 400288 408922 400344
rect 408406 389680 408462 389736
rect 408406 327800 408462 327856
rect 408406 259936 408462 259992
rect 408406 239808 408462 239864
rect 409050 319640 409106 319696
rect 408958 249600 409014 249656
rect 409326 430480 409382 430536
rect 409418 428440 409474 428496
rect 409510 399200 409566 399256
rect 409326 393080 409382 393136
rect 409602 377440 409658 377496
rect 409694 364520 409750 364576
rect 409418 342760 409474 342816
rect 409326 300600 409382 300656
rect 409326 293936 409382 293992
rect 409234 279520 409290 279576
rect 409694 339360 409750 339416
rect 409602 289720 409658 289776
rect 409510 241188 409566 241224
rect 409510 241168 409512 241188
rect 409512 241168 409564 241188
rect 409564 241168 409566 241188
rect 409510 240760 409566 240816
rect 425794 684528 425850 684584
rect 424506 683440 424562 683496
rect 416594 682896 416650 682952
rect 415490 681944 415546 682000
rect 427818 680720 427874 680776
rect 433844 680040 433900 680096
rect 445114 683712 445170 683768
rect 442538 683168 442594 683224
rect 442262 682760 442318 682816
rect 440330 681128 440386 681184
rect 441894 682216 441950 682272
rect 441250 680720 441306 680776
rect 476578 686024 476634 686080
rect 447690 682624 447746 682680
rect 454774 684800 454830 684856
rect 458638 682488 458694 682544
rect 462502 682352 462558 682408
rect 467010 681128 467066 681184
rect 472162 680992 472218 681048
rect 481178 680992 481234 681048
rect 488722 680856 488778 680912
rect 499854 683576 499910 683632
rect 500498 680584 500554 680640
rect 507582 682624 507638 682680
rect 505098 681808 505154 681864
rect 518990 680448 519046 680504
rect 528742 682352 528798 682408
rect 524970 682080 525026 682136
rect 526258 682080 526314 682136
rect 534078 682760 534134 682816
rect 531226 682216 531282 682272
rect 535274 682488 535330 682544
rect 546958 682896 547014 682952
rect 546866 681944 546922 682000
rect 549442 681808 549498 681864
rect 550178 680312 550234 680368
rect 489734 679496 489790 679552
rect 550178 678680 550234 678736
rect 550086 378800 550142 378856
rect 409786 334600 409842 334656
rect 409786 334464 409842 334520
rect 409878 315560 409934 315616
rect 550638 622920 550694 622976
rect 550454 564440 550510 564496
rect 550454 539960 550510 540016
rect 550362 522280 550418 522336
rect 550270 507320 550326 507376
rect 550638 282240 550694 282296
rect 550270 266600 550326 266656
rect 550178 242800 550234 242856
rect 550086 240760 550142 240816
rect 409050 152632 409106 152688
rect 412270 234232 412326 234288
rect 410522 151272 410578 151328
rect 427082 188536 427138 188592
rect 440606 156848 440662 156904
rect 457350 238720 457406 238776
rect 458178 238312 458234 238368
rect 453486 192616 453542 192672
rect 458178 180104 458234 180160
rect 470598 238312 470654 238368
rect 463790 153040 463846 153096
rect 476210 194520 476266 194576
rect 482466 152904 482522 152960
rect 488906 168952 488962 169008
rect 492770 185544 492826 185600
rect 495438 195336 495494 195392
rect 497278 184184 497334 184240
rect 498566 152768 498622 152824
rect 502430 167728 502486 167784
rect 524326 238176 524382 238232
rect 520186 238040 520242 238096
rect 528834 238448 528890 238504
rect 528742 237904 528798 237960
rect 523038 206216 523094 206272
rect 531318 195880 531374 195936
rect 538862 239536 538918 239592
rect 536102 195200 536158 195256
rect 537574 151680 537630 151736
rect 538770 150320 538826 150376
rect 538862 150184 538918 150240
rect 539046 149932 539102 149968
rect 539046 149912 539048 149932
rect 539048 149912 539100 149932
rect 539100 149912 539102 149932
rect 539322 149912 539378 149968
rect 539874 150184 539930 150240
rect 60002 29824 60058 29880
rect 60738 29688 60794 29744
rect 61290 29552 61346 29608
rect 65798 28192 65854 28248
rect 64878 23296 64934 23352
rect 66442 27512 66498 27568
rect 69662 27376 69718 27432
rect 64326 4800 64382 4856
rect 72330 28192 72386 28248
rect 70398 25336 70454 25392
rect 78034 28872 78090 28928
rect 74538 24384 74594 24440
rect 85762 29416 85818 29472
rect 91558 28328 91614 28384
rect 92478 28328 92534 28384
rect 96066 28192 96122 28248
rect 88338 25472 88394 25528
rect 84198 16904 84254 16960
rect 97354 28192 97410 28248
rect 97354 21664 97410 21720
rect 100758 24520 100814 24576
rect 107658 21800 107714 21856
rect 74998 3440 75054 3496
rect 117962 28056 118018 28112
rect 124218 21256 124274 21312
rect 127622 28872 127678 28928
rect 125690 23024 125746 23080
rect 125690 21392 125746 21448
rect 103334 3304 103390 3360
rect 138018 23024 138074 23080
rect 135258 21256 135314 21312
rect 128358 18536 128414 18592
rect 126978 3304 127034 3360
rect 132958 10240 133014 10296
rect 139490 18808 139546 18864
rect 150438 21392 150494 21448
rect 143538 15952 143594 16008
rect 151818 19896 151874 19952
rect 150530 16496 150586 16552
rect 161478 21528 161534 21584
rect 157798 15816 157854 15872
rect 155406 7520 155462 7576
rect 164238 24112 164294 24168
rect 169482 28328 169538 28384
rect 165802 24520 165858 24576
rect 175278 28464 175334 28520
rect 174634 27376 174690 27432
rect 173898 20032 173954 20088
rect 169574 3440 169630 3496
rect 173162 3576 173218 3632
rect 179418 21664 179474 21720
rect 178038 17720 178094 17776
rect 186226 28192 186282 28248
rect 179050 6160 179106 6216
rect 204258 19896 204314 19952
rect 207018 25608 207074 25664
rect 207018 24248 207074 24304
rect 201498 10376 201554 10432
rect 203890 3576 203946 3632
rect 213918 28736 213974 28792
rect 212630 17584 212686 17640
rect 218058 17176 218114 17232
rect 214470 16088 214526 16144
rect 222198 18944 222254 19000
rect 220910 15136 220966 15192
rect 234526 28736 234582 28792
rect 244186 29280 244242 29336
rect 235998 21800 236054 21856
rect 284114 29144 284170 29200
rect 274638 24384 274694 24440
rect 236550 14456 236606 14512
rect 242990 3712 243046 3768
rect 267738 18808 267794 18864
rect 282918 18944 282974 19000
rect 278778 18672 278834 18728
rect 276018 7656 276074 7712
rect 291198 19080 291254 19136
rect 300950 23976 301006 24032
rect 314382 29144 314438 29200
rect 319534 28600 319590 28656
rect 304998 22480 305054 22536
rect 300858 19080 300914 19136
rect 324410 22616 324466 22672
rect 324410 12960 324466 13016
rect 332598 25608 332654 25664
rect 335358 17312 335414 17368
rect 328734 11736 328790 11792
rect 339498 25472 339554 25528
rect 336738 19216 336794 19272
rect 339590 13640 339646 13696
rect 347870 23976 347926 24032
rect 353298 17448 353354 17504
rect 359462 29280 359518 29336
rect 358910 26832 358966 26888
rect 364430 25744 364486 25800
rect 369122 26968 369178 27024
rect 373630 29008 373686 29064
rect 373998 25744 374054 25800
rect 377494 28600 377550 28656
rect 378230 27104 378286 27160
rect 382646 26696 382702 26752
rect 389730 27240 389786 27296
rect 391938 22616 391994 22672
rect 386418 15000 386474 15056
rect 402978 17040 403034 17096
rect 408498 25880 408554 25936
rect 409878 25880 409934 25936
rect 407118 21120 407174 21176
rect 415398 22752 415454 22808
rect 416686 22788 416688 22808
rect 416688 22788 416740 22808
rect 416740 22788 416742 22808
rect 416686 22752 416742 22788
rect 421930 27240 421986 27296
rect 426530 22888 426586 22944
rect 431958 16496 432014 16552
rect 440330 16360 440386 16416
rect 438858 14864 438914 14920
rect 445850 22888 445906 22944
rect 445758 21936 445814 21992
rect 448610 25336 448666 25392
rect 452842 28464 452898 28520
rect 448518 20168 448574 20224
rect 459650 24656 459706 24712
rect 463790 20168 463846 20224
rect 468942 23160 468998 23216
rect 473450 24792 473506 24848
rect 465170 21936 465226 21992
rect 474738 28192 474794 28248
rect 478878 26016 478934 26072
rect 479062 26016 479118 26072
rect 487618 28328 487674 28384
rect 485042 26152 485098 26208
rect 484582 25200 484638 25256
rect 484490 24792 484546 24848
rect 505098 20304 505154 20360
rect 484398 12280 484454 12336
rect 485226 6296 485282 6352
rect 509514 29008 509570 29064
rect 511446 26968 511502 27024
rect 510802 26696 510858 26752
rect 504362 10240 504418 10296
rect 506478 3848 506534 3904
rect 519818 29416 519874 29472
rect 524326 26560 524382 26616
rect 525614 27512 525670 27568
rect 525798 20440 525854 20496
rect 526442 20304 526498 20360
rect 537850 29552 537906 29608
rect 531318 3984 531374 4040
rect 540058 147736 540114 147792
rect 540150 147328 540206 147384
rect 540058 143384 540114 143440
rect 538310 20576 538366 20632
rect 540702 149640 540758 149696
rect 540978 145424 541034 145480
rect 541070 133456 541126 133512
rect 540886 133184 540942 133240
rect 540978 129648 541034 129704
rect 540610 115912 540666 115968
rect 540794 99456 540850 99512
rect 541162 101496 541218 101552
rect 541070 95104 541126 95160
rect 541530 141752 541586 141808
rect 541898 147600 541954 147656
rect 541622 136584 541678 136640
rect 541806 133048 541862 133104
rect 543094 236544 543150 236600
rect 542358 197240 542414 197296
rect 541806 127608 541862 127664
rect 541530 102176 541586 102232
rect 541530 82864 541586 82920
rect 541254 43696 541310 43752
rect 541806 115912 541862 115968
rect 541714 115776 541770 115832
rect 542542 145696 542598 145752
rect 542450 136176 542506 136232
rect 542450 134136 542506 134192
rect 542450 131416 542506 131472
rect 542450 130736 542506 130792
rect 542450 129376 542506 129432
rect 542450 125332 542452 125352
rect 542452 125332 542504 125352
rect 542504 125332 542506 125352
rect 542450 125296 542506 125332
rect 542450 116456 542506 116512
rect 542450 113736 542506 113792
rect 542542 110336 542598 110392
rect 542450 109656 542506 109712
rect 543554 231376 543610 231432
rect 542910 141652 542912 141672
rect 542912 141652 542964 141672
rect 542964 141652 542966 141672
rect 542910 141616 542966 141652
rect 542818 135496 542874 135552
rect 542634 107616 542690 107672
rect 542910 129512 542966 129568
rect 544106 233824 544162 233880
rect 543646 149640 543702 149696
rect 543462 146376 543518 146432
rect 543278 142296 543334 142352
rect 543554 140936 543610 140992
rect 543554 138216 543610 138272
rect 542634 91296 542690 91352
rect 542726 88576 542782 88632
rect 542634 84496 542690 84552
rect 542634 75692 542636 75712
rect 542636 75692 542688 75712
rect 542688 75692 542690 75712
rect 542634 75656 542690 75692
rect 542818 65456 542874 65512
rect 542726 52536 542782 52592
rect 542726 49816 542782 49872
rect 542726 48456 542782 48512
rect 542542 30640 542598 30696
rect 543186 106256 543242 106312
rect 543554 128016 543610 128072
rect 543554 124616 543610 124672
rect 543646 121896 543702 121952
rect 543554 120536 543610 120592
rect 543554 117952 543610 118008
rect 543554 110472 543610 110528
rect 543554 97416 543610 97472
rect 543554 96056 543610 96112
rect 543646 95376 543702 95432
rect 543554 94016 543610 94072
rect 543554 92656 543610 92712
rect 543554 91976 543610 92032
rect 543554 82456 543610 82512
rect 543554 77696 543610 77752
rect 543554 76336 543610 76392
rect 543554 74976 543610 75032
rect 543554 71576 543610 71632
rect 543554 70216 543610 70272
rect 543554 66156 543610 66192
rect 543554 66136 543556 66156
rect 543556 66136 543608 66156
rect 543608 66136 543610 66156
rect 543554 64096 543610 64152
rect 543554 62076 543610 62112
rect 543554 62056 543556 62076
rect 543556 62056 543608 62076
rect 543608 62056 543610 62076
rect 543646 60696 543702 60752
rect 543554 56616 543610 56672
rect 543646 47776 543702 47832
rect 543554 45056 543610 45112
rect 543646 44376 543702 44432
rect 543554 40976 543610 41032
rect 543554 36216 543610 36272
rect 543646 35536 543702 35592
rect 543646 31184 543702 31240
rect 543646 30368 543702 30424
rect 544106 144744 544162 144800
rect 543922 78376 543978 78432
rect 544474 146512 544530 146568
rect 544658 146240 544714 146296
rect 544658 139440 544714 139496
rect 544566 136584 544622 136640
rect 544566 131144 544622 131200
rect 544290 114416 544346 114472
rect 544566 124072 544622 124128
rect 544566 117272 544622 117328
rect 547234 239400 547290 239456
rect 545210 138080 545266 138136
rect 545210 128424 545266 128480
rect 545118 127064 545174 127120
rect 545118 123936 545174 123992
rect 541990 3168 542046 3224
rect 546130 155488 546186 155544
rect 546038 139440 546094 139496
rect 546038 126928 546094 126984
rect 546958 146784 547014 146840
rect 547418 138080 547474 138136
rect 547418 126928 547474 126984
rect 548154 238584 548210 238640
rect 548982 238176 549038 238232
rect 547878 130464 547934 130520
rect 547786 85584 547842 85640
rect 549442 238040 549498 238096
rect 549350 137944 549406 138000
rect 549718 113192 549774 113248
rect 550086 126248 550142 126304
rect 550362 262520 550418 262576
rect 551098 524320 551154 524376
rect 551190 520920 551246 520976
rect 551374 684664 551430 684720
rect 551006 468560 551062 468616
rect 550914 431840 550970 431896
rect 551006 422320 551062 422376
rect 550914 407360 550970 407416
rect 550822 363840 550878 363896
rect 550822 287680 550878 287736
rect 550730 271360 550786 271416
rect 550730 234096 550786 234152
rect 551006 371320 551062 371376
rect 551098 365200 551154 365256
rect 551006 333920 551062 333976
rect 551190 327800 551246 327856
rect 552018 679360 552074 679416
rect 552018 678000 552074 678056
rect 552018 675960 552074 676016
rect 552294 674600 552350 674656
rect 552018 672424 552074 672480
rect 552202 661680 552258 661736
rect 552110 653520 552166 653576
rect 551558 650120 551614 650176
rect 552110 645360 552166 645416
rect 552018 641960 552074 642016
rect 552110 638288 552166 638344
rect 552018 637880 552074 637936
rect 552018 631760 552074 631816
rect 552018 625388 552074 625424
rect 552018 625368 552020 625388
rect 552020 625368 552072 625388
rect 552072 625368 552074 625388
rect 552018 624280 552074 624336
rect 552202 607300 552258 607336
rect 552202 607280 552204 607300
rect 552204 607280 552256 607300
rect 552256 607280 552258 607300
rect 552018 603916 552020 603936
rect 552020 603916 552072 603936
rect 552072 603916 552074 603936
rect 552018 603880 552074 603916
rect 552846 679768 552902 679824
rect 552570 654200 552626 654256
rect 552570 646720 552626 646776
rect 552478 642640 552534 642696
rect 552386 634480 552442 634536
rect 552570 620200 552626 620256
rect 552478 608660 552534 608696
rect 552478 608640 552480 608660
rect 552480 608640 552532 608660
rect 552532 608640 552534 608660
rect 552294 600480 552350 600536
rect 552018 598440 552074 598496
rect 552294 597488 552350 597544
rect 552018 596400 552074 596456
rect 552110 588956 552112 588976
rect 552112 588956 552164 588976
rect 552164 588956 552166 588976
rect 552110 588920 552166 588956
rect 552110 573996 552112 574016
rect 552112 573996 552164 574016
rect 552164 573996 552166 574016
rect 552110 573960 552166 573996
rect 552018 562420 552074 562456
rect 552018 562400 552020 562420
rect 552020 562400 552072 562420
rect 552072 562400 552074 562420
rect 552018 556960 552074 557016
rect 552570 586200 552626 586256
rect 552570 569880 552626 569936
rect 552478 568520 552534 568576
rect 552294 555600 552350 555656
rect 552018 553560 552074 553616
rect 552386 552880 552442 552936
rect 552110 545400 552166 545456
rect 552018 536560 552074 536616
rect 552018 532516 552020 532536
rect 552020 532516 552072 532536
rect 552072 532516 552074 532536
rect 552018 532480 552074 532516
rect 552018 530440 552074 530496
rect 552018 526360 552074 526416
rect 552018 525716 552020 525736
rect 552020 525716 552072 525736
rect 552072 525716 552074 525736
rect 552018 525680 552074 525716
rect 552018 521600 552074 521656
rect 552018 519424 552074 519480
rect 552018 518916 552020 518936
rect 552020 518916 552072 518936
rect 552072 518916 552074 518936
rect 552018 518880 552074 518916
rect 552018 516840 552074 516896
rect 552018 514820 552074 514856
rect 552018 514800 552020 514820
rect 552020 514800 552072 514820
rect 552072 514800 552074 514820
rect 552018 480120 552074 480176
rect 552018 465840 552074 465896
rect 552018 464344 552074 464400
rect 552018 463120 552074 463176
rect 552018 459720 552074 459776
rect 552018 459060 552074 459096
rect 552018 459040 552020 459060
rect 552020 459040 552072 459060
rect 552072 459040 552074 459060
rect 552018 457680 552074 457736
rect 552018 456340 552074 456376
rect 552018 456320 552020 456340
rect 552020 456320 552072 456340
rect 552072 456320 552074 456340
rect 552018 416200 552074 416256
rect 552018 415520 552074 415576
rect 552018 412820 552074 412856
rect 552018 412800 552020 412820
rect 552020 412800 552072 412820
rect 552072 412800 552074 412820
rect 552018 393760 552074 393816
rect 552018 367920 552074 367976
rect 552018 350940 552074 350976
rect 552018 350920 552020 350940
rect 552020 350920 552072 350940
rect 552072 350920 552074 350940
rect 552018 342796 552020 342816
rect 552020 342796 552072 342816
rect 552072 342796 552074 342816
rect 552018 342760 552074 342796
rect 552018 322360 552074 322416
rect 552018 307436 552020 307456
rect 552020 307436 552072 307456
rect 552072 307436 552074 307456
rect 552018 307400 552074 307436
rect 552018 293140 552074 293176
rect 552018 293120 552020 293140
rect 552020 293120 552072 293140
rect 552072 293120 552074 293140
rect 552018 290400 552074 290456
rect 551558 238720 551614 238776
rect 552018 263200 552074 263256
rect 552018 243344 552074 243400
rect 552570 540640 552626 540696
rect 552570 539280 552626 539336
rect 552386 534520 552442 534576
rect 552478 533840 552534 533896
rect 552294 515480 552350 515536
rect 552202 496440 552258 496496
rect 552202 460400 552258 460456
rect 552202 451424 552258 451480
rect 552202 432520 552258 432576
rect 552386 500520 552442 500576
rect 552662 531120 552718 531176
rect 552570 493720 552626 493776
rect 552478 492360 552534 492416
rect 552570 484200 552626 484256
rect 552570 478760 552626 478816
rect 552478 454960 552534 455016
rect 552386 454280 552442 454336
rect 552570 453600 552626 453656
rect 552386 446800 552442 446856
rect 552294 421640 552350 421696
rect 552294 420996 552296 421016
rect 552296 420996 552348 421016
rect 552348 420996 552350 421016
rect 552294 420960 552350 420996
rect 552202 413344 552258 413400
rect 552294 390360 552350 390416
rect 552202 360460 552258 360496
rect 552202 360440 552204 360460
rect 552204 360440 552256 360460
rect 552256 360440 552258 360460
rect 552294 351600 552350 351656
rect 552294 306040 552350 306096
rect 552202 291780 552258 291816
rect 552202 291760 552204 291780
rect 552204 291760 552256 291780
rect 552256 291760 552258 291780
rect 552294 274780 552350 274816
rect 552294 274760 552296 274780
rect 552296 274760 552348 274780
rect 552348 274760 552350 274780
rect 552570 445440 552626 445496
rect 552662 437280 552718 437336
rect 552662 435920 552718 435976
rect 552662 358400 552718 358456
rect 552662 347520 552718 347576
rect 552478 331200 552534 331256
rect 552570 314880 552626 314936
rect 552662 301280 552718 301336
rect 552846 665760 552902 665816
rect 553030 670520 553086 670576
rect 552938 597760 552994 597816
rect 552938 584840 552994 584896
rect 552938 561040 552994 561096
rect 552938 558320 552994 558376
rect 552846 484880 552902 484936
rect 552938 476040 552994 476096
rect 553306 667800 553362 667856
rect 553306 656940 553362 656976
rect 553306 656920 553308 656940
rect 553308 656920 553360 656940
rect 553360 656920 553362 656940
rect 553306 648760 553362 648816
rect 553214 644700 553270 644736
rect 553214 644680 553216 644700
rect 553216 644680 553268 644700
rect 553268 644680 553270 644700
rect 553306 641280 553362 641336
rect 553306 617480 553362 617536
rect 553214 613400 553270 613456
rect 553306 612720 553362 612776
rect 553306 611380 553362 611416
rect 553306 611360 553308 611380
rect 553308 611360 553360 611380
rect 553360 611360 553362 611380
rect 553306 610680 553362 610736
rect 553306 605920 553362 605976
rect 553306 603200 553362 603256
rect 553306 599800 553362 599856
rect 553306 586880 553362 586936
rect 553214 585520 553270 585576
rect 553122 547440 553178 547496
rect 553122 505280 553178 505336
rect 553122 501880 553178 501936
rect 553122 493040 553178 493096
rect 553030 449520 553086 449576
rect 552846 428440 552902 428496
rect 553030 426436 553032 426456
rect 553032 426436 553084 426456
rect 553084 426436 553086 426456
rect 553030 426400 553086 426436
rect 553030 425076 553032 425096
rect 553032 425076 553084 425096
rect 553084 425076 553086 425096
rect 553030 425040 553086 425076
rect 552938 424360 552994 424416
rect 553030 423700 553086 423736
rect 553030 423680 553032 423700
rect 553032 423680 553084 423700
rect 553084 423680 553086 423700
rect 553030 420280 553086 420336
rect 552938 405320 552994 405376
rect 552846 403960 552902 404016
rect 552938 403280 552994 403336
rect 552938 395120 552994 395176
rect 552846 391720 552902 391776
rect 552938 391040 552994 391096
rect 552938 388320 552994 388376
rect 552938 387640 552994 387696
rect 552938 385600 552994 385656
rect 552938 381520 552994 381576
rect 552938 377440 552994 377496
rect 552938 372700 552994 372736
rect 552938 372680 552940 372700
rect 552940 372680 552992 372700
rect 552992 372680 552994 372700
rect 552938 370640 552994 370696
rect 552846 369280 552902 369336
rect 552938 368620 552994 368656
rect 552938 368600 552940 368620
rect 552940 368600 552992 368620
rect 552992 368600 552994 368620
rect 552846 366424 552902 366480
rect 552938 365880 552994 365936
rect 552938 361120 552994 361176
rect 552938 357720 552994 357776
rect 552938 355680 552994 355736
rect 552938 340040 552994 340096
rect 552938 335960 552994 336016
rect 552938 326440 552994 326496
rect 552938 323720 552994 323776
rect 552938 318280 552994 318336
rect 552938 314200 552994 314256
rect 552938 311344 552994 311400
rect 552938 289720 552994 289776
rect 552938 279520 552994 279576
rect 552938 264560 552994 264616
rect 552938 260344 552994 260400
rect 552938 255040 552994 255096
rect 552938 250280 552994 250336
rect 552754 235320 552810 235376
rect 552018 81504 552074 81560
rect 552202 163512 552258 163568
rect 552294 151408 552350 151464
rect 552662 146920 552718 146976
rect 552662 133048 552718 133104
rect 553122 354320 553178 354376
rect 553122 353640 553178 353696
rect 553122 349424 553178 349480
rect 553122 346840 553178 346896
rect 553122 343440 553178 343496
rect 553122 338680 553178 338736
rect 553122 335300 553178 335336
rect 553122 335280 553124 335300
rect 553124 335280 553176 335300
rect 553176 335280 553178 335300
rect 553122 334600 553178 334656
rect 553122 327140 553178 327176
rect 553122 327120 553124 327140
rect 553124 327120 553176 327140
rect 553176 327120 553178 327140
rect 553122 325780 553178 325816
rect 553122 325760 553124 325780
rect 553124 325760 553176 325780
rect 553176 325760 553178 325780
rect 553122 317600 553178 317656
rect 553122 316240 553178 316296
rect 553122 312840 553178 312896
rect 553122 310800 553178 310856
rect 553122 310120 553178 310176
rect 553122 308760 553178 308816
rect 553122 305360 553178 305416
rect 553122 301960 553178 302016
rect 553122 300600 553178 300656
rect 553122 297900 553178 297936
rect 553122 297880 553124 297900
rect 553124 297880 553176 297900
rect 553176 297880 553178 297900
rect 553122 297200 553178 297256
rect 553122 292440 553178 292496
rect 553122 289040 553178 289096
rect 553122 286320 553178 286376
rect 553122 283620 553178 283656
rect 553122 283600 553124 283620
rect 553124 283600 553176 283620
rect 553176 283600 553178 283620
rect 553122 281560 553178 281616
rect 553122 280900 553178 280936
rect 553122 280880 553124 280900
rect 553124 280880 553176 280900
rect 553176 280880 553178 280900
rect 553122 280220 553178 280256
rect 553122 280200 553124 280220
rect 553124 280200 553176 280220
rect 553176 280200 553178 280220
rect 553122 278840 553178 278896
rect 553122 277480 553178 277536
rect 553122 276120 553178 276176
rect 553122 273400 553178 273456
rect 553122 270680 553178 270736
rect 553122 268660 553178 268696
rect 553122 268640 553124 268660
rect 553124 268640 553176 268660
rect 553176 268640 553178 268660
rect 553122 265240 553178 265296
rect 553122 263880 553178 263936
rect 553122 261840 553178 261896
rect 553122 259800 553178 259856
rect 553122 259120 553178 259176
rect 553122 257760 553178 257816
rect 553122 254360 553178 254416
rect 553122 253680 553178 253736
rect 553122 252320 553178 252376
rect 553122 249600 553178 249656
rect 553122 248240 553178 248296
rect 553122 246200 553178 246256
rect 553122 244840 553178 244896
rect 553306 578040 553362 578096
rect 553306 576000 553362 576056
rect 553306 567840 553362 567896
rect 553306 560360 553362 560416
rect 553306 557640 553362 557696
rect 553306 550860 553362 550896
rect 553306 550840 553308 550860
rect 553308 550840 553360 550860
rect 553360 550840 553362 550860
rect 553306 549480 553362 549536
rect 553306 546760 553362 546816
rect 553306 544040 553362 544096
rect 553306 535900 553362 535936
rect 553306 535880 553308 535900
rect 553308 535880 553360 535900
rect 553360 535880 553362 535900
rect 553306 535200 553362 535256
rect 553306 528400 553362 528456
rect 553306 510040 553362 510096
rect 553306 505960 553362 506016
rect 553306 504600 553362 504656
rect 553306 502444 553362 502480
rect 553306 502424 553308 502444
rect 553308 502424 553360 502444
rect 553360 502424 553362 502444
rect 553306 501200 553362 501256
rect 553306 499860 553362 499896
rect 553306 499840 553308 499860
rect 553308 499840 553360 499860
rect 553360 499840 553362 499860
rect 553306 498480 553362 498536
rect 553306 495760 553362 495816
rect 553306 488960 553362 489016
rect 553306 488280 553362 488336
rect 553306 479440 553362 479496
rect 553306 475360 553362 475416
rect 553306 470620 553362 470656
rect 553306 470600 553308 470620
rect 553308 470600 553360 470620
rect 553360 470600 553362 470620
rect 553306 469920 553362 469976
rect 553306 466520 553362 466576
rect 553306 448840 553362 448896
rect 553306 443400 553362 443456
rect 553306 438640 553362 438696
rect 553306 437960 553362 438016
rect 553306 436600 553362 436656
rect 553214 174528 553270 174584
rect 553582 679632 553638 679688
rect 553490 429800 553546 429856
rect 553582 378120 553638 378176
rect 553582 340720 553638 340776
rect 553398 258440 553454 258496
rect 552846 138624 552902 138680
rect 553490 247560 553546 247616
rect 553490 88984 553546 89040
rect 555146 681128 555202 681184
rect 554226 151000 554282 151056
rect 554226 89120 554282 89176
rect 554962 239808 555018 239864
rect 554870 25880 554926 25936
rect 555054 196560 555110 196616
rect 555514 231512 555570 231568
rect 555422 188264 555478 188320
rect 556158 150184 556214 150240
rect 556434 238312 556490 238368
rect 556434 234640 556490 234696
rect 556802 110880 556858 110936
rect 557814 197920 557870 197976
rect 558458 148552 558514 148608
rect 558274 20304 558330 20360
rect 560298 231240 560354 231296
rect 559654 137264 559710 137320
rect 559654 86128 559710 86184
rect 560482 197104 560538 197160
rect 560758 198736 560814 198792
rect 560666 196968 560722 197024
rect 560758 31048 560814 31104
rect 560298 17584 560354 17640
rect 561954 149232 562010 149288
rect 562414 199824 562470 199880
rect 564622 99456 564678 99512
rect 565174 231104 565230 231160
rect 564990 193840 565046 193896
rect 565174 149096 565230 149152
rect 565910 239536 565966 239592
rect 565818 136584 565874 136640
rect 566186 152632 566242 152688
rect 579066 697176 579122 697232
rect 566738 28328 566794 28384
rect 567658 237904 567714 237960
rect 567658 235184 567714 235240
rect 568578 240080 568634 240136
rect 568946 150320 569002 150376
rect 569498 157120 569554 157176
rect 570050 684528 570106 684584
rect 570510 173168 570566 173224
rect 570786 158072 570842 158128
rect 574098 105440 574154 105496
rect 574926 157936 574982 157992
rect 575478 29164 575534 29200
rect 575478 29144 575480 29164
rect 575480 29144 575532 29164
rect 575532 29144 575534 29164
rect 575662 156984 575718 157040
rect 575570 25472 575626 25528
rect 576306 240488 576362 240544
rect 577042 28600 577098 28656
rect 576950 26016 577006 26072
rect 577318 25744 577374 25800
rect 577686 237224 577742 237280
rect 578882 19760 578938 19816
rect 579986 644000 580042 644056
rect 580170 630808 580226 630864
rect 579802 524456 579858 524512
rect 580170 471416 580226 471472
rect 580170 431568 580226 431624
rect 580170 378392 580226 378448
rect 579894 28872 579950 28928
rect 579710 20032 579766 20088
rect 580170 325216 580226 325272
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 232328 580226 232384
rect 580906 670656 580962 670712
rect 580814 617480 580870 617536
rect 580722 590960 580778 591016
rect 580630 577632 580686 577688
rect 580538 564304 580594 564360
rect 580446 537784 580502 537840
rect 580354 484608 580410 484664
rect 580354 418240 580410 418296
rect 580446 365064 580502 365120
rect 580262 219000 580318 219056
rect 580538 312024 580594 312080
rect 580446 192480 580502 192536
rect 580722 179152 580778 179208
rect 580170 152632 580226 152688
rect 580170 152360 580226 152416
rect 580538 139340 580540 139360
rect 580540 139340 580592 139360
rect 580592 139340 580594 139360
rect 580538 139304 580594 139340
rect 580538 112784 580594 112840
rect 580446 99456 580502 99512
rect 580354 72936 580410 72992
rect 580354 59608 580410 59664
rect 580262 33108 580318 33144
rect 580262 33088 580264 33108
rect 580264 33088 580316 33108
rect 580316 33088 580318 33108
rect 581274 23296 581330 23352
rect 580998 16088 581054 16144
rect 580170 12280 580226 12336
rect 581826 200912 581882 200968
rect 583298 239944 583354 240000
rect 582470 15816 582526 15872
<< metal3 >>
rect 89161 700362 89227 700365
rect 551502 700362 551508 700364
rect 89161 700360 551508 700362
rect 89161 700304 89166 700360
rect 89222 700304 551508 700360
rect 89161 700302 551508 700304
rect 89161 700299 89227 700302
rect 551502 700300 551508 700302
rect 551572 700300 551578 700364
rect -960 697220 480 697460
rect 579061 697234 579127 697237
rect 583520 697234 584960 697324
rect 579061 697232 584960 697234
rect 579061 697176 579066 697232
rect 579122 697176 584960 697232
rect 579061 697174 584960 697176
rect 579061 697171 579127 697174
rect 583520 697084 584960 697174
rect 356646 686020 356652 686084
rect 356716 686082 356722 686084
rect 476573 686082 476639 686085
rect 356716 686080 476639 686082
rect 356716 686024 476578 686080
rect 476634 686024 476639 686080
rect 356716 686022 476639 686024
rect 356716 686020 356722 686022
rect 476573 686019 476639 686022
rect 28206 685884 28212 685948
rect 28276 685946 28282 685948
rect 552238 685946 552244 685948
rect 28276 685886 552244 685946
rect 28276 685884 28282 685886
rect 552238 685884 552244 685886
rect 552308 685884 552314 685948
rect 384297 684858 384363 684861
rect 454769 684858 454835 684861
rect 384297 684856 454835 684858
rect 384297 684800 384302 684856
rect 384358 684800 454774 684856
rect 454830 684800 454835 684856
rect 384297 684798 454835 684800
rect 384297 684795 384363 684798
rect 454769 684795 454835 684798
rect 407614 684660 407620 684724
rect 407684 684722 407690 684724
rect 551369 684722 551435 684725
rect 407684 684720 551435 684722
rect 407684 684664 551374 684720
rect 551430 684664 551435 684720
rect 407684 684662 551435 684664
rect 407684 684660 407690 684662
rect 551369 684659 551435 684662
rect 425789 684586 425855 684589
rect 570045 684586 570111 684589
rect 425789 684584 570111 684586
rect 425789 684528 425794 684584
rect 425850 684528 570050 684584
rect 570106 684528 570111 684584
rect 425789 684526 570111 684528
rect 425789 684523 425855 684526
rect 570045 684523 570111 684526
rect -960 684164 480 684404
rect 583520 683906 584960 683996
rect 583342 683846 584960 683906
rect 392526 683708 392532 683772
rect 392596 683770 392602 683772
rect 445109 683770 445175 683773
rect 392596 683768 445175 683770
rect 392596 683712 445114 683768
rect 445170 683712 445175 683768
rect 392596 683710 445175 683712
rect 583342 683770 583402 683846
rect 583520 683770 584960 683846
rect 583342 683756 584960 683770
rect 583342 683710 583586 683756
rect 392596 683708 392602 683710
rect 445109 683707 445175 683710
rect 393078 683572 393084 683636
rect 393148 683634 393154 683636
rect 499849 683634 499915 683637
rect 393148 683632 499915 683634
rect 393148 683576 499854 683632
rect 499910 683576 499915 683632
rect 393148 683574 499915 683576
rect 393148 683572 393154 683574
rect 499849 683571 499915 683574
rect 424501 683498 424567 683501
rect 568614 683498 568620 683500
rect 424501 683496 568620 683498
rect 424501 683440 424506 683496
rect 424562 683440 568620 683496
rect 424501 683438 568620 683440
rect 424501 683435 424567 683438
rect 568614 683436 568620 683438
rect 568684 683436 568690 683500
rect 409822 683300 409828 683364
rect 409892 683362 409898 683364
rect 583526 683362 583586 683710
rect 409892 683302 583586 683362
rect 409892 683300 409898 683302
rect 25446 683164 25452 683228
rect 25516 683226 25522 683228
rect 442533 683226 442599 683229
rect 25516 683224 442599 683226
rect 25516 683168 442538 683224
rect 442594 683168 442599 683224
rect 25516 683166 442599 683168
rect 25516 683164 25522 683166
rect 442533 683163 442599 683166
rect 416589 682954 416655 682957
rect 546953 682954 547019 682957
rect 416589 682952 547019 682954
rect 416589 682896 416594 682952
rect 416650 682896 546958 682952
rect 547014 682896 547019 682952
rect 416589 682894 547019 682896
rect 416589 682891 416655 682894
rect 546953 682891 547019 682894
rect 442257 682818 442323 682821
rect 534073 682818 534139 682821
rect 442257 682816 534139 682818
rect 442257 682760 442262 682816
rect 442318 682760 534078 682816
rect 534134 682760 534139 682816
rect 442257 682758 534139 682760
rect 442257 682755 442323 682758
rect 534073 682755 534139 682758
rect 403750 682620 403756 682684
rect 403820 682682 403826 682684
rect 447685 682682 447751 682685
rect 403820 682680 447751 682682
rect 403820 682624 447690 682680
rect 447746 682624 447751 682680
rect 403820 682622 447751 682624
rect 403820 682620 403826 682622
rect 447685 682619 447751 682622
rect 507577 682682 507643 682685
rect 552054 682682 552060 682684
rect 507577 682680 552060 682682
rect 507577 682624 507582 682680
rect 507638 682624 552060 682680
rect 507577 682622 552060 682624
rect 507577 682619 507643 682622
rect 552054 682620 552060 682622
rect 552124 682620 552130 682684
rect 403566 682484 403572 682548
rect 403636 682546 403642 682548
rect 458633 682546 458699 682549
rect 403636 682544 458699 682546
rect 403636 682488 458638 682544
rect 458694 682488 458699 682544
rect 403636 682486 458699 682488
rect 403636 682484 403642 682486
rect 458633 682483 458699 682486
rect 535269 682546 535335 682549
rect 560518 682546 560524 682548
rect 535269 682544 560524 682546
rect 535269 682488 535274 682544
rect 535330 682488 560524 682544
rect 535269 682486 560524 682488
rect 535269 682483 535335 682486
rect 560518 682484 560524 682486
rect 560588 682484 560594 682548
rect 395286 682348 395292 682412
rect 395356 682410 395362 682412
rect 462497 682410 462563 682413
rect 395356 682408 462563 682410
rect 395356 682352 462502 682408
rect 462558 682352 462563 682408
rect 395356 682350 462563 682352
rect 395356 682348 395362 682350
rect 462497 682347 462563 682350
rect 528737 682410 528803 682413
rect 561622 682410 561628 682412
rect 528737 682408 561628 682410
rect 528737 682352 528742 682408
rect 528798 682352 561628 682408
rect 528737 682350 561628 682352
rect 528737 682347 528803 682350
rect 561622 682348 561628 682350
rect 561692 682348 561698 682412
rect 358118 682212 358124 682276
rect 358188 682274 358194 682276
rect 441889 682274 441955 682277
rect 358188 682272 441955 682274
rect 358188 682216 441894 682272
rect 441950 682216 441955 682272
rect 358188 682214 441955 682216
rect 358188 682212 358194 682214
rect 441889 682211 441955 682214
rect 531221 682274 531287 682277
rect 565118 682274 565124 682276
rect 531221 682272 565124 682274
rect 531221 682216 531226 682272
rect 531282 682216 565124 682272
rect 531221 682214 565124 682216
rect 531221 682211 531287 682214
rect 565118 682212 565124 682214
rect 565188 682212 565194 682276
rect 399334 682076 399340 682140
rect 399404 682138 399410 682140
rect 524965 682138 525031 682141
rect 399404 682136 525031 682138
rect 399404 682080 524970 682136
rect 525026 682080 525031 682136
rect 399404 682078 525031 682080
rect 399404 682076 399410 682078
rect 524965 682075 525031 682078
rect 526253 682138 526319 682141
rect 566958 682138 566964 682140
rect 526253 682136 566964 682138
rect 526253 682080 526258 682136
rect 526314 682080 566964 682136
rect 526253 682078 566964 682080
rect 526253 682075 526319 682078
rect 566958 682076 566964 682078
rect 567028 682076 567034 682140
rect 397310 681940 397316 682004
rect 397380 682002 397386 682004
rect 415485 682002 415551 682005
rect 397380 682000 415551 682002
rect 397380 681944 415490 682000
rect 415546 681944 415551 682000
rect 397380 681942 415551 681944
rect 397380 681940 397386 681942
rect 415485 681939 415551 681942
rect 546861 682002 546927 682005
rect 574134 682002 574140 682004
rect 546861 682000 574140 682002
rect 546861 681944 546866 682000
rect 546922 681944 574140 682000
rect 546861 681942 574140 681944
rect 546861 681939 546927 681942
rect 574134 681940 574140 681942
rect 574204 681940 574210 682004
rect 356830 681804 356836 681868
rect 356900 681866 356906 681868
rect 505093 681866 505159 681869
rect 356900 681864 505159 681866
rect 356900 681808 505098 681864
rect 505154 681808 505159 681864
rect 356900 681806 505159 681808
rect 356900 681804 356906 681806
rect 505093 681803 505159 681806
rect 549437 681866 549503 681869
rect 578550 681866 578556 681868
rect 549437 681864 578556 681866
rect 549437 681808 549442 681864
rect 549498 681808 578556 681864
rect 549437 681806 578556 681808
rect 549437 681803 549503 681806
rect 578550 681804 578556 681806
rect 578620 681804 578626 681868
rect 405590 681124 405596 681188
rect 405660 681186 405666 681188
rect 440325 681186 440391 681189
rect 405660 681184 440391 681186
rect 405660 681128 440330 681184
rect 440386 681128 440391 681184
rect 405660 681126 440391 681128
rect 405660 681124 405666 681126
rect 440325 681123 440391 681126
rect 467005 681186 467071 681189
rect 555141 681186 555207 681189
rect 467005 681184 555207 681186
rect 467005 681128 467010 681184
rect 467066 681128 555146 681184
rect 555202 681128 555207 681184
rect 467005 681126 555207 681128
rect 467005 681123 467071 681126
rect 555141 681123 555207 681126
rect 400070 680988 400076 681052
rect 400140 681050 400146 681052
rect 472157 681050 472223 681053
rect 400140 681048 472223 681050
rect 400140 680992 472162 681048
rect 472218 680992 472223 681048
rect 400140 680990 472223 680992
rect 400140 680988 400146 680990
rect 472157 680987 472223 680990
rect 481173 681050 481239 681053
rect 575422 681050 575428 681052
rect 481173 681048 575428 681050
rect 481173 680992 481178 681048
rect 481234 680992 575428 681048
rect 481173 680990 575428 680992
rect 481173 680987 481239 680990
rect 575422 680988 575428 680990
rect 575492 680988 575498 681052
rect 363689 680914 363755 680917
rect 488717 680914 488783 680917
rect 363689 680912 488783 680914
rect 363689 680856 363694 680912
rect 363750 680856 488722 680912
rect 488778 680856 488783 680912
rect 363689 680854 488783 680856
rect 363689 680851 363755 680854
rect 488717 680851 488783 680854
rect 359406 680716 359412 680780
rect 359476 680778 359482 680780
rect 427813 680778 427879 680781
rect 359476 680776 427879 680778
rect 359476 680720 427818 680776
rect 427874 680720 427879 680776
rect 359476 680718 427879 680720
rect 359476 680716 359482 680718
rect 427813 680715 427879 680718
rect 441245 680778 441311 680781
rect 565854 680778 565860 680780
rect 441245 680776 565860 680778
rect 441245 680720 441250 680776
rect 441306 680720 565860 680776
rect 441245 680718 565860 680720
rect 441245 680715 441311 680718
rect 565854 680716 565860 680718
rect 565924 680716 565930 680780
rect 367686 680580 367692 680644
rect 367756 680642 367762 680644
rect 500493 680642 500559 680645
rect 367756 680640 500559 680642
rect 367756 680584 500498 680640
rect 500554 680584 500559 680640
rect 367756 680582 500559 680584
rect 367756 680580 367762 680582
rect 500493 680579 500559 680582
rect 369853 680506 369919 680509
rect 518985 680506 519051 680509
rect 369853 680504 519051 680506
rect 369853 680448 369858 680504
rect 369914 680448 518990 680504
rect 519046 680448 519051 680504
rect 369853 680446 519051 680448
rect 369853 680443 369919 680446
rect 518985 680443 519051 680446
rect 394233 680370 394299 680373
rect 550173 680370 550239 680373
rect 394233 680368 550239 680370
rect 394233 680312 394238 680368
rect 394294 680312 550178 680368
rect 550234 680312 550239 680368
rect 394233 680310 550239 680312
rect 394233 680307 394299 680310
rect 550173 680307 550239 680310
rect 9673 680098 9739 680101
rect 433839 680098 433905 680101
rect 9673 680096 433905 680098
rect 9673 680040 9678 680096
rect 9734 680040 433844 680096
rect 433900 680040 433905 680096
rect 9673 680038 433905 680040
rect 9673 680035 9739 680038
rect 433839 680035 433905 680038
rect 409638 679764 409644 679828
rect 409708 679826 409714 679828
rect 552841 679826 552907 679829
rect 409708 679824 552907 679826
rect 409708 679768 552846 679824
rect 552902 679768 552907 679824
rect 409708 679766 552907 679768
rect 409708 679764 409714 679766
rect 552841 679763 552907 679766
rect 405365 679690 405431 679693
rect 553577 679690 553643 679693
rect 405365 679688 553643 679690
rect 405365 679632 405370 679688
rect 405426 679632 553582 679688
rect 553638 679632 553643 679688
rect 405365 679630 553643 679632
rect 405365 679627 405431 679630
rect 553577 679627 553643 679630
rect 35249 679554 35315 679557
rect 489729 679554 489795 679557
rect 35249 679552 489795 679554
rect 35249 679496 35254 679552
rect 35310 679496 489734 679552
rect 489790 679496 489795 679552
rect 35249 679494 489795 679496
rect 35249 679491 35315 679494
rect 489729 679491 489795 679494
rect 408309 679418 408375 679421
rect 552013 679418 552079 679421
rect 408309 679416 410044 679418
rect 408309 679360 408314 679416
rect 408370 679360 410044 679416
rect 408309 679358 410044 679360
rect 549884 679416 552079 679418
rect 549884 679360 552018 679416
rect 552074 679360 552079 679416
rect 549884 679358 552079 679360
rect 408309 679355 408375 679358
rect 552013 679355 552079 679358
rect 550173 678738 550239 678741
rect 549884 678736 550239 678738
rect 549884 678680 550178 678736
rect 550234 678680 550239 678736
rect 549884 678678 550239 678680
rect 550173 678675 550239 678678
rect 408350 678268 408356 678332
rect 408420 678330 408426 678332
rect 409822 678330 409828 678332
rect 408420 678270 409828 678330
rect 408420 678268 408426 678270
rect 409822 678268 409828 678270
rect 409892 678268 409898 678332
rect 407113 678058 407179 678061
rect 552013 678058 552079 678061
rect 407113 678056 410044 678058
rect 407113 678000 407118 678056
rect 407174 678000 410044 678056
rect 407113 677998 410044 678000
rect 549884 678056 552079 678058
rect 549884 678000 552018 678056
rect 552074 678000 552079 678056
rect 549884 677998 552079 678000
rect 407113 677995 407179 677998
rect 552013 677995 552079 677998
rect 166758 676092 166764 676156
rect 166828 676154 166834 676156
rect 166901 676154 166967 676157
rect 166828 676152 166967 676154
rect 166828 676096 166906 676152
rect 166962 676096 166967 676152
rect 166828 676094 166967 676096
rect 166828 676092 166834 676094
rect 166901 676091 166967 676094
rect 552013 676018 552079 676021
rect 549884 676016 552079 676018
rect 549884 675960 552018 676016
rect 552074 675960 552079 676016
rect 549884 675958 552079 675960
rect 552013 675955 552079 675958
rect 155718 675004 155724 675068
rect 155788 675066 155794 675068
rect 346894 675066 346900 675068
rect 155788 675006 346900 675066
rect 155788 675004 155794 675006
rect 346894 675004 346900 675006
rect 346964 675004 346970 675068
rect 154481 674932 154547 674933
rect 328545 674932 328611 674933
rect 154430 674930 154436 674932
rect 154390 674870 154436 674930
rect 154500 674928 154547 674932
rect 328494 674930 328500 674932
rect 154542 674872 154547 674928
rect 154430 674868 154436 674870
rect 154500 674868 154547 674872
rect 328454 674870 328500 674930
rect 328564 674928 328611 674932
rect 328606 674872 328611 674928
rect 328494 674868 328500 674870
rect 328564 674868 328611 674872
rect 154481 674867 154547 674868
rect 328545 674867 328611 674868
rect 329741 674932 329807 674933
rect 340873 674932 340939 674933
rect 329741 674928 329788 674932
rect 329852 674930 329858 674932
rect 340822 674930 340828 674932
rect 329741 674872 329746 674928
rect 329741 674868 329788 674872
rect 329852 674870 329898 674930
rect 340782 674870 340828 674930
rect 340892 674928 340939 674932
rect 340934 674872 340939 674928
rect 329852 674868 329858 674870
rect 340822 674868 340828 674870
rect 340892 674868 340939 674872
rect 329741 674867 329807 674868
rect 340873 674867 340939 674868
rect 552289 674658 552355 674661
rect 549884 674656 552355 674658
rect 549884 674600 552294 674656
rect 552350 674600 552355 674656
rect 549884 674598 552355 674600
rect 552289 674595 552355 674598
rect 552238 673978 552244 673980
rect 549884 673918 552244 673978
rect 552238 673916 552244 673918
rect 552308 673916 552314 673980
rect 549884 672490 550282 672550
rect 550222 672482 550282 672490
rect 552013 672482 552079 672485
rect 550222 672480 552079 672482
rect 550222 672424 552018 672480
rect 552074 672424 552079 672480
rect 550222 672422 552079 672424
rect 552013 672419 552079 672422
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580901 670714 580967 670717
rect 583520 670714 584960 670804
rect 580901 670712 584960 670714
rect 580901 670656 580906 670712
rect 580962 670656 584960 670712
rect 580901 670654 584960 670656
rect 580901 670651 580967 670654
rect 407113 670578 407179 670581
rect 553025 670578 553091 670581
rect 407113 670576 410044 670578
rect 407113 670520 407118 670576
rect 407174 670520 410044 670576
rect 407113 670518 410044 670520
rect 549884 670576 553091 670578
rect 549884 670520 553030 670576
rect 553086 670520 553091 670576
rect 583520 670564 584960 670654
rect 549884 670518 553091 670520
rect 407113 670515 407179 670518
rect 553025 670515 553091 670518
rect 580942 669898 580948 669900
rect 549884 669838 580948 669898
rect 580942 669836 580948 669838
rect 581012 669836 581018 669900
rect 346564 669218 347146 669220
rect 349153 669218 349219 669221
rect 346564 669216 349219 669218
rect 172562 668677 172622 669190
rect 346564 669160 349158 669216
rect 349214 669160 349219 669216
rect 347086 669158 349219 669160
rect 349153 669155 349219 669158
rect 407113 669218 407179 669221
rect 407113 669216 410044 669218
rect 407113 669160 407118 669216
rect 407174 669160 410044 669216
rect 407113 669158 410044 669160
rect 407113 669155 407179 669158
rect 172562 668672 172671 668677
rect 172562 668616 172610 668672
rect 172666 668616 172671 668672
rect 172562 668614 172671 668616
rect 172605 668611 172671 668614
rect 557574 668538 557580 668540
rect 549884 668478 557580 668538
rect 557574 668476 557580 668478
rect 557644 668476 557650 668540
rect 406745 667858 406811 667861
rect 553301 667858 553367 667861
rect 406745 667856 410044 667858
rect 406745 667800 406750 667856
rect 406806 667800 410044 667856
rect 406745 667798 410044 667800
rect 549884 667856 553367 667858
rect 549884 667800 553306 667856
rect 553362 667800 553367 667856
rect 549884 667798 553367 667800
rect 406745 667795 406811 667798
rect 553301 667795 553367 667798
rect 407205 667178 407271 667181
rect 407205 667176 410044 667178
rect 407205 667120 407210 667176
rect 407266 667120 410044 667176
rect 407205 667118 410044 667120
rect 407205 667115 407271 667118
rect 407113 666498 407179 666501
rect 571374 666498 571380 666500
rect 407113 666496 410044 666498
rect 407113 666440 407118 666496
rect 407174 666440 410044 666496
rect 407113 666438 410044 666440
rect 549884 666438 571380 666498
rect 407113 666435 407179 666438
rect 571374 666436 571380 666438
rect 571444 666436 571450 666500
rect 552841 665818 552907 665821
rect 549884 665816 552907 665818
rect 549884 665760 552846 665816
rect 552902 665760 552907 665816
rect 549884 665758 552907 665760
rect 552841 665755 552907 665758
rect 408401 665138 408467 665141
rect 408401 665136 410044 665138
rect 408401 665080 408406 665136
rect 408462 665080 410044 665136
rect 408401 665078 410044 665080
rect 408401 665075 408467 665078
rect 407205 663778 407271 663781
rect 566038 663778 566044 663780
rect 407205 663776 410044 663778
rect 407205 663720 407210 663776
rect 407266 663720 410044 663776
rect 407205 663718 410044 663720
rect 549884 663718 566044 663778
rect 407205 663715 407271 663718
rect 566038 663716 566044 663718
rect 566108 663716 566114 663780
rect 407389 662418 407455 662421
rect 407389 662416 410044 662418
rect 407389 662360 407394 662416
rect 407450 662360 410044 662416
rect 407389 662358 410044 662360
rect 407389 662355 407455 662358
rect 407205 661738 407271 661741
rect 552197 661738 552263 661741
rect 407205 661736 410044 661738
rect 407205 661680 407210 661736
rect 407266 661680 410044 661736
rect 407205 661678 410044 661680
rect 549884 661736 552263 661738
rect 549884 661680 552202 661736
rect 552258 661680 552263 661736
rect 549884 661678 552263 661680
rect 407205 661675 407271 661678
rect 552197 661675 552263 661678
rect 407297 661058 407363 661061
rect 407297 661056 410044 661058
rect 407297 661000 407302 661056
rect 407358 661000 410044 661056
rect 407297 660998 410044 661000
rect 407297 660995 407363 660998
rect 407297 659018 407363 659021
rect 407297 659016 410044 659018
rect 407297 658960 407302 659016
rect 407358 658960 410044 659016
rect 407297 658958 410044 658960
rect 407297 658955 407363 658958
rect -960 658202 480 658292
rect 3325 658202 3391 658205
rect -960 658200 3391 658202
rect -960 658144 3330 658200
rect 3386 658144 3391 658200
rect -960 658142 3391 658144
rect -960 658052 480 658142
rect 3325 658139 3391 658142
rect 370446 657596 370452 657660
rect 370516 657658 370522 657660
rect 370516 657598 410044 657658
rect 370516 657596 370522 657598
rect 583520 657236 584960 657476
rect 553301 656978 553367 656981
rect 549884 656976 553367 656978
rect 549884 656920 553306 656976
rect 553362 656920 553367 656976
rect 549884 656918 553367 656920
rect 553301 656915 553367 656918
rect 407205 654938 407271 654941
rect 407205 654936 410044 654938
rect 407205 654880 407210 654936
rect 407266 654880 410044 654936
rect 407205 654878 410044 654880
rect 407205 654875 407271 654878
rect 407205 654258 407271 654261
rect 552565 654258 552631 654261
rect 407205 654256 410044 654258
rect 407205 654200 407210 654256
rect 407266 654200 410044 654256
rect 407205 654198 410044 654200
rect 549884 654256 552631 654258
rect 549884 654200 552570 654256
rect 552626 654200 552631 654256
rect 549884 654198 552631 654200
rect 407205 654195 407271 654198
rect 552565 654195 552631 654198
rect 552105 653578 552171 653581
rect 549884 653576 552171 653578
rect 549884 653520 552110 653576
rect 552166 653520 552171 653576
rect 549884 653518 552171 653520
rect 552105 653515 552171 653518
rect 407205 652898 407271 652901
rect 407205 652896 410044 652898
rect 407205 652840 407210 652896
rect 407266 652840 410044 652896
rect 407205 652838 410044 652840
rect 407205 652835 407271 652838
rect 402094 652156 402100 652220
rect 402164 652218 402170 652220
rect 402164 652158 410044 652218
rect 402164 652156 402170 652158
rect 575606 650858 575612 650860
rect 549884 650798 575612 650858
rect 575606 650796 575612 650798
rect 575676 650796 575682 650860
rect 407205 650178 407271 650181
rect 408217 650178 408283 650181
rect 551553 650178 551619 650181
rect 407205 650176 410044 650178
rect 407205 650120 407210 650176
rect 407266 650120 408222 650176
rect 408278 650120 410044 650176
rect 407205 650118 410044 650120
rect 549884 650176 551619 650178
rect 549884 650120 551558 650176
rect 551614 650120 551619 650176
rect 549884 650118 551619 650120
rect 407205 650115 407271 650118
rect 408217 650115 408283 650118
rect 551553 650115 551619 650118
rect 407205 649498 407271 649501
rect 556102 649498 556108 649500
rect 407205 649496 410044 649498
rect 407205 649440 407210 649496
rect 407266 649440 410044 649496
rect 407205 649438 410044 649440
rect 549884 649438 556108 649498
rect 407205 649435 407271 649438
rect 556102 649436 556108 649438
rect 556172 649436 556178 649500
rect 407481 648818 407547 648821
rect 553301 648818 553367 648821
rect 407481 648816 410044 648818
rect 407481 648760 407486 648816
rect 407542 648760 410044 648816
rect 407481 648758 410044 648760
rect 549884 648816 553367 648818
rect 549884 648760 553306 648816
rect 553362 648760 553367 648816
rect 549884 648758 553367 648760
rect 407481 648755 407547 648758
rect 553301 648755 553367 648758
rect 408401 646778 408467 646781
rect 552565 646778 552631 646781
rect 408401 646776 410044 646778
rect 408401 646720 408406 646776
rect 408462 646720 410044 646776
rect 408401 646718 410044 646720
rect 549884 646776 552631 646778
rect 549884 646720 552570 646776
rect 552626 646720 552631 646776
rect 549884 646718 552631 646720
rect 408401 646715 408467 646718
rect 552565 646715 552631 646718
rect 579654 646098 579660 646100
rect 549884 646038 579660 646098
rect 579654 646036 579660 646038
rect 579724 646036 579730 646100
rect 401358 645356 401364 645420
rect 401428 645418 401434 645420
rect 552105 645418 552171 645421
rect 401428 645358 410044 645418
rect 549884 645416 552171 645418
rect 549884 645360 552110 645416
rect 552166 645360 552171 645416
rect 549884 645358 552171 645360
rect 401428 645356 401434 645358
rect 552105 645355 552171 645358
rect -960 644996 480 645236
rect 407205 644738 407271 644741
rect 553209 644738 553275 644741
rect 407205 644736 410044 644738
rect 407205 644680 407210 644736
rect 407266 644680 410044 644736
rect 407205 644678 410044 644680
rect 549884 644736 553275 644738
rect 549884 644680 553214 644736
rect 553270 644680 553275 644736
rect 549884 644678 553275 644680
rect 407205 644675 407271 644678
rect 553209 644675 553275 644678
rect 407021 644058 407087 644061
rect 579981 644058 580047 644061
rect 583520 644058 584960 644148
rect 407021 644056 410044 644058
rect 407021 644000 407026 644056
rect 407082 644000 410044 644056
rect 407021 643998 410044 644000
rect 579981 644056 584960 644058
rect 579981 644000 579986 644056
rect 580042 644000 584960 644056
rect 579981 643998 584960 644000
rect 407021 643995 407087 643998
rect 579981 643995 580047 643998
rect 583520 643908 584960 643998
rect 552473 642698 552539 642701
rect 550222 642696 552539 642698
rect 550222 642640 552478 642696
rect 552534 642640 552539 642696
rect 550222 642638 552539 642640
rect 550222 642630 550282 642638
rect 552473 642635 552539 642638
rect 406377 642154 406443 642157
rect 410014 642154 410074 642600
rect 549884 642570 550282 642630
rect 406377 642152 410074 642154
rect 406377 642096 406382 642152
rect 406438 642096 410074 642152
rect 406377 642094 410074 642096
rect 406377 642091 406443 642094
rect 407205 642018 407271 642021
rect 552013 642018 552079 642021
rect 407205 642016 410044 642018
rect 407205 641960 407210 642016
rect 407266 641960 410044 642016
rect 407205 641958 410044 641960
rect 549884 642016 552079 642018
rect 549884 641960 552018 642016
rect 552074 641960 552079 642016
rect 549884 641958 552079 641960
rect 407205 641955 407271 641958
rect 552013 641955 552079 641958
rect 407205 641338 407271 641341
rect 553301 641338 553367 641341
rect 407205 641336 410044 641338
rect 407205 641280 407210 641336
rect 407266 641280 410044 641336
rect 407205 641278 410044 641280
rect 549884 641336 553367 641338
rect 549884 641280 553306 641336
rect 553362 641280 553367 641336
rect 549884 641278 553367 641280
rect 407205 641275 407271 641278
rect 553301 641275 553367 641278
rect 407297 638074 407363 638077
rect 410014 638074 410074 638520
rect 549884 638490 550282 638550
rect 550222 638482 550282 638490
rect 550222 638422 550650 638482
rect 550590 638346 550650 638422
rect 552105 638346 552171 638349
rect 550590 638344 552171 638346
rect 550590 638288 552110 638344
rect 552166 638288 552171 638344
rect 550590 638286 552171 638288
rect 552105 638283 552171 638286
rect 407297 638072 410074 638074
rect 407297 638016 407302 638072
rect 407358 638016 410074 638072
rect 407297 638014 410074 638016
rect 407297 638011 407363 638014
rect 407205 637938 407271 637941
rect 552013 637938 552079 637941
rect 407205 637936 410044 637938
rect 407205 637880 407210 637936
rect 407266 637880 410044 637936
rect 407205 637878 410044 637880
rect 549884 637936 552079 637938
rect 549884 637880 552018 637936
rect 552074 637880 552079 637936
rect 549884 637878 552079 637880
rect 407205 637875 407271 637878
rect 552013 637875 552079 637878
rect 407205 637258 407271 637261
rect 407205 637256 410044 637258
rect 407205 637200 407210 637256
rect 407266 637200 410044 637256
rect 407205 637198 410044 637200
rect 407205 637195 407271 637198
rect 368974 635836 368980 635900
rect 369044 635898 369050 635900
rect 369044 635838 410044 635898
rect 369044 635836 369050 635838
rect 552381 634538 552447 634541
rect 549884 634536 552447 634538
rect 549884 634480 552386 634536
rect 552442 634480 552447 634536
rect 549884 634478 552447 634480
rect 552381 634475 552447 634478
rect 407205 633858 407271 633861
rect 557758 633858 557764 633860
rect 407205 633856 410044 633858
rect 407205 633800 407210 633856
rect 407266 633800 410044 633856
rect 407205 633798 410044 633800
rect 549884 633798 557764 633858
rect 407205 633795 407271 633798
rect 557758 633796 557764 633798
rect 557828 633796 557834 633860
rect 407205 632498 407271 632501
rect 407205 632496 410044 632498
rect 407205 632440 407210 632496
rect 407266 632440 410044 632496
rect 407205 632438 410044 632440
rect 407205 632435 407271 632438
rect -960 631940 480 632180
rect 406929 631818 406995 631821
rect 552013 631818 552079 631821
rect 406929 631816 410044 631818
rect 406929 631760 406934 631816
rect 406990 631760 410044 631816
rect 406929 631758 410044 631760
rect 549884 631816 552079 631818
rect 549884 631760 552018 631816
rect 552074 631760 552079 631816
rect 549884 631758 552079 631760
rect 406929 631755 406995 631758
rect 552013 631755 552079 631758
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 557942 630458 557948 630460
rect 549884 630398 557948 630458
rect 557942 630396 557948 630398
rect 558012 630396 558018 630460
rect 407205 629098 407271 629101
rect 407205 629096 410044 629098
rect 407205 629040 407210 629096
rect 407266 629040 410044 629096
rect 407205 629038 410044 629040
rect 407205 629035 407271 629038
rect 404118 628356 404124 628420
rect 404188 628418 404194 628420
rect 571558 628418 571564 628420
rect 404188 628358 410044 628418
rect 549884 628358 571564 628418
rect 404188 628356 404194 628358
rect 571558 628356 571564 628358
rect 571628 628356 571634 628420
rect 406510 627676 406516 627740
rect 406580 627738 406586 627740
rect 406580 627678 410044 627738
rect 406580 627676 406586 627678
rect 560702 627058 560708 627060
rect 549884 626998 560708 627058
rect 560702 626996 560708 626998
rect 560772 626996 560778 627060
rect 35617 626922 35683 626925
rect 35850 626922 36064 626924
rect 35617 626920 36064 626922
rect 35617 626864 35622 626920
rect 35678 626864 36064 626920
rect 35617 626862 35910 626864
rect 35617 626859 35683 626862
rect 208301 626650 208367 626653
rect 210002 626650 210062 626894
rect 208301 626648 210062 626650
rect 208301 626592 208306 626648
rect 208362 626592 210062 626648
rect 208301 626590 210062 626592
rect 208301 626587 208367 626590
rect 34237 625970 34303 625973
rect 35850 625970 36064 625972
rect 34237 625968 36064 625970
rect 34237 625912 34242 625968
rect 34298 625912 36064 625968
rect 34237 625910 35910 625912
rect 34237 625907 34303 625910
rect 207657 625426 207723 625429
rect 210002 625426 210062 625942
rect 207657 625424 210062 625426
rect 207657 625368 207662 625424
rect 207718 625368 210062 625424
rect 207657 625366 210062 625368
rect 407021 625426 407087 625429
rect 410014 625426 410074 625600
rect 549884 625570 550282 625630
rect 550222 625562 550282 625570
rect 550222 625502 550650 625562
rect 407021 625424 410074 625426
rect 407021 625368 407026 625424
rect 407082 625368 410074 625424
rect 407021 625366 410074 625368
rect 550590 625426 550650 625502
rect 552013 625426 552079 625429
rect 550590 625424 552079 625426
rect 550590 625368 552018 625424
rect 552074 625368 552079 625424
rect 550590 625366 552079 625368
rect 207657 625363 207723 625366
rect 407021 625363 407087 625366
rect 552013 625363 552079 625366
rect 405406 624276 405412 624340
rect 405476 624338 405482 624340
rect 552013 624338 552079 624341
rect 405476 624278 410044 624338
rect 549884 624336 552079 624338
rect 549884 624280 552018 624336
rect 552074 624280 552079 624336
rect 549884 624278 552079 624280
rect 405476 624276 405482 624278
rect 552013 624275 552079 624278
rect 34421 623794 34487 623797
rect 35850 623794 36064 623796
rect 34421 623792 36064 623794
rect 34421 623736 34426 623792
rect 34482 623736 36064 623792
rect 207749 623794 207815 623797
rect 207749 623792 210062 623794
rect 207749 623736 207754 623792
rect 207810 623736 210062 623792
rect 34421 623734 35910 623736
rect 207749 623734 210062 623736
rect 34421 623731 34487 623734
rect 207749 623731 207815 623734
rect 378726 622916 378732 622980
rect 378796 622978 378802 622980
rect 550633 622978 550699 622981
rect 378796 622918 410044 622978
rect 549884 622976 550699 622978
rect 549884 622920 550638 622976
rect 550694 622920 550699 622976
rect 549884 622918 550699 622920
rect 378796 622916 378802 622918
rect 550633 622915 550699 622918
rect 34145 622842 34211 622845
rect 35850 622842 36064 622844
rect 34145 622840 36064 622842
rect 34145 622784 34150 622840
rect 34206 622784 36064 622840
rect 34145 622782 35910 622784
rect 34145 622779 34211 622782
rect 208209 622434 208275 622437
rect 210002 622434 210062 622814
rect 208209 622432 210062 622434
rect 208209 622376 208214 622432
rect 208270 622376 210062 622432
rect 208209 622374 210062 622376
rect 208209 622371 208275 622374
rect 35433 621074 35499 621077
rect 35850 621074 36064 621076
rect 35433 621072 36064 621074
rect 35433 621016 35438 621072
rect 35494 621016 36064 621072
rect 208117 621074 208183 621077
rect 208117 621072 210062 621074
rect 208117 621016 208122 621072
rect 208178 621016 210062 621072
rect 35433 621014 35910 621016
rect 208117 621014 210062 621016
rect 35433 621011 35499 621014
rect 208117 621011 208183 621014
rect 552565 620258 552631 620261
rect 549884 620256 552631 620258
rect 549884 620200 552570 620256
rect 552626 620200 552631 620256
rect 549884 620198 552631 620200
rect 552565 620195 552631 620198
rect 34881 619986 34947 619989
rect 209681 619988 209747 619989
rect 35850 619986 36064 619988
rect 34881 619984 36064 619986
rect 34881 619928 34886 619984
rect 34942 619928 36064 619984
rect 209681 619984 210032 619988
rect 209681 619928 209686 619984
rect 209742 619928 210032 619984
rect 34881 619926 35910 619928
rect 209681 619926 209790 619928
rect 34881 619923 34947 619926
rect 209681 619923 209747 619926
rect 407297 619578 407363 619581
rect 407297 619576 410044 619578
rect 407297 619520 407302 619576
rect 407358 619520 410044 619576
rect 407297 619518 410044 619520
rect 407297 619515 407363 619518
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 407205 618898 407271 618901
rect 407205 618896 410044 618898
rect 407205 618840 407210 618896
rect 407266 618840 410044 618896
rect 407205 618838 410044 618840
rect 407205 618835 407271 618838
rect 35525 618218 35591 618221
rect 35850 618218 36064 618220
rect 35525 618216 36064 618218
rect 35525 618160 35530 618216
rect 35586 618160 36064 618216
rect 35525 618158 35910 618160
rect 35525 618155 35591 618158
rect 208025 617674 208091 617677
rect 210002 617674 210062 618190
rect 208025 617672 210062 617674
rect 208025 617616 208030 617672
rect 208086 617616 210062 617672
rect 208025 617614 210062 617616
rect 208025 617611 208091 617614
rect 553301 617538 553367 617541
rect 549884 617536 553367 617538
rect 549884 617480 553306 617536
rect 553362 617480 553367 617536
rect 549884 617478 553367 617480
rect 553301 617475 553367 617478
rect 580809 617538 580875 617541
rect 583520 617538 584960 617628
rect 580809 617536 584960 617538
rect 580809 617480 580814 617536
rect 580870 617480 584960 617536
rect 580809 617478 584960 617480
rect 580809 617475 580875 617478
rect 583520 617388 584960 617478
rect 407297 616858 407363 616861
rect 407297 616856 410044 616858
rect 407297 616800 407302 616856
rect 407358 616800 410044 616856
rect 407297 616798 410044 616800
rect 407297 616795 407363 616798
rect 561806 616178 561812 616180
rect 549884 616118 561812 616178
rect 561806 616116 561812 616118
rect 561876 616116 561882 616180
rect 407297 614954 407363 614957
rect 410014 614954 410074 615468
rect 407297 614952 410074 614954
rect 407297 614896 407302 614952
rect 407358 614896 410074 614952
rect 407297 614894 410074 614896
rect 407297 614891 407363 614894
rect 407665 614818 407731 614821
rect 552238 614818 552244 614820
rect 407665 614816 410044 614818
rect 407665 614760 407670 614816
rect 407726 614760 410044 614816
rect 407665 614758 410044 614760
rect 549884 614758 552244 614818
rect 407665 614755 407731 614758
rect 552238 614756 552244 614758
rect 552308 614756 552314 614820
rect 553209 613458 553275 613461
rect 549884 613456 553275 613458
rect 549884 613400 553214 613456
rect 553270 613400 553275 613456
rect 549884 613398 553275 613400
rect 553209 613395 553275 613398
rect 407205 612778 407271 612781
rect 553301 612778 553367 612781
rect 407205 612776 410044 612778
rect 407205 612720 407210 612776
rect 407266 612720 410044 612776
rect 407205 612718 410044 612720
rect 549884 612776 553367 612778
rect 549884 612720 553306 612776
rect 553362 612720 553367 612776
rect 549884 612718 553367 612720
rect 407205 612715 407271 612718
rect 553301 612715 553367 612718
rect 556654 612098 556660 612100
rect 549884 612038 556660 612098
rect 556654 612036 556660 612038
rect 556724 612036 556730 612100
rect 377254 611356 377260 611420
rect 377324 611418 377330 611420
rect 553301 611418 553367 611421
rect 377324 611358 410044 611418
rect 549884 611416 553367 611418
rect 549884 611360 553306 611416
rect 553362 611360 553367 611416
rect 549884 611358 553367 611360
rect 377324 611356 377330 611358
rect 553301 611355 553367 611358
rect 553301 610738 553367 610741
rect 549884 610736 553367 610738
rect 549884 610680 553306 610736
rect 553362 610680 553367 610736
rect 549884 610678 553367 610680
rect 553301 610675 553367 610678
rect 346564 609378 347146 609380
rect 350441 609378 350507 609381
rect 346564 609376 350507 609378
rect 172562 608834 172622 609350
rect 346564 609320 350446 609376
rect 350502 609320 350507 609376
rect 347086 609318 350507 609320
rect 350441 609315 350507 609318
rect 175273 608834 175339 608837
rect 172562 608832 175339 608834
rect 172562 608776 175278 608832
rect 175334 608776 175339 608832
rect 172562 608774 175339 608776
rect 175273 608771 175339 608774
rect 407205 608698 407271 608701
rect 552473 608698 552539 608701
rect 407205 608696 410044 608698
rect 407205 608640 407210 608696
rect 407266 608640 410044 608696
rect 407205 608638 410044 608640
rect 550222 608696 552539 608698
rect 550222 608640 552478 608696
rect 552534 608640 552539 608696
rect 550222 608638 552539 608640
rect 407205 608635 407271 608638
rect 550222 608630 550282 608638
rect 552473 608635 552539 608638
rect 549884 608570 550282 608630
rect 556286 608018 556292 608020
rect 549884 607958 556292 608018
rect 556286 607956 556292 607958
rect 556356 607956 556362 608020
rect 346564 607746 347146 607748
rect 349245 607746 349311 607749
rect 346564 607744 349311 607746
rect 172562 607338 172622 607718
rect 346564 607688 349250 607744
rect 349306 607688 349311 607744
rect 347086 607686 349311 607688
rect 349245 607683 349311 607686
rect 176561 607338 176627 607341
rect 172562 607336 176627 607338
rect 172562 607280 176566 607336
rect 176622 607280 176627 607336
rect 172562 607278 176627 607280
rect 176561 607275 176627 607278
rect 399518 607276 399524 607340
rect 399588 607338 399594 607340
rect 552197 607338 552263 607341
rect 399588 607278 410044 607338
rect 549884 607336 552263 607338
rect 549884 607280 552202 607336
rect 552258 607280 552263 607336
rect 549884 607278 552263 607280
rect 399588 607276 399594 607278
rect 552197 607275 552263 607278
rect 346564 606386 347146 606388
rect 350441 606386 350507 606389
rect 346564 606384 350507 606386
rect -960 606114 480 606204
rect 3693 606114 3759 606117
rect -960 606112 3759 606114
rect -960 606056 3698 606112
rect 3754 606056 3759 606112
rect -960 606054 3759 606056
rect -960 605964 480 606054
rect 3693 606051 3759 606054
rect 172562 605978 172622 606358
rect 346564 606328 350446 606384
rect 350502 606328 350507 606384
rect 347086 606326 350507 606328
rect 350441 606323 350507 606326
rect 176561 605978 176627 605981
rect 172562 605976 176627 605978
rect 172562 605920 176566 605976
rect 176622 605920 176627 605976
rect 172562 605918 176627 605920
rect 176561 605915 176627 605918
rect 407941 605978 408007 605981
rect 553301 605978 553367 605981
rect 407941 605976 410044 605978
rect 407941 605920 407946 605976
rect 408002 605920 410044 605976
rect 407941 605918 410044 605920
rect 549884 605976 553367 605978
rect 549884 605920 553306 605976
rect 553362 605920 553367 605976
rect 549884 605918 553367 605920
rect 407941 605915 408007 605918
rect 553301 605915 553367 605918
rect 346564 604890 347146 604892
rect 350441 604890 350507 604893
rect 346564 604888 350507 604890
rect 172562 604482 172622 604862
rect 346564 604832 350446 604888
rect 350502 604832 350507 604888
rect 347086 604830 350507 604832
rect 350441 604827 350507 604830
rect 409462 604490 410044 604550
rect 175365 604482 175431 604485
rect 172562 604480 175431 604482
rect 172562 604424 175370 604480
rect 175426 604424 175431 604480
rect 172562 604422 175431 604424
rect 175365 604419 175431 604422
rect 387558 604420 387564 604484
rect 387628 604482 387634 604484
rect 409462 604482 409522 604490
rect 387628 604422 409522 604482
rect 387628 604420 387634 604422
rect 583520 604060 584960 604300
rect 552013 603938 552079 603941
rect 549884 603936 552079 603938
rect 549884 603880 552018 603936
rect 552074 603880 552079 603936
rect 549884 603878 552079 603880
rect 552013 603875 552079 603878
rect 346564 603666 347146 603668
rect 349337 603666 349403 603669
rect 346564 603664 349403 603666
rect 172562 603122 172622 603638
rect 346564 603608 349342 603664
rect 349398 603608 349403 603664
rect 347086 603606 349403 603608
rect 349337 603603 349403 603606
rect 553301 603258 553367 603261
rect 549884 603256 553367 603258
rect 549884 603200 553306 603256
rect 553362 603200 553367 603256
rect 549884 603198 553367 603200
rect 553301 603195 553367 603198
rect 175457 603122 175523 603125
rect 172562 603120 175523 603122
rect 172562 603064 175462 603120
rect 175518 603064 175523 603120
rect 172562 603062 175523 603064
rect 175457 603059 175523 603062
rect 407297 602578 407363 602581
rect 578734 602578 578740 602580
rect 407297 602576 410044 602578
rect 407297 602520 407302 602576
rect 407358 602520 410044 602576
rect 407297 602518 410044 602520
rect 549884 602518 578740 602578
rect 407297 602515 407363 602518
rect 578734 602516 578740 602518
rect 578804 602516 578810 602580
rect 407297 601898 407363 601901
rect 570086 601898 570092 601900
rect 407297 601896 410044 601898
rect 407297 601840 407302 601896
rect 407358 601840 410044 601896
rect 407297 601838 410044 601840
rect 549884 601838 570092 601898
rect 407297 601835 407363 601838
rect 570086 601836 570092 601838
rect 570156 601836 570162 601900
rect 407798 601156 407804 601220
rect 407868 601218 407874 601220
rect 407868 601158 410044 601218
rect 407868 601156 407874 601158
rect 552289 600538 552355 600541
rect 549884 600536 552355 600538
rect 549884 600480 552294 600536
rect 552350 600480 552355 600536
rect 549884 600478 552355 600480
rect 552289 600475 552355 600478
rect 35709 599994 35775 599997
rect 35850 599994 36064 599996
rect 35709 599992 36064 599994
rect 35709 599936 35714 599992
rect 35770 599936 36064 599992
rect 35709 599934 35910 599936
rect 35709 599931 35775 599934
rect 207013 599450 207079 599453
rect 210002 599450 210062 599966
rect 553301 599858 553367 599861
rect 549884 599856 553367 599858
rect 549884 599800 553306 599856
rect 553362 599800 553367 599856
rect 549884 599798 553367 599800
rect 553301 599795 553367 599798
rect 207013 599448 210062 599450
rect 207013 599392 207018 599448
rect 207074 599392 210062 599448
rect 207013 599390 210062 599392
rect 207013 599387 207079 599390
rect 407297 599178 407363 599181
rect 556470 599178 556476 599180
rect 407297 599176 410044 599178
rect 407297 599120 407302 599176
rect 407358 599120 410044 599176
rect 407297 599118 410044 599120
rect 549884 599118 556476 599178
rect 407297 599115 407363 599118
rect 556470 599116 556476 599118
rect 556540 599116 556546 599180
rect 382774 598436 382780 598500
rect 382844 598498 382850 598500
rect 552013 598498 552079 598501
rect 382844 598438 410044 598498
rect 549884 598496 552079 598498
rect 549884 598440 552018 598496
rect 552074 598440 552079 598496
rect 549884 598438 552079 598440
rect 382844 598436 382850 598438
rect 552013 598435 552079 598438
rect 34329 598362 34395 598365
rect 35850 598362 36064 598364
rect 34329 598360 36064 598362
rect 34329 598304 34334 598360
rect 34390 598304 36064 598360
rect 209129 598362 209195 598365
rect 209730 598362 210032 598364
rect 209129 598360 210032 598362
rect 209129 598304 209134 598360
rect 209190 598304 210032 598360
rect 34329 598302 35910 598304
rect 209129 598302 209790 598304
rect 34329 598299 34395 598302
rect 209129 598299 209195 598302
rect 34237 598090 34303 598093
rect 35850 598090 36064 598092
rect 34237 598088 36064 598090
rect 34237 598032 34242 598088
rect 34298 598032 36064 598088
rect 34237 598030 35910 598032
rect 34237 598027 34303 598030
rect 207933 597682 207999 597685
rect 210002 597682 210062 598062
rect 552933 597818 552999 597821
rect 549884 597816 552999 597818
rect 549884 597760 552938 597816
rect 552994 597760 552999 597816
rect 549884 597758 552999 597760
rect 552933 597755 552999 597758
rect 207933 597680 210062 597682
rect 207933 597624 207938 597680
rect 207994 597624 210062 597680
rect 207933 597622 210062 597624
rect 207933 597619 207999 597622
rect 551502 597484 551508 597548
rect 551572 597546 551578 597548
rect 552289 597546 552355 597549
rect 551572 597544 552355 597546
rect 551572 597488 552294 597544
rect 552350 597488 552355 597544
rect 551572 597486 552355 597488
rect 551572 597484 551578 597486
rect 552289 597483 552355 597486
rect 407297 597138 407363 597141
rect 407297 597136 410044 597138
rect 407297 597080 407302 597136
rect 407358 597080 410044 597136
rect 407297 597078 410044 597080
rect 407297 597075 407363 597078
rect 552013 596458 552079 596461
rect 549884 596456 552079 596458
rect 549884 596400 552018 596456
rect 552074 596400 552079 596456
rect 549884 596398 552079 596400
rect 552013 596395 552079 596398
rect 407297 595098 407363 595101
rect 407297 595096 410044 595098
rect 407297 595040 407302 595096
rect 407358 595040 410044 595096
rect 407297 595038 410044 595040
rect 407297 595035 407363 595038
rect 408401 594418 408467 594421
rect 408401 594416 410044 594418
rect 408401 594360 408406 594416
rect 408462 594360 410044 594416
rect 408401 594358 410044 594360
rect 408401 594355 408467 594358
rect 363454 593676 363460 593740
rect 363524 593738 363530 593740
rect 363524 593678 410044 593738
rect 363524 593676 363530 593678
rect -960 592908 480 593148
rect 407297 593058 407363 593061
rect 407297 593056 410044 593058
rect 407297 593000 407302 593056
rect 407358 593000 410044 593056
rect 407297 592998 410044 593000
rect 407297 592995 407363 592998
rect 550398 591630 550404 591632
rect 407389 591154 407455 591157
rect 410014 591154 410074 591600
rect 549884 591570 550404 591630
rect 550398 591568 550404 591570
rect 550468 591568 550474 591632
rect 407389 591152 410074 591154
rect 407389 591096 407394 591152
rect 407450 591096 410074 591152
rect 407389 591094 410074 591096
rect 407389 591091 407455 591094
rect 407297 591018 407363 591021
rect 558862 591018 558868 591020
rect 407297 591016 410044 591018
rect 407297 590960 407302 591016
rect 407358 590960 410044 591016
rect 407297 590958 410044 590960
rect 549884 590958 558868 591018
rect 407297 590955 407363 590958
rect 558862 590956 558868 590958
rect 558932 590956 558938 591020
rect 580717 591018 580783 591021
rect 583520 591018 584960 591108
rect 580717 591016 584960 591018
rect 580717 590960 580722 591016
rect 580778 590960 584960 591016
rect 580717 590958 584960 590960
rect 580717 590955 580783 590958
rect 583520 590868 584960 590958
rect 550398 590684 550404 590748
rect 550468 590746 550474 590748
rect 581126 590746 581132 590748
rect 550468 590686 581132 590746
rect 550468 590684 550474 590686
rect 581126 590684 581132 590686
rect 581196 590684 581202 590748
rect 84377 589524 84443 589525
rect 84326 589522 84332 589524
rect 84286 589462 84332 589522
rect 84396 589520 84443 589524
rect 84438 589464 84443 589520
rect 84326 589460 84332 589462
rect 84396 589460 84443 589464
rect 84377 589459 84443 589460
rect 407614 589114 407620 589116
rect 393270 589054 407620 589114
rect 257337 588978 257403 588981
rect 393270 588978 393330 589054
rect 407614 589052 407620 589054
rect 407684 589052 407690 589116
rect 257337 588976 393330 588978
rect 257337 588920 257342 588976
rect 257398 588920 393330 588976
rect 257337 588918 393330 588920
rect 407297 588978 407363 588981
rect 552105 588978 552171 588981
rect 407297 588976 410044 588978
rect 407297 588920 407302 588976
rect 407358 588920 410044 588976
rect 407297 588918 410044 588920
rect 549884 588976 552171 588978
rect 549884 588920 552110 588976
rect 552166 588920 552171 588976
rect 549884 588918 552171 588920
rect 257337 588915 257403 588918
rect 407297 588915 407363 588918
rect 552105 588915 552171 588918
rect 43846 588780 43852 588844
rect 43916 588842 43922 588844
rect 404813 588842 404879 588845
rect 43916 588840 404879 588842
rect 43916 588784 404818 588840
rect 404874 588784 404879 588840
rect 43916 588782 404879 588784
rect 43916 588780 43922 588782
rect 404813 588779 404879 588782
rect 44950 588644 44956 588708
rect 45020 588706 45026 588708
rect 407481 588706 407547 588709
rect 45020 588704 407547 588706
rect 45020 588648 407486 588704
rect 407542 588648 407547 588704
rect 45020 588646 407547 588648
rect 45020 588644 45026 588646
rect 407481 588643 407547 588646
rect 3693 588570 3759 588573
rect 388294 588570 388300 588572
rect 3693 588568 388300 588570
rect 3693 588512 3698 588568
rect 3754 588512 388300 588568
rect 3693 588510 388300 588512
rect 3693 588507 3759 588510
rect 388294 588508 388300 588510
rect 388364 588508 388370 588572
rect 52453 587890 52519 587893
rect 53046 587890 53052 587892
rect 52453 587888 53052 587890
rect 52453 587832 52458 587888
rect 52514 587832 53052 587888
rect 52453 587830 53052 587832
rect 52453 587827 52519 587830
rect 53046 587828 53052 587830
rect 53116 587828 53122 587892
rect 53833 587890 53899 587893
rect 56593 587892 56659 587893
rect 57881 587892 57947 587893
rect 54150 587890 54156 587892
rect 53833 587888 54156 587890
rect 53833 587832 53838 587888
rect 53894 587832 54156 587888
rect 53833 587830 54156 587832
rect 53833 587827 53899 587830
rect 54150 587828 54156 587830
rect 54220 587828 54226 587892
rect 56542 587890 56548 587892
rect 56502 587830 56548 587890
rect 56612 587888 56659 587892
rect 57830 587890 57836 587892
rect 56654 587832 56659 587888
rect 56542 587828 56548 587830
rect 56612 587828 56659 587832
rect 57790 587830 57836 587890
rect 57900 587888 57947 587892
rect 57942 587832 57947 587888
rect 57830 587828 57836 587830
rect 57900 587828 57947 587832
rect 56593 587827 56659 587828
rect 57881 587827 57947 587828
rect 58065 587890 58131 587893
rect 59118 587890 59124 587892
rect 58065 587888 59124 587890
rect 58065 587832 58070 587888
rect 58126 587832 59124 587888
rect 58065 587830 59124 587832
rect 58065 587827 58131 587830
rect 59118 587828 59124 587830
rect 59188 587828 59194 587892
rect 59353 587890 59419 587893
rect 60222 587890 60228 587892
rect 59353 587888 60228 587890
rect 59353 587832 59358 587888
rect 59414 587832 60228 587888
rect 59353 587830 60228 587832
rect 59353 587827 59419 587830
rect 60222 587828 60228 587830
rect 60292 587828 60298 587892
rect 62113 587890 62179 587893
rect 63493 587892 63559 587893
rect 62430 587890 62436 587892
rect 62113 587888 62436 587890
rect 62113 587832 62118 587888
rect 62174 587832 62436 587888
rect 62113 587830 62436 587832
rect 62113 587827 62179 587830
rect 62430 587828 62436 587830
rect 62500 587828 62506 587892
rect 63493 587890 63540 587892
rect 63448 587888 63540 587890
rect 63448 587832 63498 587888
rect 63448 587830 63540 587832
rect 63493 587828 63540 587830
rect 63604 587828 63610 587892
rect 63677 587890 63743 587893
rect 64270 587890 64276 587892
rect 63677 587888 64276 587890
rect 63677 587832 63682 587888
rect 63738 587832 64276 587888
rect 63677 587830 64276 587832
rect 63493 587827 63559 587828
rect 63677 587827 63743 587830
rect 64270 587828 64276 587830
rect 64340 587828 64346 587892
rect 64965 587890 65031 587893
rect 66110 587890 66116 587892
rect 64965 587888 66116 587890
rect 64965 587832 64970 587888
rect 65026 587832 66116 587888
rect 64965 587830 66116 587832
rect 64965 587827 65031 587830
rect 66110 587828 66116 587830
rect 66180 587828 66186 587892
rect 66345 587890 66411 587893
rect 66662 587890 66668 587892
rect 66345 587888 66668 587890
rect 66345 587832 66350 587888
rect 66406 587832 66668 587888
rect 66345 587830 66668 587832
rect 66345 587827 66411 587830
rect 66662 587828 66668 587830
rect 66732 587828 66738 587892
rect 67633 587890 67699 587893
rect 68318 587890 68324 587892
rect 67633 587888 68324 587890
rect 67633 587832 67638 587888
rect 67694 587832 68324 587888
rect 67633 587830 68324 587832
rect 67633 587827 67699 587830
rect 68318 587828 68324 587830
rect 68388 587828 68394 587892
rect 69013 587890 69079 587893
rect 69606 587890 69612 587892
rect 69013 587888 69612 587890
rect 69013 587832 69018 587888
rect 69074 587832 69612 587888
rect 69013 587830 69612 587832
rect 69013 587827 69079 587830
rect 69606 587828 69612 587830
rect 69676 587828 69682 587892
rect 70393 587890 70459 587893
rect 71773 587892 71839 587893
rect 70526 587890 70532 587892
rect 70393 587888 70532 587890
rect 70393 587832 70398 587888
rect 70454 587832 70532 587888
rect 70393 587830 70532 587832
rect 70393 587827 70459 587830
rect 70526 587828 70532 587830
rect 70596 587828 70602 587892
rect 71773 587888 71820 587892
rect 71884 587890 71890 587892
rect 72417 587890 72483 587893
rect 74625 587892 74691 587893
rect 72918 587890 72924 587892
rect 71773 587832 71778 587888
rect 71773 587828 71820 587832
rect 71884 587830 71930 587890
rect 72417 587888 72924 587890
rect 72417 587832 72422 587888
rect 72478 587832 72924 587888
rect 72417 587830 72924 587832
rect 71884 587828 71890 587830
rect 71773 587827 71839 587828
rect 72417 587827 72483 587830
rect 72918 587828 72924 587830
rect 72988 587828 72994 587892
rect 74574 587890 74580 587892
rect 74534 587830 74580 587890
rect 74644 587888 74691 587892
rect 74686 587832 74691 587888
rect 74574 587828 74580 587830
rect 74644 587828 74691 587832
rect 74625 587827 74691 587828
rect 77293 587890 77359 587893
rect 77702 587890 77708 587892
rect 77293 587888 77708 587890
rect 77293 587832 77298 587888
rect 77354 587832 77708 587888
rect 77293 587830 77708 587832
rect 77293 587827 77359 587830
rect 77702 587828 77708 587830
rect 77772 587828 77778 587892
rect 78673 587890 78739 587893
rect 78806 587890 78812 587892
rect 78673 587888 78812 587890
rect 78673 587832 78678 587888
rect 78734 587832 78812 587888
rect 78673 587830 78812 587832
rect 78673 587827 78739 587830
rect 78806 587828 78812 587830
rect 78876 587828 78882 587892
rect 79542 587828 79548 587892
rect 79612 587890 79618 587892
rect 79777 587890 79843 587893
rect 79612 587888 79843 587890
rect 79612 587832 79782 587888
rect 79838 587832 79843 587888
rect 79612 587830 79843 587832
rect 79612 587828 79618 587830
rect 79777 587827 79843 587830
rect 81157 587892 81223 587893
rect 81157 587888 81204 587892
rect 81268 587890 81274 587892
rect 81801 587890 81867 587893
rect 82302 587890 82308 587892
rect 81157 587832 81162 587888
rect 81157 587828 81204 587832
rect 81268 587830 81314 587890
rect 81801 587888 82308 587890
rect 81801 587832 81806 587888
rect 81862 587832 82308 587888
rect 81801 587830 82308 587832
rect 81268 587828 81274 587830
rect 81157 587827 81223 587828
rect 81801 587827 81867 587830
rect 82302 587828 82308 587830
rect 82372 587828 82378 587892
rect 82905 587890 82971 587893
rect 87137 587892 87203 587893
rect 83590 587890 83596 587892
rect 82905 587888 83596 587890
rect 82905 587832 82910 587888
rect 82966 587832 83596 587888
rect 82905 587830 83596 587832
rect 82905 587827 82971 587830
rect 83590 587828 83596 587830
rect 83660 587828 83666 587892
rect 87086 587890 87092 587892
rect 87046 587830 87092 587890
rect 87156 587888 87203 587892
rect 87198 587832 87203 587888
rect 87086 587828 87092 587830
rect 87156 587828 87203 587832
rect 87137 587827 87203 587828
rect 88333 587890 88399 587893
rect 89478 587890 89484 587892
rect 88333 587888 89484 587890
rect 88333 587832 88338 587888
rect 88394 587832 89484 587888
rect 88333 587830 89484 587832
rect 88333 587827 88399 587830
rect 89478 587828 89484 587830
rect 89548 587828 89554 587892
rect 91093 587890 91159 587893
rect 91686 587890 91692 587892
rect 91093 587888 91692 587890
rect 91093 587832 91098 587888
rect 91154 587832 91692 587888
rect 91093 587830 91692 587832
rect 91093 587827 91159 587830
rect 91686 587828 91692 587830
rect 91756 587828 91762 587892
rect 92974 587828 92980 587892
rect 93044 587890 93050 587892
rect 93117 587890 93183 587893
rect 93044 587888 93183 587890
rect 93044 587832 93122 587888
rect 93178 587832 93183 587888
rect 93044 587830 93183 587832
rect 93044 587828 93050 587830
rect 93117 587827 93183 587830
rect 93853 587890 93919 587893
rect 94078 587890 94084 587892
rect 93853 587888 94084 587890
rect 93853 587832 93858 587888
rect 93914 587832 94084 587888
rect 93853 587830 94084 587832
rect 93853 587827 93919 587830
rect 94078 587828 94084 587830
rect 94148 587828 94154 587892
rect 94446 587828 94452 587892
rect 94516 587890 94522 587892
rect 95141 587890 95207 587893
rect 99465 587892 99531 587893
rect 99414 587890 99420 587892
rect 94516 587888 95207 587890
rect 94516 587832 95146 587888
rect 95202 587832 95207 587888
rect 94516 587830 95207 587832
rect 99374 587830 99420 587890
rect 99484 587888 99531 587892
rect 99526 587832 99531 587888
rect 94516 587828 94522 587830
rect 95141 587827 95207 587830
rect 99414 587828 99420 587830
rect 99484 587828 99531 587832
rect 99465 587827 99531 587828
rect 101949 587892 102015 587893
rect 106917 587892 106983 587893
rect 101949 587888 101996 587892
rect 102060 587890 102066 587892
rect 101949 587832 101954 587888
rect 101949 587828 101996 587832
rect 102060 587830 102106 587890
rect 106917 587888 106964 587892
rect 107028 587890 107034 587892
rect 109033 587890 109099 587893
rect 109350 587890 109356 587892
rect 106917 587832 106922 587888
rect 102060 587828 102066 587830
rect 106917 587828 106964 587832
rect 107028 587830 107074 587890
rect 109033 587888 109356 587890
rect 109033 587832 109038 587888
rect 109094 587832 109356 587888
rect 109033 587830 109356 587832
rect 107028 587828 107034 587830
rect 101949 587827 102015 587828
rect 106917 587827 106983 587828
rect 109033 587827 109099 587830
rect 109350 587828 109356 587830
rect 109420 587828 109426 587892
rect 111793 587890 111859 587893
rect 111926 587890 111932 587892
rect 111793 587888 111932 587890
rect 111793 587832 111798 587888
rect 111854 587832 111932 587888
rect 111793 587830 111932 587832
rect 111793 587827 111859 587830
rect 111926 587828 111932 587830
rect 111996 587828 112002 587892
rect 114502 587828 114508 587892
rect 114572 587890 114578 587892
rect 115197 587890 115263 587893
rect 114572 587888 115263 587890
rect 114572 587832 115202 587888
rect 115258 587832 115263 587888
rect 114572 587830 115263 587832
rect 114572 587828 114578 587830
rect 115197 587827 115263 587830
rect 118693 587890 118759 587893
rect 124397 587892 124463 587893
rect 119470 587890 119476 587892
rect 118693 587888 119476 587890
rect 118693 587832 118698 587888
rect 118754 587832 119476 587888
rect 118693 587830 119476 587832
rect 118693 587827 118759 587830
rect 119470 587828 119476 587830
rect 119540 587828 119546 587892
rect 124397 587888 124444 587892
rect 124508 587890 124514 587892
rect 128353 587890 128419 587893
rect 131757 587892 131823 587893
rect 129406 587890 129412 587892
rect 124397 587832 124402 587888
rect 124397 587828 124444 587832
rect 124508 587830 124554 587890
rect 128353 587888 129412 587890
rect 128353 587832 128358 587888
rect 128414 587832 129412 587888
rect 128353 587830 129412 587832
rect 124508 587828 124514 587830
rect 124397 587827 124463 587828
rect 128353 587827 128419 587830
rect 129406 587828 129412 587830
rect 129476 587828 129482 587892
rect 131757 587888 131804 587892
rect 131868 587890 131874 587892
rect 133965 587890 134031 587893
rect 134374 587890 134380 587892
rect 131757 587832 131762 587888
rect 131757 587828 131804 587832
rect 131868 587830 131914 587890
rect 133965 587888 134380 587890
rect 133965 587832 133970 587888
rect 134026 587832 134380 587888
rect 133965 587830 134380 587832
rect 131868 587828 131874 587830
rect 131757 587827 131823 587828
rect 133965 587827 134031 587830
rect 134374 587828 134380 587830
rect 134444 587828 134450 587892
rect 136633 587890 136699 587893
rect 139393 587892 139459 587893
rect 141969 587892 142035 587893
rect 136950 587890 136956 587892
rect 136633 587888 136956 587890
rect 136633 587832 136638 587888
rect 136694 587832 136956 587888
rect 136633 587830 136956 587832
rect 136633 587827 136699 587830
rect 136950 587828 136956 587830
rect 137020 587828 137026 587892
rect 139342 587890 139348 587892
rect 139302 587830 139348 587890
rect 139412 587888 139459 587892
rect 141918 587890 141924 587892
rect 139454 587832 139459 587888
rect 139342 587828 139348 587830
rect 139412 587828 139459 587832
rect 141878 587830 141924 587890
rect 141988 587888 142035 587892
rect 142030 587832 142035 587888
rect 141918 587828 141924 587830
rect 141988 587828 142035 587832
rect 139393 587827 139459 587828
rect 141969 587827 142035 587828
rect 159081 587890 159147 587893
rect 159398 587890 159404 587892
rect 159081 587888 159404 587890
rect 159081 587832 159086 587888
rect 159142 587832 159404 587888
rect 159081 587830 159404 587832
rect 159081 587827 159147 587830
rect 159398 587828 159404 587830
rect 159468 587828 159474 587892
rect 224953 587890 225019 587893
rect 226006 587890 226012 587892
rect 224953 587888 226012 587890
rect 224953 587832 224958 587888
rect 225014 587832 226012 587888
rect 224953 587830 226012 587832
rect 224953 587827 225019 587830
rect 226006 587828 226012 587830
rect 226076 587828 226082 587892
rect 227805 587890 227871 587893
rect 228214 587890 228220 587892
rect 227805 587888 228220 587890
rect 227805 587832 227810 587888
rect 227866 587832 228220 587888
rect 227805 587830 228220 587832
rect 227805 587827 227871 587830
rect 228214 587828 228220 587830
rect 228284 587828 228290 587892
rect 230606 587828 230612 587892
rect 230676 587890 230682 587892
rect 231669 587890 231735 587893
rect 230676 587888 231735 587890
rect 230676 587832 231674 587888
rect 231730 587832 231735 587888
rect 230676 587830 231735 587832
rect 230676 587828 230682 587830
rect 231669 587827 231735 587830
rect 234286 587828 234292 587892
rect 234356 587890 234362 587892
rect 234521 587890 234587 587893
rect 234356 587888 234587 587890
rect 234356 587832 234526 587888
rect 234582 587832 234587 587888
rect 234356 587830 234587 587832
rect 234356 587828 234362 587830
rect 234521 587827 234587 587830
rect 235993 587890 236059 587893
rect 236494 587890 236500 587892
rect 235993 587888 236500 587890
rect 235993 587832 235998 587888
rect 236054 587832 236500 587888
rect 235993 587830 236500 587832
rect 235993 587827 236059 587830
rect 236494 587828 236500 587830
rect 236564 587828 236570 587892
rect 237373 587890 237439 587893
rect 237598 587890 237604 587892
rect 237373 587888 237604 587890
rect 237373 587832 237378 587888
rect 237434 587832 237604 587888
rect 237373 587830 237604 587832
rect 237373 587827 237439 587830
rect 237598 587828 237604 587830
rect 237668 587828 237674 587892
rect 238334 587828 238340 587892
rect 238404 587890 238410 587892
rect 238661 587890 238727 587893
rect 238404 587888 238727 587890
rect 238404 587832 238666 587888
rect 238722 587832 238727 587888
rect 238404 587830 238727 587832
rect 238404 587828 238410 587830
rect 238661 587827 238727 587830
rect 238845 587890 238911 587893
rect 239990 587890 239996 587892
rect 238845 587888 239996 587890
rect 238845 587832 238850 587888
rect 238906 587832 239996 587888
rect 238845 587830 239996 587832
rect 238845 587827 238911 587830
rect 239990 587828 239996 587830
rect 240060 587828 240066 587892
rect 240501 587890 240567 587893
rect 242433 587892 242499 587893
rect 241278 587890 241284 587892
rect 240501 587888 241284 587890
rect 240501 587832 240506 587888
rect 240562 587832 241284 587888
rect 240501 587830 241284 587832
rect 240501 587827 240567 587830
rect 241278 587828 241284 587830
rect 241348 587828 241354 587892
rect 242382 587890 242388 587892
rect 242342 587830 242388 587890
rect 242452 587888 242499 587892
rect 242494 587832 242499 587888
rect 242382 587828 242388 587830
rect 242452 587828 242499 587832
rect 243302 587828 243308 587892
rect 243372 587890 243378 587892
rect 243537 587890 243603 587893
rect 243372 587888 243603 587890
rect 243372 587832 243542 587888
rect 243598 587832 243603 587888
rect 243372 587830 243603 587832
rect 243372 587828 243378 587830
rect 242433 587827 242499 587828
rect 243537 587827 243603 587830
rect 244590 587828 244596 587892
rect 244660 587890 244666 587892
rect 245561 587890 245627 587893
rect 244660 587888 245627 587890
rect 244660 587832 245566 587888
rect 245622 587832 245627 587888
rect 244660 587830 245627 587832
rect 244660 587828 244666 587830
rect 245561 587827 245627 587830
rect 245837 587892 245903 587893
rect 247033 587892 247099 587893
rect 248137 587892 248203 587893
rect 245837 587888 245884 587892
rect 245948 587890 245954 587892
rect 246982 587890 246988 587892
rect 245837 587832 245842 587888
rect 245837 587828 245884 587832
rect 245948 587830 245994 587890
rect 246942 587830 246988 587890
rect 247052 587888 247099 587892
rect 248086 587890 248092 587892
rect 247094 587832 247099 587888
rect 245948 587828 245954 587830
rect 246982 587828 246988 587830
rect 247052 587828 247099 587832
rect 248046 587830 248092 587890
rect 248156 587888 248203 587892
rect 248198 587832 248203 587888
rect 248086 587828 248092 587830
rect 248156 587828 248203 587832
rect 245837 587827 245903 587828
rect 247033 587827 247099 587828
rect 248137 587827 248203 587828
rect 248413 587892 248479 587893
rect 248413 587888 248460 587892
rect 248524 587890 248530 587892
rect 248413 587832 248418 587888
rect 248413 587828 248460 587832
rect 248524 587830 248570 587890
rect 248524 587828 248530 587830
rect 249558 587828 249564 587892
rect 249628 587890 249634 587892
rect 249701 587890 249767 587893
rect 249628 587888 249767 587890
rect 249628 587832 249706 587888
rect 249762 587832 249767 587888
rect 249628 587830 249767 587832
rect 249628 587828 249634 587830
rect 248413 587827 248479 587828
rect 249701 587827 249767 587830
rect 252645 587890 252711 587893
rect 253933 587892 253999 587893
rect 252870 587890 252876 587892
rect 252645 587888 252876 587890
rect 252645 587832 252650 587888
rect 252706 587832 252876 587888
rect 252645 587830 252876 587832
rect 252645 587827 252711 587830
rect 252870 587828 252876 587830
rect 252940 587828 252946 587892
rect 253933 587888 253980 587892
rect 254044 587890 254050 587892
rect 255313 587890 255379 587893
rect 255998 587890 256004 587892
rect 253933 587832 253938 587888
rect 253933 587828 253980 587832
rect 254044 587830 254090 587890
rect 255313 587888 256004 587890
rect 255313 587832 255318 587888
rect 255374 587832 256004 587888
rect 255313 587830 256004 587832
rect 254044 587828 254050 587830
rect 253933 587827 253999 587828
rect 255313 587827 255379 587830
rect 255998 587828 256004 587830
rect 256068 587828 256074 587892
rect 256366 587828 256372 587892
rect 256436 587890 256442 587892
rect 256601 587890 256667 587893
rect 256436 587888 256667 587890
rect 256436 587832 256606 587888
rect 256662 587832 256667 587888
rect 256436 587830 256667 587832
rect 256436 587828 256442 587830
rect 256601 587827 256667 587830
rect 257654 587828 257660 587892
rect 257724 587890 257730 587892
rect 257981 587890 258047 587893
rect 257724 587888 258047 587890
rect 257724 587832 257986 587888
rect 258042 587832 258047 587888
rect 257724 587830 258047 587832
rect 257724 587828 257730 587830
rect 257981 587827 258047 587830
rect 259862 587828 259868 587892
rect 259932 587890 259938 587892
rect 260649 587890 260715 587893
rect 261017 587892 261083 587893
rect 260966 587890 260972 587892
rect 259932 587888 260715 587890
rect 259932 587832 260654 587888
rect 260710 587832 260715 587888
rect 259932 587830 260715 587832
rect 260926 587830 260972 587890
rect 261036 587888 261083 587892
rect 261078 587832 261083 587888
rect 259932 587828 259938 587830
rect 260649 587827 260715 587830
rect 260966 587828 260972 587830
rect 261036 587828 261083 587832
rect 261150 587828 261156 587892
rect 261220 587890 261226 587892
rect 262029 587890 262095 587893
rect 261220 587888 262095 587890
rect 261220 587832 262034 587888
rect 262090 587832 262095 587888
rect 261220 587830 262095 587832
rect 261220 587828 261226 587830
rect 261017 587827 261083 587828
rect 262029 587827 262095 587830
rect 262213 587892 262279 587893
rect 262213 587888 262260 587892
rect 262324 587890 262330 587892
rect 262213 587832 262218 587888
rect 262213 587828 262260 587832
rect 262324 587830 262370 587890
rect 262324 587828 262330 587830
rect 263542 587828 263548 587892
rect 263612 587890 263618 587892
rect 264881 587890 264947 587893
rect 263612 587888 264947 587890
rect 263612 587832 264886 587888
rect 264942 587832 264947 587888
rect 263612 587830 264947 587832
rect 263612 587828 263618 587830
rect 262213 587827 262279 587828
rect 264881 587827 264947 587830
rect 265750 587828 265756 587892
rect 265820 587890 265826 587892
rect 266261 587890 266327 587893
rect 265820 587888 266327 587890
rect 265820 587832 266266 587888
rect 266322 587832 266327 587888
rect 265820 587830 266327 587832
rect 265820 587828 265826 587830
rect 266261 587827 266327 587830
rect 268510 587828 268516 587892
rect 268580 587890 268586 587892
rect 268929 587890 268995 587893
rect 268580 587888 268995 587890
rect 268580 587832 268934 587888
rect 268990 587832 268995 587888
rect 268580 587830 268995 587832
rect 268580 587828 268586 587830
rect 268929 587827 268995 587830
rect 269246 587828 269252 587892
rect 269316 587890 269322 587892
rect 269757 587890 269823 587893
rect 269316 587888 269823 587890
rect 269316 587832 269762 587888
rect 269818 587832 269823 587888
rect 269316 587830 269823 587832
rect 269316 587828 269322 587830
rect 269757 587827 269823 587830
rect 270493 587890 270559 587893
rect 273529 587892 273595 587893
rect 270902 587890 270908 587892
rect 270493 587888 270908 587890
rect 270493 587832 270498 587888
rect 270554 587832 270908 587888
rect 270493 587830 270908 587832
rect 270493 587827 270559 587830
rect 270902 587828 270908 587830
rect 270972 587828 270978 587892
rect 273478 587890 273484 587892
rect 273438 587830 273484 587890
rect 273548 587888 273595 587892
rect 273590 587832 273595 587888
rect 273478 587828 273484 587830
rect 273548 587828 273595 587832
rect 273529 587827 273595 587828
rect 274633 587890 274699 587893
rect 281073 587892 281139 587893
rect 275870 587890 275876 587892
rect 274633 587888 275876 587890
rect 274633 587832 274638 587888
rect 274694 587832 275876 587888
rect 274633 587830 275876 587832
rect 274633 587827 274699 587830
rect 275870 587828 275876 587830
rect 275940 587828 275946 587892
rect 281022 587890 281028 587892
rect 280982 587830 281028 587890
rect 281092 587888 281139 587892
rect 281134 587832 281139 587888
rect 281022 587828 281028 587830
rect 281092 587828 281139 587832
rect 281073 587827 281139 587828
rect 282913 587890 282979 587893
rect 283414 587890 283420 587892
rect 282913 587888 283420 587890
rect 282913 587832 282918 587888
rect 282974 587832 283420 587888
rect 282913 587830 283420 587832
rect 282913 587827 282979 587830
rect 283414 587828 283420 587830
rect 283484 587828 283490 587892
rect 285990 587828 285996 587892
rect 286060 587890 286066 587892
rect 286317 587890 286383 587893
rect 288433 587892 288499 587893
rect 291009 587892 291075 587893
rect 288382 587890 288388 587892
rect 286060 587888 286383 587890
rect 286060 587832 286322 587888
rect 286378 587832 286383 587888
rect 286060 587830 286383 587832
rect 288342 587830 288388 587890
rect 288452 587888 288499 587892
rect 290958 587890 290964 587892
rect 288494 587832 288499 587888
rect 286060 587828 286066 587830
rect 286317 587827 286383 587830
rect 288382 587828 288388 587830
rect 288452 587828 288499 587832
rect 290918 587830 290964 587890
rect 291028 587888 291075 587892
rect 291070 587832 291075 587888
rect 290958 587828 290964 587830
rect 291028 587828 291075 587832
rect 288433 587827 288499 587828
rect 291009 587827 291075 587828
rect 298093 587890 298159 587893
rect 300853 587892 300919 587893
rect 298502 587890 298508 587892
rect 298093 587888 298508 587890
rect 298093 587832 298098 587888
rect 298154 587832 298508 587888
rect 298093 587830 298508 587832
rect 298093 587827 298159 587830
rect 298502 587828 298508 587830
rect 298572 587828 298578 587892
rect 300853 587888 300900 587892
rect 300964 587890 300970 587892
rect 302233 587890 302299 587893
rect 303470 587890 303476 587892
rect 300853 587832 300858 587888
rect 300853 587828 300900 587832
rect 300964 587830 301010 587890
rect 302233 587888 303476 587890
rect 302233 587832 302238 587888
rect 302294 587832 303476 587888
rect 302233 587830 303476 587832
rect 300964 587828 300970 587830
rect 300853 587827 300919 587828
rect 302233 587827 302299 587830
rect 303470 587828 303476 587830
rect 303540 587828 303546 587892
rect 305085 587890 305151 587893
rect 308489 587892 308555 587893
rect 305862 587890 305868 587892
rect 305085 587888 305868 587890
rect 305085 587832 305090 587888
rect 305146 587832 305868 587888
rect 305085 587830 305868 587832
rect 305085 587827 305151 587830
rect 305862 587828 305868 587830
rect 305932 587828 305938 587892
rect 308438 587890 308444 587892
rect 308398 587830 308444 587890
rect 308508 587888 308555 587892
rect 308550 587832 308555 587888
rect 308438 587828 308444 587830
rect 308508 587828 308555 587832
rect 308489 587827 308555 587828
rect 310513 587890 310579 587893
rect 310830 587890 310836 587892
rect 310513 587888 310836 587890
rect 310513 587832 310518 587888
rect 310574 587832 310836 587888
rect 310513 587830 310836 587832
rect 310513 587827 310579 587830
rect 310830 587828 310836 587830
rect 310900 587828 310906 587892
rect 313273 587890 313339 587893
rect 316033 587892 316099 587893
rect 313406 587890 313412 587892
rect 313273 587888 313412 587890
rect 313273 587832 313278 587888
rect 313334 587832 313412 587888
rect 313273 587830 313412 587832
rect 313273 587827 313339 587830
rect 313406 587828 313412 587830
rect 313476 587828 313482 587892
rect 315982 587828 315988 587892
rect 316052 587890 316099 587892
rect 316052 587888 316144 587890
rect 316094 587832 316144 587888
rect 316052 587830 316144 587832
rect 316052 587828 316099 587830
rect 333462 587828 333468 587892
rect 333532 587890 333538 587892
rect 333881 587890 333947 587893
rect 333532 587888 333947 587890
rect 333532 587832 333886 587888
rect 333942 587832 333947 587888
rect 333532 587830 333947 587832
rect 333532 587828 333538 587830
rect 316033 587827 316099 587828
rect 333881 587827 333947 587830
rect 55622 587692 55628 587756
rect 55692 587754 55698 587756
rect 56501 587754 56567 587757
rect 55692 587752 56567 587754
rect 55692 587696 56506 587752
rect 56562 587696 56567 587752
rect 55692 587694 56567 587696
rect 55692 587692 55698 587694
rect 56501 587691 56567 587694
rect 61510 587692 61516 587756
rect 61580 587754 61586 587756
rect 62021 587754 62087 587757
rect 61580 587752 62087 587754
rect 61580 587696 62026 587752
rect 62082 587696 62087 587752
rect 61580 587694 62087 587696
rect 61580 587692 61586 587694
rect 62021 587691 62087 587694
rect 63585 587754 63651 587757
rect 64638 587754 64644 587756
rect 63585 587752 64644 587754
rect 63585 587696 63590 587752
rect 63646 587696 64644 587752
rect 63585 587694 64644 587696
rect 63585 587691 63651 587694
rect 64638 587692 64644 587694
rect 64708 587692 64714 587756
rect 69422 587692 69428 587756
rect 69492 587754 69498 587756
rect 70301 587754 70367 587757
rect 69492 587752 70367 587754
rect 69492 587696 70306 587752
rect 70362 587696 70367 587752
rect 69492 587694 70367 587696
rect 69492 587692 69498 587694
rect 70301 587691 70367 587694
rect 72182 587692 72188 587756
rect 72252 587754 72258 587756
rect 73061 587754 73127 587757
rect 72252 587752 73127 587754
rect 72252 587696 73066 587752
rect 73122 587696 73127 587752
rect 72252 587694 73127 587696
rect 72252 587692 72258 587694
rect 73061 587691 73127 587694
rect 74533 587754 74599 587757
rect 77201 587756 77267 587757
rect 75494 587754 75500 587756
rect 74533 587752 75500 587754
rect 74533 587696 74538 587752
rect 74594 587696 75500 587752
rect 74533 587694 75500 587696
rect 74533 587691 74599 587694
rect 75494 587692 75500 587694
rect 75564 587692 75570 587756
rect 77150 587754 77156 587756
rect 77110 587694 77156 587754
rect 77220 587752 77267 587756
rect 77262 587696 77267 587752
rect 77150 587692 77156 587694
rect 77220 587692 77267 587696
rect 77201 587691 77267 587692
rect 78765 587754 78831 587757
rect 81893 587756 81959 587757
rect 79910 587754 79916 587756
rect 78765 587752 79916 587754
rect 78765 587696 78770 587752
rect 78826 587696 79916 587752
rect 78765 587694 79916 587696
rect 78765 587691 78831 587694
rect 79910 587692 79916 587694
rect 79980 587692 79986 587756
rect 81893 587752 81940 587756
rect 82004 587754 82010 587756
rect 86953 587754 87019 587757
rect 95233 587756 95299 587757
rect 88190 587754 88196 587756
rect 81893 587696 81898 587752
rect 81893 587692 81940 587696
rect 82004 587694 82050 587754
rect 86953 587752 88196 587754
rect 86953 587696 86958 587752
rect 87014 587696 88196 587752
rect 86953 587694 88196 587696
rect 82004 587692 82010 587694
rect 81893 587691 81959 587692
rect 86953 587691 87019 587694
rect 88190 587692 88196 587694
rect 88260 587692 88266 587756
rect 95182 587754 95188 587756
rect 95142 587694 95188 587754
rect 95252 587752 95299 587756
rect 95294 587696 95299 587752
rect 95182 587692 95188 587694
rect 95252 587692 95299 587696
rect 127014 587692 127020 587756
rect 127084 587754 127090 587756
rect 128261 587754 128327 587757
rect 127084 587752 128327 587754
rect 127084 587696 128266 587752
rect 128322 587696 128327 587752
rect 127084 587694 128327 587696
rect 127084 587692 127090 587694
rect 95233 587691 95299 587692
rect 128261 587691 128327 587694
rect 234613 587754 234679 587757
rect 240777 587756 240843 587757
rect 235390 587754 235396 587756
rect 234613 587752 235396 587754
rect 234613 587696 234618 587752
rect 234674 587696 235396 587752
rect 234613 587694 235396 587696
rect 234613 587691 234679 587694
rect 235390 587692 235396 587694
rect 235460 587692 235466 587756
rect 240726 587754 240732 587756
rect 240686 587694 240732 587754
rect 240796 587752 240843 587756
rect 240838 587696 240843 587752
rect 240726 587692 240732 587694
rect 240796 587692 240843 587696
rect 246062 587692 246068 587756
rect 246132 587754 246138 587756
rect 246941 587754 247007 587757
rect 246132 587752 247007 587754
rect 246132 587696 246946 587752
rect 247002 587696 247007 587752
rect 246132 587694 247007 587696
rect 246132 587692 246138 587694
rect 240777 587691 240843 587692
rect 246941 587691 247007 587694
rect 249793 587754 249859 587757
rect 251030 587754 251036 587756
rect 249793 587752 251036 587754
rect 249793 587696 249798 587752
rect 249854 587696 251036 587752
rect 249793 587694 251036 587696
rect 249793 587691 249859 587694
rect 251030 587692 251036 587694
rect 251100 587692 251106 587756
rect 252553 587754 252619 587757
rect 264421 587756 264487 587757
rect 253422 587754 253428 587756
rect 252553 587752 253428 587754
rect 252553 587696 252558 587752
rect 252614 587696 253428 587752
rect 252553 587694 253428 587696
rect 252553 587691 252619 587694
rect 253422 587692 253428 587694
rect 253492 587692 253498 587756
rect 264421 587752 264468 587756
rect 264532 587754 264538 587756
rect 264973 587754 265039 587757
rect 265934 587754 265940 587756
rect 264421 587696 264426 587752
rect 264421 587692 264468 587696
rect 264532 587694 264578 587754
rect 264973 587752 265940 587754
rect 264973 587696 264978 587752
rect 265034 587696 265940 587752
rect 264973 587694 265940 587696
rect 264532 587692 264538 587694
rect 264421 587691 264487 587692
rect 264973 587691 265039 587694
rect 265934 587692 265940 587694
rect 266004 587692 266010 587756
rect 74022 587556 74028 587620
rect 74092 587618 74098 587620
rect 74441 587618 74507 587621
rect 74092 587616 74507 587618
rect 74092 587560 74446 587616
rect 74502 587560 74507 587616
rect 74092 587558 74507 587560
rect 74092 587556 74098 587558
rect 74441 587555 74507 587558
rect 25773 587482 25839 587485
rect 227110 587482 227116 587484
rect 25773 587480 227116 587482
rect 25773 587424 25778 587480
rect 25834 587424 227116 587480
rect 25773 587422 227116 587424
rect 25773 587419 25839 587422
rect 227110 587420 227116 587422
rect 227180 587420 227186 587484
rect 25865 587346 25931 587349
rect 229502 587346 229508 587348
rect 25865 587344 229508 587346
rect 25865 587288 25870 587344
rect 25926 587288 229508 587344
rect 25865 587286 229508 587288
rect 25865 587283 25931 587286
rect 229502 587284 229508 587286
rect 229572 587284 229578 587348
rect 250662 587284 250668 587348
rect 250732 587346 250738 587348
rect 348366 587346 348372 587348
rect 250732 587286 348372 587346
rect 250732 587284 250738 587286
rect 348366 587284 348372 587286
rect 348436 587284 348442 587348
rect 35617 587210 35683 587213
rect 255262 587210 255268 587212
rect 35617 587208 255268 587210
rect 35617 587152 35622 587208
rect 35678 587152 255268 587208
rect 35617 587150 255268 587152
rect 35617 587147 35683 587150
rect 255262 587148 255268 587150
rect 255332 587148 255338 587212
rect 407297 586938 407363 586941
rect 553301 586938 553367 586941
rect 407297 586936 410044 586938
rect 407297 586880 407302 586936
rect 407358 586880 410044 586936
rect 407297 586878 410044 586880
rect 549884 586936 553367 586938
rect 549884 586880 553306 586936
rect 553362 586880 553367 586936
rect 549884 586878 553367 586880
rect 407297 586875 407363 586878
rect 553301 586875 553367 586878
rect 238518 586740 238524 586804
rect 238588 586802 238594 586804
rect 238753 586802 238819 586805
rect 238588 586800 238819 586802
rect 238588 586744 238758 586800
rect 238814 586744 238819 586800
rect 238588 586742 238819 586744
rect 238588 586740 238594 586742
rect 238753 586739 238819 586742
rect 257838 586740 257844 586804
rect 257908 586802 257914 586804
rect 258165 586802 258231 586805
rect 257908 586800 258231 586802
rect 257908 586744 258170 586800
rect 258226 586744 258231 586800
rect 257908 586742 258231 586744
rect 257908 586740 257914 586742
rect 258165 586739 258231 586742
rect 51942 586666 51948 586668
rect 51030 586606 51948 586666
rect 48446 586332 48452 586396
rect 48516 586394 48522 586396
rect 51030 586394 51090 586606
rect 51942 586604 51948 586606
rect 52012 586604 52018 586668
rect 67214 586666 67220 586668
rect 66486 586606 67220 586666
rect 48516 586334 51090 586394
rect 66486 586394 66546 586606
rect 67214 586604 67220 586606
rect 67284 586604 67290 586668
rect 76598 586666 76604 586668
rect 75870 586606 76604 586666
rect 67541 586394 67607 586397
rect 66486 586392 67607 586394
rect 66486 586336 67546 586392
rect 67602 586336 67607 586392
rect 66486 586334 67607 586336
rect 75870 586394 75930 586606
rect 76598 586604 76604 586606
rect 76668 586604 76674 586668
rect 86902 586604 86908 586668
rect 86972 586666 86978 586668
rect 89294 586666 89300 586668
rect 86972 586606 87706 586666
rect 86972 586604 86978 586606
rect 84142 586468 84148 586532
rect 84212 586468 84218 586532
rect 85614 586468 85620 586532
rect 85684 586468 85690 586532
rect 77109 586394 77175 586397
rect 75870 586392 77175 586394
rect 75870 586336 77114 586392
rect 77170 586336 77175 586392
rect 75870 586334 77175 586336
rect 84150 586394 84210 586468
rect 85481 586394 85547 586397
rect 84150 586392 85547 586394
rect 84150 586336 85486 586392
rect 85542 586336 85547 586392
rect 84150 586334 85547 586336
rect 85622 586394 85682 586468
rect 86861 586394 86927 586397
rect 85622 586392 86927 586394
rect 85622 586336 86866 586392
rect 86922 586336 86927 586392
rect 85622 586334 86927 586336
rect 48516 586332 48522 586334
rect 67541 586331 67607 586334
rect 77109 586331 77175 586334
rect 85481 586331 85547 586334
rect 86861 586331 86927 586334
rect 87045 586394 87111 586397
rect 87646 586394 87706 586606
rect 87045 586392 87706 586394
rect 87045 586336 87050 586392
rect 87106 586336 87706 586392
rect 87045 586334 87706 586336
rect 88566 586606 89300 586666
rect 88566 586394 88626 586606
rect 89294 586604 89300 586606
rect 89364 586604 89370 586668
rect 90398 586666 90404 586668
rect 89854 586606 90404 586666
rect 89621 586394 89687 586397
rect 88566 586392 89687 586394
rect 88566 586336 89626 586392
rect 89682 586336 89687 586392
rect 88566 586334 89687 586336
rect 89854 586394 89914 586606
rect 90398 586604 90404 586606
rect 90468 586604 90474 586668
rect 92054 586666 92060 586668
rect 91142 586606 92060 586666
rect 91001 586394 91067 586397
rect 89854 586392 91067 586394
rect 89854 586336 91006 586392
rect 91062 586336 91067 586392
rect 89854 586334 91067 586336
rect 91142 586394 91202 586606
rect 92054 586604 92060 586606
rect 92124 586604 92130 586668
rect 96838 586666 96844 586668
rect 96662 586606 96844 586666
rect 92381 586394 92447 586397
rect 91142 586392 92447 586394
rect 91142 586336 92386 586392
rect 92442 586336 92447 586392
rect 91142 586334 92447 586336
rect 96662 586394 96722 586606
rect 96838 586604 96844 586606
rect 96908 586604 96914 586668
rect 116894 586666 116900 586668
rect 115982 586606 116900 586666
rect 103462 586468 103468 586532
rect 103532 586468 103538 586532
rect 97901 586394 97967 586397
rect 96662 586392 97967 586394
rect 96662 586336 97906 586392
rect 97962 586336 97967 586392
rect 96662 586334 97967 586336
rect 103470 586394 103530 586468
rect 104801 586394 104867 586397
rect 103470 586392 104867 586394
rect 103470 586336 104806 586392
rect 104862 586336 104867 586392
rect 103470 586334 104867 586336
rect 115982 586394 116042 586606
rect 116894 586604 116900 586606
rect 116964 586604 116970 586668
rect 121862 586666 121868 586668
rect 121502 586606 121868 586666
rect 117221 586394 117287 586397
rect 115982 586392 117287 586394
rect 115982 586336 117226 586392
rect 117282 586336 117287 586392
rect 115982 586334 117287 586336
rect 121502 586394 121562 586606
rect 121862 586604 121868 586606
rect 121932 586604 121938 586668
rect 159214 586666 159220 586668
rect 158670 586606 159220 586666
rect 122741 586394 122807 586397
rect 121502 586392 122807 586394
rect 121502 586336 122746 586392
rect 122802 586336 122807 586392
rect 121502 586334 122807 586336
rect 158670 586394 158730 586606
rect 159214 586604 159220 586606
rect 159284 586604 159290 586668
rect 231710 586666 231716 586668
rect 230798 586606 231716 586666
rect 160001 586394 160067 586397
rect 158670 586392 160067 586394
rect 158670 586336 160006 586392
rect 160062 586336 160067 586392
rect 158670 586334 160067 586336
rect 230798 586394 230858 586606
rect 231710 586604 231716 586606
rect 231780 586604 231786 586668
rect 233182 586666 233188 586668
rect 231902 586606 233188 586666
rect 231761 586394 231827 586397
rect 230798 586392 231827 586394
rect 230798 586336 231766 586392
rect 231822 586336 231827 586392
rect 230798 586334 231827 586336
rect 231902 586394 231962 586606
rect 233182 586604 233188 586606
rect 233252 586604 233258 586668
rect 243670 586666 243676 586668
rect 242942 586606 243676 586666
rect 233141 586394 233207 586397
rect 231902 586392 233207 586394
rect 231902 586336 233146 586392
rect 233202 586336 233207 586392
rect 231902 586334 233207 586336
rect 242942 586394 243002 586606
rect 243670 586604 243676 586606
rect 243740 586604 243746 586668
rect 251766 586666 251772 586668
rect 251222 586606 251772 586666
rect 244181 586394 244247 586397
rect 242942 586392 244247 586394
rect 242942 586336 244186 586392
rect 244242 586336 244247 586392
rect 242942 586334 244247 586336
rect 251222 586394 251282 586606
rect 251766 586604 251772 586606
rect 251836 586604 251842 586668
rect 263358 586666 263364 586668
rect 262446 586606 263364 586666
rect 258574 586468 258580 586532
rect 258644 586468 258650 586532
rect 252461 586394 252527 586397
rect 251222 586392 252527 586394
rect 251222 586336 252466 586392
rect 252522 586336 252527 586392
rect 251222 586334 252527 586336
rect 87045 586331 87111 586334
rect 89621 586331 89687 586334
rect 91001 586331 91067 586334
rect 92381 586331 92447 586334
rect 97901 586331 97967 586334
rect 104801 586331 104867 586334
rect 117221 586331 117287 586334
rect 122741 586331 122807 586334
rect 160001 586331 160067 586334
rect 231761 586331 231827 586334
rect 233141 586331 233207 586334
rect 244181 586331 244247 586334
rect 252461 586331 252527 586334
rect 258073 586394 258139 586397
rect 258582 586394 258642 586468
rect 258073 586392 258642 586394
rect 258073 586336 258078 586392
rect 258134 586336 258642 586392
rect 258073 586334 258642 586336
rect 262446 586394 262506 586606
rect 263358 586604 263364 586606
rect 263428 586604 263434 586668
rect 267038 586666 267044 586668
rect 266310 586606 267044 586666
rect 263501 586394 263567 586397
rect 262446 586392 263567 586394
rect 262446 586336 263506 586392
rect 263562 586336 263567 586392
rect 262446 586334 263567 586336
rect 266310 586394 266370 586606
rect 267038 586604 267044 586606
rect 267108 586604 267114 586668
rect 293534 586666 293540 586668
rect 292622 586606 293540 586666
rect 267958 586468 267964 586532
rect 268028 586468 268034 586532
rect 277342 586468 277348 586532
rect 277412 586530 277418 586532
rect 277485 586530 277551 586533
rect 277412 586528 277551 586530
rect 277412 586472 277490 586528
rect 277546 586472 277551 586528
rect 277412 586470 277551 586472
rect 277412 586468 277418 586470
rect 267641 586394 267707 586397
rect 266310 586392 267707 586394
rect 266310 586336 267646 586392
rect 267702 586336 267707 586392
rect 266310 586334 267707 586336
rect 267966 586394 268026 586468
rect 277485 586467 277551 586470
rect 269021 586394 269087 586397
rect 267966 586392 269087 586394
rect 267966 586336 269026 586392
rect 269082 586336 269087 586392
rect 267966 586334 269087 586336
rect 292622 586394 292682 586606
rect 293534 586604 293540 586606
rect 293604 586604 293610 586668
rect 295926 586666 295932 586668
rect 295382 586606 295932 586666
rect 293861 586394 293927 586397
rect 292622 586392 293927 586394
rect 292622 586336 293866 586392
rect 293922 586336 293927 586392
rect 292622 586334 293927 586336
rect 295382 586394 295442 586606
rect 295926 586604 295932 586606
rect 295996 586604 296002 586668
rect 333094 586666 333100 586668
rect 332550 586606 333100 586666
rect 296621 586394 296687 586397
rect 295382 586392 296687 586394
rect 295382 586336 296626 586392
rect 296682 586336 296687 586392
rect 295382 586334 296687 586336
rect 332550 586394 332610 586606
rect 333094 586604 333100 586606
rect 333164 586604 333170 586668
rect 333789 586394 333855 586397
rect 332550 586392 333855 586394
rect 332550 586336 333794 586392
rect 333850 586336 333855 586392
rect 332550 586334 333855 586336
rect 258073 586331 258139 586334
rect 263501 586331 263567 586334
rect 267641 586331 267707 586334
rect 269021 586331 269087 586334
rect 293861 586331 293927 586334
rect 296621 586331 296687 586334
rect 333789 586331 333855 586334
rect 408401 586258 408467 586261
rect 552565 586258 552631 586261
rect 408401 586256 410044 586258
rect 408401 586200 408406 586256
rect 408462 586200 410044 586256
rect 408401 586198 410044 586200
rect 549884 586256 552631 586258
rect 549884 586200 552570 586256
rect 552626 586200 552631 586256
rect 549884 586198 552631 586200
rect 408401 586195 408467 586198
rect 552565 586195 552631 586198
rect 407665 585578 407731 585581
rect 553209 585578 553275 585581
rect 407665 585576 410044 585578
rect 407665 585520 407670 585576
rect 407726 585520 410044 585576
rect 407665 585518 410044 585520
rect 549884 585576 553275 585578
rect 549884 585520 553214 585576
rect 553270 585520 553275 585576
rect 549884 585518 553275 585520
rect 407665 585515 407731 585518
rect 553209 585515 553275 585518
rect 407297 584898 407363 584901
rect 552933 584898 552999 584901
rect 407297 584896 410044 584898
rect 407297 584840 407302 584896
rect 407358 584840 410044 584896
rect 407297 584838 410044 584840
rect 549884 584896 552999 584898
rect 549884 584840 552938 584896
rect 552994 584840 552999 584896
rect 549884 584838 552999 584840
rect 407297 584835 407363 584838
rect 552933 584835 552999 584838
rect 17861 584354 17927 584357
rect 407798 584354 407804 584356
rect 17861 584352 407804 584354
rect 17861 584296 17866 584352
rect 17922 584296 407804 584352
rect 17861 584294 407804 584296
rect 17861 584291 17927 584294
rect 407798 584292 407804 584294
rect 407868 584292 407874 584356
rect 46974 583068 46980 583132
rect 47044 583130 47050 583132
rect 288433 583130 288499 583133
rect 47044 583128 288499 583130
rect 47044 583072 288438 583128
rect 288494 583072 288499 583128
rect 47044 583070 288499 583072
rect 47044 583068 47050 583070
rect 288433 583067 288499 583070
rect 93117 582994 93183 582997
rect 346342 582994 346348 582996
rect 93117 582992 346348 582994
rect 93117 582936 93122 582992
rect 93178 582936 346348 582992
rect 93117 582934 346348 582936
rect 93117 582931 93183 582934
rect 346342 582932 346348 582934
rect 346412 582932 346418 582996
rect 570086 582178 570092 582180
rect 549884 582118 570092 582178
rect 570086 582116 570092 582118
rect 570156 582116 570162 582180
rect 72417 581634 72483 581637
rect 351126 581634 351132 581636
rect 72417 581632 351132 581634
rect 72417 581576 72422 581632
rect 72478 581576 351132 581632
rect 72417 581574 351132 581576
rect 72417 581571 72483 581574
rect 351126 581572 351132 581574
rect 351196 581572 351202 581636
rect 391238 581436 391244 581500
rect 391308 581498 391314 581500
rect 391308 581438 410044 581498
rect 391308 581436 391314 581438
rect 387006 580756 387012 580820
rect 387076 580818 387082 580820
rect 567326 580818 567332 580820
rect 387076 580758 410044 580818
rect 549884 580758 567332 580818
rect 387076 580756 387082 580758
rect 567326 580756 567332 580758
rect 567396 580756 567402 580820
rect 407297 580138 407363 580141
rect 407297 580136 410044 580138
rect -960 579852 480 580092
rect 407297 580080 407302 580136
rect 407358 580080 410044 580136
rect 407297 580078 410044 580080
rect 407297 580075 407363 580078
rect 563094 579458 563100 579460
rect 549884 579398 563100 579458
rect 563094 579396 563100 579398
rect 563164 579396 563170 579460
rect 56501 578914 56567 578917
rect 349102 578914 349108 578916
rect 56501 578912 349108 578914
rect 56501 578856 56506 578912
rect 56562 578856 349108 578912
rect 56501 578854 349108 578856
rect 56501 578851 56567 578854
rect 349102 578852 349108 578854
rect 349172 578852 349178 578916
rect 371734 578716 371740 578780
rect 371804 578778 371810 578780
rect 371804 578718 410044 578778
rect 371804 578716 371810 578718
rect 408953 578098 409019 578101
rect 553301 578098 553367 578101
rect 408953 578096 410044 578098
rect 408953 578040 408958 578096
rect 409014 578040 410044 578096
rect 408953 578038 410044 578040
rect 549884 578096 553367 578098
rect 549884 578040 553306 578096
rect 553362 578040 553367 578096
rect 549884 578038 553367 578040
rect 408953 578035 409019 578038
rect 553301 578035 553367 578038
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 46790 577492 46796 577556
rect 46860 577554 46866 577556
rect 270493 577554 270559 577557
rect 46860 577552 270559 577554
rect 46860 577496 270498 577552
rect 270554 577496 270559 577552
rect 583520 577540 584960 577630
rect 46860 577494 270559 577496
rect 46860 577492 46866 577494
rect 270493 577491 270559 577494
rect 407297 577418 407363 577421
rect 407297 577416 410044 577418
rect 407297 577360 407302 577416
rect 407358 577360 410044 577416
rect 407297 577358 410044 577360
rect 407297 577355 407363 577358
rect 407297 576738 407363 576741
rect 561990 576738 561996 576740
rect 407297 576736 410044 576738
rect 407297 576680 407302 576736
rect 407358 576680 410044 576736
rect 407297 576678 410044 576680
rect 549884 576678 561996 576738
rect 407297 576675 407363 576678
rect 561990 576676 561996 576678
rect 562060 576676 562066 576740
rect 92381 576058 92447 576061
rect 347814 576058 347820 576060
rect 92381 576056 347820 576058
rect 92381 576000 92386 576056
rect 92442 576000 347820 576056
rect 92381 575998 347820 576000
rect 92381 575995 92447 575998
rect 347814 575996 347820 575998
rect 347884 575996 347890 576060
rect 553301 576058 553367 576061
rect 549884 576056 553367 576058
rect 549884 576000 553306 576056
rect 553362 576000 553367 576056
rect 549884 575998 553367 576000
rect 553301 575995 553367 575998
rect 46606 574636 46612 574700
rect 46676 574698 46682 574700
rect 305085 574698 305151 574701
rect 46676 574696 305151 574698
rect 46676 574640 305090 574696
rect 305146 574640 305151 574696
rect 46676 574638 305151 574640
rect 46676 574636 46682 574638
rect 305085 574635 305151 574638
rect 549884 574570 550466 574630
rect 550406 574562 550466 574570
rect 550406 574502 557550 574562
rect 557490 574154 557550 574502
rect 559046 574154 559052 574156
rect 557490 574094 559052 574154
rect 559046 574092 559052 574094
rect 559116 574092 559122 574156
rect 407297 574018 407363 574021
rect 552105 574018 552171 574021
rect 407297 574016 410044 574018
rect 407297 573960 407302 574016
rect 407358 573960 410044 574016
rect 407297 573958 410044 573960
rect 549884 574016 552171 574018
rect 549884 573960 552110 574016
rect 552166 573960 552171 574016
rect 549884 573958 552171 573960
rect 407297 573955 407363 573958
rect 552105 573955 552171 573958
rect 407297 573338 407363 573341
rect 407297 573336 410044 573338
rect 407297 573280 407302 573336
rect 407358 573280 410044 573336
rect 407297 573278 410044 573280
rect 407297 573275 407363 573278
rect 407297 572658 407363 572661
rect 407297 572656 410044 572658
rect 407297 572600 407302 572656
rect 407358 572600 410044 572656
rect 407297 572598 410044 572600
rect 407297 572595 407363 572598
rect 70301 571978 70367 571981
rect 350942 571978 350948 571980
rect 70301 571976 350948 571978
rect 70301 571920 70306 571976
rect 70362 571920 350948 571976
rect 70301 571918 350948 571920
rect 70301 571915 70367 571918
rect 350942 571916 350948 571918
rect 351012 571916 351018 571980
rect 47342 570692 47348 570756
rect 47412 570754 47418 570756
rect 277485 570754 277551 570757
rect 47412 570752 277551 570754
rect 47412 570696 277490 570752
rect 277546 570696 277551 570752
rect 47412 570694 277551 570696
rect 47412 570692 47418 570694
rect 277485 570691 277551 570694
rect 34421 570618 34487 570621
rect 347998 570618 348004 570620
rect 34421 570616 348004 570618
rect 34421 570560 34426 570616
rect 34482 570560 348004 570616
rect 34421 570558 348004 570560
rect 34421 570555 34487 570558
rect 347998 570556 348004 570558
rect 348068 570556 348074 570620
rect 407941 570618 408007 570621
rect 407941 570616 410044 570618
rect 407941 570560 407946 570616
rect 408002 570560 410044 570616
rect 407941 570558 410044 570560
rect 407941 570555 408007 570558
rect 407297 569938 407363 569941
rect 552565 569938 552631 569941
rect 407297 569936 410044 569938
rect 407297 569880 407302 569936
rect 407358 569880 410044 569936
rect 407297 569878 410044 569880
rect 549884 569936 552631 569938
rect 549884 569880 552570 569936
rect 552626 569880 552631 569936
rect 549884 569878 552631 569880
rect 407297 569875 407363 569878
rect 552565 569875 552631 569878
rect 47158 569196 47164 569260
rect 47228 569258 47234 569260
rect 252645 569258 252711 569261
rect 47228 569256 252711 569258
rect 47228 569200 252650 569256
rect 252706 569200 252711 569256
rect 47228 569198 252711 569200
rect 47228 569196 47234 569198
rect 252645 569195 252711 569198
rect 289169 568850 289235 568853
rect 353518 568850 353524 568852
rect 289169 568848 353524 568850
rect 289169 568792 289174 568848
rect 289230 568792 353524 568848
rect 289169 568790 353524 568792
rect 289169 568787 289235 568790
rect 353518 568788 353524 568790
rect 353588 568788 353594 568852
rect 77753 568714 77819 568717
rect 396574 568714 396580 568716
rect 77753 568712 396580 568714
rect 77753 568656 77758 568712
rect 77814 568656 396580 568712
rect 77753 568654 396580 568656
rect 77753 568651 77819 568654
rect 396574 568652 396580 568654
rect 396644 568652 396650 568716
rect 552473 568578 552539 568581
rect 549884 568576 552539 568578
rect 549884 568520 552478 568576
rect 552534 568520 552539 568576
rect 549884 568518 552539 568520
rect 552473 568515 552539 568518
rect 46238 567836 46244 567900
rect 46308 567898 46314 567900
rect 313273 567898 313339 567901
rect 46308 567896 313339 567898
rect 46308 567840 313278 567896
rect 313334 567840 313339 567896
rect 46308 567838 313339 567840
rect 46308 567836 46314 567838
rect 313273 567835 313339 567838
rect 407297 567898 407363 567901
rect 553301 567898 553367 567901
rect 407297 567896 410044 567898
rect 407297 567840 407302 567896
rect 407358 567840 410044 567896
rect 407297 567838 410044 567840
rect 549884 567896 553367 567898
rect 549884 567840 553306 567896
rect 553362 567840 553367 567896
rect 549884 567838 553367 567840
rect 407297 567835 407363 567838
rect 553301 567835 553367 567838
rect 335353 567490 335419 567493
rect 347630 567490 347636 567492
rect 335353 567488 347636 567490
rect 335353 567432 335358 567488
rect 335414 567432 347636 567488
rect 335353 567430 347636 567432
rect 335353 567427 335419 567430
rect 347630 567428 347636 567430
rect 347700 567428 347706 567492
rect 106089 567354 106155 567357
rect 391054 567354 391060 567356
rect 106089 567352 391060 567354
rect 106089 567296 106094 567352
rect 106150 567296 391060 567352
rect 106089 567294 391060 567296
rect 106089 567291 106155 567294
rect 391054 567292 391060 567294
rect 391124 567292 391130 567356
rect 85481 567218 85547 567221
rect 398598 567218 398604 567220
rect 85481 567216 398604 567218
rect 85481 567160 85486 567216
rect 85542 567160 398604 567216
rect 85481 567158 398604 567160
rect 85481 567155 85547 567158
rect 398598 567156 398604 567158
rect 398668 567156 398674 567220
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 553342 566538 553348 566540
rect 549884 566478 553348 566538
rect 553342 566476 553348 566478
rect 553412 566476 553418 566540
rect 241421 566402 241487 566405
rect 363638 566402 363644 566404
rect 241421 566400 363644 566402
rect 241421 566344 241426 566400
rect 241482 566344 363644 566400
rect 241421 566342 363644 566344
rect 241421 566339 241487 566342
rect 363638 566340 363644 566342
rect 363708 566340 363714 566404
rect 190361 566266 190427 566269
rect 389766 566266 389772 566268
rect 190361 566264 389772 566266
rect 190361 566208 190366 566264
rect 190422 566208 389772 566264
rect 190361 566206 389772 566208
rect 190361 566203 190427 566206
rect 389766 566204 389772 566206
rect 389836 566204 389842 566268
rect 157793 566130 157859 566133
rect 359590 566130 359596 566132
rect 157793 566128 359596 566130
rect 157793 566072 157798 566128
rect 157854 566072 359596 566128
rect 157793 566070 359596 566072
rect 157793 566067 157859 566070
rect 359590 566068 359596 566070
rect 359660 566068 359666 566132
rect 109585 565994 109651 565997
rect 351862 565994 351868 565996
rect 109585 565992 351868 565994
rect 109585 565936 109590 565992
rect 109646 565936 351868 565992
rect 109585 565934 351868 565936
rect 109585 565931 109651 565934
rect 351862 565932 351868 565934
rect 351932 565932 351938 565996
rect 24669 565858 24735 565861
rect 352046 565858 352052 565860
rect 24669 565856 352052 565858
rect 24669 565800 24674 565856
rect 24730 565800 352052 565856
rect 24669 565798 352052 565800
rect 24669 565795 24735 565798
rect 352046 565796 352052 565798
rect 352116 565796 352122 565860
rect 373206 565796 373212 565860
rect 373276 565858 373282 565860
rect 373276 565798 410044 565858
rect 373276 565796 373282 565798
rect 408033 565178 408099 565181
rect 563278 565178 563284 565180
rect 408033 565176 410044 565178
rect 408033 565120 408038 565176
rect 408094 565120 410044 565176
rect 408033 565118 410044 565120
rect 549884 565118 563284 565178
rect 408033 565115 408099 565118
rect 563278 565116 563284 565118
rect 563348 565116 563354 565180
rect 322105 564906 322171 564909
rect 356094 564906 356100 564908
rect 322105 564904 356100 564906
rect 322105 564848 322110 564904
rect 322166 564848 356100 564904
rect 322105 564846 356100 564848
rect 322105 564843 322171 564846
rect 356094 564844 356100 564846
rect 356164 564844 356170 564908
rect 297633 564770 297699 564773
rect 387149 564770 387215 564773
rect 297633 564768 387215 564770
rect 297633 564712 297638 564768
rect 297694 564712 387154 564768
rect 387210 564712 387215 564768
rect 297633 564710 387215 564712
rect 297633 564707 297699 564710
rect 387149 564707 387215 564710
rect 195881 564634 195947 564637
rect 373349 564634 373415 564637
rect 195881 564632 373415 564634
rect 195881 564576 195886 564632
rect 195942 564576 373354 564632
rect 373410 564576 373415 564632
rect 195881 564574 373415 564576
rect 195881 564571 195947 564574
rect 373349 564571 373415 564574
rect 59813 564498 59879 564501
rect 394049 564498 394115 564501
rect 59813 564496 394115 564498
rect 59813 564440 59818 564496
rect 59874 564440 394054 564496
rect 394110 564440 394115 564496
rect 59813 564438 394115 564440
rect 59813 564435 59879 564438
rect 394049 564435 394115 564438
rect 407389 564498 407455 564501
rect 550449 564498 550515 564501
rect 407389 564496 410044 564498
rect 407389 564440 407394 564496
rect 407450 564440 410044 564496
rect 407389 564438 410044 564440
rect 549884 564496 550515 564498
rect 549884 564440 550454 564496
rect 550510 564440 550515 564496
rect 549884 564438 550515 564440
rect 407389 564435 407455 564438
rect 550449 564435 550515 564438
rect 580533 564362 580599 564365
rect 583520 564362 584960 564452
rect 580533 564360 584960 564362
rect 580533 564304 580538 564360
rect 580594 564304 584960 564360
rect 580533 564302 584960 564304
rect 580533 564299 580599 564302
rect 583520 564212 584960 564302
rect 46422 563620 46428 563684
rect 46492 563682 46498 563684
rect 153837 563682 153903 563685
rect 46492 563680 153903 563682
rect 46492 563624 153842 563680
rect 153898 563624 153903 563680
rect 46492 563622 153903 563624
rect 46492 563620 46498 563622
rect 153837 563619 153903 563622
rect 328361 563682 328427 563685
rect 368933 563682 368999 563685
rect 328361 563680 368999 563682
rect 328361 563624 328366 563680
rect 328422 563624 368938 563680
rect 368994 563624 368999 563680
rect 328361 563622 368999 563624
rect 328361 563619 328427 563622
rect 368933 563619 368999 563622
rect 260741 563546 260807 563549
rect 349286 563546 349292 563548
rect 260741 563544 349292 563546
rect 260741 563488 260746 563544
rect 260802 563488 349292 563544
rect 260741 563486 349292 563488
rect 260741 563483 260807 563486
rect 349286 563484 349292 563486
rect 349356 563484 349362 563548
rect 188705 563410 188771 563413
rect 381486 563410 381492 563412
rect 188705 563408 381492 563410
rect 188705 563352 188710 563408
rect 188766 563352 381492 563408
rect 188705 563350 381492 563352
rect 188705 563347 188771 563350
rect 381486 563348 381492 563350
rect 381556 563348 381562 563412
rect 83089 563274 83155 563277
rect 390001 563274 390067 563277
rect 83089 563272 390067 563274
rect 83089 563216 83094 563272
rect 83150 563216 390006 563272
rect 390062 563216 390067 563272
rect 83089 563214 390067 563216
rect 83089 563211 83155 563214
rect 390001 563211 390067 563214
rect 43989 563138 44055 563141
rect 391422 563138 391428 563140
rect 43989 563136 391428 563138
rect 43989 563080 43994 563136
rect 44050 563080 391428 563136
rect 43989 563078 391428 563080
rect 43989 563075 44055 563078
rect 391422 563076 391428 563078
rect 391492 563076 391498 563140
rect 39614 562668 39620 562732
rect 39684 562730 39690 562732
rect 294321 562730 294387 562733
rect 39684 562728 294387 562730
rect 39684 562672 294326 562728
rect 294382 562672 294387 562728
rect 39684 562670 294387 562672
rect 39684 562668 39690 562670
rect 294321 562667 294387 562670
rect 48446 562532 48452 562596
rect 48516 562594 48522 562596
rect 164325 562594 164391 562597
rect 48516 562592 164391 562594
rect 48516 562536 164330 562592
rect 164386 562536 164391 562592
rect 48516 562534 164391 562536
rect 48516 562532 48522 562534
rect 164325 562531 164391 562534
rect 274449 562594 274515 562597
rect 384573 562594 384639 562597
rect 274449 562592 384639 562594
rect 274449 562536 274454 562592
rect 274510 562536 384578 562592
rect 384634 562536 384639 562592
rect 274449 562534 384639 562536
rect 274449 562531 274515 562534
rect 384573 562531 384639 562534
rect 48630 562396 48636 562460
rect 48700 562458 48706 562460
rect 86309 562458 86375 562461
rect 48700 562456 86375 562458
rect 48700 562400 86314 562456
rect 86370 562400 86375 562456
rect 48700 562398 86375 562400
rect 48700 562396 48706 562398
rect 86309 562395 86375 562398
rect 308029 562458 308095 562461
rect 371969 562458 372035 562461
rect 552013 562458 552079 562461
rect 308029 562456 372035 562458
rect 308029 562400 308034 562456
rect 308090 562400 371974 562456
rect 372030 562400 372035 562456
rect 308029 562398 372035 562400
rect 549884 562456 552079 562458
rect 549884 562400 552018 562456
rect 552074 562400 552079 562456
rect 549884 562398 552079 562400
rect 308029 562395 308095 562398
rect 371969 562395 372035 562398
rect 552013 562395 552079 562398
rect 44766 562260 44772 562324
rect 44836 562322 44842 562324
rect 89713 562322 89779 562325
rect 44836 562320 89779 562322
rect 44836 562264 89718 562320
rect 89774 562264 89779 562320
rect 44836 562262 89779 562264
rect 44836 562260 44842 562262
rect 89713 562259 89779 562262
rect 240041 562322 240107 562325
rect 387057 562322 387123 562325
rect 240041 562320 387123 562322
rect 240041 562264 240046 562320
rect 240102 562264 387062 562320
rect 387118 562264 387123 562320
rect 240041 562262 387123 562264
rect 240041 562259 240107 562262
rect 387057 562259 387123 562262
rect 30097 562186 30163 562189
rect 57421 562186 57487 562189
rect 30097 562184 57487 562186
rect 30097 562128 30102 562184
rect 30158 562128 57426 562184
rect 57482 562128 57487 562184
rect 30097 562126 57487 562128
rect 30097 562123 30163 562126
rect 57421 562123 57487 562126
rect 59169 562186 59235 562189
rect 125685 562186 125751 562189
rect 59169 562184 125751 562186
rect 59169 562128 59174 562184
rect 59230 562128 125690 562184
rect 125746 562128 125751 562184
rect 59169 562126 125751 562128
rect 59169 562123 59235 562126
rect 125685 562123 125751 562126
rect 192569 562186 192635 562189
rect 364374 562186 364380 562188
rect 192569 562184 364380 562186
rect 192569 562128 192574 562184
rect 192630 562128 364380 562184
rect 192569 562126 364380 562128
rect 192569 562123 192635 562126
rect 364374 562124 364380 562126
rect 364444 562124 364450 562188
rect 26049 562050 26115 562053
rect 57973 562050 58039 562053
rect 26049 562048 58039 562050
rect 26049 561992 26054 562048
rect 26110 561992 57978 562048
rect 58034 561992 58039 562048
rect 26049 561990 58039 561992
rect 26049 561987 26115 561990
rect 57973 561987 58039 561990
rect 59261 562050 59327 562053
rect 170765 562050 170831 562053
rect 59261 562048 170831 562050
rect 59261 561992 59266 562048
rect 59322 561992 170770 562048
rect 170826 561992 170831 562048
rect 59261 561990 170831 561992
rect 59261 561987 59327 561990
rect 170765 561987 170831 561990
rect 189441 562050 189507 562053
rect 372153 562050 372219 562053
rect 189441 562048 372219 562050
rect 189441 561992 189446 562048
rect 189502 561992 372158 562048
rect 372214 561992 372219 562048
rect 189441 561990 372219 561992
rect 189441 561987 189507 561990
rect 372153 561987 372219 561990
rect 27470 561852 27476 561916
rect 27540 561914 27546 561916
rect 59905 561914 59971 561917
rect 27540 561912 59971 561914
rect 27540 561856 59910 561912
rect 59966 561856 59971 561912
rect 27540 561854 59971 561856
rect 27540 561852 27546 561854
rect 59905 561851 59971 561854
rect 174537 561914 174603 561917
rect 360142 561914 360148 561916
rect 174537 561912 360148 561914
rect 174537 561856 174542 561912
rect 174598 561856 360148 561912
rect 174537 561854 360148 561856
rect 174537 561851 174603 561854
rect 360142 561852 360148 561854
rect 360212 561852 360218 561916
rect 28809 561778 28875 561781
rect 48957 561778 49023 561781
rect 28809 561776 49023 561778
rect 28809 561720 28814 561776
rect 28870 561720 48962 561776
rect 49018 561720 49023 561776
rect 28809 561718 49023 561720
rect 28809 561715 28875 561718
rect 48957 561715 49023 561718
rect 341977 561778 342043 561781
rect 360326 561778 360332 561780
rect 341977 561776 360332 561778
rect 341977 561720 341982 561776
rect 342038 561720 360332 561776
rect 341977 561718 360332 561720
rect 341977 561715 342043 561718
rect 360326 561716 360332 561718
rect 360396 561716 360402 561780
rect 44909 561370 44975 561373
rect 407849 561370 407915 561373
rect 44909 561368 407915 561370
rect 44909 561312 44914 561368
rect 44970 561312 407854 561368
rect 407910 561312 407915 561368
rect 44909 561310 407915 561312
rect 44909 561307 44975 561310
rect 407849 561307 407915 561310
rect 41270 561172 41276 561236
rect 41340 561234 41346 561236
rect 59261 561234 59327 561237
rect 41340 561232 59327 561234
rect 41340 561176 59266 561232
rect 59322 561176 59327 561232
rect 41340 561174 59327 561176
rect 41340 561172 41346 561174
rect 59261 561171 59327 561174
rect 34145 561098 34211 561101
rect 64965 561098 65031 561101
rect 34145 561096 65031 561098
rect 34145 561040 34150 561096
rect 34206 561040 64970 561096
rect 65026 561040 65031 561096
rect 34145 561038 65031 561040
rect 34145 561035 34211 561038
rect 64965 561035 65031 561038
rect 336365 561098 336431 561101
rect 376201 561098 376267 561101
rect 336365 561096 376267 561098
rect 336365 561040 336370 561096
rect 336426 561040 376206 561096
rect 376262 561040 376267 561096
rect 336365 561038 376267 561040
rect 336365 561035 336431 561038
rect 376201 561035 376267 561038
rect 407297 561098 407363 561101
rect 552933 561098 552999 561101
rect 407297 561096 410044 561098
rect 407297 561040 407302 561096
rect 407358 561040 410044 561096
rect 407297 561038 410044 561040
rect 549884 561096 552999 561098
rect 549884 561040 552938 561096
rect 552994 561040 552999 561096
rect 549884 561038 552999 561040
rect 407297 561035 407363 561038
rect 552933 561035 552999 561038
rect 27245 560962 27311 560965
rect 58065 560962 58131 560965
rect 27245 560960 58131 560962
rect 27245 560904 27250 560960
rect 27306 560904 58070 560960
rect 58126 560904 58131 560960
rect 27245 560902 58131 560904
rect 27245 560899 27311 560902
rect 58065 560899 58131 560902
rect 207473 560962 207539 560965
rect 395470 560962 395476 560964
rect 207473 560960 395476 560962
rect 207473 560904 207478 560960
rect 207534 560904 395476 560960
rect 207473 560902 395476 560904
rect 207473 560899 207539 560902
rect 395470 560900 395476 560902
rect 395540 560900 395546 560964
rect 34421 560826 34487 560829
rect 268009 560826 268075 560829
rect 34421 560824 268075 560826
rect 34421 560768 34426 560824
rect 34482 560768 268014 560824
rect 268070 560768 268075 560824
rect 34421 560766 268075 560768
rect 34421 560763 34487 560766
rect 268009 560763 268075 560766
rect 31661 560690 31727 560693
rect 330477 560690 330543 560693
rect 31661 560688 330543 560690
rect 31661 560632 31666 560688
rect 31722 560632 330482 560688
rect 330538 560632 330543 560688
rect 31661 560630 330543 560632
rect 31661 560627 31727 560630
rect 330477 560627 330543 560630
rect 63217 560554 63283 560557
rect 400806 560554 400812 560556
rect 63217 560552 400812 560554
rect 63217 560496 63222 560552
rect 63278 560496 400812 560552
rect 63217 560494 400812 560496
rect 63217 560491 63283 560494
rect 400806 560492 400812 560494
rect 400876 560492 400882 560556
rect 339401 560418 339467 560421
rect 347630 560418 347636 560420
rect 339401 560416 347636 560418
rect 339401 560360 339406 560416
rect 339462 560360 347636 560416
rect 339401 560358 347636 560360
rect 339401 560355 339467 560358
rect 347630 560356 347636 560358
rect 347700 560356 347706 560420
rect 553301 560418 553367 560421
rect 549884 560416 553367 560418
rect 549884 560360 553306 560416
rect 553362 560360 553367 560416
rect 549884 560358 553367 560360
rect 553301 560355 553367 560358
rect 30281 560282 30347 560285
rect 49601 560282 49667 560285
rect 30281 560280 49667 560282
rect 30281 560224 30286 560280
rect 30342 560224 49606 560280
rect 49662 560224 49667 560280
rect 30281 560222 49667 560224
rect 30281 560219 30347 560222
rect 49601 560219 49667 560222
rect 39573 560146 39639 560149
rect 51625 560146 51691 560149
rect 39573 560144 51691 560146
rect 39573 560088 39578 560144
rect 39634 560088 51630 560144
rect 51686 560088 51691 560144
rect 39573 560086 51691 560088
rect 39573 560083 39639 560086
rect 51625 560083 51691 560086
rect 346342 560084 346348 560148
rect 346412 560146 346418 560148
rect 347262 560146 347268 560148
rect 346412 560086 347268 560146
rect 346412 560084 346418 560086
rect 347262 560084 347268 560086
rect 347332 560084 347338 560148
rect 38009 560010 38075 560013
rect 51073 560010 51139 560013
rect 38009 560008 51139 560010
rect 38009 559952 38014 560008
rect 38070 559952 51078 560008
rect 51134 559952 51139 560008
rect 38009 559950 51139 559952
rect 38009 559947 38075 559950
rect 51073 559947 51139 559950
rect 315573 560010 315639 560013
rect 398189 560010 398255 560013
rect 315573 560008 398255 560010
rect 315573 559952 315578 560008
rect 315634 559952 398194 560008
rect 398250 559952 398255 560008
rect 315573 559950 398255 559952
rect 315573 559947 315639 559950
rect 398189 559947 398255 559950
rect 408033 559058 408099 559061
rect 408033 559056 410044 559058
rect 408033 559000 408038 559056
rect 408094 559000 410044 559056
rect 408033 558998 410044 559000
rect 408033 558995 408099 558998
rect 33869 558786 33935 558789
rect 48078 558786 48084 558788
rect 33869 558784 48084 558786
rect 33869 558728 33874 558784
rect 33930 558728 48084 558784
rect 33869 558726 48084 558728
rect 33869 558723 33935 558726
rect 48078 558724 48084 558726
rect 48148 558724 48154 558788
rect 552933 558378 552999 558381
rect 549884 558376 552999 558378
rect 549884 558320 552938 558376
rect 552994 558320 552999 558376
rect 549884 558318 552999 558320
rect 552933 558315 552999 558318
rect 347630 558180 347636 558244
rect 347700 558242 347706 558244
rect 402145 558242 402211 558245
rect 347700 558240 402211 558242
rect 347700 558184 402150 558240
rect 402206 558184 402211 558240
rect 347700 558182 402211 558184
rect 347700 558180 347706 558182
rect 402145 558179 402211 558182
rect 39246 558044 39252 558108
rect 39316 558106 39322 558108
rect 48262 558106 48268 558108
rect 39316 558046 48268 558106
rect 39316 558044 39322 558046
rect 48262 558044 48268 558046
rect 48332 558044 48338 558108
rect 389950 557636 389956 557700
rect 390020 557698 390026 557700
rect 553301 557698 553367 557701
rect 390020 557638 410044 557698
rect 549884 557696 553367 557698
rect 549884 557640 553306 557696
rect 553362 557640 553367 557696
rect 549884 557638 553367 557640
rect 390020 557636 390026 557638
rect 553301 557635 553367 557638
rect 347630 557364 347636 557428
rect 347700 557426 347706 557428
rect 348550 557426 348556 557428
rect 347700 557366 348556 557426
rect 347700 557364 347706 557366
rect 348550 557364 348556 557366
rect 348620 557364 348626 557428
rect 347630 557228 347636 557292
rect 347700 557228 347706 557292
rect 347638 557124 347698 557228
rect 46289 556610 46355 556613
rect 48086 556610 48146 557056
rect 407941 557018 408007 557021
rect 552013 557018 552079 557021
rect 407941 557016 410044 557018
rect 407941 556960 407946 557016
rect 408002 556960 410044 557016
rect 407941 556958 410044 556960
rect 549884 557016 552079 557018
rect 549884 556960 552018 557016
rect 552074 556960 552079 557016
rect 549884 556958 552079 556960
rect 407941 556955 408007 556958
rect 552013 556955 552079 556958
rect 46289 556608 48146 556610
rect 46289 556552 46294 556608
rect 46350 556552 48146 556608
rect 46289 556550 48146 556552
rect 46289 556547 46355 556550
rect 406745 556338 406811 556341
rect 558126 556338 558132 556340
rect 406745 556336 410044 556338
rect 406745 556280 406750 556336
rect 406806 556280 410044 556336
rect 406745 556278 410044 556280
rect 549884 556278 558132 556338
rect 406745 556275 406811 556278
rect 558126 556276 558132 556278
rect 558196 556276 558202 556340
rect 46105 556202 46171 556205
rect 48262 556202 48268 556204
rect 46105 556200 48268 556202
rect 46105 556144 46110 556200
rect 46166 556144 48268 556200
rect 46105 556142 48268 556144
rect 46105 556139 46171 556142
rect 48262 556140 48268 556142
rect 48332 556140 48338 556204
rect 347630 556140 347636 556204
rect 347700 556202 347706 556204
rect 349470 556202 349476 556204
rect 347700 556142 349476 556202
rect 347700 556140 347706 556142
rect 349470 556140 349476 556142
rect 349540 556140 349546 556204
rect 407573 555658 407639 555661
rect 552289 555658 552355 555661
rect 407573 555656 410044 555658
rect 407573 555600 407578 555656
rect 407634 555600 410044 555656
rect 407573 555598 410044 555600
rect 549884 555656 552355 555658
rect 549884 555600 552294 555656
rect 552350 555600 552355 555656
rect 549884 555598 552355 555600
rect 407573 555595 407639 555598
rect 552289 555595 552355 555598
rect 349429 554434 349495 554437
rect 347852 554432 349495 554434
rect 347852 554376 349434 554432
rect 349490 554376 349495 554432
rect 347852 554374 349495 554376
rect 349429 554371 349495 554374
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 552013 553618 552079 553621
rect 550222 553616 552079 553618
rect 550222 553560 552018 553616
rect 552074 553560 552079 553616
rect 550222 553558 552079 553560
rect 550222 553550 550282 553558
rect 552013 553555 552079 553558
rect 549884 553490 550282 553550
rect 407297 552938 407363 552941
rect 552381 552938 552447 552941
rect 407297 552936 410044 552938
rect 407297 552880 407302 552936
rect 407358 552880 410044 552936
rect 407297 552878 410044 552880
rect 549884 552936 552447 552938
rect 549884 552880 552386 552936
rect 552442 552880 552447 552936
rect 549884 552878 552447 552880
rect 407297 552875 407363 552878
rect 552381 552875 552447 552878
rect 566222 552258 566228 552260
rect 549884 552198 566228 552258
rect 566222 552196 566228 552198
rect 566292 552196 566298 552260
rect 46289 551442 46355 551445
rect 48086 551442 48146 551616
rect 46289 551440 48146 551442
rect 46289 551384 46294 551440
rect 46350 551384 48146 551440
rect 46289 551382 48146 551384
rect 46289 551379 46355 551382
rect 347822 551170 347882 551616
rect 407389 551578 407455 551581
rect 566406 551578 566412 551580
rect 407389 551576 410044 551578
rect 407389 551520 407394 551576
rect 407450 551520 410044 551576
rect 407389 551518 410044 551520
rect 549884 551518 566412 551578
rect 407389 551515 407455 551518
rect 566406 551516 566412 551518
rect 566476 551516 566482 551580
rect 350441 551170 350507 551173
rect 347822 551168 350507 551170
rect 347822 551112 350446 551168
rect 350502 551112 350507 551168
rect 347822 551110 350507 551112
rect 350441 551107 350507 551110
rect 583520 551020 584960 551260
rect 46289 550898 46355 550901
rect 48086 550898 48146 550936
rect 46289 550896 48146 550898
rect 46289 550840 46294 550896
rect 46350 550840 48146 550896
rect 46289 550838 48146 550840
rect 407297 550898 407363 550901
rect 553301 550898 553367 550901
rect 407297 550896 410044 550898
rect 407297 550840 407302 550896
rect 407358 550840 410044 550896
rect 407297 550838 410044 550840
rect 549884 550896 553367 550898
rect 549884 550840 553306 550896
rect 553362 550840 553367 550896
rect 549884 550838 553367 550840
rect 46289 550835 46355 550838
rect 407297 550835 407363 550838
rect 553301 550835 553367 550838
rect 46289 549810 46355 549813
rect 48086 549810 48146 550256
rect 407297 550218 407363 550221
rect 407297 550216 410044 550218
rect 407297 550160 407302 550216
rect 407358 550160 410044 550216
rect 407297 550158 410044 550160
rect 407297 550155 407363 550158
rect 46289 549808 48146 549810
rect 46289 549752 46294 549808
rect 46350 549752 48146 549808
rect 46289 549750 48146 549752
rect 46289 549747 46355 549750
rect 553301 549538 553367 549541
rect 549884 549536 553367 549538
rect 549884 549480 553306 549536
rect 553362 549480 553367 549536
rect 549884 549478 553367 549480
rect 553301 549475 553367 549478
rect 352046 548994 352052 548996
rect 347852 548934 352052 548994
rect 352046 548932 352052 548934
rect 352116 548932 352122 548996
rect 45318 548252 45324 548316
rect 45388 548314 45394 548316
rect 48086 548314 48146 548896
rect 407849 548858 407915 548861
rect 407849 548856 410044 548858
rect 407849 548800 407854 548856
rect 407910 548800 410044 548856
rect 407849 548798 410044 548800
rect 407849 548795 407915 548798
rect 45388 548254 48146 548314
rect 45388 548252 45394 548254
rect 347822 547090 347882 547536
rect 407297 547498 407363 547501
rect 553117 547498 553183 547501
rect 407297 547496 410044 547498
rect 407297 547440 407302 547496
rect 407358 547440 410044 547496
rect 407297 547438 410044 547440
rect 549884 547496 553183 547498
rect 549884 547440 553122 547496
rect 553178 547440 553183 547496
rect 549884 547438 553183 547440
rect 407297 547435 407363 547438
rect 553117 547435 553183 547438
rect 350165 547090 350231 547093
rect 347822 547088 350231 547090
rect 347822 547032 350170 547088
rect 350226 547032 350231 547088
rect 347822 547030 350231 547032
rect 350165 547027 350231 547030
rect 46105 546546 46171 546549
rect 48086 546546 48146 546856
rect 46105 546544 48146 546546
rect 46105 546488 46110 546544
rect 46166 546488 48146 546544
rect 46105 546486 48146 546488
rect 347822 546546 347882 546856
rect 553301 546818 553367 546821
rect 549884 546816 553367 546818
rect 549884 546760 553306 546816
rect 553362 546760 553367 546816
rect 549884 546758 553367 546760
rect 553301 546755 553367 546758
rect 350441 546546 350507 546549
rect 347822 546544 350507 546546
rect 347822 546488 350446 546544
rect 350502 546488 350507 546544
rect 347822 546486 350507 546488
rect 46105 546483 46171 546486
rect 350441 546483 350507 546486
rect 46013 545730 46079 545733
rect 48086 545730 48146 546176
rect 407757 546138 407823 546141
rect 407757 546136 410044 546138
rect 407757 546080 407762 546136
rect 407818 546080 410044 546136
rect 407757 546078 410044 546080
rect 407757 546075 407823 546078
rect 46013 545728 48146 545730
rect 46013 545672 46018 545728
rect 46074 545672 48146 545728
rect 46013 545670 48146 545672
rect 46013 545667 46079 545670
rect 552105 545458 552171 545461
rect 549884 545456 552171 545458
rect 549884 545400 552110 545456
rect 552166 545400 552171 545456
rect 549884 545398 552171 545400
rect 552105 545395 552171 545398
rect 46105 544370 46171 544373
rect 48086 544370 48146 544816
rect 407297 544778 407363 544781
rect 574318 544778 574324 544780
rect 407297 544776 410044 544778
rect 407297 544720 407302 544776
rect 407358 544720 410044 544776
rect 407297 544718 410044 544720
rect 549884 544718 574324 544778
rect 407297 544715 407363 544718
rect 574318 544716 574324 544718
rect 574388 544716 574394 544780
rect 46105 544368 48146 544370
rect 46105 544312 46110 544368
rect 46166 544312 48146 544368
rect 46105 544310 48146 544312
rect 46105 544307 46171 544310
rect 45921 544234 45987 544237
rect 45921 544232 48116 544234
rect 45921 544176 45926 544232
rect 45982 544176 48116 544232
rect 45921 544174 48116 544176
rect 45921 544171 45987 544174
rect 407389 544098 407455 544101
rect 553301 544098 553367 544101
rect 407389 544096 410044 544098
rect 407389 544040 407394 544096
rect 407450 544040 410044 544096
rect 407389 544038 410044 544040
rect 549884 544096 553367 544098
rect 549884 544040 553306 544096
rect 553362 544040 553367 544096
rect 549884 544038 553367 544040
rect 407389 544035 407455 544038
rect 553301 544035 553367 544038
rect 347822 543010 347882 543456
rect 350441 543010 350507 543013
rect 347822 543008 350507 543010
rect 347822 542952 350446 543008
rect 350502 542952 350507 543008
rect 347822 542950 350507 542952
rect 350441 542947 350507 542950
rect 407297 542058 407363 542061
rect 407297 542056 410044 542058
rect 407297 542000 407302 542056
rect 407358 542000 410044 542056
rect 407297 541998 410044 542000
rect 407297 541995 407363 541998
rect 349153 541514 349219 541517
rect 347852 541512 349219 541514
rect 347852 541456 349158 541512
rect 349214 541456 349219 541512
rect 347852 541454 349219 541456
rect 349153 541451 349219 541454
rect 46105 541106 46171 541109
rect 48086 541106 48146 541416
rect 46105 541104 48146 541106
rect 46105 541048 46110 541104
rect 46166 541048 48146 541104
rect 46105 541046 48146 541048
rect 46105 541043 46171 541046
rect -960 540684 480 540924
rect 552565 540698 552631 540701
rect 549884 540696 552631 540698
rect 549884 540640 552570 540696
rect 552626 540640 552631 540696
rect 549884 540638 552631 540640
rect 552565 540635 552631 540638
rect 550449 540018 550515 540021
rect 549884 540016 550515 540018
rect 549884 539960 550454 540016
rect 550510 539960 550515 540016
rect 549884 539958 550515 539960
rect 550449 539955 550515 539958
rect 552565 539338 552631 539341
rect 549884 539336 552631 539338
rect 549884 539280 552570 539336
rect 552626 539280 552631 539336
rect 549884 539278 552631 539280
rect 552565 539275 552631 539278
rect 347822 538386 347882 538696
rect 350441 538386 350507 538389
rect 347822 538384 350507 538386
rect 347822 538328 350446 538384
rect 350502 538328 350507 538384
rect 347822 538326 350507 538328
rect 350441 538323 350507 538326
rect 46105 538114 46171 538117
rect 46105 538112 48116 538114
rect 46105 538056 46110 538112
rect 46166 538056 48116 538112
rect 46105 538054 48116 538056
rect 46105 538051 46171 538054
rect 407757 537978 407823 537981
rect 407757 537976 410044 537978
rect 407757 537920 407762 537976
rect 407818 537920 410044 537976
rect 407757 537918 410044 537920
rect 407757 537915 407823 537918
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect 347822 536890 347882 537336
rect 350441 536890 350507 536893
rect 347822 536888 350507 536890
rect 347822 536832 350446 536888
rect 350502 536832 350507 536888
rect 347822 536830 350507 536832
rect 350441 536827 350507 536830
rect 552013 536618 552079 536621
rect 550222 536616 552079 536618
rect 550222 536560 552018 536616
rect 552074 536560 552079 536616
rect 550222 536558 552079 536560
rect 550222 536550 550282 536558
rect 552013 536555 552079 536558
rect 549884 536490 550282 536550
rect 553301 535938 553367 535941
rect 549884 535936 553367 535938
rect 549884 535880 553306 535936
rect 553362 535880 553367 535936
rect 549884 535878 553367 535880
rect 553301 535875 553367 535878
rect 347822 534714 347882 535296
rect 407297 535258 407363 535261
rect 553301 535258 553367 535261
rect 407297 535256 410044 535258
rect 407297 535200 407302 535256
rect 407358 535200 410044 535256
rect 407297 535198 410044 535200
rect 549884 535256 553367 535258
rect 549884 535200 553306 535256
rect 553362 535200 553367 535256
rect 549884 535198 553367 535200
rect 407297 535195 407363 535198
rect 553301 535195 553367 535198
rect 350441 534714 350507 534717
rect 347822 534712 350507 534714
rect 347822 534656 350446 534712
rect 350502 534656 350507 534712
rect 347822 534654 350507 534656
rect 350441 534651 350507 534654
rect 38510 534108 38516 534172
rect 38580 534170 38586 534172
rect 48086 534170 48146 534616
rect 552381 534578 552447 534581
rect 549884 534576 552447 534578
rect 549884 534520 552386 534576
rect 552442 534520 552447 534576
rect 549884 534518 552447 534520
rect 552381 534515 552447 534518
rect 38580 534110 48146 534170
rect 38580 534108 38586 534110
rect 41822 533292 41828 533356
rect 41892 533354 41898 533356
rect 48086 533354 48146 533936
rect 347822 533490 347882 533936
rect 407614 533836 407620 533900
rect 407684 533898 407690 533900
rect 552473 533898 552539 533901
rect 407684 533838 410044 533898
rect 549884 533896 552539 533898
rect 549884 533840 552478 533896
rect 552534 533840 552539 533896
rect 549884 533838 552539 533840
rect 407684 533836 407690 533838
rect 552473 533835 552539 533838
rect 350165 533490 350231 533493
rect 347822 533488 350231 533490
rect 347822 533432 350170 533488
rect 350226 533432 350231 533488
rect 347822 533430 350231 533432
rect 350165 533427 350231 533430
rect 41892 533294 48146 533354
rect 41892 533292 41898 533294
rect 347822 532810 347882 533256
rect 350441 532810 350507 532813
rect 347822 532808 350507 532810
rect 347822 532752 350446 532808
rect 350502 532752 350507 532808
rect 347822 532750 350507 532752
rect 350441 532747 350507 532750
rect 46013 532266 46079 532269
rect 48086 532266 48146 532576
rect 46013 532264 48146 532266
rect 46013 532208 46018 532264
rect 46074 532208 48146 532264
rect 46013 532206 48146 532208
rect 46013 532203 46079 532206
rect 347822 532130 347882 532576
rect 552013 532538 552079 532541
rect 549884 532536 552079 532538
rect 549884 532480 552018 532536
rect 552074 532480 552079 532536
rect 549884 532478 552079 532480
rect 552013 532475 552079 532478
rect 349429 532130 349495 532133
rect 347822 532128 349495 532130
rect 347822 532072 349434 532128
rect 349490 532072 349495 532128
rect 347822 532070 349495 532072
rect 349429 532067 349495 532070
rect 406561 531858 406627 531861
rect 560886 531858 560892 531860
rect 406561 531856 410044 531858
rect 406561 531800 406566 531856
rect 406622 531800 410044 531856
rect 406561 531798 410044 531800
rect 549884 531798 560892 531858
rect 406561 531795 406627 531798
rect 560886 531796 560892 531798
rect 560956 531796 560962 531860
rect 44030 530708 44036 530772
rect 44100 530770 44106 530772
rect 48086 530770 48146 531216
rect 44100 530710 48146 530770
rect 347822 530770 347882 531216
rect 552657 531178 552723 531181
rect 549884 531176 552723 531178
rect 549884 531120 552662 531176
rect 552718 531120 552723 531176
rect 549884 531118 552723 531120
rect 552657 531115 552723 531118
rect 350441 530770 350507 530773
rect 347822 530768 350507 530770
rect 347822 530712 350446 530768
rect 350502 530712 350507 530768
rect 347822 530710 350507 530712
rect 44100 530708 44106 530710
rect 350441 530707 350507 530710
rect 552013 530498 552079 530501
rect 549884 530496 552079 530498
rect 549884 530440 552018 530496
rect 552074 530440 552079 530496
rect 549884 530438 552079 530440
rect 552013 530435 552079 530438
rect 46105 529954 46171 529957
rect 46105 529952 48116 529954
rect 46105 529896 46110 529952
rect 46166 529896 48116 529952
rect 46105 529894 48116 529896
rect 46105 529891 46171 529894
rect 45829 529002 45895 529005
rect 48086 529002 48146 529176
rect 407297 529138 407363 529141
rect 407297 529136 410044 529138
rect 407297 529080 407302 529136
rect 407358 529080 410044 529136
rect 407297 529078 410044 529080
rect 407297 529075 407363 529078
rect 45829 529000 48146 529002
rect 45829 528944 45834 529000
rect 45890 528944 48146 529000
rect 45829 528942 48146 528944
rect 45829 528939 45895 528942
rect 553301 528458 553367 528461
rect 549884 528456 553367 528458
rect 549884 528400 553306 528456
rect 553362 528400 553367 528456
rect 549884 528398 553367 528400
rect 553301 528395 553367 528398
rect -960 527764 480 528004
rect 37038 527308 37044 527372
rect 37108 527370 37114 527372
rect 48086 527370 48146 527816
rect 37108 527310 48146 527370
rect 37108 527308 37114 527310
rect 36854 527172 36860 527236
rect 36924 527234 36930 527236
rect 350441 527234 350507 527237
rect 36924 527174 48116 527234
rect 347852 527232 350507 527234
rect 347852 527176 350446 527232
rect 350502 527176 350507 527232
rect 347852 527174 350507 527176
rect 36924 527172 36930 527174
rect 350441 527171 350507 527174
rect 378910 527036 378916 527100
rect 378980 527098 378986 527100
rect 378980 527038 410044 527098
rect 378980 527036 378986 527038
rect 46197 526554 46263 526557
rect 46197 526552 48116 526554
rect 46197 526496 46202 526552
rect 46258 526496 48116 526552
rect 46197 526494 48116 526496
rect 46197 526491 46263 526494
rect 347822 526010 347882 526456
rect 552013 526418 552079 526421
rect 549884 526416 552079 526418
rect 549884 526360 552018 526416
rect 552074 526360 552079 526416
rect 549884 526358 552079 526360
rect 552013 526355 552079 526358
rect 350441 526010 350507 526013
rect 347822 526008 350507 526010
rect 347822 525952 350446 526008
rect 350502 525952 350507 526008
rect 347822 525950 350507 525952
rect 350441 525947 350507 525950
rect 407389 525738 407455 525741
rect 552013 525738 552079 525741
rect 407389 525736 410044 525738
rect 407389 525680 407394 525736
rect 407450 525680 410044 525736
rect 407389 525678 410044 525680
rect 549884 525736 552079 525738
rect 549884 525680 552018 525736
rect 552074 525680 552079 525736
rect 549884 525678 552079 525680
rect 407389 525675 407455 525678
rect 552013 525675 552079 525678
rect 45645 525194 45711 525197
rect 45645 525192 48116 525194
rect 45645 525136 45650 525192
rect 45706 525136 48116 525192
rect 45645 525134 48116 525136
rect 45645 525131 45711 525134
rect 407297 525058 407363 525061
rect 407297 525056 410044 525058
rect 407297 525000 407302 525056
rect 407358 525000 410044 525056
rect 407297 524998 410044 525000
rect 407297 524995 407363 524998
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 551093 524378 551159 524381
rect 549884 524376 551159 524378
rect 549884 524320 551098 524376
rect 551154 524320 551159 524376
rect 583520 524364 584960 524454
rect 549884 524318 551159 524320
rect 551093 524315 551159 524318
rect 347822 523290 347882 523736
rect 407297 523698 407363 523701
rect 407297 523696 410044 523698
rect 407297 523640 407302 523696
rect 407358 523640 410044 523696
rect 407297 523638 410044 523640
rect 407297 523635 407363 523638
rect 347998 523500 348004 523564
rect 348068 523562 348074 523564
rect 348325 523562 348391 523565
rect 348068 523560 348391 523562
rect 348068 523504 348330 523560
rect 348386 523504 348391 523560
rect 348068 523502 348391 523504
rect 348068 523500 348074 523502
rect 348325 523499 348391 523502
rect 350441 523290 350507 523293
rect 347822 523288 350507 523290
rect 347822 523232 350446 523288
rect 350502 523232 350507 523288
rect 347822 523230 350507 523232
rect 350441 523227 350507 523230
rect 347822 522885 347882 523056
rect 348918 522956 348924 523020
rect 348988 523018 348994 523020
rect 350533 523018 350599 523021
rect 348988 523016 350599 523018
rect 348988 522960 350538 523016
rect 350594 522960 350599 523016
rect 348988 522958 350599 522960
rect 348988 522956 348994 522958
rect 350533 522955 350599 522958
rect 407389 523018 407455 523021
rect 407389 523016 410044 523018
rect 407389 522960 407394 523016
rect 407450 522960 410044 523016
rect 407389 522958 410044 522960
rect 407389 522955 407455 522958
rect 347822 522880 347931 522885
rect 347822 522824 347870 522880
rect 347926 522824 347931 522880
rect 347822 522822 347931 522824
rect 347865 522819 347931 522822
rect 407297 522338 407363 522341
rect 550357 522338 550423 522341
rect 407297 522336 410044 522338
rect 407297 522280 407302 522336
rect 407358 522280 410044 522336
rect 407297 522278 410044 522280
rect 549884 522336 550423 522338
rect 549884 522280 550362 522336
rect 550418 522280 550423 522336
rect 549884 522278 550423 522280
rect 407297 522275 407363 522278
rect 550357 522275 550423 522278
rect 47485 521794 47551 521797
rect 349889 521794 349955 521797
rect 47485 521792 48116 521794
rect 47485 521736 47490 521792
rect 47546 521736 48116 521792
rect 47485 521734 48116 521736
rect 347852 521792 349955 521794
rect 347852 521736 349894 521792
rect 349950 521736 349955 521792
rect 347852 521734 349955 521736
rect 47485 521731 47551 521734
rect 349889 521731 349955 521734
rect 407297 521658 407363 521661
rect 552013 521658 552079 521661
rect 407297 521656 410044 521658
rect 407297 521600 407302 521656
rect 407358 521600 410044 521656
rect 407297 521598 410044 521600
rect 549884 521656 552079 521658
rect 549884 521600 552018 521656
rect 552074 521600 552079 521656
rect 549884 521598 552079 521600
rect 407297 521595 407363 521598
rect 552013 521595 552079 521598
rect 48086 520570 48146 521016
rect 551185 520978 551251 520981
rect 549884 520976 551251 520978
rect 549884 520920 551190 520976
rect 551246 520920 551251 520976
rect 549884 520918 551251 520920
rect 551185 520915 551251 520918
rect 40726 520510 48146 520570
rect 35750 520372 35756 520436
rect 35820 520434 35826 520436
rect 40726 520434 40786 520510
rect 35820 520374 40786 520434
rect 46197 520434 46263 520437
rect 46197 520432 48116 520434
rect 46197 520376 46202 520432
rect 46258 520376 48116 520432
rect 46197 520374 48116 520376
rect 35820 520372 35826 520374
rect 46197 520371 46263 520374
rect 347822 520298 347882 520336
rect 350574 520298 350580 520300
rect 347822 520238 350580 520298
rect 350574 520236 350580 520238
rect 350644 520236 350650 520300
rect 549884 519490 550282 519550
rect 550222 519482 550282 519490
rect 552013 519482 552079 519485
rect 550222 519480 552079 519482
rect 550222 519424 552018 519480
rect 552074 519424 552079 519480
rect 550222 519422 552079 519424
rect 552013 519419 552079 519422
rect 347822 518938 347882 518976
rect 367134 518938 367140 518940
rect 347822 518878 367140 518938
rect 367134 518876 367140 518878
rect 367204 518876 367210 518940
rect 552013 518938 552079 518941
rect 549884 518936 552079 518938
rect 549884 518880 552018 518936
rect 552074 518880 552079 518936
rect 549884 518878 552079 518880
rect 552013 518875 552079 518878
rect 407389 518258 407455 518261
rect 407389 518256 410044 518258
rect 407389 518200 407394 518256
rect 407450 518200 410044 518256
rect 407389 518198 410044 518200
rect 407389 518195 407455 518198
rect 347822 517578 347882 517616
rect 350441 517578 350507 517581
rect 347822 517576 350507 517578
rect 347822 517520 350446 517576
rect 350502 517520 350507 517576
rect 347822 517518 350507 517520
rect 350441 517515 350507 517518
rect 407297 517578 407363 517581
rect 407297 517576 410044 517578
rect 407297 517520 407302 517576
rect 407358 517520 410044 517576
rect 407297 517518 410044 517520
rect 407297 517515 407363 517518
rect 46013 516626 46079 516629
rect 48086 516626 48146 516936
rect 46013 516624 48146 516626
rect 46013 516568 46018 516624
rect 46074 516568 48146 516624
rect 46013 516566 48146 516568
rect 347822 516626 347882 516936
rect 407389 516898 407455 516901
rect 552013 516898 552079 516901
rect 407389 516896 410044 516898
rect 407389 516840 407394 516896
rect 407450 516840 410044 516896
rect 407389 516838 410044 516840
rect 549884 516896 552079 516898
rect 549884 516840 552018 516896
rect 552074 516840 552079 516896
rect 549884 516838 552079 516840
rect 407389 516835 407455 516838
rect 552013 516835 552079 516838
rect 350073 516626 350139 516629
rect 347822 516624 350139 516626
rect 347822 516568 350078 516624
rect 350134 516568 350139 516624
rect 347822 516566 350139 516568
rect 46013 516563 46079 516566
rect 350073 516563 350139 516566
rect 350441 516354 350507 516357
rect 347852 516352 350507 516354
rect 347852 516296 350446 516352
rect 350502 516296 350507 516352
rect 347852 516294 350507 516296
rect 350441 516291 350507 516294
rect 407297 516218 407363 516221
rect 407297 516216 410044 516218
rect 407297 516160 407302 516216
rect 407358 516160 410044 516216
rect 407297 516158 410044 516160
rect 407297 516155 407363 516158
rect 42006 515068 42012 515132
rect 42076 515130 42082 515132
rect 48086 515130 48146 515576
rect 552289 515538 552355 515541
rect 549884 515536 552355 515538
rect 549884 515480 552294 515536
rect 552350 515480 552355 515536
rect 549884 515478 552355 515480
rect 552289 515475 552355 515478
rect 42076 515070 48146 515130
rect 42076 515068 42082 515070
rect -960 514858 480 514948
rect 30966 514858 30972 514860
rect -960 514798 30972 514858
rect -960 514708 480 514798
rect 30966 514796 30972 514798
rect 31036 514796 31042 514860
rect 34278 514796 34284 514860
rect 34348 514858 34354 514860
rect 48086 514858 48146 514896
rect 34348 514798 48146 514858
rect 407665 514858 407731 514861
rect 552013 514858 552079 514861
rect 407665 514856 410044 514858
rect 407665 514800 407670 514856
rect 407726 514800 410044 514856
rect 407665 514798 410044 514800
rect 549884 514856 552079 514858
rect 549884 514800 552018 514856
rect 552074 514800 552079 514856
rect 549884 514798 552079 514800
rect 34348 514796 34354 514798
rect 407665 514795 407731 514798
rect 552013 514795 552079 514798
rect 45921 513906 45987 513909
rect 48086 513906 48146 514216
rect 45921 513904 48146 513906
rect 45921 513848 45926 513904
rect 45982 513848 48146 513904
rect 45921 513846 48146 513848
rect 45921 513843 45987 513846
rect 347822 513770 347882 514216
rect 350441 513770 350507 513773
rect 347822 513768 350507 513770
rect 347822 513712 350446 513768
rect 350502 513712 350507 513768
rect 347822 513710 350507 513712
rect 350441 513707 350507 513710
rect 347822 513498 347882 513536
rect 350073 513498 350139 513501
rect 347822 513496 350139 513498
rect 347822 513440 350078 513496
rect 350134 513440 350139 513496
rect 347822 513438 350139 513440
rect 350073 513435 350139 513438
rect 407297 512818 407363 512821
rect 407297 512816 410044 512818
rect 407297 512760 407302 512816
rect 407358 512760 410044 512816
rect 407297 512758 410044 512760
rect 407297 512755 407363 512758
rect 407297 512138 407363 512141
rect 407297 512136 410044 512138
rect 407297 512080 407302 512136
rect 407358 512080 410044 512136
rect 407297 512078 410044 512080
rect 407297 512075 407363 512078
rect 350441 511594 350507 511597
rect 347852 511592 350507 511594
rect 347852 511536 350446 511592
rect 350502 511536 350507 511592
rect 347852 511534 350507 511536
rect 350441 511531 350507 511534
rect 583520 511172 584960 511412
rect 45737 510914 45803 510917
rect 45737 510912 48116 510914
rect 45737 510856 45742 510912
rect 45798 510856 48116 510912
rect 45737 510854 48116 510856
rect 45737 510851 45803 510854
rect 395654 510716 395660 510780
rect 395724 510778 395730 510780
rect 395724 510718 410044 510778
rect 395724 510716 395730 510718
rect 40769 510506 40835 510509
rect 41270 510506 41276 510508
rect 40769 510504 41276 510506
rect 40769 510448 40774 510504
rect 40830 510448 41276 510504
rect 40769 510446 41276 510448
rect 40769 510443 40835 510446
rect 41270 510444 41276 510446
rect 41340 510444 41346 510508
rect 409045 510098 409111 510101
rect 553301 510098 553367 510101
rect 409045 510096 410044 510098
rect 409045 510040 409050 510096
rect 409106 510040 410044 510096
rect 409045 510038 410044 510040
rect 549884 510096 553367 510098
rect 549884 510040 553306 510096
rect 553362 510040 553367 510096
rect 549884 510038 553367 510040
rect 409045 510035 409111 510038
rect 553301 510035 553367 510038
rect 46105 509554 46171 509557
rect 46105 509552 48116 509554
rect 46105 509496 46110 509552
rect 46166 509496 48116 509552
rect 46105 509494 48116 509496
rect 46105 509491 46171 509494
rect 407297 509418 407363 509421
rect 407297 509416 410044 509418
rect 407297 509360 407302 509416
rect 407358 509360 410044 509416
rect 407297 509358 410044 509360
rect 407297 509355 407363 509358
rect 350441 508874 350507 508877
rect 347852 508872 350507 508874
rect 347852 508816 350446 508872
rect 350502 508816 350507 508872
rect 347852 508814 350507 508816
rect 350441 508811 350507 508814
rect 347822 507922 347882 508096
rect 407297 508058 407363 508061
rect 407297 508056 410044 508058
rect 407297 508000 407302 508056
rect 407358 508000 410044 508056
rect 407297 507998 410044 508000
rect 407297 507995 407363 507998
rect 350758 507922 350764 507924
rect 347822 507862 350764 507922
rect 350758 507860 350764 507862
rect 350828 507860 350834 507924
rect 46105 506970 46171 506973
rect 48086 506970 48146 507416
rect 46105 506968 48146 506970
rect 46105 506912 46110 506968
rect 46166 506912 48146 506968
rect 46105 506910 48146 506912
rect 347822 506970 347882 507416
rect 550265 507378 550331 507381
rect 549884 507376 550331 507378
rect 549884 507320 550270 507376
rect 550326 507320 550331 507376
rect 549884 507318 550331 507320
rect 550265 507315 550331 507318
rect 349981 506970 350047 506973
rect 347822 506968 350047 506970
rect 347822 506912 349986 506968
rect 350042 506912 350047 506968
rect 347822 506910 350047 506912
rect 46105 506907 46171 506910
rect 349981 506907 350047 506910
rect 407297 506698 407363 506701
rect 407297 506696 410044 506698
rect 407297 506640 407302 506696
rect 407358 506640 410044 506696
rect 407297 506638 410044 506640
rect 407297 506635 407363 506638
rect 347822 505610 347882 506056
rect 553301 506018 553367 506021
rect 549884 506016 553367 506018
rect 549884 505960 553306 506016
rect 553362 505960 553367 506016
rect 549884 505958 553367 505960
rect 553301 505955 553367 505958
rect 350073 505610 350139 505613
rect 347822 505608 350139 505610
rect 347822 505552 350078 505608
rect 350134 505552 350139 505608
rect 347822 505550 350139 505552
rect 350073 505547 350139 505550
rect 350441 505474 350507 505477
rect 347852 505472 350507 505474
rect 347852 505416 350446 505472
rect 350502 505416 350507 505472
rect 347852 505414 350507 505416
rect 350441 505411 350507 505414
rect 46105 505202 46171 505205
rect 48086 505202 48146 505376
rect 553117 505338 553183 505341
rect 549884 505336 553183 505338
rect 549884 505280 553122 505336
rect 553178 505280 553183 505336
rect 549884 505278 553183 505280
rect 553117 505275 553183 505278
rect 46105 505200 48146 505202
rect 46105 505144 46110 505200
rect 46166 505144 48146 505200
rect 46105 505142 48146 505144
rect 46105 505139 46171 505142
rect 553301 504658 553367 504661
rect 549884 504656 553367 504658
rect 549884 504600 553306 504656
rect 553362 504600 553367 504656
rect 549884 504598 553367 504600
rect 553301 504595 553367 504598
rect 47393 504114 47459 504117
rect 47393 504112 48116 504114
rect 47393 504056 47398 504112
rect 47454 504056 48116 504112
rect 47393 504054 48116 504056
rect 47393 504051 47459 504054
rect 347822 503842 347882 504016
rect 350441 503842 350507 503845
rect 347822 503840 350507 503842
rect 347822 503784 350446 503840
rect 350502 503784 350507 503840
rect 347822 503782 350507 503784
rect 350441 503779 350507 503782
rect 409462 502490 410044 502550
rect 549884 502490 550282 502550
rect 374494 502420 374500 502484
rect 374564 502482 374570 502484
rect 409462 502482 409522 502490
rect 374564 502422 409522 502482
rect 550222 502482 550282 502490
rect 553301 502482 553367 502485
rect 550222 502480 553367 502482
rect 550222 502424 553306 502480
rect 553362 502424 553367 502480
rect 550222 502422 553367 502424
rect 374564 502420 374570 502422
rect 553301 502419 553367 502422
rect 553117 501938 553183 501941
rect 549884 501936 553183 501938
rect -960 501802 480 501892
rect 549884 501880 553122 501936
rect 553178 501880 553183 501936
rect 549884 501878 553183 501880
rect 553117 501875 553183 501878
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 46105 501394 46171 501397
rect 46105 501392 48116 501394
rect 46105 501336 46110 501392
rect 46166 501336 48116 501392
rect 46105 501334 48116 501336
rect 46105 501331 46171 501334
rect 407297 501258 407363 501261
rect 553301 501258 553367 501261
rect 407297 501256 410044 501258
rect 407297 501200 407302 501256
rect 407358 501200 410044 501256
rect 407297 501198 410044 501200
rect 549884 501256 553367 501258
rect 549884 501200 553306 501256
rect 553362 501200 553367 501256
rect 549884 501198 553367 501200
rect 407297 501195 407363 501198
rect 553301 501195 553367 501198
rect 45645 500714 45711 500717
rect 45645 500712 48116 500714
rect 45645 500656 45650 500712
rect 45706 500656 48116 500712
rect 45645 500654 48116 500656
rect 45645 500651 45711 500654
rect 347822 500170 347882 500616
rect 407389 500578 407455 500581
rect 552381 500578 552447 500581
rect 407389 500576 410044 500578
rect 407389 500520 407394 500576
rect 407450 500520 410044 500576
rect 407389 500518 410044 500520
rect 549884 500576 552447 500578
rect 549884 500520 552386 500576
rect 552442 500520 552447 500576
rect 549884 500518 552447 500520
rect 407389 500515 407455 500518
rect 552381 500515 552447 500518
rect 350441 500170 350507 500173
rect 347822 500168 350507 500170
rect 347822 500112 350446 500168
rect 350502 500112 350507 500168
rect 347822 500110 350507 500112
rect 350441 500107 350507 500110
rect 349613 500034 349679 500037
rect 347852 500032 349679 500034
rect 347852 499976 349618 500032
rect 349674 499976 349679 500032
rect 347852 499974 349679 499976
rect 349613 499971 349679 499974
rect 32990 499700 32996 499764
rect 33060 499762 33066 499764
rect 48086 499762 48146 499936
rect 553301 499898 553367 499901
rect 549884 499896 553367 499898
rect 549884 499840 553306 499896
rect 553362 499840 553367 499896
rect 549884 499838 553367 499840
rect 553301 499835 553367 499838
rect 33060 499702 48146 499762
rect 33060 499700 33066 499702
rect 41270 498748 41276 498812
rect 41340 498810 41346 498812
rect 48086 498810 48146 499256
rect 41340 498750 48146 498810
rect 41340 498748 41346 498750
rect 347822 498266 347882 498576
rect 553301 498538 553367 498541
rect 549884 498536 553367 498538
rect 549884 498480 553306 498536
rect 553362 498480 553367 498536
rect 549884 498478 553367 498480
rect 553301 498475 553367 498478
rect 350441 498266 350507 498269
rect 347822 498264 350507 498266
rect 347822 498208 350446 498264
rect 350502 498208 350507 498264
rect 347822 498206 350507 498208
rect 350441 498203 350507 498206
rect 583520 497844 584960 498084
rect 46473 497314 46539 497317
rect 46473 497312 48116 497314
rect 46473 497256 46478 497312
rect 46534 497256 48116 497312
rect 46473 497254 48116 497256
rect 46473 497251 46539 497254
rect 385534 497116 385540 497180
rect 385604 497178 385610 497180
rect 550766 497178 550772 497180
rect 385604 497118 410044 497178
rect 549884 497118 550772 497178
rect 385604 497116 385610 497118
rect 550766 497116 550772 497118
rect 550836 497116 550842 497180
rect 46105 496090 46171 496093
rect 48086 496090 48146 496536
rect 552197 496498 552263 496501
rect 549884 496496 552263 496498
rect 549884 496440 552202 496496
rect 552258 496440 552263 496496
rect 549884 496438 552263 496440
rect 552197 496435 552263 496438
rect 46105 496088 48146 496090
rect 46105 496032 46110 496088
rect 46166 496032 48146 496088
rect 46105 496030 48146 496032
rect 46105 496027 46171 496030
rect 46473 495954 46539 495957
rect 46473 495952 48116 495954
rect 46473 495896 46478 495952
rect 46534 495896 48116 495952
rect 46473 495894 48116 495896
rect 46473 495891 46539 495894
rect 347822 495546 347882 495856
rect 407297 495818 407363 495821
rect 553301 495818 553367 495821
rect 407297 495816 410044 495818
rect 407297 495760 407302 495816
rect 407358 495760 410044 495816
rect 407297 495758 410044 495760
rect 549884 495816 553367 495818
rect 549884 495760 553306 495816
rect 553362 495760 553367 495816
rect 549884 495758 553367 495760
rect 407297 495755 407363 495758
rect 553301 495755 553367 495758
rect 350441 495546 350507 495549
rect 347822 495544 350507 495546
rect 347822 495488 350446 495544
rect 350502 495488 350507 495544
rect 347822 495486 350507 495488
rect 350441 495483 350507 495486
rect 46473 495274 46539 495277
rect 46473 495272 48116 495274
rect 46473 495216 46478 495272
rect 46534 495216 48116 495272
rect 46473 495214 48116 495216
rect 46473 495211 46539 495214
rect 45921 494594 45987 494597
rect 347822 494594 347882 495176
rect 350441 494594 350507 494597
rect 45921 494592 48116 494594
rect 45921 494536 45926 494592
rect 45982 494536 48116 494592
rect 45921 494534 48116 494536
rect 347822 494592 350507 494594
rect 347822 494536 350446 494592
rect 350502 494536 350507 494592
rect 347822 494534 350507 494536
rect 45921 494531 45987 494534
rect 350441 494531 350507 494534
rect 554814 494458 554820 494460
rect 549884 494398 554820 494458
rect 554814 494396 554820 494398
rect 554884 494396 554890 494460
rect 350349 493914 350415 493917
rect 347852 493912 350415 493914
rect 347852 493856 350354 493912
rect 350410 493856 350415 493912
rect 347852 493854 350415 493856
rect 350349 493851 350415 493854
rect 46473 493234 46539 493237
rect 48086 493234 48146 493816
rect 552565 493778 552631 493781
rect 549884 493776 552631 493778
rect 549884 493720 552570 493776
rect 552626 493720 552631 493776
rect 549884 493718 552631 493720
rect 552565 493715 552631 493718
rect 46473 493232 48146 493234
rect 46473 493176 46478 493232
rect 46534 493176 48146 493232
rect 46473 493174 48146 493176
rect 46473 493171 46539 493174
rect 407297 493098 407363 493101
rect 553117 493098 553183 493101
rect 407297 493096 410044 493098
rect 407297 493040 407302 493096
rect 407358 493040 410044 493096
rect 407297 493038 410044 493040
rect 549884 493096 553183 493098
rect 549884 493040 553122 493096
rect 553178 493040 553183 493096
rect 549884 493038 553183 493040
rect 407297 493035 407363 493038
rect 553117 493035 553183 493038
rect 347822 492010 347882 492456
rect 552473 492418 552539 492421
rect 549884 492416 552539 492418
rect 549884 492360 552478 492416
rect 552534 492360 552539 492416
rect 549884 492358 552539 492360
rect 552473 492355 552539 492358
rect 350349 492010 350415 492013
rect 347822 492008 350415 492010
rect 347822 491952 350354 492008
rect 350410 491952 350415 492008
rect 347822 491950 350415 491952
rect 350349 491947 350415 491950
rect 347822 491466 347882 491776
rect 553526 491738 553532 491740
rect 549884 491678 553532 491738
rect 553526 491676 553532 491678
rect 553596 491676 553602 491740
rect 350441 491466 350507 491469
rect 347822 491464 350507 491466
rect 347822 491408 350446 491464
rect 350502 491408 350507 491464
rect 347822 491406 350507 491408
rect 350441 491403 350507 491406
rect 41086 490588 41092 490652
rect 41156 490650 41162 490652
rect 48086 490650 48146 491096
rect 41156 490590 48146 490650
rect 347822 490650 347882 491096
rect 407297 491058 407363 491061
rect 407297 491056 410044 491058
rect 407297 491000 407302 491056
rect 407358 491000 410044 491056
rect 407297 490998 410044 491000
rect 407297 490995 407363 490998
rect 352046 490650 352052 490652
rect 347822 490590 352052 490650
rect 41156 490588 41162 490590
rect 352046 490588 352052 490590
rect 352116 490588 352122 490652
rect 46473 489970 46539 489973
rect 48086 489970 48146 490416
rect 347822 490106 347882 490416
rect 350441 490106 350507 490109
rect 347822 490104 350507 490106
rect 347822 490048 350446 490104
rect 350502 490048 350507 490104
rect 347822 490046 350507 490048
rect 350441 490043 350507 490046
rect 46473 489968 48146 489970
rect 46473 489912 46478 489968
rect 46534 489912 48146 489968
rect 46473 489910 48146 489912
rect 46473 489907 46539 489910
rect 46289 489834 46355 489837
rect 349153 489834 349219 489837
rect 46289 489832 48116 489834
rect 46289 489776 46294 489832
rect 46350 489776 48116 489832
rect 46289 489774 48116 489776
rect 347852 489832 349219 489834
rect 347852 489776 349158 489832
rect 349214 489776 349219 489832
rect 347852 489774 349219 489776
rect 46289 489771 46355 489774
rect 349153 489771 349219 489774
rect 407297 489698 407363 489701
rect 407297 489696 410044 489698
rect 407297 489640 407302 489696
rect 407358 489640 410044 489696
rect 407297 489638 410044 489640
rect 407297 489635 407363 489638
rect 407798 488956 407804 489020
rect 407868 489018 407874 489020
rect 553301 489018 553367 489021
rect 407868 488958 410044 489018
rect 549884 489016 553367 489018
rect 549884 488960 553306 489016
rect 553362 488960 553367 489016
rect 549884 488958 553367 488960
rect 407868 488956 407874 488958
rect 553301 488955 553367 488958
rect -960 488596 480 488836
rect 553301 488338 553367 488341
rect 549884 488336 553367 488338
rect 549884 488280 553306 488336
rect 553362 488280 553367 488336
rect 549884 488278 553367 488280
rect 553301 488275 553367 488278
rect 350441 487794 350507 487797
rect 347852 487792 350507 487794
rect 347852 487736 350446 487792
rect 350502 487736 350507 487792
rect 347852 487734 350507 487736
rect 350441 487731 350507 487734
rect 407297 487658 407363 487661
rect 407297 487656 410044 487658
rect 407297 487600 407302 487656
rect 407358 487600 410044 487656
rect 407297 487598 410044 487600
rect 407297 487595 407363 487598
rect 45134 486508 45140 486572
rect 45204 486570 45210 486572
rect 48086 486570 48146 487016
rect 407297 486978 407363 486981
rect 407297 486976 410044 486978
rect 407297 486920 407302 486976
rect 407358 486920 410044 486976
rect 407297 486918 410044 486920
rect 407297 486915 407363 486918
rect 45204 486510 48146 486570
rect 45204 486508 45210 486510
rect 46749 485890 46815 485893
rect 48086 485890 48146 486336
rect 46749 485888 48146 485890
rect 46749 485832 46754 485888
rect 46810 485832 48146 485888
rect 46749 485830 48146 485832
rect 46749 485827 46815 485830
rect 46749 485210 46815 485213
rect 48086 485210 48146 485656
rect 46749 485208 48146 485210
rect 46749 485152 46754 485208
rect 46810 485152 48146 485208
rect 46749 485150 48146 485152
rect 347822 485210 347882 485656
rect 407481 485618 407547 485621
rect 407481 485616 410044 485618
rect 407481 485560 407486 485616
rect 407542 485560 410044 485616
rect 407481 485558 410044 485560
rect 407481 485555 407547 485558
rect 349981 485210 350047 485213
rect 347822 485208 350047 485210
rect 347822 485152 349986 485208
rect 350042 485152 350047 485208
rect 347822 485150 350047 485152
rect 46749 485147 46815 485150
rect 349981 485147 350047 485150
rect 45829 484530 45895 484533
rect 48086 484530 48146 484976
rect 407297 484938 407363 484941
rect 552841 484938 552907 484941
rect 407297 484936 410044 484938
rect 407297 484880 407302 484936
rect 407358 484880 410044 484936
rect 407297 484878 410044 484880
rect 549884 484936 552907 484938
rect 549884 484880 552846 484936
rect 552902 484880 552907 484936
rect 549884 484878 552907 484880
rect 407297 484875 407363 484878
rect 552841 484875 552907 484878
rect 580349 484666 580415 484669
rect 583520 484666 584960 484756
rect 580349 484664 584960 484666
rect 580349 484608 580354 484664
rect 580410 484608 584960 484664
rect 580349 484606 584960 484608
rect 580349 484603 580415 484606
rect 45829 484528 48146 484530
rect 45829 484472 45834 484528
rect 45890 484472 48146 484528
rect 583520 484516 584960 484606
rect 45829 484470 48146 484472
rect 45829 484467 45895 484470
rect 407297 484258 407363 484261
rect 552565 484258 552631 484261
rect 407297 484256 410044 484258
rect 407297 484200 407302 484256
rect 407358 484200 410044 484256
rect 407297 484198 410044 484200
rect 549884 484256 552631 484258
rect 549884 484200 552570 484256
rect 552626 484200 552631 484256
rect 549884 484198 552631 484200
rect 407297 484195 407363 484198
rect 552565 484195 552631 484198
rect 37590 482972 37596 483036
rect 37660 483034 37666 483036
rect 48086 483034 48146 483616
rect 347822 483170 347882 483616
rect 407849 483578 407915 483581
rect 407849 483576 410044 483578
rect 407849 483520 407854 483576
rect 407910 483520 410044 483576
rect 407849 483518 410044 483520
rect 407849 483515 407915 483518
rect 350441 483170 350507 483173
rect 347822 483168 350507 483170
rect 347822 483112 350446 483168
rect 350502 483112 350507 483168
rect 347822 483110 350507 483112
rect 350441 483107 350507 483110
rect 349102 483034 349108 483036
rect 37660 482974 48146 483034
rect 347852 482974 349108 483034
rect 37660 482972 37666 482974
rect 349102 482972 349108 482974
rect 349172 482972 349178 483036
rect 46473 482354 46539 482357
rect 46473 482352 48116 482354
rect 46473 482296 46478 482352
rect 46534 482296 48116 482352
rect 46473 482294 48116 482296
rect 46473 482291 46539 482294
rect 407297 482218 407363 482221
rect 407297 482216 410044 482218
rect 407297 482160 407302 482216
rect 407358 482160 410044 482216
rect 407297 482158 410044 482160
rect 407297 482155 407363 482158
rect 350441 481674 350507 481677
rect 347852 481672 350507 481674
rect 347852 481616 350446 481672
rect 350502 481616 350507 481672
rect 347852 481614 350507 481616
rect 350441 481611 350507 481614
rect 46749 480586 46815 480589
rect 48086 480586 48146 480896
rect 347822 480722 347882 480896
rect 350073 480722 350139 480725
rect 347822 480720 350139 480722
rect 347822 480664 350078 480720
rect 350134 480664 350139 480720
rect 347822 480662 350139 480664
rect 350073 480659 350139 480662
rect 46749 480584 48146 480586
rect 46749 480528 46754 480584
rect 46810 480528 48146 480584
rect 46749 480526 48146 480528
rect 46749 480523 46815 480526
rect 46381 480314 46447 480317
rect 350441 480314 350507 480317
rect 46381 480312 48116 480314
rect 46381 480256 46386 480312
rect 46442 480256 48116 480312
rect 46381 480254 48116 480256
rect 347852 480312 350507 480314
rect 347852 480256 350446 480312
rect 350502 480256 350507 480312
rect 347852 480254 350507 480256
rect 46381 480251 46447 480254
rect 350441 480251 350507 480254
rect 392710 480116 392716 480180
rect 392780 480178 392786 480180
rect 552013 480178 552079 480181
rect 392780 480118 410044 480178
rect 549884 480176 552079 480178
rect 549884 480120 552018 480176
rect 552074 480120 552079 480176
rect 549884 480118 552079 480120
rect 392780 480116 392786 480118
rect 552013 480115 552079 480118
rect 409137 479498 409203 479501
rect 553301 479498 553367 479501
rect 409137 479496 410044 479498
rect 409137 479440 409142 479496
rect 409198 479440 410044 479496
rect 409137 479438 410044 479440
rect 549884 479496 553367 479498
rect 549884 479440 553306 479496
rect 553362 479440 553367 479496
rect 549884 479438 553367 479440
rect 409137 479435 409203 479438
rect 553301 479435 553367 479438
rect 552565 478818 552631 478821
rect 549884 478816 552631 478818
rect 549884 478760 552570 478816
rect 552626 478760 552631 478816
rect 549884 478758 552631 478760
rect 552565 478755 552631 478758
rect 407297 478138 407363 478141
rect 407297 478136 410044 478138
rect 407297 478080 407302 478136
rect 407358 478080 410044 478136
rect 407297 478078 410044 478080
rect 407297 478075 407363 478078
rect 347773 478002 347839 478005
rect 347773 478000 347882 478002
rect 347773 477944 347778 478000
rect 347834 477944 347882 478000
rect 347773 477939 347882 477944
rect 347822 477564 347882 477939
rect 39798 476308 39804 476372
rect 39868 476370 39874 476372
rect 48086 476370 48146 476816
rect 347822 476506 347882 476816
rect 409229 476778 409295 476781
rect 409229 476776 410044 476778
rect 409229 476720 409234 476776
rect 409290 476720 410044 476776
rect 409229 476718 410044 476720
rect 409229 476715 409295 476718
rect 350073 476506 350139 476509
rect 347822 476504 350139 476506
rect 347822 476448 350078 476504
rect 350134 476448 350139 476504
rect 347822 476446 350139 476448
rect 350073 476443 350139 476446
rect 39868 476310 48146 476370
rect 39868 476308 39874 476310
rect 43846 476172 43852 476236
rect 43916 476234 43922 476236
rect 350441 476234 350507 476237
rect 43916 476174 48116 476234
rect 347852 476232 350507 476234
rect 347852 476176 350446 476232
rect 350502 476176 350507 476232
rect 347852 476174 350507 476176
rect 43916 476172 43922 476174
rect 350441 476171 350507 476174
rect 408217 476234 408283 476237
rect 408534 476234 408540 476236
rect 408217 476232 408540 476234
rect 408217 476176 408222 476232
rect 408278 476176 408540 476232
rect 408217 476174 408540 476176
rect 408217 476171 408283 476174
rect 408534 476172 408540 476174
rect 408604 476172 408610 476236
rect 408217 476098 408283 476101
rect 552933 476098 552999 476101
rect 408217 476096 410044 476098
rect 408217 476040 408222 476096
rect 408278 476040 410044 476096
rect 408217 476038 410044 476040
rect 549884 476096 552999 476098
rect 549884 476040 552938 476096
rect 552994 476040 552999 476096
rect 549884 476038 552999 476040
rect 408217 476035 408283 476038
rect 552933 476035 552999 476038
rect -960 475540 480 475780
rect 46657 475554 46723 475557
rect 46657 475552 48116 475554
rect 46657 475496 46662 475552
rect 46718 475496 48116 475552
rect 46657 475494 48116 475496
rect 46657 475491 46723 475494
rect 347822 475013 347882 475456
rect 407297 475418 407363 475421
rect 553301 475418 553367 475421
rect 407297 475416 410044 475418
rect 407297 475360 407302 475416
rect 407358 475360 410044 475416
rect 407297 475358 410044 475360
rect 549884 475416 553367 475418
rect 549884 475360 553306 475416
rect 553362 475360 553367 475416
rect 549884 475358 553367 475360
rect 407297 475355 407363 475358
rect 553301 475355 553367 475358
rect 347773 475008 347882 475013
rect 347773 474952 347778 475008
rect 347834 474952 347882 475008
rect 347773 474950 347882 474952
rect 347773 474947 347839 474950
rect 407389 474738 407455 474741
rect 407389 474736 410044 474738
rect 407389 474680 407394 474736
rect 407450 474680 410044 474736
rect 407389 474678 410044 474680
rect 407389 474675 407455 474678
rect 46565 474194 46631 474197
rect 46565 474192 48116 474194
rect 46565 474136 46570 474192
rect 46626 474136 48116 474192
rect 46565 474134 48116 474136
rect 46565 474131 46631 474134
rect 407297 474058 407363 474061
rect 407297 474056 410044 474058
rect 407297 474000 407302 474056
rect 407358 474000 410044 474056
rect 407297 473998 410044 474000
rect 407297 473995 407363 473998
rect 46749 473514 46815 473517
rect 350441 473514 350507 473517
rect 46749 473512 48116 473514
rect 46749 473456 46754 473512
rect 46810 473456 48116 473512
rect 46749 473454 48116 473456
rect 347852 473512 350507 473514
rect 347852 473456 350446 473512
rect 350502 473456 350507 473512
rect 347852 473454 350507 473456
rect 46749 473451 46815 473454
rect 350441 473451 350507 473454
rect 347822 472290 347882 472736
rect 565302 472698 565308 472700
rect 549884 472638 565308 472698
rect 565302 472636 565308 472638
rect 565372 472636 565378 472700
rect 353702 472290 353708 472292
rect 347822 472230 353708 472290
rect 353702 472228 353708 472230
rect 353772 472228 353778 472292
rect 407297 472018 407363 472021
rect 407297 472016 410044 472018
rect 407297 471960 407302 472016
rect 407358 471960 410044 472016
rect 407297 471958 410044 471960
rect 407297 471955 407363 471958
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 35566 470868 35572 470932
rect 35636 470930 35642 470932
rect 48086 470930 48146 471376
rect 583520 471324 584960 471414
rect 35636 470870 48146 470930
rect 35636 470868 35642 470870
rect 349705 470794 349771 470797
rect 347852 470792 349771 470794
rect 347852 470736 349710 470792
rect 349766 470736 349771 470792
rect 347852 470734 349771 470736
rect 349705 470731 349771 470734
rect 553301 470658 553367 470661
rect 549884 470656 553367 470658
rect 549884 470600 553306 470656
rect 553362 470600 553367 470656
rect 549884 470598 553367 470600
rect 553301 470595 553367 470598
rect 46749 469706 46815 469709
rect 48086 469706 48146 470016
rect 407297 469978 407363 469981
rect 553301 469978 553367 469981
rect 407297 469976 410044 469978
rect 407297 469920 407302 469976
rect 407358 469920 410044 469976
rect 407297 469918 410044 469920
rect 549884 469976 553367 469978
rect 549884 469920 553306 469976
rect 553362 469920 553367 469976
rect 549884 469918 553367 469920
rect 407297 469915 407363 469918
rect 553301 469915 553367 469918
rect 46749 469704 48146 469706
rect 46749 469648 46754 469704
rect 46810 469648 48146 469704
rect 46749 469646 48146 469648
rect 46749 469643 46815 469646
rect 46657 468346 46723 468349
rect 48086 468346 48146 468656
rect 551001 468618 551067 468621
rect 550222 468616 551067 468618
rect 550222 468560 551006 468616
rect 551062 468560 551067 468616
rect 550222 468558 551067 468560
rect 550222 468550 550282 468558
rect 551001 468555 551067 468558
rect 46657 468344 48146 468346
rect 46657 468288 46662 468344
rect 46718 468288 48146 468344
rect 46657 468286 48146 468288
rect 46657 468283 46723 468286
rect 407297 468210 407363 468213
rect 410014 468210 410074 468520
rect 549884 468490 550282 468550
rect 407297 468208 410074 468210
rect 407297 468152 407302 468208
rect 407358 468152 410074 468208
rect 407297 468150 410074 468152
rect 407297 468147 407363 468150
rect 46749 468074 46815 468077
rect 46749 468072 48116 468074
rect 46749 468016 46754 468072
rect 46810 468016 48116 468072
rect 46749 468014 48116 468016
rect 46749 468011 46815 468014
rect 406837 467938 406903 467941
rect 406837 467936 410044 467938
rect 406837 467880 406842 467936
rect 406898 467880 410044 467936
rect 406837 467878 410044 467880
rect 406837 467875 406903 467878
rect 409229 467258 409295 467261
rect 409229 467256 410044 467258
rect 409229 467200 409234 467256
rect 409290 467200 410044 467256
rect 409229 467198 410044 467200
rect 409229 467195 409295 467198
rect 41638 466516 41644 466580
rect 41708 466578 41714 466580
rect 48086 466578 48146 466616
rect 41708 466518 48146 466578
rect 347822 466578 347882 466616
rect 350441 466578 350507 466581
rect 347822 466576 350507 466578
rect 347822 466520 350446 466576
rect 350502 466520 350507 466576
rect 347822 466518 350507 466520
rect 41708 466516 41714 466518
rect 350441 466515 350507 466518
rect 408350 466516 408356 466580
rect 408420 466578 408426 466580
rect 553301 466578 553367 466581
rect 408420 466518 410044 466578
rect 549884 466576 553367 466578
rect 549884 466520 553306 466576
rect 553362 466520 553367 466576
rect 549884 466518 553367 466520
rect 408420 466516 408426 466518
rect 553301 466515 553367 466518
rect 350073 466034 350139 466037
rect 347852 466032 350139 466034
rect 347852 465976 350078 466032
rect 350134 465976 350139 466032
rect 347852 465974 350139 465976
rect 350073 465971 350139 465974
rect 407297 465898 407363 465901
rect 552013 465898 552079 465901
rect 407297 465896 410044 465898
rect 407297 465840 407302 465896
rect 407358 465840 410044 465896
rect 407297 465838 410044 465840
rect 549884 465896 552079 465898
rect 549884 465840 552018 465896
rect 552074 465840 552079 465896
rect 549884 465838 552079 465840
rect 407297 465835 407363 465838
rect 552013 465835 552079 465838
rect 40902 465156 40908 465220
rect 40972 465218 40978 465220
rect 48086 465218 48146 465256
rect 40972 465158 48146 465218
rect 347822 465218 347882 465256
rect 350441 465218 350507 465221
rect 347822 465216 350507 465218
rect 347822 465160 350446 465216
rect 350502 465160 350507 465216
rect 347822 465158 350507 465160
rect 40972 465156 40978 465158
rect 350441 465155 350507 465158
rect 46749 464266 46815 464269
rect 48086 464266 48146 464576
rect 46749 464264 48146 464266
rect 46749 464208 46754 464264
rect 46810 464208 48146 464264
rect 46749 464206 48146 464208
rect 46749 464203 46815 464206
rect 347822 463994 347882 464576
rect 549884 464410 550282 464470
rect 550222 464402 550282 464410
rect 552013 464402 552079 464405
rect 550222 464400 552079 464402
rect 550222 464344 552018 464400
rect 552074 464344 552079 464400
rect 550222 464342 552079 464344
rect 552013 464339 552079 464342
rect 349102 463994 349108 463996
rect 347822 463934 349108 463994
rect 349102 463932 349108 463934
rect 349172 463932 349178 463996
rect 46749 463858 46815 463861
rect 48086 463858 48146 463896
rect 46749 463856 48146 463858
rect 46749 463800 46754 463856
rect 46810 463800 48146 463856
rect 46749 463798 48146 463800
rect 407297 463858 407363 463861
rect 407297 463856 410044 463858
rect 407297 463800 407302 463856
rect 407358 463800 410044 463856
rect 407297 463798 410044 463800
rect 46749 463795 46815 463798
rect 407297 463795 407363 463798
rect 46657 463314 46723 463317
rect 46657 463312 48116 463314
rect 46657 463256 46662 463312
rect 46718 463256 48116 463312
rect 46657 463254 48116 463256
rect 46657 463251 46723 463254
rect 347822 462906 347882 463216
rect 407389 463178 407455 463181
rect 552013 463178 552079 463181
rect 407389 463176 410044 463178
rect 407389 463120 407394 463176
rect 407450 463120 410044 463176
rect 407389 463118 410044 463120
rect 549884 463176 552079 463178
rect 549884 463120 552018 463176
rect 552074 463120 552079 463176
rect 549884 463118 552079 463120
rect 407389 463115 407455 463118
rect 552013 463115 552079 463118
rect 350073 462906 350139 462909
rect 347822 462904 350139 462906
rect 347822 462848 350078 462904
rect 350134 462848 350139 462904
rect 347822 462846 350139 462848
rect 350073 462843 350139 462846
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 347822 462498 347882 462536
rect 350441 462498 350507 462501
rect 347822 462496 350507 462498
rect 347822 462440 350446 462496
rect 350502 462440 350507 462496
rect 347822 462438 350507 462440
rect 350441 462435 350507 462438
rect 407297 462498 407363 462501
rect 407297 462496 410044 462498
rect 407297 462440 407302 462496
rect 407358 462440 410044 462496
rect 407297 462438 410044 462440
rect 407297 462435 407363 462438
rect 347822 461410 347882 461856
rect 355174 461756 355180 461820
rect 355244 461818 355250 461820
rect 355244 461758 410044 461818
rect 355244 461756 355250 461758
rect 350073 461410 350139 461413
rect 347822 461408 350139 461410
rect 347822 461352 350078 461408
rect 350134 461352 350139 461408
rect 347822 461350 350139 461352
rect 350073 461347 350139 461350
rect 46749 461002 46815 461005
rect 48086 461002 48146 461176
rect 347822 461138 347882 461176
rect 350441 461138 350507 461141
rect 347822 461136 350507 461138
rect 347822 461080 350446 461136
rect 350502 461080 350507 461136
rect 347822 461078 350507 461080
rect 350441 461075 350507 461078
rect 408125 461138 408191 461141
rect 408125 461136 410044 461138
rect 408125 461080 408130 461136
rect 408186 461080 410044 461136
rect 408125 461078 410044 461080
rect 408125 461075 408191 461078
rect 46749 461000 48146 461002
rect 46749 460944 46754 461000
rect 46810 460944 48146 461000
rect 46749 460942 48146 460944
rect 46749 460939 46815 460942
rect 552197 460458 552263 460461
rect 549884 460456 552263 460458
rect 549884 460400 552202 460456
rect 552258 460400 552263 460456
rect 549884 460398 552263 460400
rect 552197 460395 552263 460398
rect 46657 459914 46723 459917
rect 46657 459912 48116 459914
rect 46657 459856 46662 459912
rect 46718 459856 48116 459912
rect 46657 459854 48116 459856
rect 46657 459851 46723 459854
rect 347822 459642 347882 459816
rect 406469 459778 406535 459781
rect 552013 459778 552079 459781
rect 406469 459776 410044 459778
rect 406469 459720 406474 459776
rect 406530 459720 410044 459776
rect 406469 459718 410044 459720
rect 549884 459776 552079 459778
rect 549884 459720 552018 459776
rect 552074 459720 552079 459776
rect 549884 459718 552079 459720
rect 406469 459715 406535 459718
rect 552013 459715 552079 459718
rect 350441 459642 350507 459645
rect 347822 459640 350507 459642
rect 347822 459584 350446 459640
rect 350502 459584 350507 459640
rect 347822 459582 350507 459584
rect 350441 459579 350507 459582
rect 407297 459098 407363 459101
rect 552013 459098 552079 459101
rect 407297 459096 410044 459098
rect 407297 459040 407302 459096
rect 407358 459040 410044 459096
rect 407297 459038 410044 459040
rect 549884 459096 552079 459098
rect 549884 459040 552018 459096
rect 552074 459040 552079 459096
rect 549884 459038 552079 459040
rect 407297 459035 407363 459038
rect 552013 459035 552079 459038
rect 36670 458220 36676 458284
rect 36740 458282 36746 458284
rect 48086 458282 48146 458456
rect 36740 458222 48146 458282
rect 36740 458220 36746 458222
rect 583520 457996 584960 458236
rect 347822 457330 347882 457776
rect 408309 457738 408375 457741
rect 552013 457738 552079 457741
rect 408309 457736 410044 457738
rect 408309 457680 408314 457736
rect 408370 457680 410044 457736
rect 408309 457678 410044 457680
rect 549884 457736 552079 457738
rect 549884 457680 552018 457736
rect 552074 457680 552079 457736
rect 549884 457678 552079 457680
rect 408309 457675 408375 457678
rect 552013 457675 552079 457678
rect 350441 457330 350507 457333
rect 347822 457328 350507 457330
rect 347822 457272 350446 457328
rect 350502 457272 350507 457328
rect 347822 457270 350507 457272
rect 350441 457267 350507 457270
rect 43846 456860 43852 456924
rect 43916 456922 43922 456924
rect 48086 456922 48146 457096
rect 347822 457058 347882 457096
rect 364558 457058 364564 457060
rect 347822 456998 364564 457058
rect 364558 456996 364564 456998
rect 364628 456996 364634 457060
rect 407297 457058 407363 457061
rect 407297 457056 410044 457058
rect 407297 457000 407302 457056
rect 407358 457000 410044 457056
rect 407297 456998 410044 457000
rect 407297 456995 407363 456998
rect 43916 456862 48146 456922
rect 43916 456860 43922 456862
rect 348366 456860 348372 456924
rect 348436 456922 348442 456924
rect 349705 456922 349771 456925
rect 348436 456920 349771 456922
rect 348436 456864 349710 456920
rect 349766 456864 349771 456920
rect 348436 456862 349771 456864
rect 348436 456860 348442 456862
rect 349705 456859 349771 456862
rect 348366 456724 348372 456788
rect 348436 456786 348442 456788
rect 355409 456786 355475 456789
rect 348436 456784 355475 456786
rect 348436 456728 355414 456784
rect 355470 456728 355475 456784
rect 348436 456726 355475 456728
rect 348436 456724 348442 456726
rect 355409 456723 355475 456726
rect 46749 456514 46815 456517
rect 348233 456514 348299 456517
rect 46749 456512 48116 456514
rect 46749 456456 46754 456512
rect 46810 456456 48116 456512
rect 46749 456454 48116 456456
rect 347852 456512 348299 456514
rect 347852 456456 348238 456512
rect 348294 456456 348299 456512
rect 347852 456454 348299 456456
rect 46749 456451 46815 456454
rect 348233 456451 348299 456454
rect 552013 456378 552079 456381
rect 549884 456376 552079 456378
rect 549884 456320 552018 456376
rect 552074 456320 552079 456376
rect 549884 456318 552079 456320
rect 552013 456315 552079 456318
rect 46657 455834 46723 455837
rect 349797 455834 349863 455837
rect 46657 455832 48116 455834
rect 46657 455776 46662 455832
rect 46718 455776 48116 455832
rect 46657 455774 48116 455776
rect 347852 455832 349863 455834
rect 347852 455776 349802 455832
rect 349858 455776 349863 455832
rect 347852 455774 349863 455776
rect 46657 455771 46723 455774
rect 349797 455771 349863 455774
rect 407389 455698 407455 455701
rect 407389 455696 410044 455698
rect 407389 455640 407394 455696
rect 407450 455640 410044 455696
rect 407389 455638 410044 455640
rect 407389 455635 407455 455638
rect 407297 455018 407363 455021
rect 552473 455018 552539 455021
rect 407297 455016 410044 455018
rect 407297 454960 407302 455016
rect 407358 454960 410044 455016
rect 407297 454958 410044 454960
rect 549884 455016 552539 455018
rect 549884 454960 552478 455016
rect 552534 454960 552539 455016
rect 549884 454958 552539 454960
rect 407297 454955 407363 454958
rect 552473 454955 552539 454958
rect 347822 454202 347882 454376
rect 407389 454338 407455 454341
rect 552381 454338 552447 454341
rect 407389 454336 410044 454338
rect 407389 454280 407394 454336
rect 407450 454280 410044 454336
rect 407389 454278 410044 454280
rect 549884 454336 552447 454338
rect 549884 454280 552386 454336
rect 552442 454280 552447 454336
rect 549884 454278 552447 454280
rect 407389 454275 407455 454278
rect 552381 454275 552447 454278
rect 350441 454202 350507 454205
rect 347822 454200 350507 454202
rect 347822 454144 350446 454200
rect 350502 454144 350507 454200
rect 347822 454142 350507 454144
rect 350441 454139 350507 454142
rect 377438 453596 377444 453660
rect 377508 453658 377514 453660
rect 552565 453658 552631 453661
rect 377508 453598 410044 453658
rect 549884 453656 552631 453658
rect 549884 453600 552570 453656
rect 552626 453600 552631 453656
rect 549884 453598 552631 453600
rect 377508 453596 377514 453598
rect 552565 453595 552631 453598
rect 407665 452978 407731 452981
rect 407665 452976 410044 452978
rect 407665 452920 407670 452976
rect 407726 452920 410044 452976
rect 407665 452918 410044 452920
rect 407665 452915 407731 452918
rect 347822 451890 347882 452336
rect 350441 451890 350507 451893
rect 347822 451888 350507 451890
rect 347822 451832 350446 451888
rect 350502 451832 350507 451888
rect 347822 451830 350507 451832
rect 350441 451827 350507 451830
rect 349337 451754 349403 451757
rect 347852 451752 349403 451754
rect 347852 451696 349342 451752
rect 349398 451696 349403 451752
rect 347852 451694 349403 451696
rect 349337 451691 349403 451694
rect 407297 451618 407363 451621
rect 407297 451616 410044 451618
rect 407297 451560 407302 451616
rect 407358 451560 410044 451616
rect 407297 451558 410044 451560
rect 407297 451555 407363 451558
rect 549884 451490 550282 451550
rect 550222 451482 550282 451490
rect 552197 451482 552263 451485
rect 550222 451480 552263 451482
rect 550222 451424 552202 451480
rect 552258 451424 552263 451480
rect 550222 451422 552263 451424
rect 552197 451419 552263 451422
rect 350441 451074 350507 451077
rect 347852 451072 350507 451074
rect 347852 451016 350446 451072
rect 350502 451016 350507 451072
rect 347852 451014 350507 451016
rect 350441 451011 350507 451014
rect 39430 450468 39436 450532
rect 39500 450530 39506 450532
rect 48086 450530 48146 450976
rect 39500 450470 48146 450530
rect 39500 450468 39506 450470
rect 46749 450394 46815 450397
rect 46749 450392 48116 450394
rect 46749 450336 46754 450392
rect 46810 450336 48116 450392
rect 46749 450334 48116 450336
rect 46749 450331 46815 450334
rect 347822 449986 347882 450296
rect 561070 450258 561076 450260
rect 549884 450198 561076 450258
rect 561070 450196 561076 450198
rect 561140 450196 561146 450260
rect 350441 449986 350507 449989
rect 347822 449984 350507 449986
rect 347822 449928 350446 449984
rect 350502 449928 350507 449984
rect 347822 449926 350507 449928
rect 350441 449923 350507 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 43662 449108 43668 449172
rect 43732 449170 43738 449172
rect 48086 449170 48146 449616
rect 407297 449578 407363 449581
rect 553025 449578 553091 449581
rect 407297 449576 410044 449578
rect 407297 449520 407302 449576
rect 407358 449520 410044 449576
rect 407297 449518 410044 449520
rect 549884 449576 553091 449578
rect 549884 449520 553030 449576
rect 553086 449520 553091 449576
rect 549884 449518 553091 449520
rect 407297 449515 407363 449518
rect 553025 449515 553091 449518
rect 43732 449110 48146 449170
rect 43732 449108 43738 449110
rect 553301 448898 553367 448901
rect 549884 448896 553367 448898
rect 549884 448840 553306 448896
rect 553362 448840 553367 448896
rect 549884 448838 553367 448840
rect 553301 448835 553367 448838
rect 347822 447810 347882 448256
rect 350441 447810 350507 447813
rect 347822 447808 350507 447810
rect 347822 447752 350446 447808
rect 350502 447752 350507 447808
rect 347822 447750 350507 447752
rect 350441 447747 350507 447750
rect 407297 447266 407363 447269
rect 410014 447266 410074 447440
rect 407297 447264 410074 447266
rect 407297 447208 407302 447264
rect 407358 447208 410074 447264
rect 407297 447206 410074 447208
rect 407297 447203 407363 447206
rect 347822 446450 347882 446896
rect 552381 446858 552447 446861
rect 549884 446856 552447 446858
rect 549884 446800 552386 446856
rect 552442 446800 552447 446856
rect 549884 446798 552447 446800
rect 552381 446795 552447 446798
rect 350441 446450 350507 446453
rect 347822 446448 350507 446450
rect 347822 446392 350446 446448
rect 350502 446392 350507 446448
rect 347822 446390 350507 446392
rect 350441 446387 350507 446390
rect 46473 446042 46539 446045
rect 48086 446042 48146 446216
rect 46473 446040 48146 446042
rect 46473 445984 46478 446040
rect 46534 445984 48146 446040
rect 46473 445982 48146 445984
rect 46473 445979 46539 445982
rect 347822 445906 347882 446216
rect 407389 446178 407455 446181
rect 407389 446176 410044 446178
rect 407389 446120 407394 446176
rect 407450 446120 410044 446176
rect 407389 446118 410044 446120
rect 407389 446115 407455 446118
rect 350073 445906 350139 445909
rect 347822 445904 350139 445906
rect 347822 445848 350078 445904
rect 350134 445848 350139 445904
rect 347822 445846 350139 445848
rect 350073 445843 350139 445846
rect 350441 445634 350507 445637
rect 347852 445632 350507 445634
rect 347852 445576 350446 445632
rect 350502 445576 350507 445632
rect 347852 445574 350507 445576
rect 350441 445571 350507 445574
rect 45921 445090 45987 445093
rect 48086 445090 48146 445536
rect 552565 445498 552631 445501
rect 549884 445496 552631 445498
rect 549884 445440 552570 445496
rect 552626 445440 552631 445496
rect 549884 445438 552631 445440
rect 552565 445435 552631 445438
rect 45921 445088 48146 445090
rect 45921 445032 45926 445088
rect 45982 445032 48146 445088
rect 45921 445030 48146 445032
rect 45921 445027 45987 445030
rect 407297 444818 407363 444821
rect 407297 444816 410044 444818
rect 407297 444760 407302 444816
rect 407358 444760 410044 444816
rect 407297 444758 410044 444760
rect 407297 444755 407363 444758
rect 583520 444668 584960 444908
rect 46749 443322 46815 443325
rect 48086 443322 48146 443496
rect 553301 443458 553367 443461
rect 549884 443456 553367 443458
rect 549884 443400 553306 443456
rect 553362 443400 553367 443456
rect 549884 443398 553367 443400
rect 553301 443395 553367 443398
rect 46749 443320 48146 443322
rect 46749 443264 46754 443320
rect 46810 443264 48146 443320
rect 46749 443262 48146 443264
rect 46749 443259 46815 443262
rect 46565 442914 46631 442917
rect 46565 442912 48116 442914
rect 46565 442856 46570 442912
rect 46626 442856 48116 442912
rect 46565 442854 48116 442856
rect 46565 442851 46631 442854
rect 347822 441690 347882 442136
rect 407297 442098 407363 442101
rect 407297 442096 410044 442098
rect 407297 442040 407302 442096
rect 407358 442040 410044 442096
rect 407297 442038 410044 442040
rect 407297 442035 407363 442038
rect 350441 441690 350507 441693
rect 347822 441688 350507 441690
rect 347822 441632 350446 441688
rect 350502 441632 350507 441688
rect 347822 441630 350507 441632
rect 350441 441627 350507 441630
rect 407389 441418 407455 441421
rect 551502 441418 551508 441420
rect 407389 441416 410044 441418
rect 407389 441360 407394 441416
rect 407450 441360 410044 441416
rect 407389 441358 410044 441360
rect 549884 441358 551508 441418
rect 407389 441355 407455 441358
rect 551502 441356 551508 441358
rect 551572 441356 551578 441420
rect 347822 440330 347882 440776
rect 550214 440738 550220 440740
rect 549884 440678 550220 440738
rect 550214 440676 550220 440678
rect 550284 440676 550290 440740
rect 350441 440330 350507 440333
rect 347822 440328 350507 440330
rect 347822 440272 350446 440328
rect 350502 440272 350507 440328
rect 347822 440270 350507 440272
rect 350441 440267 350507 440270
rect 45921 439650 45987 439653
rect 48086 439650 48146 440096
rect 407205 440058 407271 440061
rect 407205 440056 410044 440058
rect 407205 440000 407210 440056
rect 407266 440000 410044 440056
rect 407205 439998 410044 440000
rect 407205 439995 407271 439998
rect 45921 439648 48146 439650
rect 45921 439592 45926 439648
rect 45982 439592 48146 439648
rect 45921 439590 48146 439592
rect 45921 439587 45987 439590
rect 40718 438908 40724 438972
rect 40788 438970 40794 438972
rect 48086 438970 48146 439416
rect 40788 438910 48146 438970
rect 40788 438908 40794 438910
rect 46289 438834 46355 438837
rect 46289 438832 48116 438834
rect 46289 438776 46294 438832
rect 46350 438776 48116 438832
rect 46289 438774 48116 438776
rect 46289 438771 46355 438774
rect 407481 438698 407547 438701
rect 553301 438698 553367 438701
rect 407481 438696 410044 438698
rect 407481 438640 407486 438696
rect 407542 438640 410044 438696
rect 407481 438638 410044 438640
rect 549884 438696 553367 438698
rect 549884 438640 553306 438696
rect 553362 438640 553367 438696
rect 549884 438638 553367 438640
rect 407481 438635 407547 438638
rect 553301 438635 553367 438638
rect 347822 437882 347882 438056
rect 407205 438018 407271 438021
rect 553301 438018 553367 438021
rect 407205 438016 410044 438018
rect 407205 437960 407210 438016
rect 407266 437960 410044 438016
rect 407205 437958 410044 437960
rect 549884 438016 553367 438018
rect 549884 437960 553306 438016
rect 553362 437960 553367 438016
rect 549884 437958 553367 437960
rect 407205 437955 407271 437958
rect 553301 437955 553367 437958
rect 350073 437882 350139 437885
rect 347822 437880 350139 437882
rect 347822 437824 350078 437880
rect 350134 437824 350139 437880
rect 347822 437822 350139 437824
rect 350073 437819 350139 437822
rect 407205 437338 407271 437341
rect 552657 437338 552723 437341
rect 407205 437336 410044 437338
rect 407205 437280 407210 437336
rect 407266 437280 410044 437336
rect 407205 437278 410044 437280
rect 549884 437336 552723 437338
rect 549884 437280 552662 437336
rect 552718 437280 552723 437336
rect 549884 437278 552723 437280
rect 407205 437275 407271 437278
rect 552657 437275 552723 437278
rect 350441 436794 350507 436797
rect 347852 436792 350507 436794
rect -960 436508 480 436748
rect 347852 436736 350446 436792
rect 350502 436736 350507 436792
rect 347852 436734 350507 436736
rect 350441 436731 350507 436734
rect 46749 436522 46815 436525
rect 48086 436522 48146 436696
rect 553301 436658 553367 436661
rect 549884 436656 553367 436658
rect 549884 436600 553306 436656
rect 553362 436600 553367 436656
rect 549884 436598 553367 436600
rect 553301 436595 553367 436598
rect 46749 436520 48146 436522
rect 46749 436464 46754 436520
rect 46810 436464 48146 436520
rect 46749 436462 48146 436464
rect 46749 436459 46815 436462
rect 407205 435978 407271 435981
rect 552657 435978 552723 435981
rect 407205 435976 410044 435978
rect 407205 435920 407210 435976
rect 407266 435920 410044 435976
rect 407205 435918 410044 435920
rect 549884 435976 552723 435978
rect 549884 435920 552662 435976
rect 552718 435920 552723 435976
rect 549884 435918 552723 435920
rect 407205 435915 407271 435918
rect 552657 435915 552723 435918
rect 347822 434890 347882 435336
rect 349654 434890 349660 434892
rect 347822 434830 349660 434890
rect 349654 434828 349660 434830
rect 349724 434828 349730 434892
rect 46749 434754 46815 434757
rect 350441 434754 350507 434757
rect 46749 434752 48116 434754
rect 46749 434696 46754 434752
rect 46810 434696 48116 434752
rect 46749 434694 48116 434696
rect 347852 434752 350507 434754
rect 347852 434696 350446 434752
rect 350502 434696 350507 434752
rect 347852 434694 350507 434696
rect 46749 434691 46815 434694
rect 350441 434691 350507 434694
rect 407297 434618 407363 434621
rect 407297 434616 410044 434618
rect 407297 434560 407302 434616
rect 407358 434560 410044 434616
rect 407297 434558 410044 434560
rect 407297 434555 407363 434558
rect 46749 433666 46815 433669
rect 48086 433666 48146 433976
rect 408401 433938 408467 433941
rect 408401 433936 410044 433938
rect 408401 433880 408406 433936
rect 408462 433880 410044 433936
rect 408401 433878 410044 433880
rect 408401 433875 408467 433878
rect 46749 433664 48146 433666
rect 46749 433608 46754 433664
rect 46810 433608 48146 433664
rect 46749 433606 48146 433608
rect 46749 433603 46815 433606
rect 348141 433394 348207 433397
rect 347852 433392 348207 433394
rect 347852 433336 348146 433392
rect 348202 433336 348207 433392
rect 347852 433334 348207 433336
rect 348141 433331 348207 433334
rect 348877 433258 348943 433261
rect 349286 433258 349292 433260
rect 348877 433256 349292 433258
rect 348877 433200 348882 433256
rect 348938 433200 349292 433256
rect 348877 433198 349292 433200
rect 348877 433195 348943 433198
rect 349286 433196 349292 433198
rect 349356 433196 349362 433260
rect 407205 433258 407271 433261
rect 407205 433256 410044 433258
rect 407205 433200 407210 433256
rect 407266 433200 410044 433256
rect 407205 433198 410044 433200
rect 407205 433195 407271 433198
rect 46381 432034 46447 432037
rect 48086 432034 48146 432616
rect 552197 432578 552263 432581
rect 549884 432576 552263 432578
rect 549884 432520 552202 432576
rect 552258 432520 552263 432576
rect 549884 432518 552263 432520
rect 552197 432515 552263 432518
rect 46381 432032 48146 432034
rect 46381 431976 46386 432032
rect 46442 431976 48146 432032
rect 46381 431974 48146 431976
rect 46381 431971 46447 431974
rect 550909 431898 550975 431901
rect 549884 431896 550975 431898
rect 549884 431840 550914 431896
rect 550970 431840 550975 431896
rect 549884 431838 550975 431840
rect 550909 431835 550975 431838
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 347822 430946 347882 431256
rect 350073 430946 350139 430949
rect 347822 430944 350139 430946
rect 347822 430888 350078 430944
rect 350134 430888 350139 430944
rect 347822 430886 350139 430888
rect 350073 430883 350139 430886
rect 350441 430674 350507 430677
rect 347852 430672 350507 430674
rect 347852 430616 350446 430672
rect 350502 430616 350507 430672
rect 347852 430614 350507 430616
rect 350441 430611 350507 430614
rect 409321 430538 409387 430541
rect 409321 430536 410044 430538
rect 409321 430480 409326 430536
rect 409382 430480 410044 430536
rect 409321 430478 410044 430480
rect 409321 430475 409387 430478
rect 46381 429994 46447 429997
rect 46381 429992 48116 429994
rect 46381 429936 46386 429992
rect 46442 429936 48116 429992
rect 46381 429934 48116 429936
rect 46381 429931 46447 429934
rect 406469 429858 406535 429861
rect 553485 429858 553551 429861
rect 406469 429856 410044 429858
rect 406469 429800 406474 429856
rect 406530 429800 410044 429856
rect 406469 429798 410044 429800
rect 549884 429856 553551 429858
rect 549884 429800 553490 429856
rect 553546 429800 553551 429856
rect 549884 429798 553551 429800
rect 406469 429795 406535 429798
rect 553485 429795 553551 429798
rect 46749 429314 46815 429317
rect 46749 429312 48116 429314
rect 46749 429256 46754 429312
rect 46810 429256 48116 429312
rect 46749 429254 48116 429256
rect 46749 429251 46815 429254
rect 407205 429178 407271 429181
rect 407205 429176 410044 429178
rect 407205 429120 407210 429176
rect 407266 429120 410044 429176
rect 407205 429118 410044 429120
rect 407205 429115 407271 429118
rect 47526 428504 47532 428568
rect 47596 428566 47602 428568
rect 47596 428506 48116 428566
rect 47596 428504 47602 428506
rect 409413 428498 409479 428501
rect 552841 428498 552907 428501
rect 409413 428496 410044 428498
rect 409413 428440 409418 428496
rect 409474 428440 410044 428496
rect 409413 428438 410044 428440
rect 549884 428496 552907 428498
rect 549884 428440 552846 428496
rect 552902 428440 552907 428496
rect 549884 428438 552907 428440
rect 409413 428435 409479 428438
rect 552841 428435 552907 428438
rect 46749 427954 46815 427957
rect 350441 427954 350507 427957
rect 46749 427952 48116 427954
rect 46749 427896 46754 427952
rect 46810 427896 48116 427952
rect 46749 427894 48116 427896
rect 347852 427952 350507 427954
rect 347852 427896 350446 427952
rect 350502 427896 350507 427952
rect 347852 427894 350507 427896
rect 46749 427891 46815 427894
rect 350441 427891 350507 427894
rect 407297 427818 407363 427821
rect 407297 427816 410044 427818
rect 407297 427760 407302 427816
rect 407358 427760 410044 427816
rect 407297 427758 410044 427760
rect 407297 427755 407363 427758
rect 407205 427138 407271 427141
rect 407205 427136 410044 427138
rect 407205 427080 407210 427136
rect 407266 427080 410044 427136
rect 407205 427078 410044 427080
rect 407205 427075 407271 427078
rect 350441 426594 350507 426597
rect 347852 426592 350507 426594
rect 347852 426536 350446 426592
rect 350502 426536 350507 426592
rect 347852 426534 350507 426536
rect 350441 426531 350507 426534
rect 553025 426458 553091 426461
rect 549884 426456 553091 426458
rect 549884 426400 553030 426456
rect 553086 426400 553091 426456
rect 549884 426398 553091 426400
rect 553025 426395 553091 426398
rect 46565 425370 46631 425373
rect 48086 425370 48146 425816
rect 46565 425368 48146 425370
rect 46565 425312 46570 425368
rect 46626 425312 48146 425368
rect 46565 425310 48146 425312
rect 347822 425370 347882 425816
rect 407205 425778 407271 425781
rect 407205 425776 410044 425778
rect 407205 425720 407210 425776
rect 407266 425720 410044 425776
rect 407205 425718 410044 425720
rect 407205 425715 407271 425718
rect 350441 425370 350507 425373
rect 347822 425368 350507 425370
rect 347822 425312 350446 425368
rect 350502 425312 350507 425368
rect 347822 425310 350507 425312
rect 46565 425307 46631 425310
rect 350441 425307 350507 425310
rect 46749 425234 46815 425237
rect 46749 425232 48116 425234
rect 46749 425176 46754 425232
rect 46810 425176 48116 425232
rect 46749 425174 48116 425176
rect 46749 425171 46815 425174
rect 553025 425098 553091 425101
rect 549884 425096 553091 425098
rect 549884 425040 553030 425096
rect 553086 425040 553091 425096
rect 549884 425038 553091 425040
rect 553025 425035 553091 425038
rect 46657 424554 46723 424557
rect 46657 424552 48116 424554
rect 46657 424496 46662 424552
rect 46718 424496 48116 424552
rect 46657 424494 48116 424496
rect 46657 424491 46723 424494
rect 552933 424418 552999 424421
rect 549884 424416 552999 424418
rect 549884 424360 552938 424416
rect 552994 424360 552999 424416
rect 549884 424358 552999 424360
rect 552933 424355 552999 424358
rect 46749 423738 46815 423741
rect 48086 423738 48146 423776
rect 46749 423736 48146 423738
rect -960 423452 480 423692
rect 46749 423680 46754 423736
rect 46810 423680 48146 423736
rect 46749 423678 48146 423680
rect 407205 423738 407271 423741
rect 553025 423738 553091 423741
rect 407205 423736 410044 423738
rect 407205 423680 407210 423736
rect 407266 423680 410044 423736
rect 407205 423678 410044 423680
rect 549884 423736 553091 423738
rect 549884 423680 553030 423736
rect 553086 423680 553091 423736
rect 549884 423678 553091 423680
rect 46749 423675 46815 423678
rect 407205 423675 407271 423678
rect 553025 423675 553091 423678
rect 407205 423058 407271 423061
rect 407205 423056 410044 423058
rect 407205 423000 407210 423056
rect 407266 423000 410044 423056
rect 407205 422998 410044 423000
rect 407205 422995 407271 422998
rect 347822 422378 347882 422416
rect 350441 422378 350507 422381
rect 551001 422378 551067 422381
rect 347822 422376 350507 422378
rect 347822 422320 350446 422376
rect 350502 422320 350507 422376
rect 347822 422318 350507 422320
rect 549884 422376 551067 422378
rect 549884 422320 551006 422376
rect 551062 422320 551067 422376
rect 549884 422318 551067 422320
rect 350441 422315 350507 422318
rect 551001 422315 551067 422318
rect 46473 421290 46539 421293
rect 48086 421290 48146 421736
rect 46473 421288 48146 421290
rect 46473 421232 46478 421288
rect 46534 421232 48146 421288
rect 46473 421230 48146 421232
rect 347822 421290 347882 421736
rect 408309 421698 408375 421701
rect 552289 421698 552355 421701
rect 408309 421696 410044 421698
rect 408309 421640 408314 421696
rect 408370 421640 410044 421696
rect 408309 421638 410044 421640
rect 549884 421696 552355 421698
rect 549884 421640 552294 421696
rect 552350 421640 552355 421696
rect 549884 421638 552355 421640
rect 408309 421635 408375 421638
rect 552289 421635 552355 421638
rect 350073 421290 350139 421293
rect 347822 421288 350139 421290
rect 347822 421232 350078 421288
rect 350134 421232 350139 421288
rect 347822 421230 350139 421232
rect 46473 421227 46539 421230
rect 350073 421227 350139 421230
rect 46749 421018 46815 421021
rect 48086 421018 48146 421056
rect 46749 421016 48146 421018
rect 46749 420960 46754 421016
rect 46810 420960 48146 421016
rect 46749 420958 48146 420960
rect 347822 421018 347882 421056
rect 350441 421018 350507 421021
rect 552289 421018 552355 421021
rect 347822 421016 350507 421018
rect 347822 420960 350446 421016
rect 350502 420960 350507 421016
rect 347822 420958 350507 420960
rect 549884 421016 552355 421018
rect 549884 420960 552294 421016
rect 552350 420960 552355 421016
rect 549884 420958 552355 420960
rect 46749 420955 46815 420958
rect 350441 420955 350507 420958
rect 552289 420955 552355 420958
rect 46657 420066 46723 420069
rect 48086 420066 48146 420376
rect 407297 420338 407363 420341
rect 553025 420338 553091 420341
rect 407297 420336 410044 420338
rect 407297 420280 407302 420336
rect 407358 420280 410044 420336
rect 407297 420278 410044 420280
rect 549884 420336 553091 420338
rect 549884 420280 553030 420336
rect 553086 420280 553091 420336
rect 549884 420278 553091 420280
rect 407297 420275 407363 420278
rect 553025 420275 553091 420278
rect 46657 420064 48146 420066
rect 46657 420008 46662 420064
rect 46718 420008 48146 420064
rect 46657 420006 48146 420008
rect 46657 420003 46723 420006
rect 46749 419658 46815 419661
rect 48086 419658 48146 419696
rect 46749 419656 48146 419658
rect 46749 419600 46754 419656
rect 46810 419600 48146 419656
rect 46749 419598 48146 419600
rect 347822 419658 347882 419696
rect 350441 419658 350507 419661
rect 347822 419656 350507 419658
rect 347822 419600 350446 419656
rect 350502 419600 350507 419656
rect 347822 419598 350507 419600
rect 46749 419595 46815 419598
rect 350441 419595 350507 419598
rect 407205 419658 407271 419661
rect 407205 419656 410044 419658
rect 407205 419600 407210 419656
rect 407266 419600 410044 419656
rect 407205 419598 410044 419600
rect 407205 419595 407271 419598
rect 46657 418706 46723 418709
rect 48086 418706 48146 419016
rect 46657 418704 48146 418706
rect 46657 418648 46662 418704
rect 46718 418648 48146 418704
rect 46657 418646 48146 418648
rect 46657 418643 46723 418646
rect 347822 418434 347882 419016
rect 407205 418978 407271 418981
rect 407205 418976 410044 418978
rect 407205 418920 407210 418976
rect 407266 418920 410044 418976
rect 407205 418918 410044 418920
rect 407205 418915 407271 418918
rect 350441 418434 350507 418437
rect 347822 418432 350507 418434
rect 347822 418376 350446 418432
rect 350502 418376 350507 418432
rect 347822 418374 350507 418376
rect 350441 418371 350507 418374
rect 46749 418298 46815 418301
rect 48086 418298 48146 418336
rect 46749 418296 48146 418298
rect 46749 418240 46754 418296
rect 46810 418240 48146 418296
rect 46749 418238 48146 418240
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 46749 418235 46815 418238
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect 347822 416938 347882 416976
rect 350441 416938 350507 416941
rect 347822 416936 350507 416938
rect 347822 416880 350446 416936
rect 350502 416880 350507 416936
rect 347822 416878 350507 416880
rect 350441 416875 350507 416878
rect 46657 415986 46723 415989
rect 48086 415986 48146 416296
rect 407573 416258 407639 416261
rect 552013 416258 552079 416261
rect 407573 416256 410044 416258
rect 407573 416200 407578 416256
rect 407634 416200 410044 416256
rect 407573 416198 410044 416200
rect 549884 416256 552079 416258
rect 549884 416200 552018 416256
rect 552074 416200 552079 416256
rect 549884 416198 552079 416200
rect 407573 416195 407639 416198
rect 552013 416195 552079 416198
rect 46657 415984 48146 415986
rect 46657 415928 46662 415984
rect 46718 415928 48146 415984
rect 46657 415926 48146 415928
rect 46657 415923 46723 415926
rect 46749 415578 46815 415581
rect 48086 415578 48146 415616
rect 552013 415578 552079 415581
rect 46749 415576 48146 415578
rect 46749 415520 46754 415576
rect 46810 415520 48146 415576
rect 46749 415518 48146 415520
rect 549884 415576 552079 415578
rect 549884 415520 552018 415576
rect 552074 415520 552079 415576
rect 549884 415518 552079 415520
rect 46749 415515 46815 415518
rect 552013 415515 552079 415518
rect 347822 414490 347882 414936
rect 407205 414898 407271 414901
rect 407205 414896 410044 414898
rect 407205 414840 407210 414896
rect 407266 414840 410044 414896
rect 407205 414838 410044 414840
rect 407205 414835 407271 414838
rect 350441 414490 350507 414493
rect 347822 414488 350507 414490
rect 347822 414432 350446 414488
rect 350502 414432 350507 414488
rect 347822 414430 350507 414432
rect 350441 414427 350507 414430
rect 46749 414082 46815 414085
rect 48086 414082 48146 414256
rect 46749 414080 48146 414082
rect 46749 414024 46754 414080
rect 46810 414024 48146 414080
rect 46749 414022 48146 414024
rect 347822 414082 347882 414256
rect 350441 414082 350507 414085
rect 347822 414080 350507 414082
rect 347822 414024 350446 414080
rect 350502 414024 350507 414080
rect 347822 414022 350507 414024
rect 46749 414019 46815 414022
rect 350441 414019 350507 414022
rect 549884 413410 550466 413470
rect 550406 413402 550466 413410
rect 552197 413402 552263 413405
rect 550406 413400 552263 413402
rect 550406 413344 552202 413400
rect 552258 413344 552263 413400
rect 550406 413342 552263 413344
rect 552197 413339 552263 413342
rect 46238 412932 46244 412996
rect 46308 412994 46314 412996
rect 46308 412934 48116 412994
rect 46308 412932 46314 412934
rect 552013 412858 552079 412861
rect 549884 412856 552079 412858
rect 549884 412800 552018 412856
rect 552074 412800 552079 412856
rect 549884 412798 552079 412800
rect 552013 412795 552079 412798
rect 407297 412178 407363 412181
rect 407297 412176 410044 412178
rect 407297 412120 407302 412176
rect 407358 412120 410044 412176
rect 407297 412118 410044 412120
rect 407297 412115 407363 412118
rect 46565 411362 46631 411365
rect 48086 411362 48146 411536
rect 46565 411360 48146 411362
rect 46565 411304 46570 411360
rect 46626 411304 48146 411360
rect 46565 411302 48146 411304
rect 347822 411362 347882 411536
rect 407205 411498 407271 411501
rect 407205 411496 410044 411498
rect 407205 411440 407210 411496
rect 407266 411440 410044 411496
rect 407205 411438 410044 411440
rect 407205 411435 407271 411438
rect 350441 411362 350507 411365
rect 347822 411360 350507 411362
rect 347822 411304 350446 411360
rect 350502 411304 350507 411360
rect 347822 411302 350507 411304
rect 46565 411299 46631 411302
rect 350441 411299 350507 411302
rect 347814 411164 347820 411228
rect 347884 411164 347890 411228
rect 347822 410924 347882 411164
rect 407205 410818 407271 410821
rect 567510 410818 567516 410820
rect 407205 410816 410044 410818
rect 407205 410760 407210 410816
rect 407266 410760 410044 410816
rect 407205 410758 410044 410760
rect 549884 410758 567516 410818
rect 407205 410755 407271 410758
rect 567510 410756 567516 410758
rect 567580 410756 567586 410820
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 349521 409594 349587 409597
rect 347852 409592 349587 409594
rect 347852 409536 349526 409592
rect 349582 409536 349587 409592
rect 347852 409534 349587 409536
rect 349521 409531 349587 409534
rect 408125 408778 408191 408781
rect 408125 408776 410044 408778
rect 408125 408720 408130 408776
rect 408186 408720 410044 408776
rect 408125 408718 410044 408720
rect 408125 408715 408191 408718
rect 46565 407690 46631 407693
rect 48086 407690 48146 408136
rect 46565 407688 48146 407690
rect 46565 407632 46570 407688
rect 46626 407632 48146 407688
rect 46565 407630 48146 407632
rect 46565 407627 46631 407630
rect 347822 407282 347882 407456
rect 407205 407418 407271 407421
rect 550909 407418 550975 407421
rect 407205 407416 410044 407418
rect 407205 407360 407210 407416
rect 407266 407360 410044 407416
rect 407205 407358 410044 407360
rect 549884 407416 550975 407418
rect 549884 407360 550914 407416
rect 550970 407360 550975 407416
rect 549884 407358 550975 407360
rect 407205 407355 407271 407358
rect 550909 407355 550975 407358
rect 350441 407282 350507 407285
rect 347822 407280 350507 407282
rect 347822 407224 350446 407280
rect 350502 407224 350507 407280
rect 347822 407222 350507 407224
rect 350441 407219 350507 407222
rect 407205 406058 407271 406061
rect 407205 406056 410044 406058
rect 407205 406000 407210 406056
rect 407266 406000 410044 406056
rect 407205 405998 410044 406000
rect 407205 405995 407271 405998
rect 347822 404970 347882 405416
rect 552933 405378 552999 405381
rect 549884 405376 552999 405378
rect 549884 405320 552938 405376
rect 552994 405320 552999 405376
rect 549884 405318 552999 405320
rect 552933 405315 552999 405318
rect 350073 404970 350139 404973
rect 347822 404968 350139 404970
rect 347822 404912 350078 404968
rect 350134 404912 350139 404968
rect 347822 404910 350139 404912
rect 350073 404907 350139 404910
rect 583520 404820 584960 405060
rect 347822 404562 347882 404736
rect 407297 404698 407363 404701
rect 554998 404698 555004 404700
rect 407297 404696 410044 404698
rect 407297 404640 407302 404696
rect 407358 404640 410044 404696
rect 407297 404638 410044 404640
rect 549884 404638 555004 404698
rect 407297 404635 407363 404638
rect 554998 404636 555004 404638
rect 555068 404636 555074 404700
rect 350441 404562 350507 404565
rect 347822 404560 350507 404562
rect 347822 404504 350446 404560
rect 350502 404504 350507 404560
rect 347822 404502 350507 404504
rect 350441 404499 350507 404502
rect 45921 403610 45987 403613
rect 48086 403610 48146 404056
rect 552841 404018 552907 404021
rect 549884 404016 552907 404018
rect 549884 403960 552846 404016
rect 552902 403960 552907 404016
rect 549884 403958 552907 403960
rect 552841 403955 552907 403958
rect 45921 403608 48146 403610
rect 45921 403552 45926 403608
rect 45982 403552 48146 403608
rect 45921 403550 48146 403552
rect 45921 403547 45987 403550
rect 552933 403338 552999 403341
rect 549884 403336 552999 403338
rect 549884 403280 552938 403336
rect 552994 403280 552999 403336
rect 549884 403278 552999 403280
rect 552933 403275 552999 403278
rect 46238 402052 46244 402116
rect 46308 402114 46314 402116
rect 48086 402114 48146 402696
rect 46308 402054 48146 402114
rect 46308 402052 46314 402054
rect 407205 401978 407271 401981
rect 407205 401976 410044 401978
rect 407205 401920 407210 401976
rect 407266 401920 410044 401976
rect 407205 401918 410044 401920
rect 407205 401915 407271 401918
rect 32806 400828 32812 400892
rect 32876 400890 32882 400892
rect 48086 400890 48146 401336
rect 32876 400830 48146 400890
rect 32876 400828 32882 400830
rect 46105 400346 46171 400349
rect 48086 400346 48146 400656
rect 46105 400344 48146 400346
rect 46105 400288 46110 400344
rect 46166 400288 48146 400344
rect 46105 400286 48146 400288
rect 347822 400346 347882 400656
rect 350441 400346 350507 400349
rect 347822 400344 350507 400346
rect 347822 400288 350446 400344
rect 350502 400288 350507 400344
rect 347822 400286 350507 400288
rect 46105 400283 46171 400286
rect 350441 400283 350507 400286
rect 408861 400346 408927 400349
rect 410014 400346 410074 400520
rect 549884 400490 550466 400550
rect 550406 400482 550466 400490
rect 550406 400422 557550 400482
rect 408861 400344 410074 400346
rect 408861 400288 408866 400344
rect 408922 400288 410074 400344
rect 408861 400286 410074 400288
rect 557490 400346 557550 400422
rect 565486 400346 565492 400348
rect 557490 400286 565492 400346
rect 408861 400283 408927 400286
rect 565486 400284 565492 400286
rect 565556 400284 565562 400348
rect 46565 399530 46631 399533
rect 48086 399530 48146 399976
rect 46565 399528 48146 399530
rect 46565 399472 46570 399528
rect 46626 399472 48146 399528
rect 46565 399470 48146 399472
rect 347822 399530 347882 399976
rect 350441 399530 350507 399533
rect 347822 399528 350507 399530
rect 347822 399472 350446 399528
rect 350502 399472 350507 399528
rect 347822 399470 350507 399472
rect 46565 399467 46631 399470
rect 350441 399467 350507 399470
rect 409505 399258 409571 399261
rect 409505 399256 410044 399258
rect 409505 399200 409510 399256
rect 409566 399200 410044 399256
rect 409505 399198 410044 399200
rect 409505 399195 409571 399198
rect 347822 397626 347882 397936
rect 407205 397898 407271 397901
rect 407205 397896 410044 397898
rect 407205 397840 407210 397896
rect 407266 397840 410044 397896
rect 407205 397838 410044 397840
rect 407205 397835 407271 397838
rect 350441 397626 350507 397629
rect 347822 397624 350507 397626
rect -960 397490 480 397580
rect 347822 397568 350446 397624
rect 350502 397568 350507 397624
rect 347822 397566 350507 397568
rect 350441 397563 350507 397566
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 46473 396674 46539 396677
rect 48086 396674 48146 397256
rect 347822 396810 347882 397256
rect 350441 396810 350507 396813
rect 347822 396808 350507 396810
rect 347822 396752 350446 396808
rect 350502 396752 350507 396808
rect 347822 396750 350507 396752
rect 350441 396747 350507 396750
rect 348141 396674 348207 396677
rect 46473 396672 48146 396674
rect 46473 396616 46478 396672
rect 46534 396616 48146 396672
rect 46473 396614 48146 396616
rect 347852 396672 348207 396674
rect 347852 396616 348146 396672
rect 348202 396616 348207 396672
rect 347852 396614 348207 396616
rect 46473 396611 46539 396614
rect 348141 396611 348207 396614
rect 347822 395450 347882 395896
rect 407205 395858 407271 395861
rect 407205 395856 410044 395858
rect 407205 395800 407210 395856
rect 407266 395800 410044 395856
rect 407205 395798 410044 395800
rect 407205 395795 407271 395798
rect 350073 395450 350139 395453
rect 347822 395448 350139 395450
rect 347822 395392 350078 395448
rect 350134 395392 350139 395448
rect 347822 395390 350139 395392
rect 350073 395387 350139 395390
rect 46565 395042 46631 395045
rect 48086 395042 48146 395216
rect 46565 395040 48146 395042
rect 46565 394984 46570 395040
rect 46626 394984 48146 395040
rect 46565 394982 48146 394984
rect 46565 394979 46631 394982
rect 347822 394906 347882 395216
rect 407941 395178 408007 395181
rect 552933 395178 552999 395181
rect 407941 395176 410044 395178
rect 407941 395120 407946 395176
rect 408002 395120 410044 395176
rect 407941 395118 410044 395120
rect 549884 395176 552999 395178
rect 549884 395120 552938 395176
rect 552994 395120 552999 395176
rect 549884 395118 552999 395120
rect 407941 395115 408007 395118
rect 552933 395115 552999 395118
rect 349797 394906 349863 394909
rect 347822 394904 349863 394906
rect 347822 394848 349802 394904
rect 349858 394848 349863 394904
rect 347822 394846 349863 394848
rect 349797 394843 349863 394846
rect 350441 394634 350507 394637
rect 347852 394632 350507 394634
rect 347852 394576 350446 394632
rect 350502 394576 350507 394632
rect 347852 394574 350507 394576
rect 350441 394571 350507 394574
rect 46565 393682 46631 393685
rect 48086 393682 48146 393856
rect 407205 393818 407271 393821
rect 552013 393818 552079 393821
rect 407205 393816 410044 393818
rect 407205 393760 407210 393816
rect 407266 393760 410044 393816
rect 407205 393758 410044 393760
rect 549884 393816 552079 393818
rect 549884 393760 552018 393816
rect 552074 393760 552079 393816
rect 549884 393758 552079 393760
rect 407205 393755 407271 393758
rect 552013 393755 552079 393758
rect 46565 393680 48146 393682
rect 46565 393624 46570 393680
rect 46626 393624 48146 393680
rect 46565 393622 48146 393624
rect 46565 393619 46631 393622
rect 46473 392730 46539 392733
rect 48086 392730 48146 393176
rect 409321 393138 409387 393141
rect 409321 393136 410044 393138
rect 409321 393080 409326 393136
rect 409382 393080 410044 393136
rect 409321 393078 410044 393080
rect 409321 393075 409387 393078
rect 46473 392728 48146 392730
rect 46473 392672 46478 392728
rect 46534 392672 48146 392728
rect 46473 392670 48146 392672
rect 46473 392667 46539 392670
rect 46565 392186 46631 392189
rect 48086 392186 48146 392496
rect 46565 392184 48146 392186
rect 46565 392128 46570 392184
rect 46626 392128 48146 392184
rect 46565 392126 48146 392128
rect 46565 392123 46631 392126
rect 347822 392050 347882 392496
rect 350441 392050 350507 392053
rect 347822 392048 350507 392050
rect 347822 391992 350446 392048
rect 350502 391992 350507 392048
rect 347822 391990 350507 391992
rect 350441 391987 350507 391990
rect 347822 391370 347882 391816
rect 407297 391778 407363 391781
rect 552841 391778 552907 391781
rect 407297 391776 410044 391778
rect 407297 391720 407302 391776
rect 407358 391720 410044 391776
rect 407297 391718 410044 391720
rect 549884 391776 552907 391778
rect 549884 391720 552846 391776
rect 552902 391720 552907 391776
rect 549884 391718 552907 391720
rect 407297 391715 407363 391718
rect 552841 391715 552907 391718
rect 583520 391628 584960 391868
rect 350073 391370 350139 391373
rect 347822 391368 350139 391370
rect 347822 391312 350078 391368
rect 350134 391312 350139 391368
rect 347822 391310 350139 391312
rect 350073 391307 350139 391310
rect 46473 390962 46539 390965
rect 48086 390962 48146 391136
rect 46473 390960 48146 390962
rect 46473 390904 46478 390960
rect 46534 390904 48146 390960
rect 46473 390902 48146 390904
rect 46473 390899 46539 390902
rect 347822 390690 347882 391136
rect 407205 391098 407271 391101
rect 552933 391098 552999 391101
rect 407205 391096 410044 391098
rect 407205 391040 407210 391096
rect 407266 391040 410044 391096
rect 407205 391038 410044 391040
rect 549884 391096 552999 391098
rect 549884 391040 552938 391096
rect 552994 391040 552999 391096
rect 549884 391038 552999 391040
rect 407205 391035 407271 391038
rect 552933 391035 552999 391038
rect 348049 390690 348115 390693
rect 347822 390688 348115 390690
rect 347822 390632 348054 390688
rect 348110 390632 348115 390688
rect 347822 390630 348115 390632
rect 348049 390627 348115 390630
rect 46565 390554 46631 390557
rect 46565 390552 48116 390554
rect 46565 390496 46570 390552
rect 46626 390496 48116 390552
rect 46565 390494 48116 390496
rect 46565 390491 46631 390494
rect 347822 390010 347882 390456
rect 552289 390418 552355 390421
rect 549884 390416 552355 390418
rect 549884 390360 552294 390416
rect 552350 390360 552355 390416
rect 549884 390358 552355 390360
rect 552289 390355 552355 390358
rect 350349 390010 350415 390013
rect 347822 390008 350415 390010
rect 347822 389952 350354 390008
rect 350410 389952 350415 390008
rect 347822 389950 350415 389952
rect 350349 389947 350415 389950
rect 350441 389874 350507 389877
rect 347852 389872 350507 389874
rect 347852 389816 350446 389872
rect 350502 389816 350507 389872
rect 347852 389814 350507 389816
rect 350441 389811 350507 389814
rect 46565 389602 46631 389605
rect 48086 389602 48146 389776
rect 408401 389738 408467 389741
rect 408401 389736 410044 389738
rect 408401 389680 408406 389736
rect 408462 389680 410044 389736
rect 408401 389678 410044 389680
rect 408401 389675 408467 389678
rect 46565 389600 48146 389602
rect 46565 389544 46570 389600
rect 46626 389544 48146 389600
rect 46565 389542 48146 389544
rect 46565 389539 46631 389542
rect 552933 388378 552999 388381
rect 549884 388376 552999 388378
rect 549884 388320 552938 388376
rect 552994 388320 552999 388376
rect 549884 388318 552999 388320
rect 552933 388315 552999 388318
rect 350441 387834 350507 387837
rect 347852 387832 350507 387834
rect 347852 387776 350446 387832
rect 350502 387776 350507 387832
rect 347852 387774 350507 387776
rect 350441 387771 350507 387774
rect 552933 387698 552999 387701
rect 549884 387696 552999 387698
rect 549884 387640 552938 387696
rect 552994 387640 552999 387696
rect 549884 387638 552999 387640
rect 552933 387635 552999 387638
rect 350349 387154 350415 387157
rect 347852 387152 350415 387154
rect 347852 387096 350354 387152
rect 350410 387096 350415 387152
rect 347852 387094 350415 387096
rect 350349 387091 350415 387094
rect 46565 386474 46631 386477
rect 46565 386472 48116 386474
rect 46565 386416 46570 386472
rect 46626 386416 48116 386472
rect 46565 386414 48116 386416
rect 46565 386411 46631 386414
rect 46473 385794 46539 385797
rect 349470 385794 349476 385796
rect 46473 385792 48116 385794
rect 46473 385736 46478 385792
rect 46534 385736 48116 385792
rect 46473 385734 48116 385736
rect 347852 385734 349476 385794
rect 46473 385731 46539 385734
rect 349470 385732 349476 385734
rect 349540 385732 349546 385796
rect 407205 385658 407271 385661
rect 552933 385658 552999 385661
rect 407205 385656 410044 385658
rect 407205 385600 407210 385656
rect 407266 385600 410044 385656
rect 407205 385598 410044 385600
rect 549884 385656 552999 385658
rect 549884 385600 552938 385656
rect 552994 385600 552999 385656
rect 549884 385598 552999 385600
rect 407205 385595 407271 385598
rect 552933 385595 552999 385598
rect 46565 385114 46631 385117
rect 350901 385114 350967 385117
rect 46565 385112 48116 385114
rect 46565 385056 46570 385112
rect 46626 385056 48116 385112
rect 46565 385054 48116 385056
rect 347852 385112 350967 385114
rect 347852 385056 350906 385112
rect 350962 385056 350967 385112
rect 347852 385054 350967 385056
rect 46565 385051 46631 385054
rect 350901 385051 350967 385054
rect 407205 384978 407271 384981
rect 407205 384976 410044 384978
rect 407205 384920 407210 384976
rect 407266 384920 410044 384976
rect 407205 384918 410044 384920
rect 407205 384915 407271 384918
rect -960 384284 480 384524
rect 351085 383754 351151 383757
rect 347852 383752 351151 383754
rect 347852 383696 351090 383752
rect 351146 383696 351151 383752
rect 347852 383694 351151 383696
rect 351085 383691 351151 383694
rect 44950 383012 44956 383076
rect 45020 383074 45026 383076
rect 407941 383074 408007 383077
rect 410014 383074 410074 383520
rect 45020 383014 48116 383074
rect 407941 383072 410074 383074
rect 407941 383016 407946 383072
rect 408002 383016 410074 383072
rect 407941 383014 410074 383016
rect 45020 383012 45026 383014
rect 407941 383011 408007 383014
rect 408125 382938 408191 382941
rect 408125 382936 410044 382938
rect 408125 382880 408130 382936
rect 408186 382880 410044 382936
rect 408125 382878 410044 382880
rect 408125 382875 408191 382878
rect 46565 382394 46631 382397
rect 350441 382394 350507 382397
rect 46565 382392 48116 382394
rect 46565 382336 46570 382392
rect 46626 382336 48116 382392
rect 46565 382334 48116 382336
rect 347852 382392 350507 382394
rect 347852 382336 350446 382392
rect 350502 382336 350507 382392
rect 347852 382334 350507 382336
rect 46565 382331 46631 382334
rect 350441 382331 350507 382334
rect 347822 381442 347882 381616
rect 407205 381578 407271 381581
rect 552933 381578 552999 381581
rect 407205 381576 410044 381578
rect 407205 381520 407210 381576
rect 407266 381520 410044 381576
rect 407205 381518 410044 381520
rect 549884 381576 552999 381578
rect 549884 381520 552938 381576
rect 552994 381520 552999 381576
rect 549884 381518 552999 381520
rect 407205 381515 407271 381518
rect 552933 381515 552999 381518
rect 350349 381442 350415 381445
rect 347822 381440 350415 381442
rect 347822 381384 350354 381440
rect 350410 381384 350415 381440
rect 347822 381382 350415 381384
rect 350349 381379 350415 381382
rect 46473 381034 46539 381037
rect 350441 381034 350507 381037
rect 46473 381032 48116 381034
rect 46473 380976 46478 381032
rect 46534 380976 48116 381032
rect 46473 380974 48116 380976
rect 347852 381032 350507 381034
rect 347852 380976 350446 381032
rect 350502 380976 350507 381032
rect 347852 380974 350507 380976
rect 46473 380971 46539 380974
rect 350441 380971 350507 380974
rect 46565 379946 46631 379949
rect 48086 379946 48146 380256
rect 46565 379944 48146 379946
rect 46565 379888 46570 379944
rect 46626 379888 48146 379944
rect 46565 379886 48146 379888
rect 46565 379883 46631 379886
rect 347822 379810 347882 380256
rect 351085 379810 351151 379813
rect 347822 379808 351151 379810
rect 347822 379752 351090 379808
rect 351146 379752 351151 379808
rect 347822 379750 351151 379752
rect 351085 379747 351151 379750
rect 407205 378858 407271 378861
rect 550081 378858 550147 378861
rect 407205 378856 410044 378858
rect 407205 378800 407210 378856
rect 407266 378800 410044 378856
rect 407205 378798 410044 378800
rect 549884 378856 550147 378858
rect 549884 378800 550086 378856
rect 550142 378800 550147 378856
rect 549884 378798 550147 378800
rect 407205 378795 407271 378798
rect 550081 378795 550147 378798
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 46565 378314 46631 378317
rect 46565 378312 48116 378314
rect 46565 378256 46570 378312
rect 46626 378256 48116 378312
rect 583520 378300 584960 378390
rect 46565 378254 48116 378256
rect 46565 378251 46631 378254
rect 407982 378116 407988 378180
rect 408052 378178 408058 378180
rect 553577 378178 553643 378181
rect 408052 378118 410044 378178
rect 549884 378176 553643 378178
rect 549884 378120 553582 378176
rect 553638 378120 553643 378176
rect 549884 378118 553643 378120
rect 408052 378116 408058 378118
rect 553577 378115 553643 378118
rect 347822 377226 347882 377536
rect 409597 377498 409663 377501
rect 552933 377498 552999 377501
rect 409597 377496 410044 377498
rect 409597 377440 409602 377496
rect 409658 377440 410044 377496
rect 409597 377438 410044 377440
rect 549884 377496 552999 377498
rect 549884 377440 552938 377496
rect 552994 377440 552999 377496
rect 549884 377438 552999 377440
rect 409597 377435 409663 377438
rect 552933 377435 552999 377438
rect 350441 377226 350507 377229
rect 347822 377224 350507 377226
rect 347822 377168 350446 377224
rect 350502 377168 350507 377224
rect 347822 377166 350507 377168
rect 350441 377163 350507 377166
rect 347957 377090 348023 377093
rect 347822 377088 348023 377090
rect 347822 377032 347962 377088
rect 348018 377032 348023 377088
rect 347822 377030 348023 377032
rect 347822 376924 347882 377030
rect 347957 377027 348023 377030
rect 47209 376274 47275 376277
rect 47209 376272 48116 376274
rect 47209 376216 47214 376272
rect 47270 376216 48116 376272
rect 47209 376214 48116 376216
rect 47209 376211 47275 376214
rect 347822 375866 347882 376176
rect 350349 375866 350415 375869
rect 347822 375864 350415 375866
rect 347822 375808 350354 375864
rect 350410 375808 350415 375864
rect 347822 375806 350415 375808
rect 350349 375803 350415 375806
rect 350441 374914 350507 374917
rect 347852 374912 350507 374914
rect 347852 374856 350446 374912
rect 350502 374856 350507 374912
rect 347852 374854 350507 374856
rect 350441 374851 350507 374854
rect 46473 374098 46539 374101
rect 48086 374098 48146 374136
rect 46473 374096 48146 374098
rect 46473 374040 46478 374096
rect 46534 374040 48146 374096
rect 46473 374038 48146 374040
rect 407205 374098 407271 374101
rect 407205 374096 410044 374098
rect 407205 374040 407210 374096
rect 407266 374040 410044 374096
rect 407205 374038 410044 374040
rect 46473 374035 46539 374038
rect 407205 374035 407271 374038
rect 46105 373146 46171 373149
rect 48086 373146 48146 373456
rect 46105 373144 48146 373146
rect 46105 373088 46110 373144
rect 46166 373088 48146 373144
rect 46105 373086 48146 373088
rect 46105 373083 46171 373086
rect 347822 372874 347882 373456
rect 407205 373418 407271 373421
rect 407205 373416 410044 373418
rect 407205 373360 407210 373416
rect 407266 373360 410044 373416
rect 407205 373358 410044 373360
rect 407205 373355 407271 373358
rect 350441 372874 350507 372877
rect 347822 372872 350507 372874
rect 347822 372816 350446 372872
rect 350502 372816 350507 372872
rect 347822 372814 350507 372816
rect 350441 372811 350507 372814
rect 46473 372738 46539 372741
rect 48086 372738 48146 372776
rect 552933 372738 552999 372741
rect 46473 372736 48146 372738
rect 46473 372680 46478 372736
rect 46534 372680 48146 372736
rect 46473 372678 48146 372680
rect 549884 372736 552999 372738
rect 549884 372680 552938 372736
rect 552994 372680 552999 372736
rect 549884 372678 552999 372680
rect 46473 372675 46539 372678
rect 552933 372675 552999 372678
rect 46473 371514 46539 371517
rect 48086 371514 48146 372096
rect 406653 372058 406719 372061
rect 406653 372056 410044 372058
rect 406653 372000 406658 372056
rect 406714 372000 410044 372056
rect 406653 371998 410044 372000
rect 406653 371995 406719 371998
rect 46473 371512 48146 371514
rect -960 371228 480 371468
rect 46473 371456 46478 371512
rect 46534 371456 48146 371512
rect 46473 371454 48146 371456
rect 46473 371451 46539 371454
rect 347822 371378 347882 371416
rect 350441 371378 350507 371381
rect 551001 371378 551067 371381
rect 347822 371376 350507 371378
rect 347822 371320 350446 371376
rect 350502 371320 350507 371376
rect 347822 371318 350507 371320
rect 549884 371376 551067 371378
rect 549884 371320 551006 371376
rect 551062 371320 551067 371376
rect 549884 371318 551067 371320
rect 350441 371315 350507 371318
rect 551001 371315 551067 371318
rect 407205 370698 407271 370701
rect 552933 370698 552999 370701
rect 407205 370696 410044 370698
rect 407205 370640 407210 370696
rect 407266 370640 410044 370696
rect 407205 370638 410044 370640
rect 549884 370696 552999 370698
rect 549884 370640 552938 370696
rect 552994 370640 552999 370696
rect 549884 370638 552999 370640
rect 407205 370635 407271 370638
rect 552933 370635 552999 370638
rect 350993 370154 351059 370157
rect 347852 370152 351059 370154
rect 347852 370096 350998 370152
rect 351054 370096 351059 370152
rect 347852 370094 351059 370096
rect 350993 370091 351059 370094
rect 46473 369066 46539 369069
rect 48086 369066 48146 369376
rect 407205 369338 407271 369341
rect 552841 369338 552907 369341
rect 407205 369336 410044 369338
rect 407205 369280 407210 369336
rect 407266 369280 410044 369336
rect 407205 369278 410044 369280
rect 549884 369336 552907 369338
rect 549884 369280 552846 369336
rect 552902 369280 552907 369336
rect 549884 369278 552907 369280
rect 407205 369275 407271 369278
rect 552841 369275 552907 369278
rect 46473 369064 48146 369066
rect 46473 369008 46478 369064
rect 46534 369008 48146 369064
rect 46473 369006 48146 369008
rect 46473 369003 46539 369006
rect 347822 368522 347882 368696
rect 552933 368658 552999 368661
rect 549884 368656 552999 368658
rect 549884 368600 552938 368656
rect 552994 368600 552999 368656
rect 549884 368598 552999 368600
rect 552933 368595 552999 368598
rect 347957 368522 348023 368525
rect 347822 368520 348023 368522
rect 347822 368464 347962 368520
rect 348018 368464 348023 368520
rect 347822 368462 348023 368464
rect 347957 368459 348023 368462
rect 46381 367706 46447 367709
rect 48086 367706 48146 368016
rect 552013 367978 552079 367981
rect 549884 367976 552079 367978
rect 549884 367920 552018 367976
rect 552074 367920 552079 367976
rect 549884 367918 552079 367920
rect 552013 367915 552079 367918
rect 46381 367704 48146 367706
rect 46381 367648 46386 367704
rect 46442 367648 48146 367704
rect 46381 367646 48146 367648
rect 46381 367643 46447 367646
rect 549884 366490 550282 366550
rect 550222 366482 550282 366490
rect 552841 366482 552907 366485
rect 550222 366480 552907 366482
rect 550222 366424 552846 366480
rect 552902 366424 552907 366480
rect 550222 366422 552907 366424
rect 552841 366419 552907 366422
rect 46473 366074 46539 366077
rect 46473 366072 48116 366074
rect 46473 366016 46478 366072
rect 46534 366016 48116 366072
rect 46473 366014 48116 366016
rect 46473 366011 46539 366014
rect 552933 365938 552999 365941
rect 549884 365936 552999 365938
rect 549884 365880 552938 365936
rect 552994 365880 552999 365936
rect 549884 365878 552999 365880
rect 552933 365875 552999 365878
rect 350441 365394 350507 365397
rect 347852 365392 350507 365394
rect 347852 365336 350446 365392
rect 350502 365336 350507 365392
rect 347852 365334 350507 365336
rect 350441 365331 350507 365334
rect 551093 365258 551159 365261
rect 549884 365256 551159 365258
rect 549884 365200 551098 365256
rect 551154 365200 551159 365256
rect 549884 365198 551159 365200
rect 551093 365195 551159 365198
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect 347822 364442 347882 364616
rect 409689 364578 409755 364581
rect 409689 364576 410044 364578
rect 409689 364520 409694 364576
rect 409750 364520 410044 364576
rect 409689 364518 410044 364520
rect 409689 364515 409755 364518
rect 350441 364442 350507 364445
rect 347822 364440 350507 364442
rect 347822 364384 350446 364440
rect 350502 364384 350507 364440
rect 347822 364382 350507 364384
rect 350441 364379 350507 364382
rect 46473 363490 46539 363493
rect 48086 363490 48146 363936
rect 46473 363488 48146 363490
rect 46473 363432 46478 363488
rect 46534 363432 48146 363488
rect 46473 363430 48146 363432
rect 46473 363427 46539 363430
rect 347822 363354 347882 363936
rect 550817 363898 550883 363901
rect 549884 363896 550883 363898
rect 549884 363840 550822 363896
rect 550878 363840 550883 363896
rect 549884 363838 550883 363840
rect 550817 363835 550883 363838
rect 350993 363354 351059 363357
rect 347822 363352 351059 363354
rect 347822 363296 350998 363352
rect 351054 363296 351059 363352
rect 347822 363294 351059 363296
rect 350993 363291 351059 363294
rect 408033 362538 408099 362541
rect 408033 362536 410044 362538
rect 408033 362480 408038 362536
rect 408094 362480 410044 362536
rect 408033 362478 410044 362480
rect 408033 362475 408099 362478
rect 407205 361178 407271 361181
rect 552933 361178 552999 361181
rect 407205 361176 410044 361178
rect 407205 361120 407210 361176
rect 407266 361120 410044 361176
rect 407205 361118 410044 361120
rect 549884 361176 552999 361178
rect 549884 361120 552938 361176
rect 552994 361120 552999 361176
rect 549884 361118 552999 361120
rect 407205 361115 407271 361118
rect 552933 361115 552999 361118
rect 407205 360498 407271 360501
rect 552197 360498 552263 360501
rect 407205 360496 410044 360498
rect 407205 360440 407210 360496
rect 407266 360440 410044 360496
rect 407205 360438 410044 360440
rect 549884 360496 552263 360498
rect 549884 360440 552202 360496
rect 552258 360440 552263 360496
rect 549884 360438 552263 360440
rect 407205 360435 407271 360438
rect 552197 360435 552263 360438
rect 45001 359410 45067 359413
rect 48086 359410 48146 359856
rect 45001 359408 48146 359410
rect 45001 359352 45006 359408
rect 45062 359352 48146 359408
rect 45001 359350 48146 359352
rect 45001 359347 45067 359350
rect 347822 358866 347882 359176
rect 349470 358866 349476 358868
rect 347822 358806 349476 358866
rect 349470 358804 349476 358806
rect 349540 358804 349546 358868
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 347822 358050 347882 358496
rect 552657 358458 552723 358461
rect 549884 358456 552723 358458
rect 549884 358400 552662 358456
rect 552718 358400 552723 358456
rect 549884 358398 552723 358400
rect 552657 358395 552723 358398
rect 350441 358050 350507 358053
rect 347822 358048 350507 358050
rect 347822 357992 350446 358048
rect 350502 357992 350507 358048
rect 347822 357990 350507 357992
rect 350441 357987 350507 357990
rect 46473 357914 46539 357917
rect 46473 357912 48116 357914
rect 46473 357856 46478 357912
rect 46534 357856 48116 357912
rect 46473 357854 48116 357856
rect 46473 357851 46539 357854
rect 407205 357778 407271 357781
rect 552933 357778 552999 357781
rect 407205 357776 410044 357778
rect 407205 357720 407210 357776
rect 407266 357720 410044 357776
rect 407205 357718 410044 357720
rect 549884 357776 552999 357778
rect 549884 357720 552938 357776
rect 552994 357720 552999 357776
rect 549884 357718 552999 357720
rect 407205 357715 407271 357718
rect 552933 357715 552999 357718
rect 347822 356690 347882 357136
rect 407205 357098 407271 357101
rect 407205 357096 410044 357098
rect 407205 357040 407210 357096
rect 407266 357040 410044 357096
rect 407205 357038 410044 357040
rect 407205 357035 407271 357038
rect 349981 356690 350047 356693
rect 347822 356688 350047 356690
rect 347822 356632 349986 356688
rect 350042 356632 350047 356688
rect 347822 356630 350047 356632
rect 349981 356627 350047 356630
rect 406653 356418 406719 356421
rect 406653 356416 410044 356418
rect 406653 356360 406658 356416
rect 406714 356360 410044 356416
rect 406653 356358 410044 356360
rect 406653 356355 406719 356358
rect 350441 355874 350507 355877
rect 347852 355872 350507 355874
rect 347852 355816 350446 355872
rect 350502 355816 350507 355872
rect 347852 355814 350507 355816
rect 350441 355811 350507 355814
rect 552933 355738 552999 355741
rect 549884 355736 552999 355738
rect 549884 355680 552938 355736
rect 552994 355680 552999 355736
rect 549884 355678 552999 355680
rect 552933 355675 552999 355678
rect 46473 354786 46539 354789
rect 48086 354786 48146 355096
rect 46473 354784 48146 354786
rect 46473 354728 46478 354784
rect 46534 354728 48146 354784
rect 46473 354726 48146 354728
rect 347822 354786 347882 355096
rect 350441 354786 350507 354789
rect 347822 354784 350507 354786
rect 347822 354728 350446 354784
rect 350502 354728 350507 354784
rect 347822 354726 350507 354728
rect 46473 354723 46539 354726
rect 350441 354723 350507 354726
rect 553117 354378 553183 354381
rect 549884 354376 553183 354378
rect 549884 354320 553122 354376
rect 553178 354320 553183 354376
rect 549884 354318 553183 354320
rect 553117 354315 553183 354318
rect 407205 353698 407271 353701
rect 553117 353698 553183 353701
rect 407205 353696 410044 353698
rect 407205 353640 407210 353696
rect 407266 353640 410044 353696
rect 407205 353638 410044 353640
rect 549884 353696 553183 353698
rect 549884 353640 553122 353696
rect 553178 353640 553183 353696
rect 549884 353638 553183 353640
rect 407205 353635 407271 353638
rect 553117 353635 553183 353638
rect 46473 353154 46539 353157
rect 46473 353152 48116 353154
rect 46473 353096 46478 353152
rect 46534 353096 48116 353152
rect 46473 353094 48116 353096
rect 46473 353091 46539 353094
rect 407297 353018 407363 353021
rect 407297 353016 410044 353018
rect 407297 352960 407302 353016
rect 407358 352960 410044 353016
rect 407297 352958 410044 352960
rect 407297 352955 407363 352958
rect 407205 352338 407271 352341
rect 407205 352336 410044 352338
rect 407205 352280 407210 352336
rect 407266 352280 410044 352336
rect 407205 352278 410044 352280
rect 407205 352275 407271 352278
rect 583520 351780 584960 352020
rect 407205 351658 407271 351661
rect 552289 351658 552355 351661
rect 407205 351656 410044 351658
rect 407205 351600 407210 351656
rect 407266 351600 410044 351656
rect 407205 351598 410044 351600
rect 549884 351656 552355 351658
rect 549884 351600 552294 351656
rect 552350 351600 552355 351656
rect 549884 351598 552355 351600
rect 407205 351595 407271 351598
rect 552289 351595 552355 351598
rect 347822 350706 347882 351016
rect 552013 350978 552079 350981
rect 549884 350976 552079 350978
rect 549884 350920 552018 350976
rect 552074 350920 552079 350976
rect 549884 350918 552079 350920
rect 552013 350915 552079 350918
rect 350441 350706 350507 350709
rect 347822 350704 350507 350706
rect 347822 350648 350446 350704
rect 350502 350648 350507 350704
rect 347822 350646 350507 350648
rect 350441 350643 350507 350646
rect 347822 349890 347882 350336
rect 350349 349890 350415 349893
rect 347822 349888 350415 349890
rect 347822 349832 350354 349888
rect 350410 349832 350415 349888
rect 347822 349830 350415 349832
rect 350349 349827 350415 349830
rect 46473 349482 46539 349485
rect 48086 349482 48146 349656
rect 46473 349480 48146 349482
rect 46473 349424 46478 349480
rect 46534 349424 48146 349480
rect 46473 349422 48146 349424
rect 46473 349419 46539 349422
rect 347822 349346 347882 349656
rect 350441 349346 350507 349349
rect 347822 349344 350507 349346
rect 347822 349288 350446 349344
rect 350502 349288 350507 349344
rect 347822 349286 350507 349288
rect 350441 349283 350507 349286
rect 407205 349346 407271 349349
rect 410014 349346 410074 349520
rect 549884 349490 550282 349550
rect 550222 349482 550282 349490
rect 553117 349482 553183 349485
rect 550222 349480 553183 349482
rect 550222 349424 553122 349480
rect 553178 349424 553183 349480
rect 550222 349422 553183 349424
rect 553117 349419 553183 349422
rect 407205 349344 410074 349346
rect 407205 349288 407210 349344
rect 407266 349288 410074 349344
rect 407205 349286 410074 349288
rect 407205 349283 407271 349286
rect 46473 347170 46539 347173
rect 48086 347170 48146 347616
rect 552657 347578 552723 347581
rect 549884 347576 552723 347578
rect 549884 347520 552662 347576
rect 552718 347520 552723 347576
rect 549884 347518 552723 347520
rect 552657 347515 552723 347518
rect 46473 347168 48146 347170
rect 46473 347112 46478 347168
rect 46534 347112 48146 347168
rect 46473 347110 48146 347112
rect 46473 347107 46539 347110
rect 349245 347034 349311 347037
rect 347852 347032 349311 347034
rect 347852 346976 349250 347032
rect 349306 346976 349311 347032
rect 347852 346974 349311 346976
rect 349245 346971 349311 346974
rect 408033 346898 408099 346901
rect 553117 346898 553183 346901
rect 408033 346896 410044 346898
rect 408033 346840 408038 346896
rect 408094 346840 410044 346896
rect 408033 346838 410044 346840
rect 549884 346896 553183 346898
rect 549884 346840 553122 346896
rect 553178 346840 553183 346896
rect 549884 346838 553183 346840
rect 408033 346835 408099 346838
rect 553117 346835 553183 346838
rect 347822 345810 347882 346256
rect 350349 345810 350415 345813
rect 347822 345808 350415 345810
rect 347822 345752 350354 345808
rect 350410 345752 350415 345808
rect 347822 345750 350415 345752
rect 350349 345747 350415 345750
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 45921 345402 45987 345405
rect 48086 345402 48146 345576
rect 407205 345538 407271 345541
rect 407205 345536 410044 345538
rect 407205 345480 407210 345536
rect 407266 345480 410044 345536
rect 407205 345478 410044 345480
rect 407205 345475 407271 345478
rect 45921 345400 48146 345402
rect 45921 345344 45926 345400
rect 45982 345344 48146 345400
rect 45921 345342 48146 345344
rect 45921 345339 45987 345342
rect 347822 344450 347882 344896
rect 407205 344858 407271 344861
rect 407205 344856 410044 344858
rect 407205 344800 407210 344856
rect 407266 344800 410044 344856
rect 407205 344798 410044 344800
rect 407205 344795 407271 344798
rect 350349 344450 350415 344453
rect 347822 344448 350415 344450
rect 347822 344392 350354 344448
rect 350410 344392 350415 344448
rect 347822 344390 350415 344392
rect 350349 344387 350415 344390
rect 347822 344042 347882 344216
rect 350165 344042 350231 344045
rect 347822 344040 350231 344042
rect 347822 343984 350170 344040
rect 350226 343984 350231 344040
rect 347822 343982 350231 343984
rect 350165 343979 350231 343982
rect 407205 343498 407271 343501
rect 553117 343498 553183 343501
rect 407205 343496 410044 343498
rect 407205 343440 407210 343496
rect 407266 343440 410044 343496
rect 407205 343438 410044 343440
rect 549884 343496 553183 343498
rect 549884 343440 553122 343496
rect 553178 343440 553183 343496
rect 549884 343438 553183 343440
rect 407205 343435 407271 343438
rect 553117 343435 553183 343438
rect 409413 342818 409479 342821
rect 552013 342818 552079 342821
rect 409413 342816 410044 342818
rect 409413 342760 409418 342816
rect 409474 342760 410044 342816
rect 409413 342758 410044 342760
rect 549884 342816 552079 342818
rect 549884 342760 552018 342816
rect 552074 342760 552079 342816
rect 549884 342758 552079 342760
rect 409413 342755 409479 342758
rect 552013 342755 552079 342758
rect 350349 342274 350415 342277
rect 347852 342272 350415 342274
rect 347852 342216 350354 342272
rect 350410 342216 350415 342272
rect 347852 342214 350415 342216
rect 350349 342211 350415 342214
rect 348734 341396 348740 341460
rect 348804 341458 348810 341460
rect 368933 341458 368999 341461
rect 348804 341456 368999 341458
rect 348804 341400 368938 341456
rect 368994 341400 368999 341456
rect 348804 341398 368999 341400
rect 348804 341396 348810 341398
rect 368933 341395 368999 341398
rect 407205 340778 407271 340781
rect 553577 340778 553643 340781
rect 407205 340776 410044 340778
rect 407205 340720 407210 340776
rect 407266 340720 410044 340776
rect 407205 340718 410044 340720
rect 549884 340776 553643 340778
rect 549884 340720 553582 340776
rect 553638 340720 553643 340776
rect 549884 340718 553643 340720
rect 407205 340715 407271 340718
rect 553577 340715 553643 340718
rect 552933 340098 552999 340101
rect 549884 340096 552999 340098
rect 549884 340040 552938 340096
rect 552994 340040 552999 340096
rect 549884 340038 552999 340040
rect 552933 340035 552999 340038
rect 45185 339554 45251 339557
rect 45185 339552 48116 339554
rect 45185 339496 45190 339552
rect 45246 339496 48116 339552
rect 45185 339494 48116 339496
rect 45185 339491 45251 339494
rect 409689 339418 409755 339421
rect 409689 339416 410044 339418
rect 409689 339360 409694 339416
rect 409750 339360 410044 339416
rect 409689 339358 410044 339360
rect 409689 339355 409755 339358
rect 553117 338738 553183 338741
rect 549884 338736 553183 338738
rect 549884 338680 553122 338736
rect 553178 338680 553183 338736
rect 549884 338678 553183 338680
rect 553117 338675 553183 338678
rect 583520 338452 584960 338692
rect 350349 338194 350415 338197
rect 347852 338192 350415 338194
rect 347852 338136 350354 338192
rect 350410 338136 350415 338192
rect 347852 338134 350415 338136
rect 350349 338131 350415 338134
rect 46473 336834 46539 336837
rect 46473 336832 48116 336834
rect 46473 336776 46478 336832
rect 46534 336776 48116 336832
rect 46473 336774 48116 336776
rect 46473 336771 46539 336774
rect 407205 336698 407271 336701
rect 559230 336698 559236 336700
rect 407205 336696 410044 336698
rect 407205 336640 407210 336696
rect 407266 336640 410044 336696
rect 407205 336638 410044 336640
rect 549884 336638 559236 336698
rect 407205 336635 407271 336638
rect 559230 336636 559236 336638
rect 559300 336636 559306 336700
rect 349613 336154 349679 336157
rect 347852 336152 349679 336154
rect 347852 336096 349618 336152
rect 349674 336096 349679 336152
rect 347852 336094 349679 336096
rect 349613 336091 349679 336094
rect 552933 336018 552999 336021
rect 549884 336016 552999 336018
rect 549884 335960 552938 336016
rect 552994 335960 552999 336016
rect 549884 335958 552999 335960
rect 552933 335955 552999 335958
rect 47209 335474 47275 335477
rect 47209 335472 48116 335474
rect 47209 335416 47214 335472
rect 47270 335416 48116 335472
rect 47209 335414 48116 335416
rect 47209 335411 47275 335414
rect 553117 335338 553183 335341
rect 549884 335336 553183 335338
rect 410014 334794 410074 335308
rect 549884 335280 553122 335336
rect 553178 335280 553183 335336
rect 549884 335278 553183 335280
rect 553117 335275 553183 335278
rect 409646 334734 410074 334794
rect 409646 334522 409706 334734
rect 409781 334658 409847 334661
rect 553117 334658 553183 334661
rect 409781 334656 410044 334658
rect 409781 334600 409786 334656
rect 409842 334600 410044 334656
rect 409781 334598 410044 334600
rect 549884 334656 553183 334658
rect 549884 334600 553122 334656
rect 553178 334600 553183 334656
rect 549884 334598 553183 334600
rect 409781 334595 409847 334598
rect 553117 334595 553183 334598
rect 409781 334522 409847 334525
rect 409646 334520 409847 334522
rect 409646 334464 409786 334520
rect 409842 334464 409847 334520
rect 409646 334462 409847 334464
rect 409781 334459 409847 334462
rect 350349 334114 350415 334117
rect 347852 334112 350415 334114
rect 347852 334056 350354 334112
rect 350410 334056 350415 334112
rect 347852 334054 350415 334056
rect 350349 334051 350415 334054
rect 551001 333978 551067 333981
rect 549884 333976 551067 333978
rect 549884 333920 551006 333976
rect 551062 333920 551067 333976
rect 549884 333918 551067 333920
rect 551001 333915 551067 333918
rect 347822 332754 347882 333336
rect 350349 332754 350415 332757
rect 347822 332752 350415 332754
rect 347822 332696 350354 332752
rect 350410 332696 350415 332752
rect 347822 332694 350415 332696
rect 350349 332691 350415 332694
rect 407297 332618 407363 332621
rect 407297 332616 410044 332618
rect 407297 332560 407302 332616
rect 407358 332560 410044 332616
rect 407297 332558 410044 332560
rect 407297 332555 407363 332558
rect -960 332196 480 332436
rect 347822 331258 347882 331296
rect 349889 331258 349955 331261
rect 347822 331256 349955 331258
rect 347822 331200 349894 331256
rect 349950 331200 349955 331256
rect 347822 331198 349955 331200
rect 349889 331195 349955 331198
rect 407205 331258 407271 331261
rect 552473 331258 552539 331261
rect 407205 331256 410044 331258
rect 407205 331200 407210 331256
rect 407266 331200 410044 331256
rect 407205 331198 410044 331200
rect 549884 331256 552539 331258
rect 549884 331200 552478 331256
rect 552534 331200 552539 331256
rect 549884 331198 552539 331200
rect 407205 331195 407271 331198
rect 552473 331195 552539 331198
rect 46841 330714 46907 330717
rect 350717 330714 350783 330717
rect 46841 330712 48116 330714
rect 46841 330656 46846 330712
rect 46902 330656 48116 330712
rect 46841 330654 48116 330656
rect 347852 330712 350783 330714
rect 347852 330656 350722 330712
rect 350778 330656 350783 330712
rect 347852 330654 350783 330656
rect 46841 330651 46907 330654
rect 350717 330651 350783 330654
rect 407205 330578 407271 330581
rect 407205 330576 410044 330578
rect 407205 330520 407210 330576
rect 407266 330520 410044 330576
rect 407205 330518 410044 330520
rect 407205 330515 407271 330518
rect 46381 329898 46447 329901
rect 48086 329898 48146 329936
rect 46381 329896 48146 329898
rect 46381 329840 46386 329896
rect 46442 329840 48146 329896
rect 46381 329838 48146 329840
rect 347822 329898 347882 329936
rect 350349 329898 350415 329901
rect 347822 329896 350415 329898
rect 347822 329840 350354 329896
rect 350410 329840 350415 329896
rect 347822 329838 350415 329840
rect 46381 329835 46447 329838
rect 350349 329835 350415 329838
rect 45829 328810 45895 328813
rect 48086 328810 48146 329256
rect 347822 328946 347882 329256
rect 350349 328946 350415 328949
rect 347822 328944 350415 328946
rect 347822 328888 350354 328944
rect 350410 328888 350415 328944
rect 347822 328886 350415 328888
rect 350349 328883 350415 328886
rect 45829 328808 48146 328810
rect 45829 328752 45834 328808
rect 45890 328752 48146 328808
rect 45829 328750 48146 328752
rect 45829 328747 45895 328750
rect 407205 328538 407271 328541
rect 407205 328536 410044 328538
rect 407205 328480 407210 328536
rect 407266 328480 410044 328536
rect 407205 328478 410044 328480
rect 407205 328475 407271 328478
rect 46841 327994 46907 327997
rect 46841 327992 48116 327994
rect 46841 327936 46846 327992
rect 46902 327936 48116 327992
rect 46841 327934 48116 327936
rect 46841 327931 46907 327934
rect 408401 327858 408467 327861
rect 551185 327858 551251 327861
rect 408401 327856 410044 327858
rect 408401 327800 408406 327856
rect 408462 327800 410044 327856
rect 408401 327798 410044 327800
rect 549884 327856 551251 327858
rect 549884 327800 551190 327856
rect 551246 327800 551251 327856
rect 549884 327798 551251 327800
rect 408401 327795 408467 327798
rect 551185 327795 551251 327798
rect 553117 327178 553183 327181
rect 549884 327176 553183 327178
rect 549884 327120 553122 327176
rect 553178 327120 553183 327176
rect 549884 327118 553183 327120
rect 553117 327115 553183 327118
rect 552933 326498 552999 326501
rect 549884 326496 552999 326498
rect 549884 326440 552938 326496
rect 552994 326440 552999 326496
rect 549884 326438 552999 326440
rect 552933 326435 552999 326438
rect 347822 325818 347882 325856
rect 350349 325818 350415 325821
rect 347822 325816 350415 325818
rect 347822 325760 350354 325816
rect 350410 325760 350415 325816
rect 347822 325758 350415 325760
rect 350349 325755 350415 325758
rect 360694 325756 360700 325820
rect 360764 325818 360770 325820
rect 553117 325818 553183 325821
rect 360764 325758 410044 325818
rect 549884 325816 553183 325818
rect 549884 325760 553122 325816
rect 553178 325760 553183 325816
rect 549884 325758 553183 325760
rect 360764 325756 360770 325758
rect 553117 325755 553183 325758
rect 46841 325274 46907 325277
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 46841 325272 48116 325274
rect 46841 325216 46846 325272
rect 46902 325216 48116 325272
rect 46841 325214 48116 325216
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 46841 325211 46907 325214
rect 580165 325211 580231 325214
rect 407205 325138 407271 325141
rect 407205 325136 410044 325138
rect 407205 325080 407210 325136
rect 407266 325080 410044 325136
rect 583520 325124 584960 325214
rect 407205 325078 410044 325080
rect 407205 325075 407271 325078
rect 350809 324594 350875 324597
rect 347852 324592 350875 324594
rect 347852 324536 350814 324592
rect 350870 324536 350875 324592
rect 347852 324534 350875 324536
rect 350809 324531 350875 324534
rect 407205 323778 407271 323781
rect 552933 323778 552999 323781
rect 407205 323776 410044 323778
rect 407205 323720 407210 323776
rect 407266 323720 410044 323776
rect 407205 323718 410044 323720
rect 549884 323776 552999 323778
rect 549884 323720 552938 323776
rect 552994 323720 552999 323776
rect 549884 323718 552999 323720
rect 407205 323715 407271 323718
rect 552933 323715 552999 323718
rect 46841 323098 46907 323101
rect 48086 323098 48146 323136
rect 46841 323096 48146 323098
rect 46841 323040 46846 323096
rect 46902 323040 48146 323096
rect 46841 323038 48146 323040
rect 407113 323098 407179 323101
rect 407113 323096 410044 323098
rect 407113 323040 407118 323096
rect 407174 323040 410044 323096
rect 407113 323038 410044 323040
rect 46841 323035 46907 323038
rect 407113 323035 407179 323038
rect 407113 322418 407179 322421
rect 552013 322418 552079 322421
rect 407113 322416 410044 322418
rect 407113 322360 407118 322416
rect 407174 322360 410044 322416
rect 407113 322358 410044 322360
rect 549884 322416 552079 322418
rect 549884 322360 552018 322416
rect 552074 322360 552079 322416
rect 549884 322358 552079 322360
rect 407113 322355 407179 322358
rect 552013 322355 552079 322358
rect 46841 321738 46907 321741
rect 48086 321738 48146 321776
rect 46841 321736 48146 321738
rect 46841 321680 46846 321736
rect 46902 321680 48146 321736
rect 46841 321678 48146 321680
rect 347822 321738 347882 321776
rect 350349 321738 350415 321741
rect 347822 321736 350415 321738
rect 347822 321680 350354 321736
rect 350410 321680 350415 321736
rect 347822 321678 350415 321680
rect 46841 321675 46907 321678
rect 350349 321675 350415 321678
rect 407205 321738 407271 321741
rect 407205 321736 410044 321738
rect 407205 321680 407210 321736
rect 407266 321680 410044 321736
rect 407205 321678 410044 321680
rect 407205 321675 407271 321678
rect 347822 320650 347882 321096
rect 407113 321058 407179 321061
rect 407113 321056 410044 321058
rect 407113 321000 407118 321056
rect 407174 321000 410044 321056
rect 407113 320998 410044 321000
rect 407113 320995 407179 320998
rect 350349 320650 350415 320653
rect 347822 320648 350415 320650
rect 347822 320592 350354 320648
rect 350410 320592 350415 320648
rect 347822 320590 350415 320592
rect 350349 320587 350415 320590
rect 46841 320242 46907 320245
rect 48086 320242 48146 320416
rect 46841 320240 48146 320242
rect 46841 320184 46846 320240
rect 46902 320184 48146 320240
rect 46841 320182 48146 320184
rect 46841 320179 46907 320182
rect -960 319140 480 319380
rect 347822 319290 347882 319736
rect 409045 319698 409111 319701
rect 409045 319696 410044 319698
rect 409045 319640 409050 319696
rect 409106 319640 410044 319696
rect 409045 319638 410044 319640
rect 409045 319635 409111 319638
rect 350349 319290 350415 319293
rect 347822 319288 350415 319290
rect 347822 319232 350354 319288
rect 350410 319232 350415 319288
rect 347822 319230 350415 319232
rect 350349 319227 350415 319230
rect 350165 319154 350231 319157
rect 347852 319152 350231 319154
rect 347852 319096 350170 319152
rect 350226 319096 350231 319152
rect 347852 319094 350231 319096
rect 350165 319091 350231 319094
rect 46841 319018 46907 319021
rect 48086 319018 48146 319056
rect 46841 319016 48146 319018
rect 46841 318960 46846 319016
rect 46902 318960 48146 319016
rect 46841 318958 48146 318960
rect 407389 319018 407455 319021
rect 407389 319016 410044 319018
rect 407389 318960 407394 319016
rect 407450 318960 410044 319016
rect 407389 318958 410044 318960
rect 46841 318955 46907 318958
rect 407389 318955 407455 318958
rect 46841 318474 46907 318477
rect 46841 318472 48116 318474
rect 46841 318416 46846 318472
rect 46902 318416 48116 318472
rect 46841 318414 48116 318416
rect 46841 318411 46907 318414
rect 347822 317794 347882 318376
rect 407113 318338 407179 318341
rect 552933 318338 552999 318341
rect 407113 318336 410044 318338
rect 407113 318280 407118 318336
rect 407174 318280 410044 318336
rect 407113 318278 410044 318280
rect 549884 318336 552999 318338
rect 549884 318280 552938 318336
rect 552994 318280 552999 318336
rect 549884 318278 552999 318280
rect 407113 318275 407179 318278
rect 552933 318275 552999 318278
rect 350349 317794 350415 317797
rect 347822 317792 350415 317794
rect 347822 317736 350354 317792
rect 350410 317736 350415 317792
rect 347822 317734 350415 317736
rect 350349 317731 350415 317734
rect 553117 317658 553183 317661
rect 549884 317656 553183 317658
rect 549884 317600 553122 317656
rect 553178 317600 553183 317656
rect 549884 317598 553183 317600
rect 553117 317595 553183 317598
rect 43437 317386 43503 317389
rect 44950 317386 44956 317388
rect 43437 317384 44956 317386
rect 43437 317328 43442 317384
rect 43498 317328 44956 317384
rect 43437 317326 44956 317328
rect 43437 317323 43503 317326
rect 44950 317324 44956 317326
rect 45020 317324 45026 317388
rect 409454 316916 409460 316980
rect 409524 316978 409530 316980
rect 409524 316918 410044 316978
rect 409524 316916 409530 316918
rect 553117 316298 553183 316301
rect 549884 316296 553183 316298
rect 549884 316240 553122 316296
rect 553178 316240 553183 316296
rect 549884 316238 553183 316240
rect 553117 316235 553183 316238
rect 347822 315210 347882 315656
rect 409873 315618 409939 315621
rect 553710 315618 553716 315620
rect 409873 315616 410044 315618
rect 409873 315560 409878 315616
rect 409934 315560 410044 315616
rect 409873 315558 410044 315560
rect 549884 315558 553716 315618
rect 409873 315555 409939 315558
rect 553710 315556 553716 315558
rect 553780 315556 553786 315620
rect 350165 315210 350231 315213
rect 347822 315208 350231 315210
rect 347822 315152 350170 315208
rect 350226 315152 350231 315208
rect 347822 315150 350231 315152
rect 350165 315147 350231 315150
rect 350349 315074 350415 315077
rect 347852 315072 350415 315074
rect 347852 315016 350354 315072
rect 350410 315016 350415 315072
rect 347852 315014 350415 315016
rect 350349 315011 350415 315014
rect 46841 314802 46907 314805
rect 48086 314802 48146 314976
rect 552565 314938 552631 314941
rect 549884 314936 552631 314938
rect 549884 314880 552570 314936
rect 552626 314880 552631 314936
rect 549884 314878 552631 314880
rect 552565 314875 552631 314878
rect 46841 314800 48146 314802
rect 46841 314744 46846 314800
rect 46902 314744 48146 314800
rect 46841 314742 48146 314744
rect 46841 314739 46907 314742
rect 552933 314258 552999 314261
rect 549884 314256 552999 314258
rect 549884 314200 552938 314256
rect 552994 314200 552999 314256
rect 549884 314198 552999 314200
rect 552933 314195 552999 314198
rect 43478 313244 43484 313308
rect 43548 313306 43554 313308
rect 44766 313306 44772 313308
rect 43548 313246 44772 313306
rect 43548 313244 43554 313246
rect 44766 313244 44772 313246
rect 44836 313244 44842 313308
rect 347822 312354 347882 312936
rect 407113 312898 407179 312901
rect 553117 312898 553183 312901
rect 407113 312896 410044 312898
rect 407113 312840 407118 312896
rect 407174 312840 410044 312896
rect 407113 312838 410044 312840
rect 549884 312896 553183 312898
rect 549884 312840 553122 312896
rect 553178 312840 553183 312896
rect 549884 312838 553183 312840
rect 407113 312835 407179 312838
rect 553117 312835 553183 312838
rect 350349 312354 350415 312357
rect 347822 312352 350415 312354
rect 347822 312296 350354 312352
rect 350410 312296 350415 312352
rect 347822 312294 350415 312296
rect 350349 312291 350415 312294
rect 580533 312082 580599 312085
rect 583520 312082 584960 312172
rect 580533 312080 584960 312082
rect 580533 312024 580538 312080
rect 580594 312024 584960 312080
rect 580533 312022 584960 312024
rect 580533 312019 580599 312022
rect 387742 311884 387748 311948
rect 387812 311946 387818 311948
rect 389081 311946 389147 311949
rect 387812 311944 389147 311946
rect 387812 311888 389086 311944
rect 389142 311888 389147 311944
rect 583520 311932 584960 312022
rect 387812 311886 389147 311888
rect 387812 311884 387818 311886
rect 389081 311883 389147 311886
rect 46841 310994 46907 310997
rect 48086 310994 48146 311576
rect 347822 311130 347882 311576
rect 350349 311130 350415 311133
rect 347822 311128 350415 311130
rect 347822 311072 350354 311128
rect 350410 311072 350415 311128
rect 347822 311070 350415 311072
rect 350349 311067 350415 311070
rect 407205 311130 407271 311133
rect 410014 311130 410074 311440
rect 549884 311410 550282 311470
rect 550222 311402 550282 311410
rect 552933 311402 552999 311405
rect 550222 311400 552999 311402
rect 550222 311344 552938 311400
rect 552994 311344 552999 311400
rect 550222 311342 552999 311344
rect 552933 311339 552999 311342
rect 407205 311128 410074 311130
rect 407205 311072 407210 311128
rect 407266 311072 410074 311128
rect 407205 311070 410074 311072
rect 407205 311067 407271 311070
rect 46841 310992 48146 310994
rect 46841 310936 46846 310992
rect 46902 310936 48146 310992
rect 46841 310934 48146 310936
rect 46841 310931 46907 310934
rect 407113 310858 407179 310861
rect 553117 310858 553183 310861
rect 407113 310856 410044 310858
rect 407113 310800 407118 310856
rect 407174 310800 410044 310856
rect 407113 310798 410044 310800
rect 549884 310856 553183 310858
rect 549884 310800 553122 310856
rect 553178 310800 553183 310856
rect 549884 310798 553183 310800
rect 407113 310795 407179 310798
rect 553117 310795 553183 310798
rect 44909 310314 44975 310317
rect 44909 310312 48116 310314
rect 44909 310256 44914 310312
rect 44970 310256 48116 310312
rect 44909 310254 48116 310256
rect 44909 310251 44975 310254
rect 407113 310178 407179 310181
rect 553117 310178 553183 310181
rect 407113 310176 410044 310178
rect 407113 310120 407118 310176
rect 407174 310120 410044 310176
rect 407113 310118 410044 310120
rect 549884 310176 553183 310178
rect 549884 310120 553122 310176
rect 553178 310120 553183 310176
rect 549884 310118 553183 310120
rect 407113 310115 407179 310118
rect 553117 310115 553183 310118
rect 46841 309226 46907 309229
rect 48086 309226 48146 309536
rect 46841 309224 48146 309226
rect 46841 309168 46846 309224
rect 46902 309168 48146 309224
rect 46841 309166 48146 309168
rect 46841 309163 46907 309166
rect 347822 308410 347882 308856
rect 553117 308818 553183 308821
rect 549884 308816 553183 308818
rect 549884 308760 553122 308816
rect 553178 308760 553183 308816
rect 549884 308758 553183 308760
rect 553117 308755 553183 308758
rect 350349 308410 350415 308413
rect 347822 308408 350415 308410
rect 347822 308352 350354 308408
rect 350410 308352 350415 308408
rect 347822 308350 350415 308352
rect 350349 308347 350415 308350
rect 407113 308138 407179 308141
rect 407113 308136 410044 308138
rect 407113 308080 407118 308136
rect 407174 308080 410044 308136
rect 407113 308078 410044 308080
rect 407113 308075 407179 308078
rect 552013 307458 552079 307461
rect 549884 307456 552079 307458
rect 549884 307400 552018 307456
rect 552074 307400 552079 307456
rect 549884 307398 552079 307400
rect 552013 307395 552079 307398
rect 407205 306778 407271 306781
rect 407205 306776 410044 306778
rect 407205 306720 407210 306776
rect 407266 306720 410044 306776
rect 407205 306718 410044 306720
rect 407205 306715 407271 306718
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 406142 306036 406148 306100
rect 406212 306098 406218 306100
rect 552289 306098 552355 306101
rect 406212 306038 410044 306098
rect 549884 306096 552355 306098
rect 549884 306040 552294 306096
rect 552350 306040 552355 306096
rect 549884 306038 552355 306040
rect 406212 306036 406218 306038
rect 552289 306035 552355 306038
rect 407113 305418 407179 305421
rect 553117 305418 553183 305421
rect 407113 305416 410044 305418
rect 407113 305360 407118 305416
rect 407174 305360 410044 305416
rect 407113 305358 410044 305360
rect 549884 305416 553183 305418
rect 549884 305360 553122 305416
rect 553178 305360 553183 305416
rect 549884 305358 553183 305360
rect 407113 305355 407179 305358
rect 553117 305355 553183 305358
rect 352649 305010 352715 305013
rect 354438 305010 354444 305012
rect 352649 305008 354444 305010
rect 352649 304952 352654 305008
rect 352710 304952 354444 305008
rect 352649 304950 354444 304952
rect 352649 304947 352715 304950
rect 354438 304948 354444 304950
rect 354508 304948 354514 305012
rect 347822 304330 347882 304776
rect 350349 304330 350415 304333
rect 347822 304328 350415 304330
rect 347822 304272 350354 304328
rect 350410 304272 350415 304328
rect 347822 304270 350415 304272
rect 350349 304267 350415 304270
rect 46841 303786 46907 303789
rect 48086 303786 48146 304096
rect 407113 304058 407179 304061
rect 407113 304056 410044 304058
rect 407113 304000 407118 304056
rect 407174 304000 410044 304056
rect 407113 303998 410044 304000
rect 407113 303995 407179 303998
rect 46841 303784 48146 303786
rect 46841 303728 46846 303784
rect 46902 303728 48146 303784
rect 46841 303726 48146 303728
rect 46841 303723 46907 303726
rect 46473 302970 46539 302973
rect 48086 302970 48146 303416
rect 46473 302968 48146 302970
rect 46473 302912 46478 302968
rect 46534 302912 48146 302968
rect 46473 302910 48146 302912
rect 347822 302970 347882 303416
rect 349889 302970 349955 302973
rect 347822 302968 349955 302970
rect 347822 302912 349894 302968
rect 349950 302912 349955 302968
rect 347822 302910 349955 302912
rect 46473 302907 46539 302910
rect 349889 302907 349955 302910
rect 347822 302426 347882 302736
rect 407389 302698 407455 302701
rect 407389 302696 410044 302698
rect 407389 302640 407394 302696
rect 407450 302640 410044 302696
rect 407389 302638 410044 302640
rect 407389 302635 407455 302638
rect 350349 302426 350415 302429
rect 347822 302424 350415 302426
rect 347822 302368 350354 302424
rect 350410 302368 350415 302424
rect 347822 302366 350415 302368
rect 350349 302363 350415 302366
rect 372654 302228 372660 302292
rect 372724 302290 372730 302292
rect 373901 302290 373967 302293
rect 372724 302288 373967 302290
rect 372724 302232 373906 302288
rect 373962 302232 373967 302288
rect 372724 302230 373967 302232
rect 372724 302228 372730 302230
rect 373901 302227 373967 302230
rect 46841 302154 46907 302157
rect 46841 302152 48116 302154
rect 46841 302096 46846 302152
rect 46902 302096 48116 302152
rect 46841 302094 48116 302096
rect 46841 302091 46907 302094
rect 407205 302018 407271 302021
rect 553117 302018 553183 302021
rect 407205 302016 410044 302018
rect 407205 301960 407210 302016
rect 407266 301960 410044 302016
rect 407205 301958 410044 301960
rect 549884 302016 553183 302018
rect 549884 301960 553122 302016
rect 553178 301960 553183 302016
rect 549884 301958 553183 301960
rect 407205 301955 407271 301958
rect 553117 301955 553183 301958
rect 46841 300930 46907 300933
rect 48086 300930 48146 301376
rect 46841 300928 48146 300930
rect 46841 300872 46846 300928
rect 46902 300872 48146 300928
rect 46841 300870 48146 300872
rect 347822 300930 347882 301376
rect 407113 301338 407179 301341
rect 552657 301338 552723 301341
rect 407113 301336 410044 301338
rect 407113 301280 407118 301336
rect 407174 301280 410044 301336
rect 407113 301278 410044 301280
rect 549884 301336 552723 301338
rect 549884 301280 552662 301336
rect 552718 301280 552723 301336
rect 549884 301278 552723 301280
rect 407113 301275 407179 301278
rect 552657 301275 552723 301278
rect 350349 300930 350415 300933
rect 347822 300928 350415 300930
rect 347822 300872 350354 300928
rect 350410 300872 350415 300928
rect 347822 300870 350415 300872
rect 46841 300867 46907 300870
rect 350349 300867 350415 300870
rect 347822 300250 347882 300696
rect 409321 300658 409387 300661
rect 553117 300658 553183 300661
rect 409321 300656 410044 300658
rect 409321 300600 409326 300656
rect 409382 300600 410044 300656
rect 409321 300598 410044 300600
rect 549884 300656 553183 300658
rect 549884 300600 553122 300656
rect 553178 300600 553183 300656
rect 549884 300598 553183 300600
rect 409321 300595 409387 300598
rect 553117 300595 553183 300598
rect 350349 300250 350415 300253
rect 347822 300248 350415 300250
rect 347822 300192 350354 300248
rect 350410 300192 350415 300248
rect 347822 300190 350415 300192
rect 350349 300187 350415 300190
rect 407113 299978 407179 299981
rect 407113 299976 410044 299978
rect 407113 299920 407118 299976
rect 407174 299920 410044 299976
rect 407113 299918 410044 299920
rect 407113 299915 407179 299918
rect 348550 299372 348556 299436
rect 348620 299434 348626 299436
rect 349153 299434 349219 299437
rect 348620 299432 349219 299434
rect 348620 299376 349158 299432
rect 349214 299376 349219 299432
rect 348620 299374 349219 299376
rect 348620 299372 348626 299374
rect 349153 299371 349219 299374
rect 347822 298890 347882 299336
rect 350349 298890 350415 298893
rect 347822 298888 350415 298890
rect 347822 298832 350354 298888
rect 350410 298832 350415 298888
rect 347822 298830 350415 298832
rect 350349 298827 350415 298830
rect 46841 298210 46907 298213
rect 48086 298210 48146 298656
rect 407665 298618 407731 298621
rect 407665 298616 410044 298618
rect 407665 298560 407670 298616
rect 407726 298560 410044 298616
rect 583520 298604 584960 298844
rect 407665 298558 410044 298560
rect 407665 298555 407731 298558
rect 46841 298208 48146 298210
rect 46841 298152 46846 298208
rect 46902 298152 48146 298208
rect 46841 298150 48146 298152
rect 46841 298147 46907 298150
rect 47301 298074 47367 298077
rect 47301 298072 48116 298074
rect 47301 298016 47306 298072
rect 47362 298016 48116 298072
rect 47301 298014 48116 298016
rect 47301 298011 47367 298014
rect 553117 297938 553183 297941
rect 549884 297936 553183 297938
rect 549884 297880 553122 297936
rect 553178 297880 553183 297936
rect 549884 297878 553183 297880
rect 553117 297875 553183 297878
rect 46841 296850 46907 296853
rect 48086 296850 48146 297296
rect 553117 297258 553183 297261
rect 549884 297256 553183 297258
rect 549884 297200 553122 297256
rect 553178 297200 553183 297256
rect 549884 297198 553183 297200
rect 553117 297195 553183 297198
rect 46841 296848 48146 296850
rect 46841 296792 46846 296848
rect 46902 296792 48146 296848
rect 46841 296790 48146 296792
rect 46841 296787 46907 296790
rect 349429 296714 349495 296717
rect 347852 296712 349495 296714
rect 347852 296656 349434 296712
rect 349490 296656 349495 296712
rect 347852 296654 349495 296656
rect 349429 296651 349495 296654
rect 348325 296034 348391 296037
rect 347852 296032 348391 296034
rect 347852 295976 348330 296032
rect 348386 295976 348391 296032
rect 347852 295974 348391 295976
rect 348325 295971 348391 295974
rect 407113 295898 407179 295901
rect 407113 295896 410044 295898
rect 407113 295840 407118 295896
rect 407174 295840 410044 295896
rect 407113 295838 410044 295840
rect 407113 295835 407179 295838
rect 350257 295354 350323 295357
rect 347852 295352 350323 295354
rect 347852 295296 350262 295352
rect 350318 295296 350323 295352
rect 347852 295294 350323 295296
rect 350257 295291 350323 295294
rect 350257 293994 350323 293997
rect 347852 293992 350323 293994
rect 347852 293936 350262 293992
rect 350318 293936 350323 293992
rect 347852 293934 350323 293936
rect 350257 293931 350323 293934
rect 409321 293994 409387 293997
rect 410014 293994 410074 294440
rect 409321 293992 410074 293994
rect 409321 293936 409326 293992
rect 409382 293936 410074 293992
rect 409321 293934 410074 293936
rect 409321 293931 409387 293934
rect 407205 293858 407271 293861
rect 407205 293856 410044 293858
rect 407205 293800 407210 293856
rect 407266 293800 410044 293856
rect 407205 293798 410044 293800
rect 407205 293795 407271 293798
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 46841 292906 46907 292909
rect 48086 292906 48146 293216
rect 407113 293178 407179 293181
rect 552013 293178 552079 293181
rect 407113 293176 410044 293178
rect 407113 293120 407118 293176
rect 407174 293120 410044 293176
rect 407113 293118 410044 293120
rect 549884 293176 552079 293178
rect 549884 293120 552018 293176
rect 552074 293120 552079 293176
rect 549884 293118 552079 293120
rect 407113 293115 407179 293118
rect 552013 293115 552079 293118
rect 46841 292904 48146 292906
rect 46841 292848 46846 292904
rect 46902 292848 48146 292904
rect 46841 292846 48146 292848
rect 46841 292843 46907 292846
rect 46473 292634 46539 292637
rect 46473 292632 48116 292634
rect 46473 292576 46478 292632
rect 46534 292576 48116 292632
rect 46473 292574 48116 292576
rect 46473 292571 46539 292574
rect 407113 292498 407179 292501
rect 553117 292498 553183 292501
rect 407113 292496 410044 292498
rect 407113 292440 407118 292496
rect 407174 292440 410044 292496
rect 407113 292438 410044 292440
rect 549884 292496 553183 292498
rect 549884 292440 553122 292496
rect 553178 292440 553183 292496
rect 549884 292438 553183 292440
rect 407113 292435 407179 292438
rect 553117 292435 553183 292438
rect 46841 291546 46907 291549
rect 48086 291546 48146 291856
rect 407205 291818 407271 291821
rect 552197 291818 552263 291821
rect 407205 291816 410044 291818
rect 407205 291760 407210 291816
rect 407266 291760 410044 291816
rect 407205 291758 410044 291760
rect 549884 291816 552263 291818
rect 549884 291760 552202 291816
rect 552258 291760 552263 291816
rect 549884 291758 552263 291760
rect 407205 291755 407271 291758
rect 552197 291755 552263 291758
rect 46841 291544 48146 291546
rect 46841 291488 46846 291544
rect 46902 291488 48146 291544
rect 46841 291486 48146 291488
rect 46841 291483 46907 291486
rect 552013 290458 552079 290461
rect 549884 290456 552079 290458
rect 549884 290400 552018 290456
rect 552074 290400 552079 290456
rect 549884 290398 552079 290400
rect 552013 290395 552079 290398
rect 409597 289778 409663 289781
rect 552933 289778 552999 289781
rect 409597 289776 410044 289778
rect 409597 289720 409602 289776
rect 409658 289720 410044 289776
rect 409597 289718 410044 289720
rect 549884 289776 552999 289778
rect 549884 289720 552938 289776
rect 552994 289720 552999 289776
rect 549884 289718 552999 289720
rect 409597 289715 409663 289718
rect 552933 289715 552999 289718
rect 347822 288690 347882 289136
rect 407113 289098 407179 289101
rect 553117 289098 553183 289101
rect 407113 289096 410044 289098
rect 407113 289040 407118 289096
rect 407174 289040 410044 289096
rect 407113 289038 410044 289040
rect 549884 289096 553183 289098
rect 549884 289040 553122 289096
rect 553178 289040 553183 289096
rect 549884 289038 553183 289040
rect 407113 289035 407179 289038
rect 553117 289035 553183 289038
rect 350257 288690 350323 288693
rect 347822 288688 350323 288690
rect 347822 288632 350262 288688
rect 350318 288632 350323 288688
rect 347822 288630 350323 288632
rect 350257 288627 350323 288630
rect 46841 288554 46907 288557
rect 350073 288554 350139 288557
rect 46841 288552 48116 288554
rect 46841 288496 46846 288552
rect 46902 288496 48116 288552
rect 46841 288494 48116 288496
rect 347852 288552 350139 288554
rect 347852 288496 350078 288552
rect 350134 288496 350139 288552
rect 347852 288494 350139 288496
rect 46841 288491 46907 288494
rect 350073 288491 350139 288494
rect 407113 288418 407179 288421
rect 407113 288416 410044 288418
rect 407113 288360 407118 288416
rect 407174 288360 410044 288416
rect 407113 288358 410044 288360
rect 407113 288355 407179 288358
rect 347822 287194 347882 287776
rect 407205 287738 407271 287741
rect 550817 287738 550883 287741
rect 407205 287736 410044 287738
rect 407205 287680 407210 287736
rect 407266 287680 410044 287736
rect 407205 287678 410044 287680
rect 549884 287736 550883 287738
rect 549884 287680 550822 287736
rect 550878 287680 550883 287736
rect 549884 287678 550883 287680
rect 407205 287675 407271 287678
rect 550817 287675 550883 287678
rect 350257 287194 350323 287197
rect 347822 287192 350323 287194
rect 347822 287136 350262 287192
rect 350318 287136 350323 287192
rect 347822 287134 350323 287136
rect 350257 287131 350323 287134
rect 407113 287058 407179 287061
rect 407113 287056 410044 287058
rect 407113 287000 407118 287056
rect 407174 287000 410044 287056
rect 407113 286998 410044 287000
rect 407113 286995 407179 286998
rect 350257 286514 350323 286517
rect 347852 286512 350323 286514
rect 347852 286456 350262 286512
rect 350318 286456 350323 286512
rect 347852 286454 350323 286456
rect 350257 286451 350323 286454
rect 46841 285834 46907 285837
rect 48086 285834 48146 286416
rect 553117 286378 553183 286381
rect 549884 286376 553183 286378
rect 549884 286320 553122 286376
rect 553178 286320 553183 286376
rect 549884 286318 553183 286320
rect 553117 286315 553183 286318
rect 355501 285834 355567 285837
rect 46841 285832 48146 285834
rect 46841 285776 46846 285832
rect 46902 285776 48146 285832
rect 46841 285774 48146 285776
rect 347852 285832 355567 285834
rect 347852 285776 355506 285832
rect 355562 285776 355567 285832
rect 347852 285774 355567 285776
rect 46841 285771 46907 285774
rect 355501 285771 355567 285774
rect 44950 285228 44956 285292
rect 45020 285290 45026 285292
rect 46933 285290 46999 285293
rect 45020 285288 46999 285290
rect 45020 285232 46938 285288
rect 46994 285232 46999 285288
rect 583520 285276 584960 285516
rect 45020 285230 46999 285232
rect 45020 285228 45026 285230
rect 46933 285227 46999 285230
rect 350257 285154 350323 285157
rect 347852 285152 350323 285154
rect 347852 285096 350262 285152
rect 350318 285096 350323 285152
rect 347852 285094 350323 285096
rect 350257 285091 350323 285094
rect 407205 285018 407271 285021
rect 407205 285016 410044 285018
rect 407205 284960 407210 285016
rect 407266 284960 410044 285016
rect 407205 284958 410044 284960
rect 407205 284955 407271 284958
rect 46473 284338 46539 284341
rect 48086 284338 48146 284376
rect 46473 284336 48146 284338
rect 46473 284280 46478 284336
rect 46534 284280 48146 284336
rect 46473 284278 48146 284280
rect 347822 284338 347882 284376
rect 350625 284338 350691 284341
rect 347822 284336 350691 284338
rect 347822 284280 350630 284336
rect 350686 284280 350691 284336
rect 347822 284278 350691 284280
rect 46473 284275 46539 284278
rect 350625 284275 350691 284278
rect 407113 284338 407179 284341
rect 407113 284336 410044 284338
rect 407113 284280 407118 284336
rect 407174 284280 410044 284336
rect 407113 284278 410044 284280
rect 407113 284275 407179 284278
rect 44817 283250 44883 283253
rect 48086 283250 48146 283696
rect 407205 283658 407271 283661
rect 553117 283658 553183 283661
rect 407205 283656 410044 283658
rect 407205 283600 407210 283656
rect 407266 283600 410044 283656
rect 407205 283598 410044 283600
rect 549884 283656 553183 283658
rect 549884 283600 553122 283656
rect 553178 283600 553183 283656
rect 549884 283598 553183 283600
rect 407205 283595 407271 283598
rect 553117 283595 553183 283598
rect 44817 283248 48146 283250
rect 44817 283192 44822 283248
rect 44878 283192 48146 283248
rect 44817 283190 48146 283192
rect 44817 283187 44883 283190
rect 407113 282978 407179 282981
rect 407113 282976 410044 282978
rect 407113 282920 407118 282976
rect 407174 282920 410044 282976
rect 407113 282918 410044 282920
rect 407113 282915 407179 282918
rect 47393 281890 47459 281893
rect 48086 281890 48146 282336
rect 550633 282298 550699 282301
rect 549884 282296 550699 282298
rect 549884 282240 550638 282296
rect 550694 282240 550699 282296
rect 549884 282238 550699 282240
rect 550633 282235 550699 282238
rect 47393 281888 48146 281890
rect 47393 281832 47398 281888
rect 47454 281832 48146 281888
rect 47393 281830 48146 281832
rect 47393 281827 47459 281830
rect 46841 281618 46907 281621
rect 48086 281618 48146 281656
rect 553117 281618 553183 281621
rect 46841 281616 48146 281618
rect 46841 281560 46846 281616
rect 46902 281560 48146 281616
rect 46841 281558 48146 281560
rect 549884 281616 553183 281618
rect 549884 281560 553122 281616
rect 553178 281560 553183 281616
rect 549884 281558 553183 281560
rect 46841 281555 46907 281558
rect 553117 281555 553183 281558
rect 347822 280530 347882 280976
rect 553117 280938 553183 280941
rect 549884 280936 553183 280938
rect 549884 280880 553122 280936
rect 553178 280880 553183 280936
rect 549884 280878 553183 280880
rect 553117 280875 553183 280878
rect 349613 280530 349679 280533
rect 347822 280528 349679 280530
rect 347822 280472 349618 280528
rect 349674 280472 349679 280528
rect 347822 280470 349679 280472
rect 349613 280467 349679 280470
rect 553117 280258 553183 280261
rect 549884 280256 553183 280258
rect -960 279972 480 280212
rect 549884 280200 553122 280256
rect 553178 280200 553183 280256
rect 549884 280198 553183 280200
rect 553117 280195 553183 280198
rect 349337 279714 349403 279717
rect 347852 279712 349403 279714
rect 347852 279656 349342 279712
rect 349398 279656 349403 279712
rect 347852 279654 349403 279656
rect 349337 279651 349403 279654
rect 409229 279578 409295 279581
rect 552933 279578 552999 279581
rect 409229 279576 410044 279578
rect 409229 279520 409234 279576
rect 409290 279520 410044 279576
rect 409229 279518 410044 279520
rect 549884 279576 552999 279578
rect 549884 279520 552938 279576
rect 552994 279520 552999 279576
rect 549884 279518 552999 279520
rect 409229 279515 409295 279518
rect 552933 279515 552999 279518
rect 407113 278898 407179 278901
rect 553117 278898 553183 278901
rect 407113 278896 410044 278898
rect 407113 278840 407118 278896
rect 407174 278840 410044 278896
rect 407113 278838 410044 278840
rect 549884 278896 553183 278898
rect 549884 278840 553122 278896
rect 553178 278840 553183 278896
rect 549884 278838 553183 278840
rect 407113 278835 407179 278838
rect 553117 278835 553183 278838
rect 351126 278354 351132 278356
rect 347852 278294 351132 278354
rect 351126 278292 351132 278294
rect 351196 278292 351202 278356
rect 46841 277810 46907 277813
rect 48086 277810 48146 278256
rect 46841 277808 48146 277810
rect 46841 277752 46846 277808
rect 46902 277752 48146 277808
rect 46841 277750 48146 277752
rect 46841 277747 46907 277750
rect 347822 277538 347882 277576
rect 350257 277538 350323 277541
rect 347822 277536 350323 277538
rect 347822 277480 350262 277536
rect 350318 277480 350323 277536
rect 347822 277478 350323 277480
rect 350257 277475 350323 277478
rect 409638 277476 409644 277540
rect 409708 277538 409714 277540
rect 553117 277538 553183 277541
rect 409708 277478 410044 277538
rect 550222 277536 553183 277538
rect 550222 277480 553122 277536
rect 553178 277480 553183 277536
rect 550222 277478 553183 277480
rect 409708 277476 409714 277478
rect 550222 277470 550282 277478
rect 553117 277475 553183 277478
rect 549884 277410 550282 277470
rect 408033 276858 408099 276861
rect 408033 276856 410044 276858
rect 408033 276800 408038 276856
rect 408094 276800 410044 276856
rect 408033 276798 410044 276800
rect 408033 276795 408099 276798
rect 347822 276045 347882 276216
rect 407113 276178 407179 276181
rect 553117 276178 553183 276181
rect 407113 276176 410044 276178
rect 407113 276120 407118 276176
rect 407174 276120 410044 276176
rect 407113 276118 410044 276120
rect 549884 276176 553183 276178
rect 549884 276120 553122 276176
rect 553178 276120 553183 276176
rect 549884 276118 553183 276120
rect 407113 276115 407179 276118
rect 553117 276115 553183 276118
rect 40769 276042 40835 276045
rect 44766 276042 44772 276044
rect 40769 276040 44772 276042
rect 40769 275984 40774 276040
rect 40830 275984 44772 276040
rect 40769 275982 44772 275984
rect 40769 275979 40835 275982
rect 44766 275980 44772 275982
rect 44836 275980 44842 276044
rect 347822 276040 347931 276045
rect 347822 275984 347870 276040
rect 347926 275984 347931 276040
rect 347822 275982 347931 275984
rect 347865 275979 347931 275982
rect 350257 275634 350323 275637
rect 347852 275632 350323 275634
rect 347852 275576 350262 275632
rect 350318 275576 350323 275632
rect 347852 275574 350323 275576
rect 350257 275571 350323 275574
rect 407113 275498 407179 275501
rect 407113 275496 410044 275498
rect 407113 275440 407118 275496
rect 407174 275440 410044 275496
rect 407113 275438 410044 275440
rect 407113 275435 407179 275438
rect 552289 274818 552355 274821
rect 549884 274816 552355 274818
rect 549884 274760 552294 274816
rect 552350 274760 552355 274816
rect 549884 274758 552355 274760
rect 552289 274755 552355 274758
rect 31518 273668 31524 273732
rect 31588 273730 31594 273732
rect 48086 273730 48146 274176
rect 347822 273866 347882 274176
rect 350165 273866 350231 273869
rect 347822 273864 350231 273866
rect 347822 273808 350170 273864
rect 350226 273808 350231 273864
rect 347822 273806 350231 273808
rect 350165 273803 350231 273806
rect 31588 273670 48146 273730
rect 31588 273668 31594 273670
rect 47301 273322 47367 273325
rect 48086 273322 48146 273496
rect 347822 273458 347882 273496
rect 350257 273458 350323 273461
rect 553117 273458 553183 273461
rect 347822 273456 350323 273458
rect 347822 273400 350262 273456
rect 350318 273400 350323 273456
rect 347822 273398 350323 273400
rect 549884 273456 553183 273458
rect 549884 273400 553122 273456
rect 553178 273400 553183 273456
rect 549884 273398 553183 273400
rect 350257 273395 350323 273398
rect 553117 273395 553183 273398
rect 47301 273320 48146 273322
rect 47301 273264 47306 273320
rect 47362 273264 48146 273320
rect 47301 273262 48146 273264
rect 47301 273259 47367 273262
rect 347822 272234 347882 272816
rect 407113 272778 407179 272781
rect 407113 272776 410044 272778
rect 407113 272720 407118 272776
rect 407174 272720 410044 272776
rect 407113 272718 410044 272720
rect 407113 272715 407179 272718
rect 350257 272234 350323 272237
rect 347822 272232 350323 272234
rect 347822 272176 350262 272232
rect 350318 272176 350323 272232
rect 347822 272174 350323 272176
rect 350257 272171 350323 272174
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 407205 271418 407271 271421
rect 550725 271418 550791 271421
rect 407205 271416 410044 271418
rect 407205 271360 407210 271416
rect 407266 271360 410044 271416
rect 407205 271358 410044 271360
rect 549884 271416 550791 271418
rect 549884 271360 550730 271416
rect 550786 271360 550791 271416
rect 549884 271358 550791 271360
rect 407205 271355 407271 271358
rect 550725 271355 550791 271358
rect 553117 270738 553183 270741
rect 549884 270736 553183 270738
rect 549884 270680 553122 270736
rect 553178 270680 553183 270736
rect 549884 270678 553183 270680
rect 553117 270675 553183 270678
rect 47117 270194 47183 270197
rect 350257 270194 350323 270197
rect 47117 270192 48116 270194
rect 47117 270136 47122 270192
rect 47178 270136 48116 270192
rect 47117 270134 48116 270136
rect 347852 270192 350323 270194
rect 347852 270136 350262 270192
rect 350318 270136 350323 270192
rect 347852 270134 350323 270136
rect 47117 270131 47183 270134
rect 350257 270131 350323 270134
rect 407113 270058 407179 270061
rect 407113 270056 410044 270058
rect 407113 270000 407118 270056
rect 407174 270000 410044 270056
rect 407113 269998 410044 270000
rect 407113 269995 407179 269998
rect 350257 268834 350323 268837
rect 347852 268832 350323 268834
rect 347852 268776 350262 268832
rect 350318 268776 350323 268832
rect 347852 268774 350323 268776
rect 350257 268771 350323 268774
rect 46841 268290 46907 268293
rect 48086 268290 48146 268736
rect 553117 268698 553183 268701
rect 549884 268696 553183 268698
rect 549884 268640 553122 268696
rect 553178 268640 553183 268696
rect 549884 268638 553183 268640
rect 553117 268635 553183 268638
rect 46841 268288 48146 268290
rect 46841 268232 46846 268288
rect 46902 268232 48146 268288
rect 46841 268230 48146 268232
rect 46841 268227 46907 268230
rect 350942 268154 350948 268156
rect 347852 268094 350948 268154
rect 350942 268092 350948 268094
rect 351012 268092 351018 268156
rect 35382 267956 35388 268020
rect 35452 268018 35458 268020
rect 48086 268018 48146 268056
rect 35452 267958 48146 268018
rect 407113 268018 407179 268021
rect 407113 268016 410044 268018
rect 407113 267960 407118 268016
rect 407174 267960 410044 268016
rect 407113 267958 410044 267960
rect 35452 267956 35458 267958
rect 407113 267955 407179 267958
rect -960 267052 480 267292
rect 347822 266794 347882 267376
rect 407757 267338 407823 267341
rect 407757 267336 410044 267338
rect 407757 267280 407762 267336
rect 407818 267280 410044 267336
rect 407757 267278 410044 267280
rect 407757 267275 407823 267278
rect 350257 266794 350323 266797
rect 347822 266792 350323 266794
rect 347822 266736 350262 266792
rect 350318 266736 350323 266792
rect 347822 266734 350323 266736
rect 350257 266731 350323 266734
rect 550265 266658 550331 266661
rect 549884 266656 550331 266658
rect 549884 266600 550270 266656
rect 550326 266600 550331 266656
rect 549884 266598 550331 266600
rect 550265 266595 550331 266598
rect 553117 265298 553183 265301
rect 549884 265296 553183 265298
rect 549884 265240 553122 265296
rect 553178 265240 553183 265296
rect 549884 265238 553183 265240
rect 553117 265235 553183 265238
rect 44173 264890 44239 264893
rect 44582 264890 44588 264892
rect 44173 264888 44588 264890
rect 44173 264832 44178 264888
rect 44234 264832 44588 264888
rect 44173 264830 44588 264832
rect 44173 264827 44239 264830
rect 44582 264828 44588 264830
rect 44652 264828 44658 264892
rect 45093 264754 45159 264757
rect 45093 264752 48116 264754
rect 45093 264696 45098 264752
rect 45154 264696 48116 264752
rect 45093 264694 48116 264696
rect 45093 264691 45159 264694
rect 43478 264556 43484 264620
rect 43548 264618 43554 264620
rect 45829 264618 45895 264621
rect 552933 264618 552999 264621
rect 43548 264616 45895 264618
rect 43548 264560 45834 264616
rect 45890 264560 45895 264616
rect 43548 264558 45895 264560
rect 549884 264616 552999 264618
rect 549884 264560 552938 264616
rect 552994 264560 552999 264616
rect 549884 264558 552999 264560
rect 43548 264556 43554 264558
rect 45829 264555 45895 264558
rect 552933 264555 552999 264558
rect 347822 263938 347882 263976
rect 350257 263938 350323 263941
rect 347822 263936 350323 263938
rect 347822 263880 350262 263936
rect 350318 263880 350323 263936
rect 347822 263878 350323 263880
rect 350257 263875 350323 263878
rect 407113 263938 407179 263941
rect 553117 263938 553183 263941
rect 407113 263936 410044 263938
rect 407113 263880 407118 263936
rect 407174 263880 410044 263936
rect 407113 263878 410044 263880
rect 549884 263936 553183 263938
rect 549884 263880 553122 263936
rect 553178 263880 553183 263936
rect 549884 263878 553183 263880
rect 407113 263875 407179 263878
rect 553117 263875 553183 263878
rect 347822 262850 347882 263296
rect 552013 263258 552079 263261
rect 549884 263256 552079 263258
rect 549884 263200 552018 263256
rect 552074 263200 552079 263256
rect 549884 263198 552079 263200
rect 552013 263195 552079 263198
rect 406561 262986 406627 262989
rect 409086 262986 409092 262988
rect 406561 262984 409092 262986
rect 406561 262928 406566 262984
rect 406622 262928 409092 262984
rect 406561 262926 409092 262928
rect 406561 262923 406627 262926
rect 409086 262924 409092 262926
rect 409156 262924 409162 262988
rect 349429 262850 349495 262853
rect 347822 262848 349495 262850
rect 347822 262792 349434 262848
rect 349490 262792 349495 262848
rect 347822 262790 349495 262792
rect 349429 262787 349495 262790
rect 349245 262714 349311 262717
rect 347852 262712 349311 262714
rect 347852 262656 349250 262712
rect 349306 262656 349311 262712
rect 347852 262654 349311 262656
rect 349245 262651 349311 262654
rect 36486 262244 36492 262308
rect 36556 262306 36562 262308
rect 48086 262306 48146 262616
rect 407113 262578 407179 262581
rect 550357 262578 550423 262581
rect 407113 262576 410044 262578
rect 407113 262520 407118 262576
rect 407174 262520 410044 262576
rect 407113 262518 410044 262520
rect 549884 262576 550423 262578
rect 549884 262520 550362 262576
rect 550418 262520 550423 262576
rect 549884 262518 550423 262520
rect 407113 262515 407179 262518
rect 550357 262515 550423 262518
rect 36556 262246 48146 262306
rect 36556 262244 36562 262246
rect 406326 262108 406332 262172
rect 406396 262170 406402 262172
rect 407481 262170 407547 262173
rect 406396 262168 407547 262170
rect 406396 262112 407486 262168
rect 407542 262112 407547 262168
rect 406396 262110 407547 262112
rect 406396 262108 406402 262110
rect 407481 262107 407547 262110
rect 407113 261898 407179 261901
rect 553117 261898 553183 261901
rect 407113 261896 410044 261898
rect 407113 261840 407118 261896
rect 407174 261840 410044 261896
rect 407113 261838 410044 261840
rect 549884 261896 553183 261898
rect 549884 261840 553122 261896
rect 553178 261840 553183 261896
rect 549884 261838 553183 261840
rect 407113 261835 407179 261838
rect 553117 261835 553183 261838
rect 350257 261354 350323 261357
rect 347852 261352 350323 261354
rect 347852 261296 350262 261352
rect 350318 261296 350323 261352
rect 347852 261294 350323 261296
rect 350257 261291 350323 261294
rect 408401 259994 408467 259997
rect 410014 259994 410074 260440
rect 549884 260410 550282 260470
rect 550222 260402 550282 260410
rect 552933 260402 552999 260405
rect 550222 260400 552999 260402
rect 550222 260344 552938 260400
rect 552994 260344 552999 260400
rect 550222 260342 552999 260344
rect 552933 260339 552999 260342
rect 408401 259992 410074 259994
rect 408401 259936 408406 259992
rect 408462 259936 410074 259992
rect 408401 259934 410074 259936
rect 408401 259931 408467 259934
rect 407113 259858 407179 259861
rect 553117 259858 553183 259861
rect 407113 259856 410044 259858
rect 407113 259800 407118 259856
rect 407174 259800 410044 259856
rect 407113 259798 410044 259800
rect 549884 259856 553183 259858
rect 549884 259800 553122 259856
rect 553178 259800 553183 259856
rect 549884 259798 553183 259800
rect 407113 259795 407179 259798
rect 553117 259795 553183 259798
rect 44766 259524 44772 259588
rect 44836 259586 44842 259588
rect 47485 259586 47551 259589
rect 44836 259584 47551 259586
rect 44836 259528 47490 259584
rect 47546 259528 47551 259584
rect 44836 259526 47551 259528
rect 44836 259524 44842 259526
rect 47485 259523 47551 259526
rect 347822 258770 347882 259216
rect 553117 259178 553183 259181
rect 549884 259176 553183 259178
rect 549884 259120 553122 259176
rect 553178 259120 553183 259176
rect 549884 259118 553183 259120
rect 553117 259115 553183 259118
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 349521 258770 349587 258773
rect 347822 258768 349587 258770
rect 347822 258712 349526 258768
rect 349582 258712 349587 258768
rect 583520 258756 584960 258846
rect 347822 258710 349587 258712
rect 349521 258707 349587 258710
rect 44950 258164 44956 258228
rect 45020 258226 45026 258228
rect 48086 258226 48146 258536
rect 553393 258498 553459 258501
rect 549884 258496 553459 258498
rect 549884 258440 553398 258496
rect 553454 258440 553459 258496
rect 549884 258438 553459 258440
rect 553393 258435 553459 258438
rect 45020 258166 48146 258226
rect 45020 258164 45026 258166
rect 45277 257954 45343 257957
rect 349705 257954 349771 257957
rect 45277 257952 48116 257954
rect 45277 257896 45282 257952
rect 45338 257896 48116 257952
rect 45277 257894 48116 257896
rect 347852 257952 349771 257954
rect 347852 257896 349710 257952
rect 349766 257896 349771 257952
rect 347852 257894 349771 257896
rect 45277 257891 45343 257894
rect 349705 257891 349771 257894
rect 407205 257818 407271 257821
rect 553117 257818 553183 257821
rect 407205 257816 410044 257818
rect 407205 257760 407210 257816
rect 407266 257760 410044 257816
rect 407205 257758 410044 257760
rect 549884 257816 553183 257818
rect 549884 257760 553122 257816
rect 553178 257760 553183 257816
rect 549884 257758 553183 257760
rect 407205 257755 407271 257758
rect 553117 257755 553183 257758
rect 45921 256730 45987 256733
rect 48086 256730 48146 257176
rect 407113 257138 407179 257141
rect 407113 257136 410044 257138
rect 407113 257080 407118 257136
rect 407174 257080 410044 257136
rect 407113 257078 410044 257080
rect 407113 257075 407179 257078
rect 45921 256728 48146 256730
rect 45921 256672 45926 256728
rect 45982 256672 48146 256728
rect 45921 256670 48146 256672
rect 45921 256667 45987 256670
rect 347822 256050 347882 256496
rect 349981 256050 350047 256053
rect 347822 256048 350047 256050
rect 347822 255992 349986 256048
rect 350042 255992 350047 256048
rect 347822 255990 350047 255992
rect 349981 255987 350047 255990
rect 347822 255370 347882 255816
rect 350441 255370 350507 255373
rect 347822 255368 350507 255370
rect 347822 255312 350446 255368
rect 350502 255312 350507 255368
rect 347822 255310 350507 255312
rect 350441 255307 350507 255310
rect 407113 255098 407179 255101
rect 552933 255098 552999 255101
rect 407113 255096 410044 255098
rect 407113 255040 407118 255096
rect 407174 255040 410044 255096
rect 407113 255038 410044 255040
rect 549884 255096 552999 255098
rect 549884 255040 552938 255096
rect 552994 255040 552999 255096
rect 549884 255038 552999 255040
rect 407113 255035 407179 255038
rect 552933 255035 552999 255038
rect 46565 254282 46631 254285
rect 48086 254282 48146 254456
rect 46565 254280 48146 254282
rect -960 254146 480 254236
rect 46565 254224 46570 254280
rect 46626 254224 48146 254280
rect 46565 254222 48146 254224
rect 46565 254219 46631 254222
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 347822 254010 347882 254456
rect 407389 254418 407455 254421
rect 553117 254418 553183 254421
rect 407389 254416 410044 254418
rect 407389 254360 407394 254416
rect 407450 254360 410044 254416
rect 407389 254358 410044 254360
rect 549884 254416 553183 254418
rect 549884 254360 553122 254416
rect 553178 254360 553183 254416
rect 549884 254358 553183 254360
rect 407389 254355 407455 254358
rect 553117 254355 553183 254358
rect 350441 254010 350507 254013
rect 347822 254008 350507 254010
rect 347822 253952 350446 254008
rect 350502 253952 350507 254008
rect 347822 253950 350507 253952
rect 350441 253947 350507 253950
rect 553117 253738 553183 253741
rect 549884 253736 553183 253738
rect 549884 253680 553122 253736
rect 553178 253680 553183 253736
rect 549884 253678 553183 253680
rect 553117 253675 553183 253678
rect 46054 252452 46060 252516
rect 46124 252514 46130 252516
rect 46381 252514 46447 252517
rect 46124 252512 46447 252514
rect 46124 252456 46386 252512
rect 46442 252456 46447 252512
rect 46124 252454 46447 252456
rect 46124 252452 46130 252454
rect 46381 252451 46447 252454
rect 553117 252378 553183 252381
rect 549884 252376 553183 252378
rect 549884 252320 553122 252376
rect 553178 252320 553183 252376
rect 549884 252318 553183 252320
rect 553117 252315 553183 252318
rect 46422 251772 46428 251836
rect 46492 251834 46498 251836
rect 376201 251834 376267 251837
rect 404854 251834 404860 251836
rect 46492 251774 48116 251834
rect 376201 251832 404860 251834
rect 376201 251776 376206 251832
rect 376262 251776 404860 251832
rect 376201 251774 404860 251776
rect 46492 251772 46498 251774
rect 376201 251771 376267 251774
rect 404854 251772 404860 251774
rect 404924 251772 404930 251836
rect 407205 251698 407271 251701
rect 407205 251696 410044 251698
rect 407205 251640 407210 251696
rect 407266 251640 410044 251696
rect 407205 251638 410044 251640
rect 407205 251635 407271 251638
rect 407205 251018 407271 251021
rect 407205 251016 410044 251018
rect 407205 250960 407210 251016
rect 407266 250960 410044 251016
rect 407205 250958 410044 250960
rect 407205 250955 407271 250958
rect 347822 249930 347882 250376
rect 407113 250338 407179 250341
rect 552933 250338 552999 250341
rect 407113 250336 410044 250338
rect 407113 250280 407118 250336
rect 407174 250280 410044 250336
rect 407113 250278 410044 250280
rect 549884 250336 552999 250338
rect 549884 250280 552938 250336
rect 552994 250280 552999 250336
rect 549884 250278 552999 250280
rect 407113 250275 407179 250278
rect 552933 250275 552999 250278
rect 350441 249930 350507 249933
rect 347822 249928 350507 249930
rect 347822 249872 350446 249928
rect 350502 249872 350507 249928
rect 347822 249870 350507 249872
rect 350441 249867 350507 249870
rect 408953 249658 409019 249661
rect 553117 249658 553183 249661
rect 408953 249656 410044 249658
rect 408953 249600 408958 249656
rect 409014 249600 410044 249656
rect 408953 249598 410044 249600
rect 549884 249656 553183 249658
rect 549884 249600 553122 249656
rect 553178 249600 553183 249656
rect 549884 249598 553183 249600
rect 408953 249595 409019 249598
rect 553117 249595 553183 249598
rect 347822 248570 347882 249016
rect 350441 248570 350507 248573
rect 347822 248568 350507 248570
rect 347822 248512 350446 248568
rect 350502 248512 350507 248568
rect 347822 248510 350507 248512
rect 350441 248507 350507 248510
rect 553117 248298 553183 248301
rect 549884 248296 553183 248298
rect 549884 248240 553122 248296
rect 553178 248240 553183 248296
rect 549884 248238 553183 248240
rect 553117 248235 553183 248238
rect 350073 247754 350139 247757
rect 347852 247752 350139 247754
rect 347852 247696 350078 247752
rect 350134 247696 350139 247752
rect 347852 247694 350139 247696
rect 350073 247691 350139 247694
rect 46422 247556 46428 247620
rect 46492 247618 46498 247620
rect 46749 247618 46815 247621
rect 46492 247616 46815 247618
rect 46492 247560 46754 247616
rect 46810 247560 46815 247616
rect 46492 247558 46815 247560
rect 46492 247556 46498 247558
rect 46749 247555 46815 247558
rect 46749 247482 46815 247485
rect 48086 247482 48146 247656
rect 553485 247618 553551 247621
rect 549884 247616 553551 247618
rect 549884 247560 553490 247616
rect 553546 247560 553551 247616
rect 549884 247558 553551 247560
rect 553485 247555 553551 247558
rect 46749 247480 48146 247482
rect 46749 247424 46754 247480
rect 46810 247424 48146 247480
rect 46749 247422 48146 247424
rect 46749 247419 46815 247422
rect 46606 247012 46612 247076
rect 46676 247074 46682 247076
rect 46676 247014 48116 247074
rect 46676 247012 46682 247014
rect 407205 246938 407271 246941
rect 563462 246938 563468 246940
rect 407205 246936 410044 246938
rect 407205 246880 407210 246936
rect 407266 246880 410044 246936
rect 407205 246878 410044 246880
rect 549884 246878 563468 246938
rect 407205 246875 407271 246878
rect 563462 246876 563468 246878
rect 563532 246876 563538 246940
rect 46749 245850 46815 245853
rect 48086 245850 48146 246296
rect 347822 246122 347882 246296
rect 407113 246258 407179 246261
rect 553117 246258 553183 246261
rect 407113 246256 410044 246258
rect 407113 246200 407118 246256
rect 407174 246200 410044 246256
rect 407113 246198 410044 246200
rect 549884 246256 553183 246258
rect 549884 246200 553122 246256
rect 553178 246200 553183 246256
rect 549884 246198 553183 246200
rect 407113 246195 407179 246198
rect 553117 246195 553183 246198
rect 350349 246122 350415 246125
rect 347822 246120 350415 246122
rect 347822 246064 350354 246120
rect 350410 246064 350415 246120
rect 347822 246062 350415 246064
rect 350349 246059 350415 246062
rect 46749 245848 48146 245850
rect 46749 245792 46754 245848
rect 46810 245792 48146 245848
rect 46749 245790 48146 245792
rect 350441 245850 350507 245853
rect 350441 245848 350642 245850
rect 350441 245792 350446 245848
rect 350502 245792 350642 245848
rect 350441 245790 350642 245792
rect 46749 245787 46815 245790
rect 350441 245787 350507 245790
rect 350441 245714 350507 245717
rect 347852 245712 350507 245714
rect 347852 245656 350446 245712
rect 350502 245656 350507 245712
rect 347852 245654 350507 245656
rect 350441 245651 350507 245654
rect 350582 245578 350642 245790
rect 350942 245578 350948 245580
rect 350582 245518 350948 245578
rect 350942 245516 350948 245518
rect 351012 245516 351018 245580
rect 407205 245578 407271 245581
rect 407205 245576 410044 245578
rect 407205 245520 407210 245576
rect 407266 245520 410044 245576
rect 407205 245518 410044 245520
rect 407205 245515 407271 245518
rect 44582 245380 44588 245444
rect 44652 245442 44658 245444
rect 46381 245442 46447 245445
rect 44652 245440 46447 245442
rect 44652 245384 46386 245440
rect 46442 245384 46447 245440
rect 583520 245428 584960 245668
rect 44652 245382 46447 245384
rect 44652 245380 44658 245382
rect 46381 245379 46447 245382
rect 347822 244490 347882 244936
rect 407113 244898 407179 244901
rect 553117 244898 553183 244901
rect 407113 244896 410044 244898
rect 407113 244840 407118 244896
rect 407174 244840 410044 244896
rect 407113 244838 410044 244840
rect 549884 244896 553183 244898
rect 549884 244840 553122 244896
rect 553178 244840 553183 244896
rect 549884 244838 553183 244840
rect 407113 244835 407179 244838
rect 553117 244835 553183 244838
rect 350533 244490 350599 244493
rect 347822 244488 350599 244490
rect 347822 244432 350538 244488
rect 350594 244432 350599 244488
rect 347822 244430 350599 244432
rect 350533 244427 350599 244430
rect 44766 244292 44772 244356
rect 44836 244354 44842 244356
rect 45093 244354 45159 244357
rect 46657 244356 46723 244357
rect 46606 244354 46612 244356
rect 44836 244352 45159 244354
rect 44836 244296 45098 244352
rect 45154 244296 45159 244352
rect 44836 244294 45159 244296
rect 46566 244294 46612 244354
rect 46676 244352 46723 244356
rect 46718 244296 46723 244352
rect 44836 244292 44842 244294
rect 45093 244291 45159 244294
rect 46606 244292 46612 244294
rect 46676 244292 46723 244296
rect 46790 244292 46796 244356
rect 46860 244354 46866 244356
rect 350073 244354 350139 244357
rect 46860 244294 48116 244354
rect 347852 244352 350139 244354
rect 347852 244296 350078 244352
rect 350134 244296 350139 244352
rect 347852 244294 350139 244296
rect 46860 244292 46866 244294
rect 46657 244291 46723 244292
rect 350073 244291 350139 244294
rect 347822 243266 347882 243576
rect 396206 243476 396212 243540
rect 396276 243538 396282 243540
rect 397361 243538 397427 243541
rect 396276 243536 397427 243538
rect 396276 243480 397366 243536
rect 397422 243480 397427 243536
rect 396276 243478 397427 243480
rect 396276 243476 396282 243478
rect 397361 243475 397427 243478
rect 350441 243266 350507 243269
rect 347822 243264 350507 243266
rect 347822 243208 350446 243264
rect 350502 243208 350507 243264
rect 347822 243206 350507 243208
rect 350441 243203 350507 243206
rect 45829 242994 45895 242997
rect 350165 242994 350231 242997
rect 45829 242992 48116 242994
rect 45829 242936 45834 242992
rect 45890 242936 48116 242992
rect 45829 242934 48116 242936
rect 347852 242992 350231 242994
rect 347852 242936 350170 242992
rect 350226 242936 350231 242992
rect 347852 242934 350231 242936
rect 45829 242931 45895 242934
rect 350165 242931 350231 242934
rect 407757 242994 407823 242997
rect 410014 242994 410074 243440
rect 549884 243410 550282 243470
rect 550222 243402 550282 243410
rect 552013 243402 552079 243405
rect 550222 243400 552079 243402
rect 550222 243344 552018 243400
rect 552074 243344 552079 243400
rect 550222 243342 552079 243344
rect 552013 243339 552079 243342
rect 407757 242992 410074 242994
rect 407757 242936 407762 242992
rect 407818 242936 410074 242992
rect 407757 242934 410074 242936
rect 407757 242931 407823 242934
rect 409822 242796 409828 242860
rect 409892 242858 409898 242860
rect 550173 242858 550239 242861
rect 409892 242798 410044 242858
rect 549884 242856 550239 242858
rect 549884 242800 550178 242856
rect 550234 242800 550239 242856
rect 549884 242798 550239 242800
rect 409892 242796 409898 242798
rect 550173 242795 550239 242798
rect 407665 242586 407731 242589
rect 410006 242586 410012 242588
rect 407665 242584 410012 242586
rect 407665 242528 407670 242584
rect 407726 242528 410012 242584
rect 407665 242526 410012 242528
rect 407665 242523 407731 242526
rect 410006 242524 410012 242526
rect 410076 242524 410082 242588
rect 407113 242178 407179 242181
rect 407113 242176 410044 242178
rect 407113 242120 407118 242176
rect 407174 242120 410044 242176
rect 407113 242118 410044 242120
rect 407113 242115 407179 242118
rect 47485 241498 47551 241501
rect 47710 241498 47716 241500
rect 47485 241496 47716 241498
rect 47485 241440 47490 241496
rect 47546 241440 47716 241496
rect 47485 241438 47716 241440
rect 47485 241435 47551 241438
rect 47710 241436 47716 241438
rect 47780 241436 47786 241500
rect 409505 241226 409571 241229
rect 410014 241226 410074 241468
rect 409505 241224 410074 241226
rect -960 241090 480 241180
rect 409505 241168 409510 241224
rect 409566 241168 410074 241224
rect 409505 241166 410074 241168
rect 409505 241163 409571 241166
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 47342 240892 47348 240956
rect 47412 240954 47418 240956
rect 47412 240894 48116 240954
rect 47412 240892 47418 240894
rect 409505 240818 409571 240821
rect 550081 240818 550147 240821
rect 409505 240816 410044 240818
rect 409505 240760 409510 240816
rect 409566 240760 410044 240816
rect 409505 240758 410044 240760
rect 549884 240816 550147 240818
rect 549884 240760 550086 240816
rect 550142 240760 550147 240816
rect 549884 240758 550147 240760
rect 409505 240755 409571 240758
rect 550081 240755 550147 240758
rect 391422 240484 391428 240548
rect 391492 240546 391498 240548
rect 576301 240546 576367 240549
rect 391492 240544 576367 240546
rect 391492 240488 576306 240544
rect 576362 240488 576367 240544
rect 391492 240486 576367 240488
rect 391492 240484 391498 240486
rect 576301 240483 576367 240486
rect 366541 240138 366607 240141
rect 568573 240138 568639 240141
rect 366541 240136 568639 240138
rect 366541 240080 366546 240136
rect 366602 240080 568578 240136
rect 568634 240080 568639 240136
rect 366541 240078 568639 240080
rect 366541 240075 366607 240078
rect 568573 240075 568639 240078
rect 396441 240002 396507 240005
rect 583293 240002 583359 240005
rect 396441 240000 583359 240002
rect 396441 239944 396446 240000
rect 396502 239944 583298 240000
rect 583354 239944 583359 240000
rect 396441 239942 583359 239944
rect 396441 239939 396507 239942
rect 583293 239939 583359 239942
rect 408401 239866 408467 239869
rect 554957 239866 555023 239869
rect 408401 239864 555023 239866
rect 408401 239808 408406 239864
rect 408462 239808 554962 239864
rect 555018 239808 555023 239864
rect 408401 239806 555023 239808
rect 408401 239803 408467 239806
rect 554957 239803 555023 239806
rect 538857 239594 538923 239597
rect 565905 239594 565971 239597
rect 538857 239592 565971 239594
rect 538857 239536 538862 239592
rect 538918 239536 565910 239592
rect 565966 239536 565971 239592
rect 538857 239534 565971 239536
rect 538857 239531 538923 239534
rect 565905 239531 565971 239534
rect 347822 239322 347882 239496
rect 393037 239458 393103 239461
rect 547229 239458 547295 239461
rect 393037 239456 547295 239458
rect 393037 239400 393042 239456
rect 393098 239400 547234 239456
rect 547290 239400 547295 239456
rect 393037 239398 547295 239400
rect 393037 239395 393103 239398
rect 547229 239395 547295 239398
rect 350349 239322 350415 239325
rect 347822 239320 350415 239322
rect 347822 239264 350354 239320
rect 350410 239264 350415 239320
rect 347822 239262 350415 239264
rect 350349 239259 350415 239262
rect 350441 238914 350507 238917
rect 347852 238912 350507 238914
rect 347852 238856 350446 238912
rect 350502 238856 350507 238912
rect 347852 238854 350507 238856
rect 350441 238851 350507 238854
rect 457345 238778 457411 238781
rect 551553 238778 551619 238781
rect 457345 238776 551619 238778
rect 457345 238720 457350 238776
rect 457406 238720 551558 238776
rect 551614 238720 551619 238776
rect 457345 238718 551619 238720
rect 457345 238715 457411 238718
rect 551553 238715 551619 238718
rect 399569 238642 399635 238645
rect 548149 238642 548215 238645
rect 399569 238640 548215 238642
rect 399569 238584 399574 238640
rect 399630 238584 548154 238640
rect 548210 238584 548215 238640
rect 399569 238582 548215 238584
rect 399569 238579 399635 238582
rect 548149 238579 548215 238582
rect 398281 238506 398347 238509
rect 528829 238506 528895 238509
rect 398281 238504 528895 238506
rect 398281 238448 398286 238504
rect 398342 238448 528834 238504
rect 528890 238448 528895 238504
rect 398281 238446 528895 238448
rect 398281 238443 398347 238446
rect 528829 238443 528895 238446
rect 388294 238308 388300 238372
rect 388364 238370 388370 238372
rect 458173 238370 458239 238373
rect 388364 238368 458239 238370
rect 388364 238312 458178 238368
rect 458234 238312 458239 238368
rect 388364 238310 458239 238312
rect 388364 238308 388370 238310
rect 458173 238307 458239 238310
rect 470593 238370 470659 238373
rect 556429 238370 556495 238373
rect 470593 238368 556495 238370
rect 470593 238312 470598 238368
rect 470654 238312 556434 238368
rect 556490 238312 556495 238368
rect 470593 238310 556495 238312
rect 470593 238307 470659 238310
rect 556429 238307 556495 238310
rect 46841 238234 46907 238237
rect 524321 238234 524387 238237
rect 548977 238234 549043 238237
rect 46841 238232 48116 238234
rect 46841 238176 46846 238232
rect 46902 238176 48116 238232
rect 46841 238174 48116 238176
rect 524321 238232 549043 238234
rect 524321 238176 524326 238232
rect 524382 238176 548982 238232
rect 549038 238176 549043 238232
rect 524321 238174 549043 238176
rect 46841 238171 46907 238174
rect 524321 238171 524387 238174
rect 548977 238171 549043 238174
rect 520181 238098 520247 238101
rect 549437 238098 549503 238101
rect 520181 238096 549503 238098
rect 520181 238040 520186 238096
rect 520242 238040 549442 238096
rect 549498 238040 549503 238096
rect 520181 238038 549503 238040
rect 520181 238035 520247 238038
rect 549437 238035 549503 238038
rect 528737 237962 528803 237965
rect 567653 237962 567719 237965
rect 528737 237960 567719 237962
rect 528737 237904 528742 237960
rect 528798 237904 567658 237960
rect 567714 237904 567719 237960
rect 528737 237902 567719 237904
rect 528737 237899 528803 237902
rect 567653 237899 567719 237902
rect 46841 237554 46907 237557
rect 46841 237552 48116 237554
rect 46841 237496 46846 237552
rect 46902 237496 48116 237552
rect 46841 237494 48116 237496
rect 46841 237491 46907 237494
rect 385953 237282 386019 237285
rect 577681 237282 577747 237285
rect 385953 237280 577747 237282
rect 385953 237224 385958 237280
rect 386014 237224 577686 237280
rect 577742 237224 577747 237280
rect 385953 237222 577747 237224
rect 385953 237219 386019 237222
rect 577681 237219 577747 237222
rect 393078 236676 393084 236740
rect 393148 236738 393154 236740
rect 547086 236738 547092 236740
rect 393148 236678 547092 236738
rect 393148 236676 393154 236678
rect 547086 236676 547092 236678
rect 547156 236676 547162 236740
rect 377213 236602 377279 236605
rect 543089 236602 543155 236605
rect 377213 236600 543155 236602
rect 377213 236544 377218 236600
rect 377274 236544 543094 236600
rect 543150 236544 543155 236600
rect 377213 236542 543155 236544
rect 377213 236539 377279 236542
rect 543089 236539 543155 236542
rect 350441 236194 350507 236197
rect 347852 236192 350507 236194
rect 347852 236136 350446 236192
rect 350502 236136 350507 236192
rect 347852 236134 350507 236136
rect 350441 236131 350507 236134
rect 46841 236058 46907 236061
rect 48086 236058 48146 236096
rect 46841 236056 48146 236058
rect 46841 236000 46846 236056
rect 46902 236000 48146 236056
rect 46841 235998 48146 236000
rect 46841 235995 46907 235998
rect 405590 235724 405596 235788
rect 405660 235786 405666 235788
rect 548006 235786 548012 235788
rect 405660 235726 548012 235786
rect 405660 235724 405666 235726
rect 548006 235724 548012 235726
rect 548076 235724 548082 235788
rect 400070 235588 400076 235652
rect 400140 235650 400146 235652
rect 544326 235650 544332 235652
rect 400140 235590 544332 235650
rect 400140 235588 400146 235590
rect 544326 235588 544332 235590
rect 544396 235588 544402 235652
rect 387558 235452 387564 235516
rect 387628 235514 387634 235516
rect 540278 235514 540284 235516
rect 387628 235454 540284 235514
rect 387628 235452 387634 235454
rect 540278 235452 540284 235454
rect 540348 235452 540354 235516
rect 347822 234970 347882 235416
rect 380433 235378 380499 235381
rect 541566 235378 541572 235380
rect 380433 235376 541572 235378
rect 380433 235320 380438 235376
rect 380494 235320 541572 235376
rect 380433 235318 541572 235320
rect 380433 235315 380499 235318
rect 541566 235316 541572 235318
rect 541636 235316 541642 235380
rect 552749 235378 552815 235381
rect 556838 235378 556844 235380
rect 552749 235376 556844 235378
rect 552749 235320 552754 235376
rect 552810 235320 556844 235376
rect 552749 235318 556844 235320
rect 552749 235315 552815 235318
rect 556838 235316 556844 235318
rect 556908 235316 556914 235380
rect 406142 235180 406148 235244
rect 406212 235242 406218 235244
rect 567653 235242 567719 235245
rect 406212 235240 567719 235242
rect 406212 235184 567658 235240
rect 567714 235184 567719 235240
rect 406212 235182 567719 235184
rect 406212 235180 406218 235182
rect 567653 235179 567719 235182
rect 350441 234970 350507 234973
rect 347822 234968 350507 234970
rect 347822 234912 350446 234968
rect 350502 234912 350507 234968
rect 347822 234910 350507 234912
rect 350441 234907 350507 234910
rect 45645 234698 45711 234701
rect 48086 234698 48146 234736
rect 45645 234696 48146 234698
rect 45645 234640 45650 234696
rect 45706 234640 48146 234696
rect 45645 234638 48146 234640
rect 556429 234698 556495 234701
rect 556654 234698 556660 234700
rect 556429 234696 556660 234698
rect 556429 234640 556434 234696
rect 556490 234640 556660 234696
rect 556429 234638 556660 234640
rect 45645 234635 45711 234638
rect 556429 234635 556495 234638
rect 556654 234636 556660 234638
rect 556724 234636 556730 234700
rect 412265 234290 412331 234293
rect 538806 234290 538812 234292
rect 412265 234288 538812 234290
rect 412265 234232 412270 234288
rect 412326 234232 538812 234288
rect 412265 234230 538812 234232
rect 412265 234227 412331 234230
rect 538806 234228 538812 234230
rect 538876 234228 538882 234292
rect 405406 234092 405412 234156
rect 405476 234154 405482 234156
rect 550725 234154 550791 234157
rect 405476 234152 550791 234154
rect 405476 234096 550730 234152
rect 550786 234096 550791 234152
rect 405476 234094 550791 234096
rect 405476 234092 405482 234094
rect 550725 234091 550791 234094
rect 404118 233956 404124 234020
rect 404188 234018 404194 234020
rect 549478 234018 549484 234020
rect 404188 233958 549484 234018
rect 404188 233956 404194 233958
rect 549478 233956 549484 233958
rect 549548 233956 549554 234020
rect 348918 233820 348924 233884
rect 348988 233882 348994 233884
rect 349153 233882 349219 233885
rect 348988 233880 349219 233882
rect 348988 233824 349158 233880
rect 349214 233824 349219 233880
rect 348988 233822 349219 233824
rect 348988 233820 348994 233822
rect 349153 233819 349219 233822
rect 388989 233882 389055 233885
rect 544101 233882 544167 233885
rect 388989 233880 544167 233882
rect 388989 233824 388994 233880
rect 389050 233824 544106 233880
rect 544162 233824 544167 233880
rect 388989 233822 544167 233824
rect 388989 233819 389055 233822
rect 544101 233819 544167 233822
rect 47025 233474 47091 233477
rect 47025 233472 48116 233474
rect 47025 233416 47030 233472
rect 47086 233416 48116 233472
rect 47025 233414 48116 233416
rect 47025 233411 47091 233414
rect 46841 232386 46907 232389
rect 48086 232386 48146 232696
rect 46841 232384 48146 232386
rect 46841 232328 46846 232384
rect 46902 232328 48146 232384
rect 46841 232326 48146 232328
rect 46841 232323 46907 232326
rect 347822 232250 347882 232696
rect 366633 232522 366699 232525
rect 538990 232522 538996 232524
rect 366633 232520 538996 232522
rect 366633 232464 366638 232520
rect 366694 232464 538996 232520
rect 366633 232462 538996 232464
rect 366633 232459 366699 232462
rect 538990 232460 538996 232462
rect 539060 232460 539066 232524
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 350441 232250 350507 232253
rect 347822 232248 350507 232250
rect 347822 232192 350446 232248
rect 350502 232192 350507 232248
rect 583520 232236 584960 232326
rect 347822 232190 350507 232192
rect 350441 232187 350507 232190
rect 400673 231706 400739 231709
rect 539174 231706 539180 231708
rect 400673 231704 539180 231706
rect 400673 231648 400678 231704
rect 400734 231648 539180 231704
rect 400673 231646 539180 231648
rect 400673 231643 400739 231646
rect 539174 231644 539180 231646
rect 539244 231644 539250 231708
rect 402094 231508 402100 231572
rect 402164 231570 402170 231572
rect 555509 231570 555575 231573
rect 402164 231568 555575 231570
rect 402164 231512 555514 231568
rect 555570 231512 555575 231568
rect 402164 231510 555575 231512
rect 402164 231508 402170 231510
rect 555509 231507 555575 231510
rect 383561 231434 383627 231437
rect 543549 231434 543615 231437
rect 383561 231432 543615 231434
rect 383561 231376 383566 231432
rect 383622 231376 543554 231432
rect 543610 231376 543615 231432
rect 383561 231374 543615 231376
rect 383561 231371 383627 231374
rect 543549 231371 543615 231374
rect 47025 230890 47091 230893
rect 48086 230890 48146 231336
rect 397310 231236 397316 231300
rect 397380 231298 397386 231300
rect 560293 231298 560359 231301
rect 397380 231296 560359 231298
rect 397380 231240 560298 231296
rect 560354 231240 560359 231296
rect 397380 231238 560359 231240
rect 397380 231236 397386 231238
rect 560293 231235 560359 231238
rect 401358 231100 401364 231164
rect 401428 231162 401434 231164
rect 565169 231162 565235 231165
rect 401428 231160 565235 231162
rect 401428 231104 565174 231160
rect 565230 231104 565235 231160
rect 401428 231102 565235 231104
rect 401428 231100 401434 231102
rect 565169 231099 565235 231102
rect 47025 230888 48146 230890
rect 47025 230832 47030 230888
rect 47086 230832 48146 230888
rect 47025 230830 48146 230832
rect 47025 230827 47091 230830
rect 46841 230618 46907 230621
rect 48086 230618 48146 230656
rect 46841 230616 48146 230618
rect 46841 230560 46846 230616
rect 46902 230560 48146 230616
rect 46841 230558 48146 230560
rect 347822 230618 347882 230656
rect 350441 230618 350507 230621
rect 347822 230616 350507 230618
rect 347822 230560 350446 230616
rect 350502 230560 350507 230616
rect 347822 230558 350507 230560
rect 46841 230555 46907 230558
rect 350441 230555 350507 230558
rect 47761 229394 47827 229397
rect 47761 229392 48116 229394
rect 47761 229336 47766 229392
rect 47822 229336 48116 229392
rect 47761 229334 48116 229336
rect 47761 229331 47827 229334
rect 347822 229258 347882 229296
rect 350441 229258 350507 229261
rect 347822 229256 350507 229258
rect 347822 229200 350446 229256
rect 350502 229200 350507 229256
rect 347822 229198 350507 229200
rect 350441 229195 350507 229198
rect -960 227884 480 228124
rect 46841 227898 46907 227901
rect 48086 227898 48146 227936
rect 46841 227896 48146 227898
rect 46841 227840 46846 227896
rect 46902 227840 48146 227896
rect 46841 227838 48146 227840
rect 46841 227835 46907 227838
rect 46565 226674 46631 226677
rect 46565 226672 48116 226674
rect 46565 226616 46570 226672
rect 46626 226616 48116 226672
rect 46565 226614 48116 226616
rect 46565 226611 46631 226614
rect 47761 226404 47827 226405
rect 47710 226402 47716 226404
rect 47670 226342 47716 226402
rect 47780 226400 47827 226404
rect 47822 226344 47827 226400
rect 47710 226340 47716 226342
rect 47780 226340 47827 226344
rect 47761 226339 47827 226340
rect 347822 225042 347882 225216
rect 350441 225042 350507 225045
rect 347822 225040 350507 225042
rect 347822 224984 350446 225040
rect 350502 224984 350507 225040
rect 347822 224982 350507 224984
rect 350441 224979 350507 224982
rect 46841 224090 46907 224093
rect 48086 224090 48146 224536
rect 46841 224088 48146 224090
rect 46841 224032 46846 224088
rect 46902 224032 48146 224088
rect 46841 224030 48146 224032
rect 46841 224027 46907 224030
rect 350441 222594 350507 222597
rect 347852 222592 350507 222594
rect 347852 222536 350446 222592
rect 350502 222536 350507 222592
rect 347852 222534 350507 222536
rect 350441 222531 350507 222534
rect 46841 222458 46907 222461
rect 48086 222458 48146 222496
rect 46841 222456 48146 222458
rect 46841 222400 46846 222456
rect 46902 222400 48146 222456
rect 46841 222398 48146 222400
rect 46841 222395 46907 222398
rect 46381 222186 46447 222189
rect 47710 222186 47716 222188
rect 46381 222184 47716 222186
rect 46381 222128 46386 222184
rect 46442 222128 47716 222184
rect 46381 222126 47716 222128
rect 46381 222123 46447 222126
rect 47710 222124 47716 222126
rect 47780 222124 47786 222188
rect 46657 221370 46723 221373
rect 48086 221370 48146 221816
rect 46657 221368 48146 221370
rect 46657 221312 46662 221368
rect 46718 221312 48146 221368
rect 46657 221310 48146 221312
rect 46657 221307 46723 221310
rect 347822 221234 347882 221816
rect 350441 221234 350507 221237
rect 347822 221232 350507 221234
rect 347822 221176 350446 221232
rect 350502 221176 350507 221232
rect 347822 221174 350507 221176
rect 350441 221171 350507 221174
rect 46841 221098 46907 221101
rect 48086 221098 48146 221136
rect 46841 221096 48146 221098
rect 46841 221040 46846 221096
rect 46902 221040 48146 221096
rect 46841 221038 48146 221040
rect 46841 221035 46907 221038
rect 37733 220826 37799 220829
rect 39246 220826 39252 220828
rect 37733 220824 39252 220826
rect 37733 220768 37738 220824
rect 37794 220768 39252 220824
rect 37733 220766 39252 220768
rect 37733 220763 37799 220766
rect 39246 220764 39252 220766
rect 39316 220764 39322 220828
rect 44173 220826 44239 220829
rect 44766 220826 44772 220828
rect 44173 220824 44772 220826
rect 44173 220768 44178 220824
rect 44234 220768 44772 220824
rect 44173 220766 44772 220768
rect 44173 220763 44239 220766
rect 44766 220764 44772 220766
rect 44836 220764 44842 220828
rect 47158 220492 47164 220556
rect 47228 220554 47234 220556
rect 47228 220494 48116 220554
rect 47228 220492 47234 220494
rect 47761 220282 47827 220285
rect 48078 220282 48084 220284
rect 47761 220280 48084 220282
rect 47761 220224 47766 220280
rect 47822 220224 48084 220280
rect 47761 220222 48084 220224
rect 47761 220219 47827 220222
rect 48078 220220 48084 220222
rect 48148 220220 48154 220284
rect 35801 220146 35867 220149
rect 44582 220146 44588 220148
rect 35801 220144 44588 220146
rect 35801 220088 35806 220144
rect 35862 220088 44588 220144
rect 35801 220086 44588 220088
rect 35801 220083 35867 220086
rect 44582 220084 44588 220086
rect 44652 220084 44658 220148
rect 347822 220010 347882 220456
rect 350349 220010 350415 220013
rect 347822 220008 350415 220010
rect 347822 219952 350354 220008
rect 350410 219952 350415 220008
rect 347822 219950 350415 219952
rect 350349 219947 350415 219950
rect 46565 218650 46631 218653
rect 48086 218650 48146 219096
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 46565 218648 48146 218650
rect 46565 218592 46570 218648
rect 46626 218592 48146 218648
rect 46565 218590 48146 218592
rect 46565 218587 46631 218590
rect 38101 218106 38167 218109
rect 39246 218106 39252 218108
rect 38101 218104 39252 218106
rect 38101 218048 38106 218104
rect 38162 218048 39252 218104
rect 38101 218046 39252 218048
rect 38101 218043 38167 218046
rect 39246 218044 39252 218046
rect 39316 218044 39322 218108
rect 46841 218106 46907 218109
rect 48086 218106 48146 218416
rect 46841 218104 48146 218106
rect 46841 218048 46846 218104
rect 46902 218048 48146 218104
rect 46841 218046 48146 218048
rect 347822 218106 347882 218416
rect 350441 218106 350507 218109
rect 347822 218104 350507 218106
rect 347822 218048 350446 218104
rect 350502 218048 350507 218104
rect 347822 218046 350507 218048
rect 46841 218043 46907 218046
rect 350441 218043 350507 218046
rect 46013 217290 46079 217293
rect 48086 217290 48146 217736
rect 347822 217562 347882 217736
rect 350441 217562 350507 217565
rect 347822 217560 350507 217562
rect 347822 217504 350446 217560
rect 350502 217504 350507 217560
rect 347822 217502 350507 217504
rect 350441 217499 350507 217502
rect 46013 217288 48146 217290
rect 46013 217232 46018 217288
rect 46074 217232 48146 217288
rect 46013 217230 48146 217232
rect 46013 217227 46079 217230
rect 350257 217154 350323 217157
rect 347852 217152 350323 217154
rect 347852 217096 350262 217152
rect 350318 217096 350323 217152
rect 347852 217094 350323 217096
rect 350257 217091 350323 217094
rect 47485 216746 47551 216749
rect 48086 216746 48146 217056
rect 47485 216744 48146 216746
rect 47485 216688 47490 216744
rect 47546 216688 48146 216744
rect 47485 216686 48146 216688
rect 47485 216683 47551 216686
rect 46841 215386 46907 215389
rect 48086 215386 48146 215696
rect 46841 215384 48146 215386
rect 46841 215328 46846 215384
rect 46902 215328 48146 215384
rect 46841 215326 48146 215328
rect 347822 215386 347882 215696
rect 350441 215386 350507 215389
rect 347822 215384 350507 215386
rect 347822 215328 350446 215384
rect 350502 215328 350507 215384
rect 347822 215326 350507 215328
rect 46841 215323 46907 215326
rect 350441 215323 350507 215326
rect -960 214828 480 215068
rect 46841 214026 46907 214029
rect 48086 214026 48146 214336
rect 46841 214024 48146 214026
rect 46841 213968 46846 214024
rect 46902 213968 48146 214024
rect 46841 213966 48146 213968
rect 46841 213963 46907 213966
rect 347822 213210 347882 213656
rect 350441 213210 350507 213213
rect 347822 213208 350507 213210
rect 347822 213152 350446 213208
rect 350502 213152 350507 213208
rect 347822 213150 350507 213152
rect 350441 213147 350507 213150
rect 46841 211306 46907 211309
rect 48086 211306 48146 211616
rect 46841 211304 48146 211306
rect 46841 211248 46846 211304
rect 46902 211248 48146 211304
rect 46841 211246 48146 211248
rect 46841 211243 46907 211246
rect 46974 210292 46980 210356
rect 47044 210354 47050 210356
rect 372153 210354 372219 210357
rect 542670 210354 542676 210356
rect 47044 210294 48116 210354
rect 372153 210352 542676 210354
rect 372153 210296 372158 210352
rect 372214 210296 542676 210352
rect 372153 210294 542676 210296
rect 47044 210292 47050 210294
rect 372153 210291 372219 210294
rect 542670 210292 542676 210294
rect 542740 210292 542746 210356
rect 347822 210082 347882 210256
rect 349521 210082 349587 210085
rect 347822 210080 349587 210082
rect 347822 210024 349526 210080
rect 349582 210024 349587 210080
rect 347822 210022 349587 210024
rect 349521 210019 349587 210022
rect 347822 209130 347882 209576
rect 350441 209130 350507 209133
rect 347822 209128 350507 209130
rect 347822 209072 350446 209128
rect 350502 209072 350507 209128
rect 347822 209070 350507 209072
rect 350441 209067 350507 209070
rect 347822 207770 347882 208216
rect 350257 207770 350323 207773
rect 347822 207768 350323 207770
rect 347822 207712 350262 207768
rect 350318 207712 350323 207768
rect 347822 207710 350323 207712
rect 350257 207707 350323 207710
rect 46841 207634 46907 207637
rect 46841 207632 48116 207634
rect 46841 207576 46846 207632
rect 46902 207576 48116 207632
rect 46841 207574 48116 207576
rect 46841 207571 46907 207574
rect 347822 207226 347882 207536
rect 350441 207226 350507 207229
rect 347822 207224 350507 207226
rect 347822 207168 350446 207224
rect 350502 207168 350507 207224
rect 347822 207166 350507 207168
rect 350441 207163 350507 207166
rect 46841 206954 46907 206957
rect 350441 206954 350507 206957
rect 46841 206952 48116 206954
rect 46841 206896 46846 206952
rect 46902 206896 48116 206952
rect 46841 206894 48116 206896
rect 347852 206952 350507 206954
rect 347852 206896 350446 206952
rect 350502 206896 350507 206952
rect 347852 206894 350507 206896
rect 46841 206891 46907 206894
rect 350441 206891 350507 206894
rect 406510 206212 406516 206276
rect 406580 206274 406586 206276
rect 523033 206274 523099 206277
rect 406580 206272 523099 206274
rect 406580 206216 523038 206272
rect 523094 206216 523099 206272
rect 406580 206214 523099 206216
rect 406580 206212 406586 206214
rect 523033 206211 523099 206214
rect 37733 205730 37799 205733
rect 39062 205730 39068 205732
rect 37733 205728 39068 205730
rect 37733 205672 37738 205728
rect 37794 205672 39068 205728
rect 37733 205670 39068 205672
rect 37733 205667 37799 205670
rect 39062 205668 39068 205670
rect 39132 205668 39138 205732
rect 39246 205668 39252 205732
rect 39316 205730 39322 205732
rect 42977 205730 43043 205733
rect 39316 205728 43043 205730
rect 39316 205672 42982 205728
rect 43038 205672 43043 205728
rect 39316 205670 43043 205672
rect 39316 205668 39322 205670
rect 42977 205667 43043 205670
rect 46841 205730 46907 205733
rect 48086 205730 48146 206176
rect 46841 205728 48146 205730
rect 46841 205672 46846 205728
rect 46902 205672 48146 205728
rect 46841 205670 48146 205672
rect 46841 205667 46907 205670
rect 583520 205580 584960 205820
rect 347822 205050 347882 205496
rect 350257 205050 350323 205053
rect 347822 205048 350323 205050
rect 347822 204992 350262 205048
rect 350318 204992 350323 205048
rect 347822 204990 350323 204992
rect 350257 204987 350323 204990
rect 39614 204852 39620 204916
rect 39684 204914 39690 204916
rect 40677 204914 40743 204917
rect 39684 204912 40743 204914
rect 39684 204856 40682 204912
rect 40738 204856 40743 204912
rect 39684 204854 40743 204856
rect 39684 204852 39690 204854
rect 40677 204851 40743 204854
rect 47526 204444 47532 204508
rect 47596 204506 47602 204508
rect 47894 204506 47900 204508
rect 47596 204446 47900 204506
rect 47596 204444 47602 204446
rect 47894 204444 47900 204446
rect 47964 204444 47970 204508
rect 46197 204370 46263 204373
rect 47526 204370 47532 204372
rect 46197 204368 47532 204370
rect 46197 204312 46202 204368
rect 46258 204312 47532 204368
rect 46197 204310 47532 204312
rect 46197 204307 46263 204310
rect 47526 204308 47532 204310
rect 47596 204308 47602 204372
rect 350441 204234 350507 204237
rect 347852 204232 350507 204234
rect 347852 204176 350446 204232
rect 350502 204176 350507 204232
rect 347852 204174 350507 204176
rect 350441 204171 350507 204174
rect 45645 203690 45711 203693
rect 48086 203690 48146 204136
rect 45645 203688 48146 203690
rect 45645 203632 45650 203688
rect 45706 203632 48146 203688
rect 45645 203630 48146 203632
rect 45645 203627 45711 203630
rect 33961 203554 34027 203557
rect 39246 203554 39252 203556
rect 33961 203552 39252 203554
rect 33961 203496 33966 203552
rect 34022 203496 39252 203552
rect 33961 203494 39252 203496
rect 33961 203491 34027 203494
rect 39246 203492 39252 203494
rect 39316 203492 39322 203556
rect 347822 203146 347882 203456
rect 350441 203146 350507 203149
rect 347822 203144 350507 203146
rect 347822 203088 350446 203144
rect 350502 203088 350507 203144
rect 347822 203086 350507 203088
rect 350441 203083 350507 203086
rect 45553 202874 45619 202877
rect 45553 202872 48116 202874
rect 45553 202816 45558 202872
rect 45614 202816 48116 202872
rect 45553 202814 48116 202816
rect 45553 202811 45619 202814
rect 347822 202330 347882 202776
rect 349337 202330 349403 202333
rect 347822 202328 349403 202330
rect 347822 202272 349342 202328
rect 349398 202272 349403 202328
rect 347822 202270 349403 202272
rect 349337 202267 349403 202270
rect -960 201922 480 202012
rect 4061 201922 4127 201925
rect -960 201920 4127 201922
rect -960 201864 4066 201920
rect 4122 201864 4127 201920
rect -960 201862 4127 201864
rect -960 201772 480 201862
rect 4061 201859 4127 201862
rect 44582 201588 44588 201652
rect 44652 201650 44658 201652
rect 46197 201650 46263 201653
rect 48270 201652 48330 202096
rect 347822 201786 347882 202096
rect 350441 201786 350507 201789
rect 347822 201784 350507 201786
rect 347822 201728 350446 201784
rect 350502 201728 350507 201784
rect 347822 201726 350507 201728
rect 350441 201723 350507 201726
rect 44652 201648 46263 201650
rect 44652 201592 46202 201648
rect 46258 201592 46263 201648
rect 44652 201590 46263 201592
rect 44652 201588 44658 201590
rect 46197 201587 46263 201590
rect 48262 201588 48268 201652
rect 48332 201588 48338 201652
rect 44766 201452 44772 201516
rect 44836 201514 44842 201516
rect 45737 201514 45803 201517
rect 44836 201512 45803 201514
rect 44836 201456 45742 201512
rect 45798 201456 45803 201512
rect 44836 201454 45803 201456
rect 44836 201452 44842 201454
rect 45737 201451 45803 201454
rect 347814 201044 347820 201108
rect 347884 201106 347890 201108
rect 353293 201106 353359 201109
rect 347884 201104 353359 201106
rect 347884 201048 353298 201104
rect 353354 201048 353359 201104
rect 347884 201046 353359 201048
rect 347884 201044 347890 201046
rect 353293 201043 353359 201046
rect 347681 200970 347747 200973
rect 581821 200970 581887 200973
rect 347681 200968 581887 200970
rect 347681 200912 347686 200968
rect 347742 200912 581826 200968
rect 581882 200912 581887 200968
rect 347681 200910 581887 200912
rect 347681 200907 347747 200910
rect 581821 200907 581887 200910
rect 45093 200562 45159 200565
rect 48262 200562 48268 200564
rect 45093 200560 48268 200562
rect 45093 200504 45098 200560
rect 45154 200504 48268 200560
rect 45093 200502 48268 200504
rect 45093 200499 45159 200502
rect 48262 200500 48268 200502
rect 48332 200500 48338 200564
rect 347630 200500 347636 200564
rect 347700 200562 347706 200564
rect 349705 200562 349771 200565
rect 347700 200560 349771 200562
rect 347700 200504 349710 200560
rect 349766 200504 349771 200560
rect 347700 200502 349771 200504
rect 347700 200500 347706 200502
rect 349705 200499 349771 200502
rect 347681 200290 347747 200293
rect 348693 200290 348759 200293
rect 347681 200288 348759 200290
rect 347681 200232 347686 200288
rect 347742 200232 348698 200288
rect 348754 200232 348759 200288
rect 347681 200230 348759 200232
rect 347681 200227 347747 200230
rect 348693 200227 348759 200230
rect 41873 200020 41939 200021
rect 41822 200018 41828 200020
rect 41782 199958 41828 200018
rect 41892 200016 41939 200020
rect 41934 199960 41939 200016
rect 41822 199956 41828 199958
rect 41892 199956 41939 199960
rect 41873 199955 41939 199956
rect 39205 199882 39271 199885
rect 562409 199882 562475 199885
rect 39205 199880 562475 199882
rect 39205 199824 39210 199880
rect 39266 199824 562414 199880
rect 562470 199824 562475 199880
rect 39205 199822 562475 199824
rect 39205 199819 39271 199822
rect 562409 199819 562475 199822
rect 37181 199746 37247 199749
rect 362401 199746 362467 199749
rect 37181 199744 362467 199746
rect 37181 199688 37186 199744
rect 37242 199688 362406 199744
rect 362462 199688 362467 199744
rect 37181 199686 362467 199688
rect 37181 199683 37247 199686
rect 362401 199683 362467 199686
rect 47853 199610 47919 199613
rect 48998 199610 49004 199612
rect 47853 199608 49004 199610
rect 47853 199552 47858 199608
rect 47914 199552 49004 199608
rect 47853 199550 49004 199552
rect 47853 199547 47919 199550
rect 48998 199548 49004 199550
rect 49068 199548 49074 199612
rect 347446 199548 347452 199612
rect 347516 199610 347522 199612
rect 347589 199610 347655 199613
rect 347516 199608 347655 199610
rect 347516 199552 347594 199608
rect 347650 199552 347655 199608
rect 347516 199550 347655 199552
rect 347516 199548 347522 199550
rect 347589 199547 347655 199550
rect 346117 199338 346183 199341
rect 382917 199338 382983 199341
rect 346117 199336 382983 199338
rect 346117 199280 346122 199336
rect 346178 199280 382922 199336
rect 382978 199280 382983 199336
rect 346117 199278 382983 199280
rect 346117 199275 346183 199278
rect 382917 199275 382983 199278
rect 35709 199066 35775 199069
rect 174905 199066 174971 199069
rect 35709 199064 174971 199066
rect 35709 199008 35714 199064
rect 35770 199008 174910 199064
rect 174966 199008 174971 199064
rect 35709 199006 174971 199008
rect 35709 199003 35775 199006
rect 174905 199003 174971 199006
rect 200021 199066 200087 199069
rect 363689 199066 363755 199069
rect 200021 199064 363755 199066
rect 200021 199008 200026 199064
rect 200082 199008 363694 199064
rect 363750 199008 363755 199064
rect 200021 199006 363755 199008
rect 200021 199003 200087 199006
rect 363689 199003 363755 199006
rect 38285 198930 38351 198933
rect 257889 198930 257955 198933
rect 38285 198928 257955 198930
rect 38285 198872 38290 198928
rect 38346 198872 257894 198928
rect 257950 198872 257955 198928
rect 38285 198870 257955 198872
rect 38285 198867 38351 198870
rect 257889 198867 257955 198870
rect 348693 198930 348759 198933
rect 350942 198930 350948 198932
rect 348693 198928 350948 198930
rect 348693 198872 348698 198928
rect 348754 198872 350948 198928
rect 348693 198870 350948 198872
rect 348693 198867 348759 198870
rect 350942 198868 350948 198870
rect 351012 198868 351018 198932
rect 83457 198794 83523 198797
rect 560753 198794 560819 198797
rect 83457 198792 560819 198794
rect 83457 198736 83462 198792
rect 83518 198736 560758 198792
rect 560814 198736 560819 198792
rect 83457 198734 560819 198736
rect 83457 198731 83523 198734
rect 560753 198731 560819 198734
rect 19977 198658 20043 198661
rect 396533 198658 396599 198661
rect 19977 198656 396599 198658
rect 19977 198600 19982 198656
rect 20038 198600 396538 198656
rect 396594 198600 396599 198656
rect 19977 198598 396599 198600
rect 19977 198595 20043 198598
rect 396533 198595 396599 198598
rect 21265 198522 21331 198525
rect 347681 198522 347747 198525
rect 21265 198520 347747 198522
rect 21265 198464 21270 198520
rect 21326 198464 347686 198520
rect 347742 198464 347747 198520
rect 21265 198462 347747 198464
rect 21265 198459 21331 198462
rect 347681 198459 347747 198462
rect 35617 198386 35683 198389
rect 82813 198386 82879 198389
rect 35617 198384 82879 198386
rect 35617 198328 35622 198384
rect 35678 198328 82818 198384
rect 82874 198328 82879 198384
rect 35617 198326 82879 198328
rect 35617 198323 35683 198326
rect 82813 198323 82879 198326
rect 94405 198386 94471 198389
rect 368974 198386 368980 198388
rect 94405 198384 368980 198386
rect 94405 198328 94410 198384
rect 94466 198328 368980 198384
rect 94405 198326 368980 198328
rect 94405 198323 94471 198326
rect 368974 198324 368980 198326
rect 369044 198324 369050 198388
rect 25865 198250 25931 198253
rect 53833 198250 53899 198253
rect 25865 198248 53899 198250
rect 25865 198192 25870 198248
rect 25926 198192 53838 198248
rect 53894 198192 53899 198248
rect 25865 198190 53899 198192
rect 25865 198187 25931 198190
rect 53833 198187 53899 198190
rect 122741 198250 122807 198253
rect 356830 198250 356836 198252
rect 122741 198248 356836 198250
rect 122741 198192 122746 198248
rect 122802 198192 356836 198248
rect 122741 198190 356836 198192
rect 122741 198187 122807 198190
rect 356830 198188 356836 198190
rect 356900 198188 356906 198252
rect 36537 198114 36603 198117
rect 153653 198114 153719 198117
rect 36537 198112 153719 198114
rect 36537 198056 36542 198112
rect 36598 198056 153658 198112
rect 153714 198056 153719 198112
rect 36537 198054 153719 198056
rect 36537 198051 36603 198054
rect 153653 198051 153719 198054
rect 170397 198114 170463 198117
rect 359406 198114 359412 198116
rect 170397 198112 359412 198114
rect 170397 198056 170402 198112
rect 170458 198056 359412 198112
rect 170397 198054 359412 198056
rect 170397 198051 170463 198054
rect 359406 198052 359412 198054
rect 359476 198052 359482 198116
rect 47526 197916 47532 197980
rect 47596 197978 47602 197980
rect 93117 197978 93183 197981
rect 47596 197976 93183 197978
rect 47596 197920 93122 197976
rect 93178 197920 93183 197976
rect 47596 197918 93183 197920
rect 47596 197916 47602 197918
rect 93117 197915 93183 197918
rect 208117 197978 208183 197981
rect 557809 197978 557875 197981
rect 208117 197976 557875 197978
rect 208117 197920 208122 197976
rect 208178 197920 557814 197976
rect 557870 197920 557875 197976
rect 208117 197918 557875 197920
rect 208117 197915 208183 197918
rect 557809 197915 557875 197918
rect 3417 197298 3483 197301
rect 542353 197298 542419 197301
rect 3417 197296 542419 197298
rect 3417 197240 3422 197296
rect 3478 197240 542358 197296
rect 542414 197240 542419 197296
rect 3417 197238 542419 197240
rect 3417 197235 3483 197238
rect 542353 197235 542419 197238
rect 58985 197162 59051 197165
rect 560477 197162 560543 197165
rect 58985 197160 560543 197162
rect 58985 197104 58990 197160
rect 59046 197104 560482 197160
rect 560538 197104 560543 197160
rect 58985 197102 560543 197104
rect 58985 197099 59051 197102
rect 560477 197099 560543 197102
rect 120165 197026 120231 197029
rect 560661 197026 560727 197029
rect 120165 197024 560727 197026
rect 120165 196968 120170 197024
rect 120226 196968 560666 197024
rect 560722 196968 560727 197024
rect 120165 196966 560727 196968
rect 120165 196963 120231 196966
rect 560661 196963 560727 196966
rect 34329 196890 34395 196893
rect 342345 196890 342411 196893
rect 34329 196888 342411 196890
rect 34329 196832 34334 196888
rect 34390 196832 342350 196888
rect 342406 196832 342411 196888
rect 34329 196830 342411 196832
rect 34329 196827 34395 196830
rect 342345 196827 342411 196830
rect 187785 196754 187851 196757
rect 367686 196754 367692 196756
rect 187785 196752 367692 196754
rect 187785 196696 187790 196752
rect 187846 196696 367692 196752
rect 187785 196694 367692 196696
rect 187785 196691 187851 196694
rect 367686 196692 367692 196694
rect 367756 196692 367762 196756
rect 47894 196556 47900 196620
rect 47964 196618 47970 196620
rect 235165 196618 235231 196621
rect 47964 196616 235231 196618
rect 47964 196560 235170 196616
rect 235226 196560 235231 196616
rect 47964 196558 235231 196560
rect 47964 196556 47970 196558
rect 235165 196555 235231 196558
rect 270585 196618 270651 196621
rect 555049 196618 555115 196621
rect 270585 196616 555115 196618
rect 270585 196560 270590 196616
rect 270646 196560 555054 196616
rect 555110 196560 555115 196616
rect 270585 196558 555115 196560
rect 270585 196555 270651 196558
rect 555049 196555 555115 196558
rect 36670 195876 36676 195940
rect 36740 195938 36746 195940
rect 531313 195938 531379 195941
rect 36740 195936 531379 195938
rect 36740 195880 531318 195936
rect 531374 195880 531379 195936
rect 36740 195878 531379 195880
rect 36740 195876 36746 195878
rect 531313 195875 531379 195878
rect 60273 195802 60339 195805
rect 403750 195802 403756 195804
rect 60273 195800 403756 195802
rect 60273 195744 60278 195800
rect 60334 195744 403756 195800
rect 60273 195742 403756 195744
rect 60273 195739 60339 195742
rect 403750 195740 403756 195742
rect 403820 195740 403826 195804
rect 56133 195530 56199 195533
rect 349102 195530 349108 195532
rect 56133 195528 349108 195530
rect 56133 195472 56138 195528
rect 56194 195472 349108 195528
rect 56133 195470 349108 195472
rect 56133 195467 56199 195470
rect 349102 195468 349108 195470
rect 349172 195468 349178 195532
rect 45921 195394 45987 195397
rect 495433 195394 495499 195397
rect 45921 195392 495499 195394
rect 45921 195336 45926 195392
rect 45982 195336 495438 195392
rect 495494 195336 495499 195392
rect 45921 195334 495499 195336
rect 45921 195331 45987 195334
rect 495433 195331 495499 195334
rect 46238 195196 46244 195260
rect 46308 195258 46314 195260
rect 536097 195258 536163 195261
rect 46308 195256 536163 195258
rect 46308 195200 536102 195256
rect 536158 195200 536163 195256
rect 46308 195198 536163 195200
rect 46308 195196 46314 195198
rect 536097 195195 536163 195198
rect 30966 194516 30972 194580
rect 31036 194578 31042 194580
rect 476205 194578 476271 194581
rect 31036 194576 476271 194578
rect 31036 194520 476210 194576
rect 476266 194520 476271 194576
rect 31036 194518 476271 194520
rect 31036 194516 31042 194518
rect 476205 194515 476271 194518
rect 4061 194442 4127 194445
rect 395654 194442 395660 194444
rect 4061 194440 395660 194442
rect 4061 194384 4066 194440
rect 4122 194384 395660 194440
rect 4061 194382 395660 194384
rect 4061 194379 4127 194382
rect 395654 194380 395660 194382
rect 395724 194380 395730 194444
rect 27245 194306 27311 194309
rect 330753 194306 330819 194309
rect 27245 194304 330819 194306
rect 27245 194248 27250 194304
rect 27306 194248 330758 194304
rect 330814 194248 330819 194304
rect 27245 194246 330819 194248
rect 27245 194243 27311 194246
rect 330753 194243 330819 194246
rect 133045 194170 133111 194173
rect 368473 194170 368539 194173
rect 133045 194168 368539 194170
rect 133045 194112 133050 194168
rect 133106 194112 368478 194168
rect 368534 194112 368539 194168
rect 133045 194110 368539 194112
rect 133045 194107 133111 194110
rect 368473 194107 368539 194110
rect 48262 193972 48268 194036
rect 48332 194034 48338 194036
rect 196801 194034 196867 194037
rect 48332 194032 196867 194034
rect 48332 193976 196806 194032
rect 196862 193976 196867 194032
rect 48332 193974 196867 193976
rect 48332 193972 48338 193974
rect 196801 193971 196867 193974
rect 53046 193836 53052 193900
rect 53116 193898 53122 193900
rect 564985 193898 565051 193901
rect 53116 193896 565051 193898
rect 53116 193840 564990 193896
rect 565046 193840 565051 193896
rect 53116 193838 565051 193840
rect 53116 193836 53122 193838
rect 564985 193835 565051 193838
rect 48998 192884 49004 192948
rect 49068 192946 49074 192948
rect 139393 192946 139459 192949
rect 49068 192944 139459 192946
rect 49068 192888 139398 192944
rect 139454 192888 139459 192944
rect 49068 192886 139459 192888
rect 49068 192884 49074 192886
rect 139393 192883 139459 192886
rect 146293 192946 146359 192949
rect 356094 192946 356100 192948
rect 146293 192944 356100 192946
rect 146293 192888 146298 192944
rect 146354 192888 356100 192944
rect 146293 192886 356100 192888
rect 146293 192883 146359 192886
rect 356094 192884 356100 192886
rect 356164 192884 356170 192948
rect 27613 192810 27679 192813
rect 374494 192810 374500 192812
rect 27613 192808 374500 192810
rect 27613 192752 27618 192808
rect 27674 192752 374500 192808
rect 27613 192750 374500 192752
rect 27613 192747 27679 192750
rect 374494 192748 374500 192750
rect 374564 192748 374570 192812
rect 45134 192612 45140 192676
rect 45204 192674 45210 192676
rect 453481 192674 453547 192677
rect 45204 192672 453547 192674
rect 45204 192616 453486 192672
rect 453542 192616 453547 192672
rect 45204 192614 453547 192616
rect 45204 192612 45210 192614
rect 453481 192611 453547 192614
rect 1393 192538 1459 192541
rect 554998 192538 555004 192540
rect 1393 192536 555004 192538
rect 1393 192480 1398 192536
rect 1454 192480 555004 192536
rect 1393 192478 555004 192480
rect 1393 192475 1459 192478
rect 554998 192476 555004 192478
rect 555068 192476 555074 192540
rect 580441 192538 580507 192541
rect 583520 192538 584960 192628
rect 580441 192536 584960 192538
rect 580441 192480 580446 192536
rect 580502 192480 584960 192536
rect 580441 192478 584960 192480
rect 580441 192475 580507 192478
rect 583520 192388 584960 192478
rect 158161 191722 158227 191725
rect 347446 191722 347452 191724
rect 158161 191720 347452 191722
rect 158161 191664 158166 191720
rect 158222 191664 347452 191720
rect 158161 191662 347452 191664
rect 158161 191659 158227 191662
rect 347446 191660 347452 191662
rect 347516 191660 347522 191724
rect 278589 191586 278655 191589
rect 347078 191586 347084 191588
rect 278589 191584 347084 191586
rect 278589 191528 278594 191584
rect 278650 191528 347084 191584
rect 278589 191526 347084 191528
rect 278589 191523 278655 191526
rect 347078 191524 347084 191526
rect 347148 191524 347154 191588
rect 55070 191252 55076 191316
rect 55140 191314 55146 191316
rect 370957 191314 371023 191317
rect 55140 191312 371023 191314
rect 55140 191256 370962 191312
rect 371018 191256 371023 191312
rect 55140 191254 371023 191256
rect 55140 191252 55146 191254
rect 370957 191251 371023 191254
rect 57830 191116 57836 191180
rect 57900 191178 57906 191180
rect 550214 191178 550220 191180
rect 57900 191118 550220 191178
rect 57900 191116 57906 191118
rect 550214 191116 550220 191118
rect 550284 191116 550290 191180
rect 2773 191042 2839 191045
rect 551502 191042 551508 191044
rect 2773 191040 551508 191042
rect 2773 190984 2778 191040
rect 2834 190984 551508 191040
rect 2773 190982 551508 190984
rect 2773 190979 2839 190982
rect 551502 190980 551508 190982
rect 551572 190980 551578 191044
rect 211981 190362 212047 190365
rect 350574 190362 350580 190364
rect 211981 190360 350580 190362
rect 211981 190304 211986 190360
rect 212042 190304 350580 190360
rect 211981 190302 350580 190304
rect 211981 190299 212047 190302
rect 350574 190300 350580 190302
rect 350644 190300 350650 190364
rect 61326 190164 61332 190228
rect 61396 190226 61402 190228
rect 365897 190226 365963 190229
rect 61396 190224 365963 190226
rect 61396 190168 365902 190224
rect 365958 190168 365963 190224
rect 61396 190166 365963 190168
rect 61396 190164 61402 190166
rect 365897 190163 365963 190166
rect 50470 190028 50476 190092
rect 50540 190090 50546 190092
rect 373717 190090 373783 190093
rect 50540 190088 373783 190090
rect 50540 190032 373722 190088
rect 373778 190032 373783 190088
rect 50540 190030 373783 190032
rect 50540 190028 50546 190030
rect 373717 190027 373783 190030
rect 41229 189954 41295 189957
rect 377254 189954 377260 189956
rect 41229 189952 377260 189954
rect 41229 189896 41234 189952
rect 41290 189896 377260 189952
rect 41229 189894 377260 189896
rect 41229 189891 41295 189894
rect 377254 189892 377260 189894
rect 377324 189892 377330 189956
rect 53598 189756 53604 189820
rect 53668 189818 53674 189820
rect 399518 189818 399524 189820
rect 53668 189758 399524 189818
rect 53668 189756 53674 189758
rect 399518 189756 399524 189758
rect 399588 189756 399594 189820
rect 55438 189620 55444 189684
rect 55508 189682 55514 189684
rect 407614 189682 407620 189684
rect 55508 189622 407620 189682
rect 55508 189620 55514 189622
rect 407614 189620 407620 189622
rect 407684 189620 407690 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 46381 188866 46447 188869
rect 378910 188866 378916 188868
rect 46381 188864 378916 188866
rect 46381 188808 46386 188864
rect 46442 188808 378916 188864
rect 46381 188806 378916 188808
rect 46381 188803 46447 188806
rect 378910 188804 378916 188806
rect 378980 188804 378986 188868
rect 47894 188668 47900 188732
rect 47964 188730 47970 188732
rect 385534 188730 385540 188732
rect 47964 188670 385540 188730
rect 47964 188668 47970 188670
rect 385534 188668 385540 188670
rect 385604 188668 385610 188732
rect 43662 188532 43668 188596
rect 43732 188594 43738 188596
rect 427077 188594 427143 188597
rect 43732 188592 427143 188594
rect 43732 188536 427082 188592
rect 427138 188536 427143 188592
rect 43732 188534 427143 188536
rect 43732 188532 43738 188534
rect 427077 188531 427143 188534
rect 55622 188396 55628 188460
rect 55692 188458 55698 188460
rect 552238 188458 552244 188460
rect 55692 188398 552244 188458
rect 55692 188396 55698 188398
rect 552238 188396 552244 188398
rect 552308 188396 552314 188460
rect 36670 188260 36676 188324
rect 36740 188322 36746 188324
rect 555417 188322 555483 188325
rect 36740 188320 555483 188322
rect 36740 188264 555422 188320
rect 555478 188264 555483 188320
rect 36740 188262 555483 188264
rect 36740 188260 36746 188262
rect 555417 188259 555483 188262
rect 61510 187580 61516 187644
rect 61580 187642 61586 187644
rect 363229 187642 363295 187645
rect 61580 187640 363295 187642
rect 61580 187584 363234 187640
rect 363290 187584 363295 187640
rect 61580 187582 363295 187584
rect 61580 187580 61586 187582
rect 363229 187579 363295 187582
rect 58566 187444 58572 187508
rect 58636 187506 58642 187508
rect 367093 187506 367159 187509
rect 58636 187504 367159 187506
rect 58636 187448 367098 187504
rect 367154 187448 367159 187504
rect 58636 187446 367159 187448
rect 58636 187444 58642 187446
rect 367093 187443 367159 187446
rect 59118 187308 59124 187372
rect 59188 187370 59194 187372
rect 368657 187370 368723 187373
rect 59188 187368 368723 187370
rect 59188 187312 368662 187368
rect 368718 187312 368723 187368
rect 59188 187310 368723 187312
rect 59188 187308 59194 187310
rect 368657 187307 368723 187310
rect 54702 187172 54708 187236
rect 54772 187234 54778 187236
rect 374913 187234 374979 187237
rect 54772 187232 374979 187234
rect 54772 187176 374918 187232
rect 374974 187176 374979 187232
rect 54772 187174 374979 187176
rect 54772 187172 54778 187174
rect 374913 187171 374979 187174
rect 48681 187098 48747 187101
rect 396206 187098 396212 187100
rect 48681 187096 396212 187098
rect 48681 187040 48686 187096
rect 48742 187040 396212 187096
rect 48681 187038 396212 187040
rect 48681 187035 48747 187038
rect 396206 187036 396212 187038
rect 396276 187036 396282 187100
rect 68001 186962 68067 186965
rect 539542 186962 539548 186964
rect 68001 186960 539548 186962
rect 68001 186904 68006 186960
rect 68062 186904 539548 186960
rect 68001 186902 539548 186904
rect 68001 186899 68067 186902
rect 539542 186900 539548 186902
rect 539612 186900 539618 186964
rect 49550 185812 49556 185876
rect 49620 185874 49626 185876
rect 360326 185874 360332 185876
rect 49620 185814 360332 185874
rect 49620 185812 49626 185814
rect 360326 185812 360332 185814
rect 360396 185812 360402 185876
rect 50654 185676 50660 185740
rect 50724 185738 50730 185740
rect 373533 185738 373599 185741
rect 50724 185736 373599 185738
rect 50724 185680 373538 185736
rect 373594 185680 373599 185736
rect 50724 185678 373599 185680
rect 50724 185676 50730 185678
rect 373533 185675 373599 185678
rect 36854 185540 36860 185604
rect 36924 185602 36930 185604
rect 492765 185602 492831 185605
rect 36924 185600 492831 185602
rect 36924 185544 492770 185600
rect 492826 185544 492831 185600
rect 36924 185542 492831 185544
rect 36924 185540 36930 185542
rect 492765 185539 492831 185542
rect 60590 184588 60596 184652
rect 60660 184650 60666 184652
rect 353518 184650 353524 184652
rect 60660 184590 353524 184650
rect 60660 184588 60666 184590
rect 353518 184588 353524 184590
rect 353588 184588 353594 184652
rect 36445 184514 36511 184517
rect 353702 184514 353708 184516
rect 36445 184512 353708 184514
rect 36445 184456 36450 184512
rect 36506 184456 353708 184512
rect 36445 184454 353708 184456
rect 36445 184451 36511 184454
rect 353702 184452 353708 184454
rect 353772 184452 353778 184516
rect 56317 184378 56383 184381
rect 407982 184378 407988 184380
rect 56317 184376 407988 184378
rect 56317 184320 56322 184376
rect 56378 184320 407988 184376
rect 56317 184318 407988 184320
rect 56317 184315 56383 184318
rect 407982 184316 407988 184318
rect 408052 184316 408058 184380
rect 37038 184180 37044 184244
rect 37108 184242 37114 184244
rect 497273 184242 497339 184245
rect 37108 184240 497339 184242
rect 37108 184184 497278 184240
rect 497334 184184 497339 184240
rect 37108 184182 497339 184184
rect 37108 184180 37114 184182
rect 497273 184179 497339 184182
rect 54886 182820 54892 182884
rect 54956 182882 54962 182884
rect 387006 182882 387012 182884
rect 54956 182822 387012 182882
rect 54956 182820 54962 182822
rect 387006 182820 387012 182822
rect 387076 182820 387082 182884
rect 147673 181658 147739 181661
rect 348366 181658 348372 181660
rect 147673 181656 348372 181658
rect 147673 181600 147678 181656
rect 147734 181600 348372 181656
rect 147673 181598 348372 181600
rect 147673 181595 147739 181598
rect 348366 181596 348372 181598
rect 348436 181596 348442 181660
rect 45369 181522 45435 181525
rect 348734 181522 348740 181524
rect 45369 181520 348740 181522
rect 45369 181464 45374 181520
rect 45430 181464 348740 181520
rect 45369 181462 348740 181464
rect 45369 181459 45435 181462
rect 348734 181460 348740 181462
rect 348804 181460 348810 181524
rect 50286 181324 50292 181388
rect 50356 181386 50362 181388
rect 367134 181386 367140 181388
rect 50356 181326 367140 181386
rect 50356 181324 50362 181326
rect 367134 181324 367140 181326
rect 367204 181324 367210 181388
rect 108297 180706 108363 180709
rect 395286 180706 395292 180708
rect 108297 180704 395292 180706
rect 108297 180648 108302 180704
rect 108358 180648 395292 180704
rect 108297 180646 395292 180648
rect 108297 180643 108363 180646
rect 395286 180644 395292 180646
rect 395356 180644 395362 180708
rect 41086 180508 41092 180572
rect 41156 180570 41162 180572
rect 329189 180570 329255 180573
rect 41156 180568 329255 180570
rect 41156 180512 329194 180568
rect 329250 180512 329255 180568
rect 41156 180510 329255 180512
rect 41156 180508 41162 180510
rect 329189 180507 329255 180510
rect 49366 180372 49372 180436
rect 49436 180434 49442 180436
rect 382774 180434 382780 180436
rect 49436 180374 382780 180434
rect 49436 180372 49442 180374
rect 382774 180372 382780 180374
rect 382844 180372 382850 180436
rect 41045 180298 41111 180301
rect 391238 180298 391244 180300
rect 41045 180296 391244 180298
rect 41045 180240 41050 180296
rect 41106 180240 391244 180296
rect 41045 180238 391244 180240
rect 41045 180235 41111 180238
rect 391238 180236 391244 180238
rect 391308 180236 391314 180300
rect 34278 180100 34284 180164
rect 34348 180162 34354 180164
rect 458173 180162 458239 180165
rect 34348 180160 458239 180162
rect 34348 180104 458178 180160
rect 458234 180104 458239 180160
rect 34348 180102 458239 180104
rect 34348 180100 34354 180102
rect 458173 180099 458239 180102
rect 77385 180026 77451 180029
rect 539726 180026 539732 180028
rect 77385 180024 539732 180026
rect 77385 179968 77390 180024
rect 77446 179968 539732 180024
rect 77385 179966 539732 179968
rect 77385 179963 77451 179966
rect 539726 179964 539732 179966
rect 539796 179964 539802 180028
rect 172053 179890 172119 179893
rect 350758 179890 350764 179892
rect 172053 179888 350764 179890
rect 172053 179832 172058 179888
rect 172114 179832 350764 179888
rect 172053 179830 350764 179832
rect 172053 179827 172119 179830
rect 350758 179828 350764 179830
rect 350828 179828 350834 179892
rect 580717 179210 580783 179213
rect 583520 179210 584960 179300
rect 580717 179208 584960 179210
rect 580717 179152 580722 179208
rect 580778 179152 584960 179208
rect 580717 179150 584960 179152
rect 580717 179147 580783 179150
rect 583520 179060 584960 179150
rect 46657 178802 46723 178805
rect 364558 178802 364564 178804
rect 46657 178800 364564 178802
rect 46657 178744 46662 178800
rect 46718 178744 364564 178800
rect 46657 178742 364564 178744
rect 46657 178739 46723 178742
rect 364558 178740 364564 178742
rect 364628 178740 364634 178804
rect 45870 178604 45876 178668
rect 45940 178666 45946 178668
rect 376385 178666 376451 178669
rect 45940 178664 376451 178666
rect 45940 178608 376390 178664
rect 376446 178608 376451 178664
rect 45940 178606 376451 178608
rect 45940 178604 45946 178606
rect 376385 178603 376451 178606
rect 61694 177788 61700 177852
rect 61764 177850 61770 177852
rect 362953 177850 363019 177853
rect 61764 177848 363019 177850
rect 61764 177792 362958 177848
rect 363014 177792 363019 177848
rect 61764 177790 363019 177792
rect 61764 177788 61770 177790
rect 362953 177787 363019 177790
rect 44633 177714 44699 177717
rect 349654 177714 349660 177716
rect 44633 177712 349660 177714
rect 44633 177656 44638 177712
rect 44694 177656 349660 177712
rect 44633 177654 349660 177656
rect 44633 177651 44699 177654
rect 349654 177652 349660 177654
rect 349724 177652 349730 177716
rect 50429 177578 50495 177581
rect 378726 177578 378732 177580
rect 50429 177576 378732 177578
rect 50429 177520 50434 177576
rect 50490 177520 378732 177576
rect 50429 177518 378732 177520
rect 50429 177515 50495 177518
rect 378726 177516 378732 177518
rect 378796 177516 378802 177580
rect 49182 177380 49188 177444
rect 49252 177442 49258 177444
rect 392526 177442 392532 177444
rect 49252 177382 392532 177442
rect 49252 177380 49258 177382
rect 392526 177380 392532 177382
rect 392596 177380 392602 177444
rect 73337 177306 73403 177309
rect 541014 177306 541020 177308
rect 73337 177304 541020 177306
rect 73337 177248 73342 177304
rect 73398 177248 541020 177304
rect 73337 177246 541020 177248
rect 73337 177243 73403 177246
rect 541014 177244 541020 177246
rect 541084 177244 541090 177308
rect -960 175796 480 176036
rect 60406 174932 60412 174996
rect 60476 174994 60482 174996
rect 372613 174994 372679 174997
rect 60476 174992 372679 174994
rect 60476 174936 372618 174992
rect 372674 174936 372679 174992
rect 60476 174934 372679 174936
rect 60476 174932 60482 174934
rect 372613 174931 372679 174934
rect 52310 174796 52316 174860
rect 52380 174858 52386 174860
rect 376017 174858 376083 174861
rect 52380 174856 376083 174858
rect 52380 174800 376022 174856
rect 376078 174800 376083 174856
rect 52380 174798 376083 174800
rect 52380 174796 52386 174798
rect 376017 174795 376083 174798
rect 46606 174660 46612 174724
rect 46676 174722 46682 174724
rect 542670 174722 542676 174724
rect 46676 174662 542676 174722
rect 46676 174660 46682 174662
rect 542670 174660 542676 174662
rect 542740 174660 542746 174724
rect 41086 174524 41092 174588
rect 41156 174586 41162 174588
rect 553209 174586 553275 174589
rect 41156 174584 553275 174586
rect 41156 174528 553214 174584
rect 553270 174528 553275 174584
rect 41156 174526 553275 174528
rect 41156 174524 41162 174526
rect 553209 174523 553275 174526
rect 41270 173300 41276 173364
rect 41340 173362 41346 173364
rect 371233 173362 371299 173365
rect 41340 173360 371299 173362
rect 41340 173304 371238 173360
rect 371294 173304 371299 173360
rect 41340 173302 371299 173304
rect 41340 173300 41346 173302
rect 371233 173299 371299 173302
rect 50838 173164 50844 173228
rect 50908 173226 50914 173228
rect 570505 173226 570571 173229
rect 50908 173224 570571 173226
rect 50908 173168 570510 173224
rect 570566 173168 570571 173224
rect 50908 173166 570571 173168
rect 50908 173164 50914 173166
rect 570505 173163 570571 173166
rect 195237 172410 195303 172413
rect 346894 172410 346900 172412
rect 195237 172408 346900 172410
rect 195237 172352 195242 172408
rect 195298 172352 346900 172408
rect 195237 172350 346900 172352
rect 195237 172347 195303 172350
rect 346894 172348 346900 172350
rect 346964 172348 346970 172412
rect 53414 172212 53420 172276
rect 53484 172274 53490 172276
rect 377438 172274 377444 172276
rect 53484 172214 377444 172274
rect 53484 172212 53490 172214
rect 377438 172212 377444 172214
rect 377508 172212 377514 172276
rect 41270 172076 41276 172140
rect 41340 172138 41346 172140
rect 373206 172138 373212 172140
rect 41340 172078 373212 172138
rect 41340 172076 41346 172078
rect 373206 172076 373212 172078
rect 373276 172076 373282 172140
rect 46238 171940 46244 172004
rect 46308 172002 46314 172004
rect 387742 172002 387748 172004
rect 46308 171942 387748 172002
rect 46308 171940 46314 171942
rect 387742 171940 387748 171942
rect 387812 171940 387818 172004
rect 31753 171866 31819 171869
rect 389950 171866 389956 171868
rect 31753 171864 389956 171866
rect 31753 171808 31758 171864
rect 31814 171808 389956 171864
rect 31753 171806 389956 171808
rect 31753 171803 31819 171806
rect 389950 171804 389956 171806
rect 390020 171804 390026 171868
rect 46054 171668 46060 171732
rect 46124 171730 46130 171732
rect 543958 171730 543964 171732
rect 46124 171670 543964 171730
rect 46124 171668 46130 171670
rect 543958 171668 543964 171670
rect 544028 171668 544034 171732
rect 43662 170444 43668 170508
rect 43732 170506 43738 170508
rect 392710 170506 392716 170508
rect 43732 170446 392716 170506
rect 43732 170444 43738 170446
rect 392710 170444 392716 170446
rect 392780 170444 392786 170508
rect 157885 170370 157951 170373
rect 563278 170370 563284 170372
rect 157885 170368 563284 170370
rect 157885 170312 157890 170368
rect 157946 170312 563284 170368
rect 157885 170310 563284 170312
rect 157885 170307 157951 170310
rect 563278 170308 563284 170310
rect 563348 170308 563354 170372
rect 41638 168948 41644 169012
rect 41708 169010 41714 169012
rect 488901 169010 488967 169013
rect 41708 169008 488967 169010
rect 41708 168952 488906 169008
rect 488962 168952 488967 169008
rect 41708 168950 488967 168952
rect 41708 168948 41714 168950
rect 488901 168947 488967 168950
rect 39430 167724 39436 167788
rect 39500 167786 39506 167788
rect 502425 167786 502491 167789
rect 39500 167784 502491 167786
rect 39500 167728 502430 167784
rect 502486 167728 502491 167784
rect 39500 167726 502491 167728
rect 39500 167724 39506 167726
rect 502425 167723 502491 167726
rect 77385 167650 77451 167653
rect 559046 167650 559052 167652
rect 77385 167648 559052 167650
rect 77385 167592 77390 167648
rect 77446 167592 559052 167648
rect 77385 167590 559052 167592
rect 77385 167587 77451 167590
rect 559046 167588 559052 167590
rect 559116 167588 559122 167652
rect 54518 166500 54524 166564
rect 54588 166562 54594 166564
rect 363454 166562 363460 166564
rect 54588 166502 363460 166562
rect 54588 166500 54594 166502
rect 363454 166500 363460 166502
rect 363524 166500 363530 166564
rect 384573 166562 384639 166565
rect 545430 166562 545436 166564
rect 384573 166560 545436 166562
rect 384573 166504 384578 166560
rect 384634 166504 545436 166560
rect 384573 166502 545436 166504
rect 384573 166499 384639 166502
rect 545430 166500 545436 166502
rect 545500 166500 545506 166564
rect 53230 166364 53236 166428
rect 53300 166426 53306 166428
rect 393957 166426 394023 166429
rect 53300 166424 394023 166426
rect 53300 166368 393962 166424
rect 394018 166368 394023 166424
rect 53300 166366 394023 166368
rect 53300 166364 53306 166366
rect 393957 166363 394023 166366
rect 404261 166426 404327 166429
rect 562174 166426 562180 166428
rect 404261 166424 562180 166426
rect 404261 166368 404266 166424
rect 404322 166368 562180 166424
rect 404261 166366 562180 166368
rect 404261 166363 404327 166366
rect 562174 166364 562180 166366
rect 562244 166364 562250 166428
rect 40718 166228 40724 166292
rect 40788 166290 40794 166292
rect 383929 166290 383995 166293
rect 40788 166288 383995 166290
rect 40788 166232 383934 166288
rect 383990 166232 383995 166288
rect 40788 166230 383995 166232
rect 40788 166228 40794 166230
rect 383929 166227 383995 166230
rect 395981 166290 396047 166293
rect 563278 166290 563284 166292
rect 395981 166288 563284 166290
rect 395981 166232 395986 166288
rect 396042 166232 563284 166288
rect 395981 166230 563284 166232
rect 395981 166227 396047 166230
rect 563278 166228 563284 166230
rect 563348 166228 563354 166292
rect 583520 165732 584960 165972
rect 321461 163706 321527 163709
rect 399334 163706 399340 163708
rect 321461 163704 399340 163706
rect 321461 163648 321466 163704
rect 321522 163648 399340 163704
rect 321461 163646 399340 163648
rect 321461 163643 321527 163646
rect 399334 163644 399340 163646
rect 399404 163644 399410 163708
rect 389766 163508 389772 163572
rect 389836 163570 389842 163572
rect 552197 163570 552263 163573
rect 389836 163568 552263 163570
rect 389836 163512 552202 163568
rect 552258 163512 552263 163568
rect 389836 163510 552263 163512
rect 389836 163508 389842 163510
rect 552197 163507 552263 163510
rect 271229 163434 271295 163437
rect 358118 163434 358124 163436
rect 271229 163432 358124 163434
rect 271229 163376 271234 163432
rect 271290 163376 358124 163432
rect 271229 163374 358124 163376
rect 271229 163371 271295 163374
rect 358118 163372 358124 163374
rect 358188 163372 358194 163436
rect 374729 163434 374795 163437
rect 541198 163434 541204 163436
rect 374729 163432 541204 163434
rect 374729 163376 374734 163432
rect 374790 163376 541204 163432
rect 374729 163374 541204 163376
rect 374729 163371 374795 163374
rect 541198 163372 541204 163374
rect 541268 163372 541274 163436
rect -960 162740 480 162980
rect 251265 162074 251331 162077
rect 403566 162074 403572 162076
rect 251265 162072 403572 162074
rect 251265 162016 251270 162072
rect 251326 162016 403572 162072
rect 251265 162014 403572 162016
rect 251265 162011 251331 162014
rect 403566 162012 403572 162014
rect 403636 162012 403642 162076
rect 402421 161258 402487 161261
rect 549846 161258 549852 161260
rect 402421 161256 549852 161258
rect 402421 161200 402426 161256
rect 402482 161200 549852 161256
rect 402421 161198 549852 161200
rect 402421 161195 402487 161198
rect 549846 161196 549852 161198
rect 549916 161196 549922 161260
rect 387149 161122 387215 161125
rect 548190 161122 548196 161124
rect 387149 161120 548196 161122
rect 387149 161064 387154 161120
rect 387210 161064 548196 161120
rect 387149 161062 548196 161064
rect 387149 161059 387215 161062
rect 548190 161060 548196 161062
rect 548260 161060 548266 161124
rect 57646 160924 57652 160988
rect 57716 160986 57722 160988
rect 371734 160986 371740 160988
rect 57716 160926 371740 160986
rect 57716 160924 57722 160926
rect 371734 160924 371740 160926
rect 371804 160924 371810 160988
rect 391054 160924 391060 160988
rect 391124 160986 391130 160988
rect 552238 160986 552244 160988
rect 391124 160926 552244 160986
rect 391124 160924 391130 160926
rect 552238 160924 552244 160926
rect 552308 160924 552314 160988
rect 110413 160850 110479 160853
rect 547454 160850 547460 160852
rect 110413 160848 547460 160850
rect 110413 160792 110418 160848
rect 110474 160792 547460 160848
rect 110413 160790 547460 160792
rect 110413 160787 110479 160790
rect 547454 160788 547460 160790
rect 547524 160788 547530 160852
rect 28809 160714 28875 160717
rect 552422 160714 552428 160716
rect 28809 160712 552428 160714
rect 28809 160656 28814 160712
rect 28870 160656 552428 160712
rect 28809 160654 552428 160656
rect 28809 160651 28875 160654
rect 552422 160652 552428 160654
rect 552492 160652 552498 160716
rect 56869 159626 56935 159629
rect 355174 159626 355180 159628
rect 56869 159624 355180 159626
rect 56869 159568 56874 159624
rect 56930 159568 355180 159624
rect 56869 159566 355180 159568
rect 56869 159563 56935 159566
rect 355174 159564 355180 159566
rect 355244 159564 355250 159628
rect 401133 159626 401199 159629
rect 543774 159626 543780 159628
rect 401133 159624 543780 159626
rect 401133 159568 401138 159624
rect 401194 159568 543780 159624
rect 401133 159566 543780 159568
rect 401133 159563 401199 159566
rect 543774 159564 543780 159566
rect 543844 159564 543850 159628
rect 57462 159428 57468 159492
rect 57532 159490 57538 159492
rect 359549 159490 359615 159493
rect 57532 159488 359615 159490
rect 57532 159432 359554 159488
rect 359610 159432 359615 159488
rect 57532 159430 359615 159432
rect 57532 159428 57538 159430
rect 359549 159427 359615 159430
rect 393221 159490 393287 159493
rect 545798 159490 545804 159492
rect 393221 159488 545804 159490
rect 393221 159432 393226 159488
rect 393282 159432 545804 159488
rect 393221 159430 545804 159432
rect 393221 159427 393287 159430
rect 545798 159428 545804 159430
rect 545868 159428 545874 159492
rect 57789 159354 57855 159357
rect 563094 159354 563100 159356
rect 57789 159352 563100 159354
rect 57789 159296 57794 159352
rect 57850 159296 563100 159352
rect 57789 159294 563100 159296
rect 57789 159291 57855 159294
rect 563094 159292 563100 159294
rect 563164 159292 563170 159356
rect 334065 158674 334131 158677
rect 539358 158674 539364 158676
rect 334065 158672 539364 158674
rect 334065 158616 334070 158672
rect 334126 158616 539364 158672
rect 334065 158614 539364 158616
rect 334065 158611 334131 158614
rect 539358 158612 539364 158614
rect 539428 158612 539434 158676
rect 56961 158538 57027 158541
rect 352046 158538 352052 158540
rect 56961 158536 352052 158538
rect 56961 158480 56966 158536
rect 57022 158480 352052 158536
rect 56961 158478 352052 158480
rect 56961 158475 57027 158478
rect 352046 158476 352052 158478
rect 352116 158476 352122 158540
rect 373349 158538 373415 158541
rect 549662 158538 549668 158540
rect 373349 158536 549668 158538
rect 373349 158480 373354 158536
rect 373410 158480 549668 158536
rect 373349 158478 549668 158480
rect 373349 158475 373415 158478
rect 549662 158476 549668 158478
rect 549732 158476 549738 158540
rect 58934 158340 58940 158404
rect 59004 158402 59010 158404
rect 373993 158402 374059 158405
rect 59004 158400 374059 158402
rect 59004 158344 373998 158400
rect 374054 158344 374059 158400
rect 59004 158342 374059 158344
rect 59004 158340 59010 158342
rect 373993 158339 374059 158342
rect 46422 158204 46428 158268
rect 46492 158266 46498 158268
rect 544142 158266 544148 158268
rect 46492 158206 544148 158266
rect 46492 158204 46498 158206
rect 544142 158204 544148 158206
rect 544212 158204 544218 158268
rect 26877 158130 26943 158133
rect 570781 158130 570847 158133
rect 26877 158128 570847 158130
rect 26877 158072 26882 158128
rect 26938 158072 570786 158128
rect 570842 158072 570847 158128
rect 26877 158070 570847 158072
rect 26877 158067 26943 158070
rect 570781 158067 570847 158070
rect 27061 157994 27127 157997
rect 574921 157994 574987 157997
rect 27061 157992 574987 157994
rect 27061 157936 27066 157992
rect 27122 157936 574926 157992
rect 574982 157936 574987 157992
rect 27061 157934 574987 157936
rect 27061 157931 27127 157934
rect 574921 157931 574987 157934
rect 398598 157252 398604 157316
rect 398668 157314 398674 157316
rect 552606 157314 552612 157316
rect 398668 157254 552612 157314
rect 398668 157252 398674 157254
rect 552606 157252 552612 157254
rect 552676 157252 552682 157316
rect 409086 157116 409092 157180
rect 409156 157178 409162 157180
rect 569493 157178 569559 157181
rect 409156 157176 569559 157178
rect 409156 157120 569498 157176
rect 569554 157120 569559 157176
rect 409156 157118 569559 157120
rect 409156 157116 409162 157118
rect 569493 157115 569559 157118
rect 40902 156980 40908 157044
rect 40972 157042 40978 157044
rect 384573 157042 384639 157045
rect 40972 157040 384639 157042
rect 40972 156984 384578 157040
rect 384634 156984 384639 157040
rect 40972 156982 384639 156984
rect 40972 156980 40978 156982
rect 384573 156979 384639 156982
rect 409454 156980 409460 157044
rect 409524 157042 409530 157044
rect 575657 157042 575723 157045
rect 409524 157040 575723 157042
rect 409524 156984 575662 157040
rect 575718 156984 575723 157040
rect 409524 156982 575723 156984
rect 409524 156980 409530 156982
rect 575657 156979 575723 156982
rect 35566 156844 35572 156908
rect 35636 156906 35642 156908
rect 440601 156906 440667 156909
rect 35636 156904 440667 156906
rect 35636 156848 440606 156904
rect 440662 156848 440667 156904
rect 35636 156846 440667 156848
rect 35636 156844 35642 156846
rect 440601 156843 440667 156846
rect 46473 156770 46539 156773
rect 539910 156770 539916 156772
rect 46473 156768 539916 156770
rect 46473 156712 46478 156768
rect 46534 156712 539916 156768
rect 46473 156710 539916 156712
rect 46473 156707 46539 156710
rect 539910 156708 539916 156710
rect 539980 156708 539986 156772
rect 19057 156634 19123 156637
rect 563094 156634 563100 156636
rect 19057 156632 563100 156634
rect 19057 156576 19062 156632
rect 19118 156576 563100 156632
rect 19057 156574 563100 156576
rect 19057 156571 19123 156574
rect 563094 156572 563100 156574
rect 563164 156572 563170 156636
rect 46381 155956 46447 155957
rect 46381 155954 46428 155956
rect 46336 155952 46428 155954
rect 46336 155896 46386 155952
rect 46336 155894 46428 155896
rect 46381 155892 46428 155894
rect 46492 155892 46498 155956
rect 46381 155891 46447 155892
rect 317597 155818 317663 155821
rect 351862 155818 351868 155820
rect 317597 155816 351868 155818
rect 317597 155760 317602 155816
rect 317658 155760 351868 155816
rect 317597 155758 351868 155760
rect 317597 155755 317663 155758
rect 351862 155756 351868 155758
rect 351932 155756 351938 155820
rect 60038 155620 60044 155684
rect 60108 155682 60114 155684
rect 365713 155682 365779 155685
rect 60108 155680 365779 155682
rect 60108 155624 365718 155680
rect 365774 155624 365779 155680
rect 60108 155622 365779 155624
rect 60108 155620 60114 155622
rect 365713 155619 365779 155622
rect 384665 155682 384731 155685
rect 543406 155682 543412 155684
rect 384665 155680 543412 155682
rect 384665 155624 384670 155680
rect 384726 155624 543412 155680
rect 384665 155622 543412 155624
rect 384665 155619 384731 155622
rect 543406 155620 543412 155622
rect 543476 155620 543482 155684
rect 51717 155546 51783 155549
rect 364374 155546 364380 155548
rect 51717 155544 364380 155546
rect 51717 155488 51722 155544
rect 51778 155488 364380 155544
rect 51717 155486 364380 155488
rect 51717 155483 51783 155486
rect 364374 155484 364380 155486
rect 364444 155484 364450 155548
rect 384205 155546 384271 155549
rect 546125 155546 546191 155549
rect 384205 155544 546191 155546
rect 384205 155488 384210 155544
rect 384266 155488 546130 155544
rect 546186 155488 546191 155544
rect 384205 155486 546191 155488
rect 384205 155483 384271 155486
rect 546125 155483 546191 155486
rect 45093 155410 45159 155413
rect 360142 155410 360148 155412
rect 45093 155408 360148 155410
rect 45093 155352 45098 155408
rect 45154 155352 360148 155408
rect 45093 155350 360148 155352
rect 45093 155347 45159 155350
rect 360142 155348 360148 155350
rect 360212 155348 360218 155412
rect 375281 155410 375347 155413
rect 545246 155410 545252 155412
rect 375281 155408 545252 155410
rect 375281 155352 375286 155408
rect 375342 155352 545252 155408
rect 375281 155350 545252 155352
rect 375281 155347 375347 155350
rect 545246 155348 545252 155350
rect 545316 155348 545322 155412
rect 58750 155212 58756 155276
rect 58820 155274 58826 155276
rect 407798 155274 407804 155276
rect 58820 155214 407804 155274
rect 58820 155212 58826 155214
rect 407798 155212 407804 155214
rect 407868 155212 407874 155276
rect 406326 154260 406332 154324
rect 406396 154322 406402 154324
rect 547822 154322 547828 154324
rect 406396 154262 547828 154322
rect 406396 154260 406402 154262
rect 547822 154260 547828 154262
rect 547892 154260 547898 154324
rect 381721 154186 381787 154189
rect 542854 154186 542860 154188
rect 381721 154184 542860 154186
rect 381721 154128 381726 154184
rect 381782 154128 542860 154184
rect 381721 154126 542860 154128
rect 381721 154123 381787 154126
rect 542854 154124 542860 154126
rect 542924 154124 542930 154188
rect 57513 154050 57579 154053
rect 360694 154050 360700 154052
rect 57513 154048 360700 154050
rect 57513 153992 57518 154048
rect 57574 153992 360700 154048
rect 57513 153990 360700 153992
rect 57513 153987 57579 153990
rect 360694 153988 360700 153990
rect 360764 153988 360770 154052
rect 363638 153988 363644 154052
rect 363708 154050 363714 154052
rect 549294 154050 549300 154052
rect 363708 153990 549300 154050
rect 363708 153988 363714 153990
rect 549294 153988 549300 153990
rect 549364 153988 549370 154052
rect 111885 153914 111951 153917
rect 545062 153914 545068 153916
rect 111885 153912 545068 153914
rect 111885 153856 111890 153912
rect 111946 153856 545068 153912
rect 111885 153854 545068 153856
rect 111885 153851 111951 153854
rect 545062 153852 545068 153854
rect 545132 153852 545138 153916
rect 24209 153778 24275 153781
rect 551502 153778 551508 153780
rect 24209 153776 551508 153778
rect 24209 153720 24214 153776
rect 24270 153720 551508 153776
rect 24209 153718 551508 153720
rect 24209 153715 24275 153718
rect 551502 153716 551508 153718
rect 551572 153716 551578 153780
rect 61929 153098 61995 153101
rect 168373 153098 168439 153101
rect 61929 153096 168439 153098
rect 61929 153040 61934 153096
rect 61990 153040 168378 153096
rect 168434 153040 168439 153096
rect 61929 153038 168439 153040
rect 61929 153035 61995 153038
rect 168373 153035 168439 153038
rect 396574 153036 396580 153100
rect 396644 153098 396650 153100
rect 463785 153098 463851 153101
rect 396644 153096 463851 153098
rect 396644 153040 463790 153096
rect 463846 153040 463851 153096
rect 396644 153038 463851 153040
rect 396644 153036 396650 153038
rect 463785 153035 463851 153038
rect 48814 152900 48820 152964
rect 48884 152962 48890 152964
rect 204897 152962 204963 152965
rect 48884 152960 204963 152962
rect 48884 152904 204902 152960
rect 204958 152904 204963 152960
rect 48884 152902 204963 152904
rect 48884 152900 48890 152902
rect 204897 152899 204963 152902
rect 341793 152962 341859 152965
rect 356646 152962 356652 152964
rect 341793 152960 356652 152962
rect 341793 152904 341798 152960
rect 341854 152904 356652 152960
rect 341793 152902 356652 152904
rect 341793 152899 341859 152902
rect 356646 152900 356652 152902
rect 356716 152900 356722 152964
rect 400806 152900 400812 152964
rect 400876 152962 400882 152964
rect 482461 152962 482527 152965
rect 400876 152960 482527 152962
rect 400876 152904 482466 152960
rect 482522 152904 482527 152960
rect 400876 152902 482527 152904
rect 400876 152900 400882 152902
rect 482461 152899 482527 152902
rect 47710 152764 47716 152828
rect 47780 152826 47786 152828
rect 170121 152826 170187 152829
rect 47780 152824 170187 152826
rect 47780 152768 170126 152824
rect 170182 152768 170187 152824
rect 47780 152766 170187 152768
rect 47780 152764 47786 152766
rect 170121 152763 170187 152766
rect 179137 152826 179203 152829
rect 377397 152826 377463 152829
rect 179137 152824 377463 152826
rect 179137 152768 179142 152824
rect 179198 152768 377402 152824
rect 377458 152768 377463 152824
rect 179137 152766 377463 152768
rect 179137 152763 179203 152766
rect 377397 152763 377463 152766
rect 395470 152764 395476 152828
rect 395540 152826 395546 152828
rect 498561 152826 498627 152829
rect 395540 152824 498627 152826
rect 395540 152768 498566 152824
rect 498622 152768 498627 152824
rect 395540 152766 498627 152768
rect 395540 152764 395546 152766
rect 498561 152763 498627 152766
rect 19149 152690 19215 152693
rect 153377 152690 153443 152693
rect 19149 152688 153443 152690
rect 19149 152632 19154 152688
rect 19210 152632 153382 152688
rect 153438 152632 153443 152688
rect 19149 152630 153443 152632
rect 19149 152627 19215 152630
rect 153377 152627 153443 152630
rect 199101 152690 199167 152693
rect 398097 152690 398163 152693
rect 199101 152688 398163 152690
rect 199101 152632 199106 152688
rect 199162 152632 398102 152688
rect 398158 152632 398163 152688
rect 199101 152630 398163 152632
rect 199101 152627 199167 152630
rect 398097 152627 398163 152630
rect 408534 152628 408540 152692
rect 408604 152690 408610 152692
rect 409045 152690 409111 152693
rect 408604 152688 409111 152690
rect 408604 152632 409050 152688
rect 409106 152632 409111 152688
rect 408604 152630 409111 152632
rect 408604 152628 408610 152630
rect 409045 152627 409111 152630
rect 409822 152628 409828 152692
rect 409892 152690 409898 152692
rect 566181 152690 566247 152693
rect 409892 152688 566247 152690
rect 409892 152632 566186 152688
rect 566242 152632 566247 152688
rect 409892 152630 566247 152632
rect 409892 152628 409898 152630
rect 566181 152627 566247 152630
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 28625 152554 28691 152557
rect 240961 152554 241027 152557
rect 28625 152552 241027 152554
rect 28625 152496 28630 152552
rect 28686 152496 240966 152552
rect 241022 152496 241027 152552
rect 28625 152494 241027 152496
rect 28625 152491 28691 152494
rect 240961 152491 241027 152494
rect 325049 152554 325115 152557
rect 354438 152554 354444 152556
rect 325049 152552 354444 152554
rect 325049 152496 325054 152552
rect 325110 152496 354444 152552
rect 325049 152494 354444 152496
rect 325049 152491 325115 152494
rect 354438 152492 354444 152494
rect 354508 152492 354514 152556
rect 381486 152492 381492 152556
rect 381556 152554 381562 152556
rect 553894 152554 553900 152556
rect 381556 152494 553900 152554
rect 381556 152492 381562 152494
rect 553894 152492 553900 152494
rect 553964 152492 553970 152556
rect 583520 152540 584960 152630
rect 72877 152418 72943 152421
rect 370446 152418 370452 152420
rect 72877 152416 370452 152418
rect 72877 152360 72882 152416
rect 72938 152360 370452 152416
rect 72877 152358 370452 152360
rect 72877 152355 72943 152358
rect 370446 152356 370452 152358
rect 370516 152356 370522 152420
rect 376109 152418 376175 152421
rect 580165 152418 580231 152421
rect 376109 152416 580231 152418
rect 376109 152360 376114 152416
rect 376170 152360 580170 152416
rect 580226 152360 580231 152416
rect 376109 152358 580231 152360
rect 376109 152355 376175 152358
rect 580165 152355 580231 152358
rect 59445 151738 59511 151741
rect 59629 151738 59695 151741
rect 59445 151736 59695 151738
rect 59445 151680 59450 151736
rect 59506 151680 59634 151736
rect 59690 151680 59695 151736
rect 59445 151678 59695 151680
rect 59445 151675 59511 151678
rect 59629 151675 59695 151678
rect 537569 151738 537635 151741
rect 541382 151738 541388 151740
rect 537569 151736 541388 151738
rect 537569 151680 537574 151736
rect 537630 151680 541388 151736
rect 537569 151678 541388 151680
rect 537569 151675 537635 151678
rect 541382 151676 541388 151678
rect 541452 151676 541458 151740
rect 59721 151466 59787 151469
rect 59997 151466 60063 151469
rect 59721 151464 60063 151466
rect 59721 151408 59726 151464
rect 59782 151408 60002 151464
rect 60058 151408 60063 151464
rect 59721 151406 60063 151408
rect 59721 151403 59787 151406
rect 59997 151403 60063 151406
rect 410190 151404 410196 151468
rect 410260 151466 410266 151468
rect 552289 151466 552355 151469
rect 410260 151464 552355 151466
rect 410260 151408 552294 151464
rect 552350 151408 552355 151464
rect 410260 151406 552355 151408
rect 410260 151404 410266 151406
rect 552289 151403 552355 151406
rect 59721 151330 59787 151333
rect 117313 151330 117379 151333
rect 59721 151328 117379 151330
rect 59721 151272 59726 151328
rect 59782 151272 117318 151328
rect 117374 151272 117379 151328
rect 59721 151270 117379 151272
rect 59721 151267 59787 151270
rect 117313 151267 117379 151270
rect 410517 151330 410583 151333
rect 559046 151330 559052 151332
rect 410517 151328 559052 151330
rect 410517 151272 410522 151328
rect 410578 151272 559052 151328
rect 410517 151270 559052 151272
rect 410517 151267 410583 151270
rect 559046 151268 559052 151270
rect 559116 151268 559122 151332
rect 55765 151194 55831 151197
rect 349470 151194 349476 151196
rect 55765 151192 349476 151194
rect 55765 151136 55770 151192
rect 55826 151136 349476 151192
rect 55765 151134 349476 151136
rect 55765 151131 55831 151134
rect 349470 151132 349476 151134
rect 349540 151132 349546 151196
rect 359590 151132 359596 151196
rect 359660 151194 359666 151196
rect 554998 151194 555004 151196
rect 359660 151134 555004 151194
rect 359660 151132 359666 151134
rect 554998 151132 555004 151134
rect 555068 151132 555074 151196
rect 57278 150996 57284 151060
rect 57348 151058 57354 151060
rect 372654 151058 372660 151060
rect 57348 150998 372660 151058
rect 57348 150996 57354 150998
rect 372654 150996 372660 150998
rect 372724 150996 372730 151060
rect 404854 150996 404860 151060
rect 404924 151058 404930 151060
rect 554221 151058 554287 151061
rect 404924 151056 554287 151058
rect 404924 151000 554226 151056
rect 554282 151000 554287 151056
rect 404924 150998 554287 151000
rect 404924 150996 404930 150998
rect 554221 150995 554287 150998
rect 539174 150452 539180 150516
rect 539244 150514 539250 150516
rect 540094 150514 540100 150516
rect 539244 150454 540100 150514
rect 539244 150452 539250 150454
rect 540094 150452 540100 150454
rect 540164 150452 540170 150516
rect 538765 150378 538831 150381
rect 568941 150378 569007 150381
rect 538765 150376 569007 150378
rect 538765 150320 538770 150376
rect 538826 150320 568946 150376
rect 569002 150320 569007 150376
rect 538765 150318 569007 150320
rect 538765 150315 538831 150318
rect 568941 150315 569007 150318
rect 538857 150242 538923 150245
rect 539869 150242 539935 150245
rect 556153 150242 556219 150245
rect 538857 150240 539794 150242
rect 538857 150184 538862 150240
rect 538918 150184 539794 150240
rect 538857 150182 539794 150184
rect 538857 150179 538923 150182
rect 59537 150106 59603 150109
rect 59997 150106 60063 150109
rect 59537 150104 60063 150106
rect 59537 150048 59542 150104
rect 59598 150048 60002 150104
rect 60058 150048 60063 150104
rect 59537 150046 60063 150048
rect 59537 150043 59603 150046
rect 59997 150043 60063 150046
rect 60222 150044 60228 150108
rect 60292 150106 60298 150108
rect 61326 150106 61332 150108
rect 60292 150046 61332 150106
rect 60292 150044 60298 150046
rect 61326 150044 61332 150046
rect 61396 150044 61402 150108
rect 399937 150106 400003 150109
rect 539734 150106 539794 150182
rect 539869 150240 556219 150242
rect 539869 150184 539874 150240
rect 539930 150184 556158 150240
rect 556214 150184 556219 150240
rect 539869 150182 556219 150184
rect 539869 150179 539935 150182
rect 556153 150179 556219 150182
rect 399937 150104 539610 150106
rect 399937 150048 399942 150104
rect 399998 150048 539610 150104
rect 399937 150046 539610 150048
rect 539734 150046 553410 150106
rect 399937 150043 400003 150046
rect 59905 149970 59971 149973
rect 61510 149970 61516 149972
rect 59905 149968 61516 149970
rect -960 149834 480 149924
rect 59905 149912 59910 149968
rect 59966 149912 61516 149968
rect 59905 149910 61516 149912
rect 59905 149907 59971 149910
rect 61510 149908 61516 149910
rect 61580 149908 61586 149972
rect 386321 149970 386387 149973
rect 539041 149970 539107 149973
rect 386321 149968 539107 149970
rect 386321 149912 386326 149968
rect 386382 149912 539046 149968
rect 539102 149912 539107 149968
rect 386321 149910 539107 149912
rect 386321 149907 386387 149910
rect 539041 149907 539107 149910
rect 539317 149970 539383 149973
rect 539550 149970 539610 150046
rect 547270 149970 547276 149972
rect 539317 149968 539426 149970
rect 539317 149912 539322 149968
rect 539378 149912 539426 149968
rect 539317 149907 539426 149912
rect 539550 149910 547276 149970
rect 547270 149908 547276 149910
rect 547340 149908 547346 149972
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect 539366 149804 539426 149907
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 540697 149698 540763 149701
rect 543641 149698 543707 149701
rect 540697 149696 543707 149698
rect 540697 149640 540702 149696
rect 540758 149640 543646 149696
rect 543702 149640 543707 149696
rect 540697 149638 543707 149640
rect 540697 149635 540763 149638
rect 543641 149635 543707 149638
rect 553350 149290 553410 150046
rect 561949 149290 562015 149293
rect 553350 149288 562015 149290
rect 553350 149232 561954 149288
rect 562010 149232 562015 149288
rect 553350 149230 562015 149232
rect 561949 149227 562015 149230
rect 48681 149154 48747 149157
rect 48998 149154 49004 149156
rect 48681 149152 49004 149154
rect 48681 149096 48686 149152
rect 48742 149096 49004 149152
rect 48681 149094 49004 149096
rect 48681 149091 48747 149094
rect 48998 149092 49004 149094
rect 49068 149092 49074 149156
rect 563646 149092 563652 149156
rect 563716 149154 563722 149156
rect 565169 149154 565235 149157
rect 563716 149152 565235 149154
rect 563716 149096 565174 149152
rect 565230 149096 565235 149152
rect 563716 149094 565235 149096
rect 563716 149092 563722 149094
rect 565169 149091 565235 149094
rect 56225 149018 56291 149021
rect 59721 149018 59787 149021
rect 56225 149016 59787 149018
rect 56225 148960 56230 149016
rect 56286 148960 59726 149016
rect 59782 148960 59787 149016
rect 56225 148958 59787 148960
rect 56225 148955 56291 148958
rect 59721 148955 59787 148958
rect 51022 148684 51028 148748
rect 51092 148746 51098 148748
rect 60222 148746 60228 148748
rect 51092 148686 60228 148746
rect 51092 148684 51098 148686
rect 60222 148684 60228 148686
rect 60292 148684 60298 148748
rect 540094 148548 540100 148612
rect 540164 148610 540170 148612
rect 558453 148610 558519 148613
rect 540164 148608 558519 148610
rect 540164 148552 558458 148608
rect 558514 148552 558519 148608
rect 540164 148550 558519 148552
rect 540164 148548 540170 148550
rect 558453 148547 558519 148550
rect 47710 147732 47716 147796
rect 47780 147794 47786 147796
rect 51717 147794 51783 147797
rect 47780 147792 51783 147794
rect 47780 147736 51722 147792
rect 51778 147736 51783 147792
rect 47780 147734 51783 147736
rect 47780 147732 47786 147734
rect 51717 147731 51783 147734
rect 540053 147794 540119 147797
rect 540053 147792 540346 147794
rect 540053 147736 540058 147792
rect 540114 147736 540346 147792
rect 540053 147734 540346 147736
rect 540053 147731 540119 147734
rect 51809 147658 51875 147661
rect 59629 147658 59695 147661
rect 51809 147656 59695 147658
rect 51809 147600 51814 147656
rect 51870 147600 59634 147656
rect 59690 147600 59695 147656
rect 51809 147598 59695 147600
rect 540286 147658 540346 147734
rect 541893 147658 541959 147661
rect 540286 147656 541959 147658
rect 540286 147600 541898 147656
rect 541954 147600 541959 147656
rect 540286 147598 541959 147600
rect 51809 147595 51875 147598
rect 59629 147595 59695 147598
rect 541893 147595 541959 147598
rect 51022 147460 51028 147524
rect 51092 147522 51098 147524
rect 52126 147522 52132 147524
rect 51092 147462 52132 147522
rect 51092 147460 51098 147462
rect 52126 147460 52132 147462
rect 52196 147460 52202 147524
rect 539358 147324 539364 147388
rect 539428 147386 539434 147388
rect 540145 147386 540211 147389
rect 539428 147384 540211 147386
rect 539428 147328 540150 147384
rect 540206 147328 540211 147384
rect 539428 147326 540211 147328
rect 539428 147324 539434 147326
rect 540145 147323 540211 147326
rect 540278 146916 540284 146980
rect 540348 146978 540354 146980
rect 552657 146978 552723 146981
rect 540348 146976 552723 146978
rect 540348 146920 552662 146976
rect 552718 146920 552723 146976
rect 540348 146918 552723 146920
rect 540348 146916 540354 146918
rect 552657 146915 552723 146918
rect 539358 146780 539364 146844
rect 539428 146842 539434 146844
rect 546953 146842 547019 146845
rect 539428 146840 547019 146842
rect 539428 146784 546958 146840
rect 547014 146784 547019 146840
rect 539428 146782 547019 146784
rect 539428 146780 539434 146782
rect 546953 146779 547019 146782
rect 52361 146570 52427 146573
rect 60038 146570 60044 146572
rect 52361 146568 60044 146570
rect 52361 146512 52366 146568
rect 52422 146512 60044 146568
rect 52361 146510 60044 146512
rect 52361 146507 52427 146510
rect 60038 146508 60044 146510
rect 60108 146508 60114 146572
rect 539358 146508 539364 146572
rect 539428 146570 539434 146572
rect 544469 146570 544535 146573
rect 539428 146568 544535 146570
rect 539428 146512 544474 146568
rect 544530 146512 544535 146568
rect 539428 146510 544535 146512
rect 539428 146508 539434 146510
rect 544469 146507 544535 146510
rect 543457 146434 543523 146437
rect 539948 146432 543523 146434
rect 539948 146376 543462 146432
rect 543518 146376 543523 146432
rect 539948 146374 543523 146376
rect 543457 146371 543523 146374
rect 544142 146236 544148 146300
rect 544212 146298 544218 146300
rect 544653 146298 544719 146301
rect 544212 146296 544719 146298
rect 544212 146240 544658 146296
rect 544714 146240 544719 146296
rect 544212 146238 544719 146240
rect 544212 146236 544218 146238
rect 544653 146235 544719 146238
rect 542854 146100 542860 146164
rect 542924 146162 542930 146164
rect 544694 146162 544700 146164
rect 542924 146102 544700 146162
rect 542924 146100 542930 146102
rect 544694 146100 544700 146102
rect 544764 146100 544770 146164
rect 57881 145754 57947 145757
rect 542537 145754 542603 145757
rect 57881 145752 60076 145754
rect 57881 145696 57886 145752
rect 57942 145696 60076 145752
rect 57881 145694 60076 145696
rect 539948 145752 542603 145754
rect 539948 145696 542542 145752
rect 542598 145696 542603 145752
rect 539948 145694 542603 145696
rect 57881 145691 57947 145694
rect 542537 145691 542603 145694
rect 539358 145420 539364 145484
rect 539428 145482 539434 145484
rect 540973 145482 541039 145485
rect 539428 145480 541039 145482
rect 539428 145424 540978 145480
rect 541034 145424 541039 145480
rect 539428 145422 541039 145424
rect 539428 145420 539434 145422
rect 540973 145419 541039 145422
rect 59077 144938 59143 144941
rect 59302 144938 59308 144940
rect 59077 144936 59308 144938
rect 59077 144880 59082 144936
rect 59138 144880 59308 144936
rect 59077 144878 59308 144880
rect 59077 144875 59143 144878
rect 59302 144876 59308 144878
rect 59372 144876 59378 144940
rect 540830 144740 540836 144804
rect 540900 144802 540906 144804
rect 544101 144802 544167 144805
rect 540900 144800 544167 144802
rect 540900 144744 544106 144800
rect 544162 144744 544167 144800
rect 540900 144742 544167 144744
rect 540900 144740 540906 144742
rect 544101 144739 544167 144742
rect 57605 143578 57671 143581
rect 58014 143578 58020 143580
rect 57605 143576 58020 143578
rect 57605 143520 57610 143576
rect 57666 143520 58020 143576
rect 57605 143518 58020 143520
rect 57605 143515 57671 143518
rect 58014 143516 58020 143518
rect 58084 143516 58090 143580
rect 58750 143516 58756 143580
rect 58820 143578 58826 143580
rect 58893 143578 58959 143581
rect 58820 143576 58959 143578
rect 58820 143520 58898 143576
rect 58954 143520 58959 143576
rect 58820 143518 58959 143520
rect 58820 143516 58826 143518
rect 58893 143515 58959 143518
rect 540053 143442 540119 143445
rect 539918 143440 540119 143442
rect 539918 143384 540058 143440
rect 540114 143384 540119 143440
rect 539918 143382 540119 143384
rect 57789 143034 57855 143037
rect 57789 143032 60076 143034
rect 57789 142976 57794 143032
rect 57850 142976 60076 143032
rect 539918 143004 539978 143382
rect 540053 143379 540119 143382
rect 57789 142974 60076 142976
rect 57789 142971 57855 142974
rect 52310 142354 52316 142356
rect 51950 142294 52316 142354
rect 51533 142082 51599 142085
rect 51950 142082 52010 142294
rect 52310 142292 52316 142294
rect 52380 142292 52386 142356
rect 543273 142354 543339 142357
rect 539948 142352 543339 142354
rect 539948 142296 543278 142352
rect 543334 142296 543339 142352
rect 539948 142294 543339 142296
rect 543273 142291 543339 142294
rect 52177 142218 52243 142221
rect 52177 142216 52378 142218
rect 52177 142160 52182 142216
rect 52238 142160 52378 142216
rect 52177 142158 52378 142160
rect 52177 142155 52243 142158
rect 52318 142084 52378 142158
rect 51533 142080 52010 142082
rect 51533 142024 51538 142080
rect 51594 142024 52010 142080
rect 51533 142022 52010 142024
rect 51533 142019 51599 142022
rect 52310 142020 52316 142084
rect 52380 142020 52386 142084
rect 59118 142020 59124 142084
rect 59188 142082 59194 142084
rect 59486 142082 59492 142084
rect 59188 142022 59492 142082
rect 59188 142020 59194 142022
rect 59486 142020 59492 142022
rect 59556 142020 59562 142084
rect 539358 141748 539364 141812
rect 539428 141810 539434 141812
rect 541525 141810 541591 141813
rect 539428 141808 541591 141810
rect 539428 141752 541530 141808
rect 541586 141752 541591 141808
rect 539428 141750 541591 141752
rect 539428 141748 539434 141750
rect 541525 141747 541591 141750
rect 56685 141674 56751 141677
rect 542905 141674 542971 141677
rect 56685 141672 60076 141674
rect 56685 141616 56690 141672
rect 56746 141616 60076 141672
rect 56685 141614 60076 141616
rect 539948 141672 542971 141674
rect 539948 141616 542910 141672
rect 542966 141616 542971 141672
rect 539948 141614 542971 141616
rect 56685 141611 56751 141614
rect 542905 141611 542971 141614
rect 543549 140994 543615 140997
rect 539948 140992 543615 140994
rect 539948 140936 543554 140992
rect 543610 140936 543615 140992
rect 539948 140934 543615 140936
rect 543549 140931 543615 140934
rect 56685 140314 56751 140317
rect 56685 140312 60076 140314
rect 56685 140256 56690 140312
rect 56746 140256 60076 140312
rect 56685 140254 60076 140256
rect 56685 140251 56751 140254
rect 57237 139634 57303 139637
rect 57237 139632 60076 139634
rect 57237 139576 57242 139632
rect 57298 139576 60076 139632
rect 57237 139574 60076 139576
rect 57237 139571 57303 139574
rect 544326 139572 544332 139636
rect 544396 139634 544402 139636
rect 545614 139634 545620 139636
rect 544396 139574 545620 139634
rect 544396 139572 544402 139574
rect 545614 139572 545620 139574
rect 545684 139572 545690 139636
rect 544510 139436 544516 139500
rect 544580 139498 544586 139500
rect 544653 139498 544719 139501
rect 544580 139496 544719 139498
rect 544580 139440 544658 139496
rect 544714 139440 544719 139496
rect 544580 139438 544719 139440
rect 544580 139436 544586 139438
rect 544653 139435 544719 139438
rect 545430 139436 545436 139500
rect 545500 139498 545506 139500
rect 546033 139498 546099 139501
rect 545500 139496 546099 139498
rect 545500 139440 546038 139496
rect 546094 139440 546099 139496
rect 545500 139438 546099 139440
rect 545500 139436 545506 139438
rect 546033 139435 546099 139438
rect 580533 139362 580599 139365
rect 583520 139362 584960 139452
rect 580533 139360 584960 139362
rect 580533 139304 580538 139360
rect 580594 139304 584960 139360
rect 580533 139302 584960 139304
rect 580533 139299 580599 139302
rect 59261 139226 59327 139229
rect 60590 139226 60596 139228
rect 59261 139224 60596 139226
rect 59261 139168 59266 139224
rect 59322 139168 60596 139224
rect 59261 139166 60596 139168
rect 59261 139163 59327 139166
rect 60590 139164 60596 139166
rect 60660 139164 60666 139228
rect 583520 139212 584960 139302
rect 547270 138620 547276 138684
rect 547340 138682 547346 138684
rect 552841 138682 552907 138685
rect 547340 138680 552907 138682
rect 547340 138624 552846 138680
rect 552902 138624 552907 138680
rect 547340 138622 552907 138624
rect 547340 138620 547346 138622
rect 552841 138619 552907 138622
rect 543549 138274 543615 138277
rect 539948 138272 543615 138274
rect 539948 138216 543554 138272
rect 543610 138216 543615 138272
rect 539948 138214 543615 138216
rect 543549 138211 543615 138214
rect 51022 138076 51028 138140
rect 51092 138138 51098 138140
rect 52126 138138 52132 138140
rect 51092 138078 52132 138138
rect 51092 138076 51098 138078
rect 52126 138076 52132 138078
rect 52196 138076 52202 138140
rect 544694 138076 544700 138140
rect 544764 138138 544770 138140
rect 545205 138138 545271 138141
rect 544764 138136 545271 138138
rect 544764 138080 545210 138136
rect 545266 138080 545271 138136
rect 544764 138078 545271 138080
rect 544764 138076 544770 138078
rect 545205 138075 545271 138078
rect 547270 138076 547276 138140
rect 547340 138138 547346 138140
rect 547413 138138 547479 138141
rect 547340 138136 547479 138138
rect 547340 138080 547418 138136
rect 547474 138080 547479 138136
rect 547340 138078 547479 138080
rect 547340 138076 547346 138078
rect 547413 138075 547479 138078
rect 544694 137940 544700 138004
rect 544764 138002 544770 138004
rect 549345 138002 549411 138005
rect 544764 138000 549411 138002
rect 544764 137944 549350 138000
rect 549406 137944 549411 138000
rect 544764 137942 549411 137944
rect 544764 137940 544770 137942
rect 549345 137939 549411 137942
rect 57605 137594 57671 137597
rect 57605 137592 60076 137594
rect 57605 137536 57610 137592
rect 57666 137536 60076 137592
rect 57605 137534 60076 137536
rect 57605 137531 57671 137534
rect 59077 137322 59143 137325
rect 59302 137322 59308 137324
rect 59077 137320 59308 137322
rect 59077 137264 59082 137320
rect 59138 137264 59308 137320
rect 59077 137262 59308 137264
rect 59077 137259 59143 137262
rect 59302 137260 59308 137262
rect 59372 137260 59378 137324
rect 559649 137322 559715 137325
rect 563646 137322 563652 137324
rect 559649 137320 563652 137322
rect 559649 137264 559654 137320
rect 559710 137264 563652 137320
rect 559649 137262 563652 137264
rect 559649 137259 559715 137262
rect 563646 137260 563652 137262
rect 563716 137260 563722 137324
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 58893 136642 58959 136645
rect 59118 136642 59124 136644
rect 58893 136640 59124 136642
rect 58893 136584 58898 136640
rect 58954 136584 59124 136640
rect 58893 136582 59124 136584
rect 58893 136579 58959 136582
rect 59118 136580 59124 136582
rect 59188 136580 59194 136644
rect 541617 136642 541683 136645
rect 544561 136644 544627 136645
rect 544326 136642 544332 136644
rect 541617 136640 544332 136642
rect 541617 136584 541622 136640
rect 541678 136584 544332 136640
rect 541617 136582 544332 136584
rect 541617 136579 541683 136582
rect 544326 136580 544332 136582
rect 544396 136580 544402 136644
rect 544510 136580 544516 136644
rect 544580 136642 544627 136644
rect 544580 136640 544672 136642
rect 544622 136584 544672 136640
rect 544580 136582 544672 136584
rect 544580 136580 544627 136582
rect 564014 136580 564020 136644
rect 564084 136642 564090 136644
rect 565813 136642 565879 136645
rect 564084 136640 565879 136642
rect 564084 136584 565818 136640
rect 565874 136584 565879 136640
rect 564084 136582 565879 136584
rect 564084 136580 564090 136582
rect 544561 136579 544627 136580
rect 565813 136579 565879 136582
rect 542445 136234 542511 136237
rect 539948 136232 542511 136234
rect 539948 136176 542450 136232
rect 542506 136176 542511 136232
rect 539948 136174 542511 136176
rect 542445 136171 542511 136174
rect 53741 135962 53807 135965
rect 58566 135962 58572 135964
rect 53741 135960 58572 135962
rect 53741 135904 53746 135960
rect 53802 135904 58572 135960
rect 53741 135902 58572 135904
rect 53741 135899 53807 135902
rect 58566 135900 58572 135902
rect 58636 135900 58642 135964
rect 542813 135554 542879 135557
rect 539948 135552 542879 135554
rect 41086 135220 41092 135284
rect 41156 135282 41162 135284
rect 60046 135282 60106 135524
rect 539948 135496 542818 135552
rect 542874 135496 542879 135552
rect 539948 135494 542879 135496
rect 542813 135491 542879 135494
rect 41156 135222 60106 135282
rect 41156 135220 41162 135222
rect 57605 134874 57671 134877
rect 57605 134872 60076 134874
rect 57605 134816 57610 134872
rect 57666 134816 60076 134872
rect 57605 134814 60076 134816
rect 57605 134811 57671 134814
rect 542445 134194 542511 134197
rect 539948 134192 542511 134194
rect 539948 134136 542450 134192
rect 542506 134136 542511 134192
rect 539948 134134 542511 134136
rect 542445 134131 542511 134134
rect 541065 133514 541131 133517
rect 539948 133512 541131 133514
rect 539948 133456 541070 133512
rect 541126 133456 541131 133512
rect 539948 133454 541131 133456
rect 541065 133451 541131 133454
rect 540881 133242 540947 133245
rect 541382 133242 541388 133244
rect 540881 133240 541388 133242
rect 540881 133184 540886 133240
rect 540942 133184 541388 133240
rect 540881 133182 541388 133184
rect 540881 133179 540947 133182
rect 541382 133180 541388 133182
rect 541452 133180 541458 133244
rect 541801 133106 541867 133109
rect 552657 133106 552723 133109
rect 541801 133104 552723 133106
rect 541801 133048 541806 133104
rect 541862 133048 552662 133104
rect 552718 133048 552723 133104
rect 541801 133046 552723 133048
rect 541801 133043 541867 133046
rect 552657 133043 552723 133046
rect 57605 132834 57671 132837
rect 57605 132832 60076 132834
rect 57605 132776 57610 132832
rect 57666 132776 60076 132832
rect 57605 132774 60076 132776
rect 57605 132771 57671 132774
rect 547270 132772 547276 132836
rect 547340 132834 547346 132836
rect 547638 132834 547644 132836
rect 547340 132774 547644 132834
rect 547340 132772 547346 132774
rect 547638 132772 547644 132774
rect 547708 132772 547714 132836
rect 57605 131474 57671 131477
rect 542445 131474 542511 131477
rect 57605 131472 60076 131474
rect 57605 131416 57610 131472
rect 57666 131416 60076 131472
rect 57605 131414 60076 131416
rect 539948 131472 542511 131474
rect 539948 131416 542450 131472
rect 542506 131416 542511 131472
rect 539948 131414 542511 131416
rect 57605 131411 57671 131414
rect 542445 131411 542511 131414
rect 541934 131276 541940 131340
rect 542004 131338 542010 131340
rect 544694 131338 544700 131340
rect 542004 131278 544700 131338
rect 542004 131276 542010 131278
rect 544694 131276 544700 131278
rect 544764 131276 544770 131340
rect 544561 131204 544627 131205
rect 544510 131202 544516 131204
rect 544470 131142 544516 131202
rect 544580 131200 544627 131204
rect 544622 131144 544627 131200
rect 544510 131140 544516 131142
rect 544580 131140 544627 131144
rect 544561 131139 544627 131140
rect 57605 130794 57671 130797
rect 542445 130794 542511 130797
rect 57605 130792 60076 130794
rect 57605 130736 57610 130792
rect 57666 130736 60076 130792
rect 57605 130734 60076 130736
rect 539948 130792 542511 130794
rect 539948 130736 542450 130792
rect 542506 130736 542511 130792
rect 539948 130734 542511 130736
rect 57605 130731 57671 130734
rect 542445 130731 542511 130734
rect 541566 130460 541572 130524
rect 541636 130522 541642 130524
rect 547873 130522 547939 130525
rect 541636 130520 547939 130522
rect 541636 130464 547878 130520
rect 547934 130464 547939 130520
rect 541636 130462 547939 130464
rect 541636 130460 541642 130462
rect 547873 130459 547939 130462
rect 542118 130324 542124 130388
rect 542188 130386 542194 130388
rect 548006 130386 548012 130388
rect 542188 130326 548012 130386
rect 542188 130324 542194 130326
rect 548006 130324 548012 130326
rect 548076 130324 548082 130388
rect 540646 129644 540652 129708
rect 540716 129706 540722 129708
rect 540973 129706 541039 129709
rect 540716 129704 541039 129706
rect 540716 129648 540978 129704
rect 541034 129648 541039 129704
rect 540716 129646 541039 129648
rect 540716 129644 540722 129646
rect 540973 129643 541039 129646
rect 542905 129570 542971 129573
rect 548374 129570 548380 129572
rect 542905 129568 548380 129570
rect 542905 129512 542910 129568
rect 542966 129512 548380 129568
rect 542905 129510 548380 129512
rect 542905 129507 542971 129510
rect 548374 129508 548380 129510
rect 548444 129508 548450 129572
rect 57605 129434 57671 129437
rect 542445 129434 542511 129437
rect 57605 129432 60076 129434
rect 57605 129376 57610 129432
rect 57666 129376 60076 129432
rect 57605 129374 60076 129376
rect 539948 129432 542511 129434
rect 539948 129376 542450 129432
rect 542506 129376 542511 129432
rect 539948 129374 542511 129376
rect 57605 129371 57671 129374
rect 542445 129371 542511 129374
rect 543038 128420 543044 128484
rect 543108 128482 543114 128484
rect 545205 128482 545271 128485
rect 543108 128480 545271 128482
rect 543108 128424 545210 128480
rect 545266 128424 545271 128480
rect 543108 128422 545271 128424
rect 543108 128420 543114 128422
rect 545205 128419 545271 128422
rect 57605 128074 57671 128077
rect 543549 128074 543615 128077
rect 57605 128072 60076 128074
rect 57605 128016 57610 128072
rect 57666 128016 60076 128072
rect 57605 128014 60076 128016
rect 539948 128072 543615 128074
rect 539948 128016 543554 128072
rect 543610 128016 543615 128072
rect 539948 128014 543615 128016
rect 57605 128011 57671 128014
rect 543549 128011 543615 128014
rect 541801 127666 541867 127669
rect 544142 127666 544148 127668
rect 541801 127664 544148 127666
rect 541801 127608 541806 127664
rect 541862 127608 544148 127664
rect 541801 127606 544148 127608
rect 541801 127603 541867 127606
rect 544142 127604 544148 127606
rect 544212 127604 544218 127668
rect 544326 127604 544332 127668
rect 544396 127666 544402 127668
rect 545430 127666 545436 127668
rect 544396 127606 545436 127666
rect 544396 127604 544402 127606
rect 545430 127604 545436 127606
rect 545500 127604 545506 127668
rect 545113 127122 545179 127125
rect 545614 127122 545620 127124
rect 545113 127120 545620 127122
rect 545113 127064 545118 127120
rect 545174 127064 545620 127120
rect 545113 127062 545620 127064
rect 545113 127059 545179 127062
rect 545614 127060 545620 127062
rect 545684 127060 545690 127124
rect 545614 126924 545620 126988
rect 545684 126986 545690 126988
rect 546033 126986 546099 126989
rect 545684 126984 546099 126986
rect 545684 126928 546038 126984
rect 546094 126928 546099 126984
rect 545684 126926 546099 126928
rect 545684 126924 545690 126926
rect 546033 126923 546099 126926
rect 547413 126986 547479 126989
rect 547638 126986 547644 126988
rect 547413 126984 547644 126986
rect 547413 126928 547418 126984
rect 547474 126928 547644 126984
rect 547413 126926 547644 126928
rect 547413 126923 547479 126926
rect 547638 126924 547644 126926
rect 547708 126924 547714 126988
rect 545798 126788 545804 126852
rect 545868 126850 545874 126852
rect 547270 126850 547276 126852
rect 545868 126790 547276 126850
rect 545868 126788 545874 126790
rect 547270 126788 547276 126790
rect 547340 126788 547346 126852
rect 57605 126714 57671 126717
rect 57605 126712 60076 126714
rect 57605 126656 57610 126712
rect 57666 126656 60076 126712
rect 57605 126654 60076 126656
rect 57605 126651 57671 126654
rect 540830 126244 540836 126308
rect 540900 126306 540906 126308
rect 550081 126306 550147 126309
rect 540900 126304 550147 126306
rect 540900 126248 550086 126304
rect 550142 126248 550147 126304
rect 540900 126246 550147 126248
rect 540900 126244 540906 126246
rect 550081 126243 550147 126246
rect 583520 125884 584960 126124
rect 59261 125490 59327 125493
rect 59486 125490 59492 125492
rect 59261 125488 59492 125490
rect 59261 125432 59266 125488
rect 59322 125432 59492 125488
rect 59261 125430 59492 125432
rect 59261 125427 59327 125430
rect 59486 125428 59492 125430
rect 59556 125428 59562 125492
rect 56685 125354 56751 125357
rect 542445 125354 542511 125357
rect 56685 125352 60076 125354
rect 56685 125296 56690 125352
rect 56746 125296 60076 125352
rect 56685 125294 60076 125296
rect 539948 125352 542511 125354
rect 539948 125296 542450 125352
rect 542506 125296 542511 125352
rect 539948 125294 542511 125296
rect 56685 125291 56751 125294
rect 542445 125291 542511 125294
rect 53741 124810 53807 124813
rect 58566 124810 58572 124812
rect 53741 124808 58572 124810
rect 53741 124752 53746 124808
rect 53802 124752 58572 124808
rect 53741 124750 58572 124752
rect 53741 124747 53807 124750
rect 58566 124748 58572 124750
rect 58636 124748 58642 124812
rect 543549 124674 543615 124677
rect 539948 124672 543615 124674
rect 539948 124616 543554 124672
rect 543610 124616 543615 124672
rect 539948 124614 543615 124616
rect 543549 124611 543615 124614
rect 58934 124266 58940 124268
rect 58206 124206 58940 124266
rect 50337 124130 50403 124133
rect 51022 124130 51028 124132
rect 50337 124128 51028 124130
rect 50337 124072 50342 124128
rect 50398 124072 51028 124128
rect 50337 124070 51028 124072
rect 50337 124067 50403 124070
rect 51022 124068 51028 124070
rect 51092 124068 51098 124132
rect 51533 124130 51599 124133
rect 52126 124130 52132 124132
rect 51533 124128 52132 124130
rect 51533 124072 51538 124128
rect 51594 124072 52132 124128
rect 51533 124070 52132 124072
rect 51533 124067 51599 124070
rect 52126 124068 52132 124070
rect 52196 124068 52202 124132
rect 58065 124130 58131 124133
rect 58206 124130 58266 124206
rect 58934 124204 58940 124206
rect 59004 124204 59010 124268
rect 544561 124132 544627 124133
rect 58065 124128 58266 124130
rect 58065 124072 58070 124128
rect 58126 124072 58266 124128
rect 58065 124070 58266 124072
rect 58065 124067 58131 124070
rect 544510 124068 544516 124132
rect 544580 124130 544627 124132
rect 544580 124128 544672 124130
rect 544622 124072 544672 124128
rect 544580 124070 544672 124072
rect 544580 124068 544627 124070
rect 544561 124067 544627 124068
rect 544326 123932 544332 123996
rect 544396 123994 544402 123996
rect 545113 123994 545179 123997
rect 544396 123992 545179 123994
rect 544396 123936 545118 123992
rect 545174 123936 545179 123992
rect 544396 123934 545179 123936
rect 544396 123932 544402 123934
rect 545113 123931 545179 123934
rect -960 123572 480 123812
rect 46422 123524 46428 123588
rect 46492 123586 46498 123588
rect 58750 123586 58756 123588
rect 46492 123526 58756 123586
rect 46492 123524 46498 123526
rect 58750 123524 58756 123526
rect 58820 123524 58826 123588
rect 46238 123388 46244 123452
rect 46308 123450 46314 123452
rect 59854 123450 59860 123452
rect 46308 123390 59860 123450
rect 46308 123388 46314 123390
rect 59854 123388 59860 123390
rect 59924 123388 59930 123452
rect 57605 123314 57671 123317
rect 57605 123312 60076 123314
rect 57605 123256 57610 123312
rect 57666 123256 60076 123312
rect 57605 123254 60076 123256
rect 57605 123251 57671 123254
rect 54661 122090 54727 122093
rect 59670 122090 59676 122092
rect 54661 122088 59676 122090
rect 54661 122032 54666 122088
rect 54722 122032 59676 122088
rect 54661 122030 59676 122032
rect 54661 122027 54727 122030
rect 59670 122028 59676 122030
rect 59740 122028 59746 122092
rect 543641 121954 543707 121957
rect 539948 121952 543707 121954
rect 539948 121896 543646 121952
rect 543702 121896 543707 121952
rect 539948 121894 543707 121896
rect 543641 121891 543707 121894
rect 57421 120594 57487 120597
rect 543549 120594 543615 120597
rect 57421 120592 60076 120594
rect 57421 120536 57426 120592
rect 57482 120536 60076 120592
rect 57421 120534 60076 120536
rect 539948 120592 543615 120594
rect 539948 120536 543554 120592
rect 543610 120536 543615 120592
rect 539948 120534 543615 120536
rect 57421 120531 57487 120534
rect 543549 120531 543615 120534
rect 59261 120188 59327 120189
rect 59261 120186 59308 120188
rect 59216 120184 59308 120186
rect 59216 120128 59266 120184
rect 59216 120126 59308 120128
rect 59261 120124 59308 120126
rect 59372 120124 59378 120188
rect 59261 120123 59327 120124
rect 56961 119914 57027 119917
rect 56961 119912 60076 119914
rect 56961 119856 56966 119912
rect 57022 119856 60076 119912
rect 56961 119854 60076 119856
rect 56961 119851 57027 119854
rect 57421 119234 57487 119237
rect 57421 119232 60076 119234
rect 57421 119176 57426 119232
rect 57482 119176 60076 119232
rect 57421 119174 60076 119176
rect 57421 119171 57487 119174
rect 56961 118010 57027 118013
rect 58014 118010 58020 118012
rect 56961 118008 58020 118010
rect 56961 117952 56966 118008
rect 57022 117952 58020 118008
rect 56961 117950 58020 117952
rect 56961 117947 57027 117950
rect 58014 117948 58020 117950
rect 58084 117948 58090 118012
rect 543549 118010 543615 118013
rect 544142 118010 544148 118012
rect 543549 118008 544148 118010
rect 543549 117952 543554 118008
rect 543610 117952 544148 118008
rect 543549 117950 544148 117952
rect 543549 117947 543615 117950
rect 544142 117948 544148 117950
rect 544212 117948 544218 118012
rect 544561 117332 544627 117333
rect 544510 117330 544516 117332
rect 544470 117270 544516 117330
rect 544580 117328 544627 117332
rect 544622 117272 544627 117328
rect 544510 117268 544516 117270
rect 544580 117268 544627 117272
rect 544561 117267 544627 117268
rect 57053 117194 57119 117197
rect 57053 117192 60076 117194
rect 57053 117136 57058 117192
rect 57114 117136 60076 117192
rect 57053 117134 60076 117136
rect 57053 117131 57119 117134
rect 542445 116514 542511 116517
rect 539948 116512 542511 116514
rect 539948 116456 542450 116512
rect 542506 116456 542511 116512
rect 539948 116454 542511 116456
rect 542445 116451 542511 116454
rect 540605 115970 540671 115973
rect 541801 115972 541867 115973
rect 541198 115970 541204 115972
rect 540605 115968 541204 115970
rect 540605 115912 540610 115968
rect 540666 115912 541204 115968
rect 540605 115910 541204 115912
rect 540605 115907 540671 115910
rect 541198 115908 541204 115910
rect 541268 115908 541274 115972
rect 541750 115970 541756 115972
rect 541710 115910 541756 115970
rect 541820 115968 541867 115972
rect 541862 115912 541867 115968
rect 541750 115908 541756 115910
rect 541820 115908 541867 115912
rect 541801 115907 541867 115908
rect 58249 115834 58315 115837
rect 541709 115834 541775 115837
rect 58249 115832 60076 115834
rect 58249 115776 58254 115832
rect 58310 115776 60076 115832
rect 58249 115774 60076 115776
rect 539948 115832 541775 115834
rect 539948 115776 541714 115832
rect 541770 115776 541775 115832
rect 539948 115774 541775 115776
rect 58249 115771 58315 115774
rect 541709 115771 541775 115774
rect 57421 115154 57487 115157
rect 57421 115152 60076 115154
rect 57421 115096 57426 115152
rect 57482 115096 60076 115152
rect 57421 115094 60076 115096
rect 57421 115091 57487 115094
rect 57421 114474 57487 114477
rect 544285 114474 544351 114477
rect 544510 114474 544516 114476
rect 57421 114472 60076 114474
rect 57421 114416 57426 114472
rect 57482 114416 60076 114472
rect 544285 114472 544516 114474
rect 57421 114414 60076 114416
rect 57421 114411 57487 114414
rect 539918 114338 539978 114444
rect 544285 114416 544290 114472
rect 544346 114416 544516 114472
rect 544285 114414 544516 114416
rect 544285 114411 544351 114414
rect 544510 114412 544516 114414
rect 544580 114412 544586 114476
rect 547454 114338 547460 114340
rect 539918 114278 547460 114338
rect 547454 114276 547460 114278
rect 547524 114276 547530 114340
rect 542445 113794 542511 113797
rect 539948 113792 542511 113794
rect 539948 113736 542450 113792
rect 542506 113736 542511 113792
rect 539948 113734 542511 113736
rect 542445 113731 542511 113734
rect 549478 113188 549484 113252
rect 549548 113250 549554 113252
rect 549713 113250 549779 113253
rect 549548 113248 549779 113250
rect 549548 113192 549718 113248
rect 549774 113192 549779 113248
rect 549548 113190 549779 113192
rect 549548 113188 549554 113190
rect 549713 113187 549779 113190
rect 56869 113114 56935 113117
rect 542486 113114 542492 113116
rect 56869 113112 60076 113114
rect 56869 113056 56874 113112
rect 56930 113056 60076 113112
rect 56869 113054 60076 113056
rect 539948 113054 542492 113114
rect 56869 113051 56935 113054
rect 542486 113052 542492 113054
rect 542556 113052 542562 113116
rect 580533 112842 580599 112845
rect 583520 112842 584960 112932
rect 580533 112840 584960 112842
rect 580533 112784 580538 112840
rect 580594 112784 584960 112840
rect 580533 112782 584960 112784
rect 580533 112779 580599 112782
rect 583520 112692 584960 112782
rect 58893 111890 58959 111893
rect 59302 111890 59308 111892
rect 58893 111888 59308 111890
rect 58893 111832 58898 111888
rect 58954 111832 59308 111888
rect 58893 111830 59308 111832
rect 58893 111827 58959 111830
rect 59302 111828 59308 111830
rect 59372 111828 59378 111892
rect 542854 110876 542860 110940
rect 542924 110938 542930 110940
rect 556797 110938 556863 110941
rect 542924 110936 556863 110938
rect 542924 110880 556802 110936
rect 556858 110880 556863 110936
rect 542924 110878 556863 110880
rect 542924 110876 542930 110878
rect 556797 110875 556863 110878
rect -960 110516 480 110756
rect 541934 110604 541940 110668
rect 542004 110666 542010 110668
rect 547454 110666 547460 110668
rect 542004 110606 547460 110666
rect 542004 110604 542010 110606
rect 547454 110604 547460 110606
rect 547524 110604 547530 110668
rect 543549 110530 543615 110533
rect 544142 110530 544148 110532
rect 543549 110528 544148 110530
rect 543549 110472 543554 110528
rect 543610 110472 544148 110528
rect 543549 110470 544148 110472
rect 543549 110467 543615 110470
rect 544142 110468 544148 110470
rect 544212 110468 544218 110532
rect 57513 110394 57579 110397
rect 542537 110394 542603 110397
rect 57513 110392 60076 110394
rect 57513 110336 57518 110392
rect 57574 110336 60076 110392
rect 57513 110334 60076 110336
rect 539948 110392 542603 110394
rect 539948 110336 542542 110392
rect 542598 110336 542603 110392
rect 539948 110334 542603 110336
rect 57513 110331 57579 110334
rect 542537 110331 542603 110334
rect 540646 110196 540652 110260
rect 540716 110258 540722 110260
rect 541198 110258 541204 110260
rect 540716 110198 541204 110258
rect 540716 110196 540722 110198
rect 541198 110196 541204 110198
rect 541268 110196 541274 110260
rect 542445 109714 542511 109717
rect 539948 109712 542511 109714
rect 539948 109656 542450 109712
rect 542506 109656 542511 109712
rect 539948 109654 542511 109656
rect 542445 109651 542511 109654
rect 57513 108354 57579 108357
rect 57513 108352 60076 108354
rect 57513 108296 57518 108352
rect 57574 108296 60076 108352
rect 57513 108294 60076 108296
rect 57513 108291 57579 108294
rect 56593 107674 56659 107677
rect 542629 107674 542695 107677
rect 56593 107672 60076 107674
rect 56593 107616 56598 107672
rect 56654 107616 60076 107672
rect 56593 107614 60076 107616
rect 539948 107672 542695 107674
rect 539948 107616 542634 107672
rect 542690 107616 542695 107672
rect 539948 107614 542695 107616
rect 56593 107611 56659 107614
rect 542629 107611 542695 107614
rect 541750 107476 541756 107540
rect 541820 107538 541826 107540
rect 542486 107538 542492 107540
rect 541820 107478 542492 107538
rect 541820 107476 541826 107478
rect 542486 107476 542492 107478
rect 542556 107476 542562 107540
rect 543181 106314 543247 106317
rect 539948 106312 543247 106314
rect 539948 106256 543186 106312
rect 543242 106256 543247 106312
rect 539948 106254 543247 106256
rect 543181 106251 543247 106254
rect 541566 105436 541572 105500
rect 541636 105498 541642 105500
rect 574093 105498 574159 105501
rect 541636 105496 574159 105498
rect 541636 105440 574098 105496
rect 574154 105440 574159 105496
rect 541636 105438 574159 105440
rect 541636 105436 541642 105438
rect 574093 105435 574159 105438
rect 56869 104274 56935 104277
rect 543406 104274 543412 104276
rect 56869 104272 60076 104274
rect 56869 104216 56874 104272
rect 56930 104216 60076 104272
rect 56869 104214 60076 104216
rect 539948 104214 543412 104274
rect 56869 104211 56935 104214
rect 543406 104212 543412 104214
rect 543476 104212 543482 104276
rect 57513 103594 57579 103597
rect 57513 103592 60076 103594
rect 57513 103536 57518 103592
rect 57574 103536 60076 103592
rect 57513 103534 60076 103536
rect 57513 103531 57579 103534
rect 57513 102914 57579 102917
rect 57513 102912 60076 102914
rect 57513 102856 57518 102912
rect 57574 102856 60076 102912
rect 57513 102854 60076 102856
rect 57513 102851 57579 102854
rect 541382 102308 541388 102372
rect 541452 102370 541458 102372
rect 543038 102370 543044 102372
rect 541452 102310 543044 102370
rect 541452 102308 541458 102310
rect 543038 102308 543044 102310
rect 543108 102308 543114 102372
rect 57881 102234 57947 102237
rect 541525 102234 541591 102237
rect 542118 102234 542124 102236
rect 57881 102232 60076 102234
rect 57881 102176 57886 102232
rect 57942 102176 60076 102232
rect 57881 102174 60076 102176
rect 541525 102232 542124 102234
rect 541525 102176 541530 102232
rect 541586 102176 542124 102232
rect 541525 102174 542124 102176
rect 57881 102171 57947 102174
rect 541525 102171 541591 102174
rect 542118 102172 542124 102174
rect 542188 102172 542194 102236
rect 57513 101554 57579 101557
rect 541157 101554 541223 101557
rect 57513 101552 60076 101554
rect 57513 101496 57518 101552
rect 57574 101496 60076 101552
rect 57513 101494 60076 101496
rect 539948 101552 541223 101554
rect 539948 101496 541162 101552
rect 541218 101496 541223 101552
rect 539948 101494 541223 101496
rect 57513 101491 57579 101494
rect 541157 101491 541223 101494
rect 40493 100058 40559 100061
rect 59302 100058 59308 100060
rect 40493 100056 59308 100058
rect 40493 100000 40498 100056
rect 40554 100000 59308 100056
rect 40493 99998 59308 100000
rect 40493 99995 40559 99998
rect 59302 99996 59308 99998
rect 59372 99996 59378 100060
rect 57513 99514 57579 99517
rect 540789 99514 540855 99517
rect 541198 99514 541204 99516
rect 57513 99512 60076 99514
rect 57513 99456 57518 99512
rect 57574 99456 60076 99512
rect 57513 99454 60076 99456
rect 540789 99512 541204 99514
rect 540789 99456 540794 99512
rect 540850 99456 541204 99512
rect 540789 99454 541204 99456
rect 57513 99451 57579 99454
rect 540789 99451 540855 99454
rect 541198 99452 541204 99454
rect 541268 99452 541274 99516
rect 564014 99452 564020 99516
rect 564084 99514 564090 99516
rect 564617 99514 564683 99517
rect 564084 99512 564683 99514
rect 564084 99456 564622 99512
rect 564678 99456 564683 99512
rect 564084 99454 564683 99456
rect 564084 99452 564090 99454
rect 564617 99451 564683 99454
rect 580441 99514 580507 99517
rect 583520 99514 584960 99604
rect 580441 99512 584960 99514
rect 580441 99456 580446 99512
rect 580502 99456 584960 99512
rect 580441 99454 584960 99456
rect 580441 99451 580507 99454
rect 583520 99364 584960 99454
rect 55857 98154 55923 98157
rect 55857 98152 60076 98154
rect 55857 98096 55862 98152
rect 55918 98096 60076 98152
rect 55857 98094 60076 98096
rect 55857 98091 55923 98094
rect -960 97610 480 97700
rect 2865 97610 2931 97613
rect -960 97608 2931 97610
rect -960 97552 2870 97608
rect 2926 97552 2931 97608
rect -960 97550 2931 97552
rect -960 97460 480 97550
rect 2865 97547 2931 97550
rect 543549 97474 543615 97477
rect 539948 97472 543615 97474
rect 539948 97416 543554 97472
rect 543610 97416 543615 97472
rect 539948 97414 543615 97416
rect 543549 97411 543615 97414
rect 59077 96794 59143 96797
rect 59077 96792 60076 96794
rect 59077 96736 59082 96792
rect 59138 96736 60076 96792
rect 59077 96734 60076 96736
rect 59077 96731 59143 96734
rect 543549 96114 543615 96117
rect 539948 96112 543615 96114
rect 539948 96056 543554 96112
rect 543610 96056 543615 96112
rect 539948 96054 543615 96056
rect 543549 96051 543615 96054
rect 543641 95434 543707 95437
rect 539948 95432 543707 95434
rect 539948 95376 543646 95432
rect 543702 95376 543707 95432
rect 539948 95374 543707 95376
rect 543641 95371 543707 95374
rect 540094 95100 540100 95164
rect 540164 95162 540170 95164
rect 541065 95162 541131 95165
rect 540164 95160 541131 95162
rect 540164 95104 541070 95160
rect 541126 95104 541131 95160
rect 540164 95102 541131 95104
rect 540164 95100 540170 95102
rect 541065 95099 541131 95102
rect 57513 94074 57579 94077
rect 543549 94074 543615 94077
rect 57513 94072 60076 94074
rect 57513 94016 57518 94072
rect 57574 94016 60076 94072
rect 57513 94014 60076 94016
rect 539948 94072 543615 94074
rect 539948 94016 543554 94072
rect 543610 94016 543615 94072
rect 539948 94014 543615 94016
rect 57513 94011 57579 94014
rect 543549 94011 543615 94014
rect 57513 92714 57579 92717
rect 543549 92714 543615 92717
rect 57513 92712 60076 92714
rect 57513 92656 57518 92712
rect 57574 92656 60076 92712
rect 57513 92654 60076 92656
rect 539948 92712 543615 92714
rect 539948 92656 543554 92712
rect 543610 92656 543615 92712
rect 539948 92654 543615 92656
rect 57513 92651 57579 92654
rect 543549 92651 543615 92654
rect 543549 92034 543615 92037
rect 539948 92032 543615 92034
rect 539948 91976 543554 92032
rect 543610 91976 543615 92032
rect 539948 91974 543615 91976
rect 543549 91971 543615 91974
rect 542629 91354 542695 91357
rect 539948 91352 542695 91354
rect 539948 91296 542634 91352
rect 542690 91296 542695 91352
rect 539948 91294 542695 91296
rect 542629 91291 542695 91294
rect 57145 90674 57211 90677
rect 57145 90672 60076 90674
rect 57145 90616 57150 90672
rect 57206 90616 60076 90672
rect 57145 90614 60076 90616
rect 57145 90611 57211 90614
rect 57605 89314 57671 89317
rect 57605 89312 60076 89314
rect 57605 89256 57610 89312
rect 57666 89256 60076 89312
rect 57605 89254 60076 89256
rect 57605 89251 57671 89254
rect 554221 89178 554287 89181
rect 547830 89176 554287 89178
rect 547830 89120 554226 89176
rect 554282 89120 554287 89176
rect 547830 89118 554287 89120
rect 543222 88980 543228 89044
rect 543292 89042 543298 89044
rect 547830 89042 547890 89118
rect 554221 89115 554287 89118
rect 543292 88982 547890 89042
rect 553485 89042 553551 89045
rect 553894 89042 553900 89044
rect 553485 89040 553900 89042
rect 553485 88984 553490 89040
rect 553546 88984 553900 89040
rect 553485 88982 553900 88984
rect 543292 88980 543298 88982
rect 553485 88979 553551 88982
rect 553894 88980 553900 88982
rect 553964 88980 553970 89044
rect 542721 88634 542787 88637
rect 539948 88632 542787 88634
rect 539948 88576 542726 88632
rect 542782 88576 542787 88632
rect 539948 88574 542787 88576
rect 542721 88571 542787 88574
rect 542302 87954 542308 87956
rect 539948 87894 542308 87954
rect 542302 87892 542308 87894
rect 542372 87892 542378 87956
rect 57605 86594 57671 86597
rect 57605 86592 60076 86594
rect 57605 86536 57610 86592
rect 57666 86536 60076 86592
rect 57605 86534 60076 86536
rect 57605 86531 57671 86534
rect 543038 86124 543044 86188
rect 543108 86186 543114 86188
rect 559649 86186 559715 86189
rect 543108 86184 559715 86186
rect 543108 86128 559654 86184
rect 559710 86128 559715 86184
rect 543108 86126 559715 86128
rect 543108 86124 543114 86126
rect 559649 86123 559715 86126
rect 583520 86036 584960 86276
rect 547781 85642 547847 85645
rect 548374 85642 548380 85644
rect 547781 85640 548380 85642
rect 547781 85584 547786 85640
rect 547842 85584 548380 85640
rect 547781 85582 548380 85584
rect 547781 85579 547847 85582
rect 548374 85580 548380 85582
rect 548444 85580 548450 85644
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect 539918 84690 539978 85204
rect 548190 84690 548196 84692
rect 539918 84630 548196 84690
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 548190 84628 548196 84630
rect 548260 84628 548266 84692
rect 542629 84554 542695 84557
rect 539948 84552 542695 84554
rect 539948 84496 542634 84552
rect 542690 84496 542695 84552
rect 539948 84494 542695 84496
rect 542629 84491 542695 84494
rect 539918 83330 539978 83844
rect 549846 83330 549852 83332
rect 539918 83270 549852 83330
rect 549846 83268 549852 83270
rect 549916 83268 549922 83332
rect 541198 82860 541204 82924
rect 541268 82922 541274 82924
rect 541525 82922 541591 82925
rect 541268 82920 541591 82922
rect 541268 82864 541530 82920
rect 541586 82864 541591 82920
rect 541268 82862 541591 82864
rect 541268 82860 541274 82862
rect 541525 82859 541591 82862
rect 57605 82514 57671 82517
rect 543549 82514 543615 82517
rect 57605 82512 60076 82514
rect 57605 82456 57610 82512
rect 57666 82456 60076 82512
rect 57605 82454 60076 82456
rect 539948 82512 543615 82514
rect 539948 82456 543554 82512
rect 543610 82456 543615 82512
rect 539948 82454 543615 82456
rect 57605 82451 57671 82454
rect 543549 82451 543615 82454
rect 57513 81834 57579 81837
rect 57513 81832 60076 81834
rect 57513 81776 57518 81832
rect 57574 81776 60076 81832
rect 57513 81774 60076 81776
rect 57513 81771 57579 81774
rect 549846 81500 549852 81564
rect 549916 81562 549922 81564
rect 552013 81562 552079 81565
rect 549916 81560 552079 81562
rect 549916 81504 552018 81560
rect 552074 81504 552079 81560
rect 549916 81502 552079 81504
rect 549916 81500 549922 81502
rect 552013 81499 552079 81502
rect 57881 81154 57947 81157
rect 57881 81152 60076 81154
rect 57881 81096 57886 81152
rect 57942 81096 60076 81152
rect 57881 81094 60076 81096
rect 57881 81091 57947 81094
rect 543917 78434 543983 78437
rect 539948 78432 543983 78434
rect 539948 78376 543922 78432
rect 543978 78376 543983 78432
rect 539948 78374 543983 78376
rect 543917 78371 543983 78374
rect 543549 77754 543615 77757
rect 539948 77752 543615 77754
rect 539948 77696 543554 77752
rect 543610 77696 543615 77752
rect 539948 77694 543615 77696
rect 543549 77691 543615 77694
rect 55949 77074 56015 77077
rect 55949 77072 60076 77074
rect 55949 77016 55954 77072
rect 56010 77016 60076 77072
rect 55949 77014 60076 77016
rect 55949 77011 56015 77014
rect 543549 76394 543615 76397
rect 539948 76392 543615 76394
rect 539948 76336 543554 76392
rect 543610 76336 543615 76392
rect 539948 76334 543615 76336
rect 543549 76331 543615 76334
rect 57605 75714 57671 75717
rect 542629 75714 542695 75717
rect 57605 75712 60076 75714
rect 57605 75656 57610 75712
rect 57666 75656 60076 75712
rect 57605 75654 60076 75656
rect 539948 75712 542695 75714
rect 539948 75656 542634 75712
rect 542690 75656 542695 75712
rect 539948 75654 542695 75656
rect 57605 75651 57671 75654
rect 542629 75651 542695 75654
rect 57278 74972 57284 75036
rect 57348 75034 57354 75036
rect 543549 75034 543615 75037
rect 57348 74974 60076 75034
rect 539948 75032 543615 75034
rect 539948 74976 543554 75032
rect 543610 74976 543615 75032
rect 539948 74974 543615 74976
rect 57348 74972 57354 74974
rect 543549 74971 543615 74974
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 539918 72314 539978 72964
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect 549662 72314 549668 72316
rect 539918 72254 549668 72314
rect 549662 72252 549668 72254
rect 549732 72252 549738 72316
rect -960 71484 480 71724
rect 543549 71634 543615 71637
rect 539948 71632 543615 71634
rect 539948 71576 543554 71632
rect 543610 71576 543615 71632
rect 539948 71574 543615 71576
rect 543549 71571 543615 71574
rect 541014 70954 541020 70956
rect 539948 70894 541020 70954
rect 541014 70892 541020 70894
rect 541084 70892 541090 70956
rect 56133 70274 56199 70277
rect 543549 70274 543615 70277
rect 56133 70272 60076 70274
rect 56133 70216 56138 70272
rect 56194 70216 60076 70272
rect 56133 70214 60076 70216
rect 539948 70272 543615 70274
rect 539948 70216 543554 70272
rect 543610 70216 543615 70272
rect 539948 70214 543615 70216
rect 56133 70211 56199 70214
rect 543549 70211 543615 70214
rect 57881 68914 57947 68917
rect 543958 68914 543964 68916
rect 57881 68912 60076 68914
rect 57881 68856 57886 68912
rect 57942 68856 60076 68912
rect 57881 68854 60076 68856
rect 539948 68854 543964 68914
rect 57881 68851 57947 68854
rect 543958 68852 543964 68854
rect 544028 68852 544034 68916
rect 57145 68234 57211 68237
rect 57145 68232 60076 68234
rect 57145 68176 57150 68232
rect 57206 68176 60076 68232
rect 57145 68174 60076 68176
rect 57145 68171 57211 68174
rect 57881 67554 57947 67557
rect 57881 67552 60076 67554
rect 57881 67496 57886 67552
rect 57942 67496 60076 67552
rect 57881 67494 60076 67496
rect 57881 67491 57947 67494
rect 543549 66194 543615 66197
rect 539948 66192 543615 66194
rect 539948 66136 543554 66192
rect 543610 66136 543615 66192
rect 539948 66134 543615 66136
rect 543549 66131 543615 66134
rect 542813 65514 542879 65517
rect 539948 65512 542879 65514
rect 539948 65456 542818 65512
rect 542874 65456 542879 65512
rect 539948 65454 542879 65456
rect 542813 65451 542879 65454
rect 57830 64772 57836 64836
rect 57900 64834 57906 64836
rect 57900 64774 60076 64834
rect 57900 64772 57906 64774
rect 57881 64154 57947 64157
rect 543549 64154 543615 64157
rect 57881 64152 60076 64154
rect 57881 64096 57886 64152
rect 57942 64096 60076 64152
rect 57881 64094 60076 64096
rect 539948 64152 543615 64154
rect 539948 64096 543554 64152
rect 543610 64096 543615 64152
rect 539948 64094 543615 64096
rect 57881 64091 57947 64094
rect 543549 64091 543615 64094
rect 57881 63474 57947 63477
rect 57881 63472 60076 63474
rect 57881 63416 57886 63472
rect 57942 63416 60076 63472
rect 57881 63414 60076 63416
rect 57881 63411 57947 63414
rect 57881 62114 57947 62117
rect 543549 62114 543615 62117
rect 57881 62112 60076 62114
rect 57881 62056 57886 62112
rect 57942 62056 60076 62112
rect 57881 62054 60076 62056
rect 539948 62112 543615 62114
rect 539948 62056 543554 62112
rect 543610 62056 543615 62112
rect 539948 62054 543615 62056
rect 57881 62051 57947 62054
rect 543549 62051 543615 62054
rect 543641 60754 543707 60757
rect 539948 60752 543707 60754
rect 539948 60696 543646 60752
rect 543702 60696 543707 60752
rect 539948 60694 543707 60696
rect 543641 60691 543707 60694
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect 57462 59332 57468 59396
rect 57532 59394 57538 59396
rect 57532 59334 60076 59394
rect 57532 59332 57538 59334
rect 57881 58714 57947 58717
rect 57881 58712 60076 58714
rect -960 58578 480 58668
rect 57881 58656 57886 58712
rect 57942 58656 60076 58712
rect 57881 58654 60076 58656
rect 57881 58651 57947 58654
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 55438 57972 55444 58036
rect 55508 58034 55514 58036
rect 55508 57974 60076 58034
rect 55508 57972 55514 57974
rect 57881 57354 57947 57357
rect 57881 57352 60076 57354
rect 57881 57296 57886 57352
rect 57942 57296 60076 57352
rect 57881 57294 60076 57296
rect 57881 57291 57947 57294
rect 543549 56674 543615 56677
rect 539948 56672 543615 56674
rect 539948 56616 543554 56672
rect 543610 56616 543615 56672
rect 539948 56614 543615 56616
rect 543549 56611 543615 56614
rect 56777 55994 56843 55997
rect 56777 55992 60076 55994
rect 56777 55936 56782 55992
rect 56838 55936 60076 55992
rect 56777 55934 60076 55936
rect 56777 55931 56843 55934
rect 539918 55450 539978 55964
rect 539918 55390 547890 55450
rect 57881 55314 57947 55317
rect 547830 55314 547890 55390
rect 563094 55314 563100 55316
rect 57881 55312 60076 55314
rect 57881 55256 57886 55312
rect 57942 55256 60076 55312
rect 57881 55254 60076 55256
rect 547830 55254 563100 55314
rect 57881 55251 57947 55254
rect 563094 55252 563100 55254
rect 563164 55252 563170 55316
rect 56317 54634 56383 54637
rect 56317 54632 60076 54634
rect 56317 54576 56322 54632
rect 56378 54576 60076 54632
rect 56317 54574 60076 54576
rect 56317 54571 56383 54574
rect 58985 53274 59051 53277
rect 58985 53272 60076 53274
rect 58985 53216 58990 53272
rect 59046 53216 60076 53272
rect 58985 53214 60076 53216
rect 58985 53211 59051 53214
rect 542721 52594 542787 52597
rect 539948 52592 542787 52594
rect 539948 52536 542726 52592
rect 542782 52536 542787 52592
rect 539948 52534 542787 52536
rect 542721 52531 542787 52534
rect 539918 51098 539978 51204
rect 552606 51098 552612 51100
rect 539918 51038 552612 51098
rect 552606 51036 552612 51038
rect 552676 51036 552682 51100
rect 542721 49874 542787 49877
rect 539948 49872 542787 49874
rect 539948 49816 542726 49872
rect 542782 49816 542787 49872
rect 539948 49814 542787 49816
rect 542721 49811 542787 49814
rect 41270 48588 41276 48652
rect 41340 48650 41346 48652
rect 60046 48650 60106 49164
rect 41340 48590 60106 48650
rect 41340 48588 41346 48590
rect 542721 48514 542787 48517
rect 539948 48512 542787 48514
rect 539948 48456 542726 48512
rect 542782 48456 542787 48512
rect 539948 48454 542787 48456
rect 542721 48451 542787 48454
rect 543641 47834 543707 47837
rect 539948 47832 543707 47834
rect 539948 47776 543646 47832
rect 543702 47776 543707 47832
rect 539948 47774 543707 47776
rect 543641 47771 543707 47774
rect 57145 47154 57211 47157
rect 57145 47152 60076 47154
rect 57145 47096 57150 47152
rect 57206 47096 60076 47152
rect 57145 47094 60076 47096
rect 57145 47091 57211 47094
rect 539726 46820 539732 46884
rect 539796 46820 539802 46884
rect 57053 46474 57119 46477
rect 57053 46472 60076 46474
rect 57053 46416 57058 46472
rect 57114 46416 60076 46472
rect 539734 46444 539794 46820
rect 57053 46414 60076 46416
rect 57053 46411 57119 46414
rect 583520 46188 584960 46428
rect 58157 45794 58223 45797
rect 58157 45792 60076 45794
rect 58157 45736 58162 45792
rect 58218 45736 60076 45792
rect 58157 45734 60076 45736
rect 58157 45731 58223 45734
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 57145 45114 57211 45117
rect 543549 45114 543615 45117
rect 57145 45112 60076 45114
rect 57145 45056 57150 45112
rect 57206 45056 60076 45112
rect 57145 45054 60076 45056
rect 539948 45112 543615 45114
rect 539948 45056 543554 45112
rect 543610 45056 543615 45112
rect 539948 45054 543615 45056
rect 57145 45051 57211 45054
rect 543549 45051 543615 45054
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 543641 44434 543707 44437
rect 539948 44432 543707 44434
rect 539948 44376 543646 44432
rect 543702 44376 543707 44432
rect 539948 44374 543707 44376
rect 543641 44371 543707 44374
rect 53046 44298 53052 44300
rect 6870 44238 53052 44298
rect 53046 44236 53052 44238
rect 53116 44236 53122 44300
rect 541249 43754 541315 43757
rect 539948 43752 541315 43754
rect 539948 43696 541254 43752
rect 541310 43696 541315 43752
rect 539948 43694 541315 43696
rect 541249 43691 541315 43694
rect 56041 41714 56107 41717
rect 539918 41714 539978 42364
rect 551502 41714 551508 41716
rect 56041 41712 60076 41714
rect 56041 41656 56046 41712
rect 56102 41656 60076 41712
rect 56041 41654 60076 41656
rect 539918 41654 551508 41714
rect 56041 41651 56107 41654
rect 551502 41652 551508 41654
rect 551572 41652 551578 41716
rect 56685 41034 56751 41037
rect 543549 41034 543615 41037
rect 56685 41032 60076 41034
rect 56685 40976 56690 41032
rect 56746 40976 60076 41032
rect 56685 40974 60076 40976
rect 539948 41032 543615 41034
rect 539948 40976 543554 41032
rect 543610 40976 543615 41032
rect 539948 40974 543615 40976
rect 56685 40971 56751 40974
rect 543549 40971 543615 40974
rect 57881 40354 57947 40357
rect 57881 40352 60076 40354
rect 57881 40296 57886 40352
rect 57942 40296 60076 40352
rect 57881 40294 60076 40296
rect 57881 40291 57947 40294
rect 57881 39674 57947 39677
rect 57881 39672 60076 39674
rect 57881 39616 57886 39672
rect 57942 39616 60076 39672
rect 57881 39614 60076 39616
rect 57881 39611 57947 39614
rect 539910 38524 539916 38588
rect 539980 38524 539986 38588
rect 539918 38284 539978 38524
rect 539918 37362 539978 37604
rect 552422 37362 552428 37364
rect 539918 37302 552428 37362
rect 552422 37300 552428 37302
rect 552492 37300 552498 37364
rect 543549 36274 543615 36277
rect 539948 36272 543615 36274
rect 539948 36216 543554 36272
rect 543610 36216 543615 36272
rect 539948 36214 543615 36216
rect 543549 36211 543615 36214
rect 55622 35532 55628 35596
rect 55692 35594 55698 35596
rect 543641 35594 543707 35597
rect 55692 35534 60076 35594
rect 539948 35592 543707 35594
rect 539948 35536 543646 35592
rect 543702 35536 543707 35592
rect 539948 35534 543707 35536
rect 55692 35532 55698 35534
rect 543641 35531 543707 35534
rect 539542 35260 539548 35324
rect 539612 35260 539618 35324
rect 57646 34852 57652 34916
rect 57716 34914 57722 34916
rect 57716 34854 60076 34914
rect 539550 34884 539610 35260
rect 57716 34852 57722 34854
rect 57881 33554 57947 33557
rect 57881 33552 60076 33554
rect 57881 33496 57886 33552
rect 57942 33496 60076 33552
rect 57881 33494 60076 33496
rect 57881 33491 57947 33494
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect 57881 32874 57947 32877
rect 57881 32872 60076 32874
rect 57881 32816 57886 32872
rect 57942 32816 60076 32872
rect 57881 32814 60076 32816
rect 57881 32811 57947 32814
rect -960 32316 480 32556
rect 56409 32194 56475 32197
rect 56409 32192 60076 32194
rect 56409 32136 56414 32192
rect 56470 32136 60076 32192
rect 56409 32134 60076 32136
rect 56409 32131 56475 32134
rect 45870 30908 45876 30972
rect 45940 30970 45946 30972
rect 60046 30970 60106 31484
rect 539918 31242 539978 31484
rect 543641 31242 543707 31245
rect 539918 31240 543707 31242
rect 539918 31184 543646 31240
rect 543702 31184 543707 31240
rect 539918 31182 543707 31184
rect 543641 31179 543707 31182
rect 539358 31044 539364 31108
rect 539428 31106 539434 31108
rect 560753 31106 560819 31109
rect 539428 31104 560819 31106
rect 539428 31048 560758 31104
rect 560814 31048 560819 31104
rect 539428 31046 560819 31048
rect 539428 31044 539434 31046
rect 560753 31043 560819 31046
rect 45940 30910 60106 30970
rect 45940 30908 45946 30910
rect 540278 30908 540284 30972
rect 540348 30970 540354 30972
rect 554998 30970 555004 30972
rect 540348 30910 555004 30970
rect 540348 30908 540354 30910
rect 554998 30908 555004 30910
rect 555068 30908 555074 30972
rect 59118 30772 59124 30836
rect 59188 30834 59194 30836
rect 59188 30774 60076 30834
rect 59188 30772 59194 30774
rect 539918 30698 539978 30804
rect 542537 30698 542603 30701
rect 539918 30696 542603 30698
rect 539918 30640 542542 30696
rect 542598 30640 542603 30696
rect 539918 30638 542603 30640
rect 542537 30635 542603 30638
rect 543641 30426 543707 30429
rect 552238 30426 552244 30428
rect 543641 30424 552244 30426
rect 543641 30368 543646 30424
rect 543702 30368 552244 30424
rect 543641 30366 552244 30368
rect 543641 30363 543707 30366
rect 552238 30364 552244 30366
rect 552308 30364 552314 30428
rect 59302 29820 59308 29884
rect 59372 29882 59378 29884
rect 59997 29882 60063 29885
rect 59372 29880 60063 29882
rect 59372 29824 60002 29880
rect 60058 29824 60063 29880
rect 59372 29822 60063 29824
rect 59372 29820 59378 29822
rect 59997 29819 60063 29822
rect 55029 29746 55095 29749
rect 60733 29746 60799 29749
rect 55029 29744 60799 29746
rect 55029 29688 55034 29744
rect 55090 29688 60738 29744
rect 60794 29688 60799 29744
rect 55029 29686 60799 29688
rect 55029 29683 55095 29686
rect 60733 29683 60799 29686
rect 50286 29548 50292 29612
rect 50356 29610 50362 29612
rect 61285 29610 61351 29613
rect 50356 29608 61351 29610
rect 50356 29552 61290 29608
rect 61346 29552 61351 29608
rect 50356 29550 61351 29552
rect 50356 29548 50362 29550
rect 61285 29547 61351 29550
rect 537845 29610 537911 29613
rect 545246 29610 545252 29612
rect 537845 29608 545252 29610
rect 537845 29552 537850 29608
rect 537906 29552 545252 29608
rect 537845 29550 545252 29552
rect 537845 29547 537911 29550
rect 545246 29548 545252 29550
rect 545316 29548 545322 29612
rect 52126 29412 52132 29476
rect 52196 29474 52202 29476
rect 85757 29474 85823 29477
rect 52196 29472 85823 29474
rect 52196 29416 85762 29472
rect 85818 29416 85823 29472
rect 52196 29414 85823 29416
rect 52196 29412 52202 29414
rect 85757 29411 85823 29414
rect 519813 29474 519879 29477
rect 547638 29474 547644 29476
rect 519813 29472 547644 29474
rect 519813 29416 519818 29472
rect 519874 29416 547644 29472
rect 519813 29414 547644 29416
rect 519813 29411 519879 29414
rect 547638 29412 547644 29414
rect 547708 29412 547714 29476
rect 31477 29338 31543 29341
rect 244181 29338 244247 29341
rect 31477 29336 244247 29338
rect 31477 29280 31482 29336
rect 31538 29280 244186 29336
rect 244242 29280 244247 29336
rect 31477 29278 244247 29280
rect 31477 29275 31543 29278
rect 244181 29275 244247 29278
rect 359457 29338 359523 29341
rect 561806 29338 561812 29340
rect 359457 29336 561812 29338
rect 359457 29280 359462 29336
rect 359518 29280 561812 29336
rect 359457 29278 561812 29280
rect 359457 29275 359523 29278
rect 561806 29276 561812 29278
rect 561876 29276 561882 29340
rect 27521 29202 27587 29205
rect 284109 29202 284175 29205
rect 27521 29200 284175 29202
rect 27521 29144 27526 29200
rect 27582 29144 284114 29200
rect 284170 29144 284175 29200
rect 27521 29142 284175 29144
rect 27521 29139 27587 29142
rect 284109 29139 284175 29142
rect 314377 29202 314443 29205
rect 561990 29202 561996 29204
rect 314377 29200 561996 29202
rect 314377 29144 314382 29200
rect 314438 29144 561996 29200
rect 314377 29142 561996 29144
rect 314377 29139 314443 29142
rect 561990 29140 561996 29142
rect 562060 29140 562066 29204
rect 575473 29202 575539 29205
rect 575606 29202 575612 29204
rect 575473 29200 575612 29202
rect 575473 29144 575478 29200
rect 575534 29144 575612 29200
rect 575473 29142 575612 29144
rect 575473 29139 575539 29142
rect 575606 29140 575612 29142
rect 575676 29140 575682 29204
rect 31293 29066 31359 29069
rect 373625 29066 373691 29069
rect 31293 29064 373691 29066
rect 31293 29008 31298 29064
rect 31354 29008 373630 29064
rect 373686 29008 373691 29064
rect 31293 29006 373691 29008
rect 31293 29003 31359 29006
rect 373625 29003 373691 29006
rect 509509 29066 509575 29069
rect 543774 29066 543780 29068
rect 509509 29064 543780 29066
rect 509509 29008 509514 29064
rect 509570 29008 543780 29064
rect 509509 29006 543780 29008
rect 509509 29003 509575 29006
rect 543774 29004 543780 29006
rect 543844 29004 543850 29068
rect 59854 28868 59860 28932
rect 59924 28930 59930 28932
rect 78029 28930 78095 28933
rect 59924 28928 78095 28930
rect 59924 28872 78034 28928
rect 78090 28872 78095 28928
rect 59924 28870 78095 28872
rect 59924 28868 59930 28870
rect 78029 28867 78095 28870
rect 127617 28930 127683 28933
rect 579889 28930 579955 28933
rect 127617 28928 579955 28930
rect 127617 28872 127622 28928
rect 127678 28872 579894 28928
rect 579950 28872 579955 28928
rect 127617 28870 579955 28872
rect 127617 28867 127683 28870
rect 579889 28867 579955 28870
rect 39798 28732 39804 28796
rect 39868 28794 39874 28796
rect 213913 28794 213979 28797
rect 39868 28792 213979 28794
rect 39868 28736 213918 28792
rect 213974 28736 213979 28792
rect 39868 28734 213979 28736
rect 39868 28732 39874 28734
rect 213913 28731 213979 28734
rect 234521 28794 234587 28797
rect 541198 28794 541204 28796
rect 234521 28792 541204 28794
rect 234521 28736 234526 28792
rect 234582 28736 541204 28792
rect 234521 28734 541204 28736
rect 234521 28731 234587 28734
rect 541198 28732 541204 28734
rect 541268 28732 541274 28796
rect 38561 28658 38627 28661
rect 319529 28658 319595 28661
rect 38561 28656 319595 28658
rect 38561 28600 38566 28656
rect 38622 28600 319534 28656
rect 319590 28600 319595 28656
rect 38561 28598 319595 28600
rect 38561 28595 38627 28598
rect 319529 28595 319595 28598
rect 377489 28658 377555 28661
rect 577037 28658 577103 28661
rect 377489 28656 577103 28658
rect 377489 28600 377494 28656
rect 377550 28600 577042 28656
rect 577098 28600 577103 28656
rect 377489 28598 577103 28600
rect 377489 28595 377555 28598
rect 577037 28595 577103 28598
rect 44030 28460 44036 28524
rect 44100 28522 44106 28524
rect 175273 28522 175339 28525
rect 44100 28520 175339 28522
rect 44100 28464 175278 28520
rect 175334 28464 175339 28520
rect 44100 28462 175339 28464
rect 44100 28460 44106 28462
rect 175273 28459 175339 28462
rect 452837 28522 452903 28525
rect 560518 28522 560524 28524
rect 452837 28520 560524 28522
rect 452837 28464 452842 28520
rect 452898 28464 560524 28520
rect 452837 28462 560524 28464
rect 452837 28459 452903 28462
rect 560518 28460 560524 28462
rect 560588 28460 560594 28524
rect 50470 28324 50476 28388
rect 50540 28386 50546 28388
rect 91553 28386 91619 28389
rect 50540 28384 91619 28386
rect 50540 28328 91558 28384
rect 91614 28328 91619 28384
rect 50540 28326 91619 28328
rect 50540 28324 50546 28326
rect 91553 28323 91619 28326
rect 92473 28386 92539 28389
rect 169477 28386 169543 28389
rect 92473 28384 169543 28386
rect 92473 28328 92478 28384
rect 92534 28328 169482 28384
rect 169538 28328 169543 28384
rect 92473 28326 169543 28328
rect 92473 28323 92539 28326
rect 169477 28323 169543 28326
rect 487613 28386 487679 28389
rect 566733 28386 566799 28389
rect 487613 28384 566799 28386
rect 487613 28328 487618 28384
rect 487674 28328 566738 28384
rect 566794 28328 566799 28384
rect 487613 28326 566799 28328
rect 487613 28323 487679 28326
rect 566733 28323 566799 28326
rect 58750 28188 58756 28252
rect 58820 28250 58826 28252
rect 65793 28250 65859 28253
rect 58820 28248 65859 28250
rect 58820 28192 65798 28248
rect 65854 28192 65859 28248
rect 58820 28190 65859 28192
rect 58820 28188 58826 28190
rect 65793 28187 65859 28190
rect 72325 28250 72391 28253
rect 96061 28250 96127 28253
rect 72325 28248 96127 28250
rect 72325 28192 72330 28248
rect 72386 28192 96066 28248
rect 96122 28192 96127 28248
rect 72325 28190 96127 28192
rect 72325 28187 72391 28190
rect 96061 28187 96127 28190
rect 97349 28250 97415 28253
rect 186221 28250 186287 28253
rect 97349 28248 186287 28250
rect 97349 28192 97354 28248
rect 97410 28192 186226 28248
rect 186282 28192 186287 28248
rect 97349 28190 186287 28192
rect 97349 28187 97415 28190
rect 186221 28187 186287 28190
rect 474733 28250 474799 28253
rect 552054 28250 552060 28252
rect 474733 28248 552060 28250
rect 474733 28192 474738 28248
rect 474794 28192 552060 28248
rect 474733 28190 552060 28192
rect 474733 28187 474799 28190
rect 552054 28188 552060 28190
rect 552124 28188 552130 28252
rect 45318 28052 45324 28116
rect 45388 28114 45394 28116
rect 117957 28114 118023 28117
rect 45388 28112 118023 28114
rect 45388 28056 117962 28112
rect 118018 28056 118023 28112
rect 45388 28054 118023 28056
rect 45388 28052 45394 28054
rect 117957 28051 118023 28054
rect 48998 27508 49004 27572
rect 49068 27570 49074 27572
rect 66437 27570 66503 27573
rect 49068 27568 66503 27570
rect 49068 27512 66442 27568
rect 66498 27512 66503 27568
rect 49068 27510 66503 27512
rect 49068 27508 49074 27510
rect 66437 27507 66503 27510
rect 525609 27570 525675 27573
rect 549294 27570 549300 27572
rect 525609 27568 549300 27570
rect 525609 27512 525614 27568
rect 525670 27512 549300 27568
rect 525609 27510 549300 27512
rect 525609 27507 525675 27510
rect 549294 27508 549300 27510
rect 549364 27508 549370 27572
rect 30189 27434 30255 27437
rect 69657 27434 69723 27437
rect 30189 27432 69723 27434
rect 30189 27376 30194 27432
rect 30250 27376 69662 27432
rect 69718 27376 69723 27432
rect 30189 27374 69723 27376
rect 30189 27371 30255 27374
rect 69657 27371 69723 27374
rect 174629 27434 174695 27437
rect 561070 27434 561076 27436
rect 174629 27432 561076 27434
rect 174629 27376 174634 27432
rect 174690 27376 561076 27432
rect 174629 27374 561076 27376
rect 174629 27371 174695 27374
rect 561070 27372 561076 27374
rect 561140 27372 561146 27436
rect 44950 27236 44956 27300
rect 45020 27298 45026 27300
rect 389725 27298 389791 27301
rect 45020 27296 389791 27298
rect 45020 27240 389730 27296
rect 389786 27240 389791 27296
rect 45020 27238 389791 27240
rect 45020 27236 45026 27238
rect 389725 27235 389791 27238
rect 421925 27298 421991 27301
rect 566038 27298 566044 27300
rect 421925 27296 566044 27298
rect 421925 27240 421930 27296
rect 421986 27240 566044 27296
rect 421925 27238 566044 27240
rect 421925 27235 421991 27238
rect 566038 27236 566044 27238
rect 566108 27236 566114 27300
rect 378225 27162 378291 27165
rect 578550 27162 578556 27164
rect 378225 27160 578556 27162
rect 378225 27104 378230 27160
rect 378286 27104 578556 27160
rect 378225 27102 578556 27104
rect 378225 27099 378291 27102
rect 578550 27100 578556 27102
rect 578620 27100 578626 27164
rect 43846 26964 43852 27028
rect 43916 27026 43922 27028
rect 369117 27026 369183 27029
rect 43916 27024 369183 27026
rect 43916 26968 369122 27024
rect 369178 26968 369183 27024
rect 43916 26966 369183 26968
rect 43916 26964 43922 26966
rect 369117 26963 369183 26966
rect 511441 27026 511507 27029
rect 545062 27026 545068 27028
rect 511441 27024 545068 27026
rect 511441 26968 511446 27024
rect 511502 26968 545068 27024
rect 511441 26966 545068 26968
rect 511441 26963 511507 26966
rect 545062 26964 545068 26966
rect 545132 26964 545138 27028
rect 358905 26890 358971 26893
rect 561622 26890 561628 26892
rect 358905 26888 561628 26890
rect 358905 26832 358910 26888
rect 358966 26832 561628 26888
rect 358905 26830 561628 26832
rect 358905 26827 358971 26830
rect 561622 26828 561628 26830
rect 561692 26828 561698 26892
rect 42006 26692 42012 26756
rect 42076 26754 42082 26756
rect 382641 26754 382707 26757
rect 42076 26752 382707 26754
rect 42076 26696 382646 26752
rect 382702 26696 382707 26752
rect 42076 26694 382707 26696
rect 42076 26692 42082 26694
rect 382641 26691 382707 26694
rect 510797 26754 510863 26757
rect 545614 26754 545620 26756
rect 510797 26752 545620 26754
rect 510797 26696 510802 26752
rect 510858 26696 545620 26752
rect 510797 26694 545620 26696
rect 510797 26691 510863 26694
rect 545614 26692 545620 26694
rect 545684 26692 545690 26756
rect 36486 26556 36492 26620
rect 36556 26618 36562 26620
rect 524321 26618 524387 26621
rect 36556 26616 524387 26618
rect 36556 26560 524326 26616
rect 524382 26560 524387 26616
rect 36556 26558 524387 26560
rect 36556 26556 36562 26558
rect 524321 26555 524387 26558
rect 485037 26210 485103 26213
rect 567142 26210 567148 26212
rect 485037 26208 567148 26210
rect 485037 26152 485042 26208
rect 485098 26152 567148 26208
rect 485037 26150 567148 26152
rect 485037 26147 485103 26150
rect 567142 26148 567148 26150
rect 567212 26148 567218 26212
rect 32990 26012 32996 26076
rect 33060 26074 33066 26076
rect 478873 26074 478939 26077
rect 33060 26072 478939 26074
rect 33060 26016 478878 26072
rect 478934 26016 478939 26072
rect 33060 26014 478939 26016
rect 33060 26012 33066 26014
rect 478873 26011 478939 26014
rect 479057 26074 479123 26077
rect 576945 26074 577011 26077
rect 479057 26072 577011 26074
rect 479057 26016 479062 26072
rect 479118 26016 576950 26072
rect 577006 26016 577011 26072
rect 479057 26014 577011 26016
rect 479057 26011 479123 26014
rect 576945 26011 577011 26014
rect 38510 25876 38516 25940
rect 38580 25938 38586 25940
rect 408493 25938 408559 25941
rect 38580 25936 408559 25938
rect 38580 25880 408498 25936
rect 408554 25880 408559 25936
rect 38580 25878 408559 25880
rect 38580 25876 38586 25878
rect 408493 25875 408559 25878
rect 409873 25938 409939 25941
rect 554865 25938 554931 25941
rect 409873 25936 554931 25938
rect 409873 25880 409878 25936
rect 409934 25880 554870 25936
rect 554926 25880 554931 25936
rect 409873 25878 554931 25880
rect 409873 25875 409939 25878
rect 554865 25875 554931 25878
rect 37590 25740 37596 25804
rect 37660 25802 37666 25804
rect 364425 25802 364491 25805
rect 37660 25800 364491 25802
rect 37660 25744 364430 25800
rect 364486 25744 364491 25800
rect 37660 25742 364491 25744
rect 37660 25740 37666 25742
rect 364425 25739 364491 25742
rect 373993 25802 374059 25805
rect 577313 25802 577379 25805
rect 373993 25800 577379 25802
rect 373993 25744 373998 25800
rect 374054 25744 577318 25800
rect 577374 25744 577379 25800
rect 373993 25742 577379 25744
rect 373993 25739 374059 25742
rect 577313 25739 577379 25742
rect 60038 25604 60044 25668
rect 60108 25666 60114 25668
rect 207013 25666 207079 25669
rect 60108 25664 207079 25666
rect 60108 25608 207018 25664
rect 207074 25608 207079 25664
rect 60108 25606 207079 25608
rect 60108 25604 60114 25606
rect 207013 25603 207079 25606
rect 332593 25666 332659 25669
rect 566406 25666 566412 25668
rect 332593 25664 566412 25666
rect 332593 25608 332598 25664
rect 332654 25608 566412 25664
rect 332593 25606 566412 25608
rect 332593 25603 332659 25606
rect 566406 25604 566412 25606
rect 566476 25604 566482 25668
rect 53230 25468 53236 25532
rect 53300 25530 53306 25532
rect 53649 25530 53715 25533
rect 53300 25528 53715 25530
rect 53300 25472 53654 25528
rect 53710 25472 53715 25528
rect 53300 25470 53715 25472
rect 53300 25468 53306 25470
rect 53649 25467 53715 25470
rect 54518 25468 54524 25532
rect 54588 25530 54594 25532
rect 88333 25530 88399 25533
rect 54588 25528 88399 25530
rect 54588 25472 88338 25528
rect 88394 25472 88399 25528
rect 54588 25470 88399 25472
rect 54588 25468 54594 25470
rect 88333 25467 88399 25470
rect 339493 25530 339559 25533
rect 575565 25530 575631 25533
rect 339493 25528 575631 25530
rect 339493 25472 339498 25528
rect 339554 25472 575570 25528
rect 575626 25472 575631 25528
rect 339493 25470 575631 25472
rect 339493 25467 339559 25470
rect 575565 25467 575631 25470
rect 53414 25332 53420 25396
rect 53484 25394 53490 25396
rect 70393 25394 70459 25397
rect 53484 25392 70459 25394
rect 53484 25336 70398 25392
rect 70454 25336 70459 25392
rect 53484 25334 70459 25336
rect 53484 25332 53490 25334
rect 70393 25331 70459 25334
rect 448605 25394 448671 25397
rect 538806 25394 538812 25396
rect 448605 25392 538812 25394
rect 448605 25336 448610 25392
rect 448666 25336 538812 25392
rect 448605 25334 538812 25336
rect 448605 25331 448671 25334
rect 538806 25332 538812 25334
rect 538876 25332 538882 25396
rect 32806 25196 32812 25260
rect 32876 25258 32882 25260
rect 484577 25258 484643 25261
rect 32876 25256 484643 25258
rect 32876 25200 484582 25256
rect 484638 25200 484643 25256
rect 32876 25198 484643 25200
rect 32876 25196 32882 25198
rect 484577 25195 484643 25198
rect 41781 24850 41847 24853
rect 473445 24850 473511 24853
rect 41781 24848 473511 24850
rect 41781 24792 41786 24848
rect 41842 24792 473450 24848
rect 473506 24792 473511 24848
rect 41781 24790 473511 24792
rect 41781 24787 41847 24790
rect 473445 24787 473511 24790
rect 484485 24850 484551 24853
rect 547270 24850 547276 24852
rect 484485 24848 547276 24850
rect 484485 24792 484490 24848
rect 484546 24792 547276 24848
rect 484485 24790 547276 24792
rect 484485 24787 484551 24790
rect 547270 24788 547276 24790
rect 547340 24788 547346 24852
rect 30281 24714 30347 24717
rect 459645 24714 459711 24717
rect 30281 24712 459711 24714
rect 30281 24656 30286 24712
rect 30342 24656 459650 24712
rect 459706 24656 459711 24712
rect 30281 24654 459711 24656
rect 30281 24651 30347 24654
rect 459645 24651 459711 24654
rect 54702 24516 54708 24580
rect 54772 24578 54778 24580
rect 100753 24578 100819 24581
rect 54772 24576 100819 24578
rect 54772 24520 100758 24576
rect 100814 24520 100819 24576
rect 54772 24518 100819 24520
rect 54772 24516 54778 24518
rect 100753 24515 100819 24518
rect 165797 24578 165863 24581
rect 556654 24578 556660 24580
rect 165797 24576 556660 24578
rect 165797 24520 165802 24576
rect 165858 24520 556660 24576
rect 165797 24518 556660 24520
rect 165797 24515 165863 24518
rect 556654 24516 556660 24518
rect 556724 24516 556730 24580
rect 52310 24380 52316 24444
rect 52380 24442 52386 24444
rect 74533 24442 74599 24445
rect 52380 24440 74599 24442
rect 52380 24384 74538 24440
rect 74594 24384 74599 24440
rect 52380 24382 74599 24384
rect 52380 24380 52386 24382
rect 74533 24379 74599 24382
rect 274633 24442 274699 24445
rect 565302 24442 565308 24444
rect 274633 24440 565308 24442
rect 274633 24384 274638 24440
rect 274694 24384 565308 24440
rect 274633 24382 565308 24384
rect 274633 24379 274699 24382
rect 565302 24380 565308 24382
rect 565372 24380 565378 24444
rect 207013 24306 207079 24309
rect 567326 24306 567332 24308
rect 207013 24304 567332 24306
rect 207013 24248 207018 24304
rect 207074 24248 567332 24304
rect 207013 24246 567332 24248
rect 207013 24243 207079 24246
rect 567326 24244 567332 24246
rect 567396 24244 567402 24308
rect 164233 24170 164299 24173
rect 553342 24170 553348 24172
rect 164233 24168 553348 24170
rect 164233 24112 164238 24168
rect 164294 24112 553348 24168
rect 164233 24110 553348 24112
rect 164233 24107 164299 24110
rect 553342 24108 553348 24110
rect 553412 24108 553418 24172
rect 39062 23972 39068 24036
rect 39132 24034 39138 24036
rect 300945 24034 301011 24037
rect 39132 24032 301011 24034
rect 39132 23976 300950 24032
rect 301006 23976 301011 24032
rect 39132 23974 301011 23976
rect 39132 23972 39138 23974
rect 300945 23971 301011 23974
rect 347865 24034 347931 24037
rect 566222 24034 566228 24036
rect 347865 24032 566228 24034
rect 347865 23976 347870 24032
rect 347926 23976 566228 24032
rect 347865 23974 566228 23976
rect 347865 23971 347931 23974
rect 566222 23972 566228 23974
rect 566292 23972 566298 24036
rect 64873 23354 64939 23357
rect 581269 23354 581335 23357
rect 64873 23352 581335 23354
rect 64873 23296 64878 23352
rect 64934 23296 581274 23352
rect 581330 23296 581335 23352
rect 64873 23294 581335 23296
rect 64873 23291 64939 23294
rect 581269 23291 581335 23294
rect 21909 23218 21975 23221
rect 468937 23218 469003 23221
rect 21909 23216 469003 23218
rect 21909 23160 21914 23216
rect 21970 23160 468942 23216
rect 468998 23160 469003 23216
rect 21909 23158 469003 23160
rect 21909 23155 21975 23158
rect 468937 23155 469003 23158
rect 53598 23020 53604 23084
rect 53668 23082 53674 23084
rect 125685 23082 125751 23085
rect 53668 23080 125751 23082
rect 53668 23024 125690 23080
rect 125746 23024 125751 23080
rect 53668 23022 125751 23024
rect 53668 23020 53674 23022
rect 125685 23019 125751 23022
rect 138013 23082 138079 23085
rect 581126 23082 581132 23084
rect 138013 23080 581132 23082
rect 138013 23024 138018 23080
rect 138074 23024 581132 23080
rect 138013 23022 581132 23024
rect 138013 23019 138079 23022
rect 581126 23020 581132 23022
rect 581196 23020 581202 23084
rect 24485 22946 24551 22949
rect 426525 22946 426591 22949
rect 24485 22944 426591 22946
rect 24485 22888 24490 22944
rect 24546 22888 426530 22944
rect 426586 22888 426591 22944
rect 24485 22886 426591 22888
rect 24485 22883 24551 22886
rect 426525 22883 426591 22886
rect 445845 22946 445911 22949
rect 548374 22946 548380 22948
rect 445845 22944 548380 22946
rect 445845 22888 445850 22944
rect 445906 22888 548380 22944
rect 445845 22886 548380 22888
rect 445845 22883 445911 22886
rect 548374 22884 548380 22886
rect 548444 22884 548450 22948
rect 23289 22810 23355 22813
rect 415393 22810 415459 22813
rect 23289 22808 415459 22810
rect 23289 22752 23294 22808
rect 23350 22752 415398 22808
rect 415454 22752 415459 22808
rect 23289 22750 415459 22752
rect 23289 22747 23355 22750
rect 415393 22747 415459 22750
rect 416681 22810 416747 22813
rect 579654 22810 579660 22812
rect 416681 22808 579660 22810
rect 416681 22752 416686 22808
rect 416742 22752 579660 22808
rect 416681 22750 579660 22752
rect 416681 22747 416747 22750
rect 579654 22748 579660 22750
rect 579724 22748 579730 22812
rect 48078 22612 48084 22676
rect 48148 22674 48154 22676
rect 324405 22674 324471 22677
rect 48148 22672 324471 22674
rect 48148 22616 324410 22672
rect 324466 22616 324471 22672
rect 48148 22614 324471 22616
rect 48148 22612 48154 22614
rect 324405 22611 324471 22614
rect 391933 22674 391999 22677
rect 547086 22674 547092 22676
rect 391933 22672 547092 22674
rect 391933 22616 391938 22672
rect 391994 22616 547092 22672
rect 391933 22614 547092 22616
rect 391933 22611 391999 22614
rect 547086 22612 547092 22614
rect 547156 22612 547162 22676
rect 304993 22538 305059 22541
rect 578734 22538 578740 22540
rect 304993 22536 578740 22538
rect 304993 22480 304998 22536
rect 305054 22480 578740 22536
rect 304993 22478 578740 22480
rect 304993 22475 305059 22478
rect 578734 22476 578740 22478
rect 578804 22476 578810 22540
rect 35750 21932 35756 21996
rect 35820 21994 35826 21996
rect 445753 21994 445819 21997
rect 35820 21992 445819 21994
rect 35820 21936 445758 21992
rect 445814 21936 445819 21992
rect 35820 21934 445819 21936
rect 35820 21932 35826 21934
rect 445753 21931 445819 21934
rect 465165 21994 465231 21997
rect 540278 21994 540284 21996
rect 465165 21992 540284 21994
rect 465165 21936 465170 21992
rect 465226 21936 540284 21992
rect 465165 21934 540284 21936
rect 465165 21931 465231 21934
rect 540278 21932 540284 21934
rect 540348 21932 540354 21996
rect 49550 21796 49556 21860
rect 49620 21858 49626 21860
rect 107653 21858 107719 21861
rect 49620 21856 107719 21858
rect 49620 21800 107658 21856
rect 107714 21800 107719 21856
rect 49620 21798 107719 21800
rect 49620 21796 49626 21798
rect 107653 21795 107719 21798
rect 235993 21858 236059 21861
rect 565486 21858 565492 21860
rect 235993 21856 565492 21858
rect 235993 21800 235998 21856
rect 236054 21800 565492 21856
rect 235993 21798 565492 21800
rect 235993 21795 236059 21798
rect 565486 21796 565492 21798
rect 565556 21796 565562 21860
rect 57513 21722 57579 21725
rect 97349 21722 97415 21725
rect 57513 21720 97415 21722
rect 57513 21664 57518 21720
rect 57574 21664 97354 21720
rect 97410 21664 97415 21720
rect 57513 21662 97415 21664
rect 57513 21659 57579 21662
rect 97349 21659 97415 21662
rect 179413 21722 179479 21725
rect 571374 21722 571380 21724
rect 179413 21720 571380 21722
rect 179413 21664 179418 21720
rect 179474 21664 571380 21720
rect 179413 21662 571380 21664
rect 179413 21659 179479 21662
rect 571374 21660 571380 21662
rect 571444 21660 571450 21724
rect 161473 21586 161539 21589
rect 565118 21586 565124 21588
rect 161473 21584 565124 21586
rect 161473 21528 161478 21584
rect 161534 21528 565124 21584
rect 161473 21526 565124 21528
rect 161473 21523 161539 21526
rect 565118 21524 565124 21526
rect 565188 21524 565194 21588
rect 50654 21388 50660 21452
rect 50724 21450 50730 21452
rect 125685 21450 125751 21453
rect 50724 21448 125751 21450
rect 50724 21392 125690 21448
rect 125746 21392 125751 21448
rect 50724 21390 125751 21392
rect 50724 21388 50730 21390
rect 125685 21387 125751 21390
rect 150433 21450 150499 21453
rect 567510 21450 567516 21452
rect 150433 21448 567516 21450
rect 150433 21392 150438 21448
rect 150494 21392 567516 21448
rect 150433 21390 567516 21392
rect 150433 21387 150499 21390
rect 567510 21388 567516 21390
rect 567580 21388 567586 21452
rect 49182 21252 49188 21316
rect 49252 21314 49258 21316
rect 124213 21314 124279 21317
rect 49252 21312 124279 21314
rect 49252 21256 124218 21312
rect 124274 21256 124279 21312
rect 49252 21254 124279 21256
rect 49252 21252 49258 21254
rect 124213 21251 124279 21254
rect 135253 21314 135319 21317
rect 570086 21314 570092 21316
rect 135253 21312 570092 21314
rect 135253 21256 135258 21312
rect 135314 21256 570092 21312
rect 135253 21254 570092 21256
rect 135253 21251 135319 21254
rect 570086 21252 570092 21254
rect 570156 21252 570162 21316
rect 407113 21178 407179 21181
rect 558862 21178 558868 21180
rect 407113 21176 558868 21178
rect 407113 21120 407118 21176
rect 407174 21120 558868 21176
rect 407113 21118 558868 21120
rect 407113 21115 407179 21118
rect 558862 21116 558868 21118
rect 558932 21116 558938 21180
rect 31518 20572 31524 20636
rect 31588 20634 31594 20636
rect 538305 20634 538371 20637
rect 31588 20632 538371 20634
rect 31588 20576 538310 20632
rect 538366 20576 538371 20632
rect 31588 20574 538371 20576
rect 31588 20572 31594 20574
rect 538305 20571 538371 20574
rect 22737 20498 22803 20501
rect 525793 20498 525859 20501
rect 22737 20496 525859 20498
rect 22737 20440 22742 20496
rect 22798 20440 525798 20496
rect 525854 20440 525859 20496
rect 22737 20438 525859 20440
rect 22737 20435 22803 20438
rect 525793 20435 525859 20438
rect 20529 20362 20595 20365
rect 505093 20362 505159 20365
rect 20529 20360 505159 20362
rect 20529 20304 20534 20360
rect 20590 20304 505098 20360
rect 505154 20304 505159 20360
rect 20529 20302 505159 20304
rect 20529 20299 20595 20302
rect 505093 20299 505159 20302
rect 526437 20362 526503 20365
rect 558269 20362 558335 20365
rect 526437 20360 558335 20362
rect 526437 20304 526442 20360
rect 526498 20304 558274 20360
rect 558330 20304 558335 20360
rect 526437 20302 558335 20304
rect 526437 20299 526503 20302
rect 558269 20299 558335 20302
rect 27470 20164 27476 20228
rect 27540 20226 27546 20228
rect 448513 20226 448579 20229
rect 27540 20224 448579 20226
rect 27540 20168 448518 20224
rect 448574 20168 448579 20224
rect 27540 20166 448579 20168
rect 27540 20164 27546 20166
rect 448513 20163 448579 20166
rect 463785 20226 463851 20229
rect 543222 20226 543228 20228
rect 463785 20224 543228 20226
rect 463785 20168 463790 20224
rect 463846 20168 543228 20224
rect 463785 20166 543228 20168
rect 463785 20163 463851 20166
rect 543222 20164 543228 20166
rect 543292 20164 543298 20228
rect 173893 20090 173959 20093
rect 579705 20090 579771 20093
rect 173893 20088 579771 20090
rect 173893 20032 173898 20088
rect 173954 20032 579710 20088
rect 579766 20032 579771 20088
rect 173893 20030 579771 20032
rect 173893 20027 173959 20030
rect 579705 20027 579771 20030
rect 49366 19892 49372 19956
rect 49436 19954 49442 19956
rect 151813 19954 151879 19957
rect 49436 19952 151879 19954
rect 49436 19896 151818 19952
rect 151874 19896 151879 19952
rect 49436 19894 151879 19896
rect 49436 19892 49442 19894
rect 151813 19891 151879 19894
rect 204253 19954 204319 19957
rect 554814 19954 554820 19956
rect 204253 19952 554820 19954
rect 204253 19896 204258 19952
rect 204314 19896 554820 19952
rect 204253 19894 554820 19896
rect 204253 19891 204319 19894
rect 554814 19892 554820 19894
rect 554884 19892 554890 19956
rect 578877 19818 578943 19821
rect 583520 19818 584960 19908
rect 578877 19816 584960 19818
rect 578877 19760 578882 19816
rect 578938 19760 584960 19816
rect 578877 19758 584960 19760
rect 578877 19755 578943 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 28206 19410 28212 19412
rect -960 19350 28212 19410
rect -960 19260 480 19350
rect 28206 19348 28212 19350
rect 28276 19348 28282 19412
rect 57237 19274 57303 19277
rect 336733 19274 336799 19277
rect 57237 19272 336799 19274
rect 57237 19216 57242 19272
rect 57298 19216 336738 19272
rect 336794 19216 336799 19272
rect 57237 19214 336799 19216
rect 57237 19211 57303 19214
rect 336733 19211 336799 19214
rect 47710 19076 47716 19140
rect 47780 19138 47786 19140
rect 291193 19138 291259 19141
rect 47780 19136 291259 19138
rect 47780 19080 291198 19136
rect 291254 19080 291259 19136
rect 47780 19078 291259 19080
rect 47780 19076 47786 19078
rect 291193 19075 291259 19078
rect 300853 19138 300919 19141
rect 544326 19138 544332 19140
rect 300853 19136 544332 19138
rect 300853 19080 300858 19136
rect 300914 19080 544332 19136
rect 300853 19078 544332 19080
rect 300853 19075 300919 19078
rect 544326 19076 544332 19078
rect 544396 19076 544402 19140
rect 58566 18940 58572 19004
rect 58636 19002 58642 19004
rect 222193 19002 222259 19005
rect 58636 19000 222259 19002
rect 58636 18944 222198 19000
rect 222254 18944 222259 19000
rect 58636 18942 222259 18944
rect 58636 18940 58642 18942
rect 222193 18939 222259 18942
rect 282913 19002 282979 19005
rect 559046 19002 559052 19004
rect 282913 19000 559052 19002
rect 282913 18944 282918 19000
rect 282974 18944 559052 19000
rect 282913 18942 559052 18944
rect 282913 18939 282979 18942
rect 559046 18940 559052 18942
rect 559116 18940 559122 19004
rect 44766 18804 44772 18868
rect 44836 18866 44842 18868
rect 139485 18866 139551 18869
rect 44836 18864 139551 18866
rect 44836 18808 139490 18864
rect 139546 18808 139551 18864
rect 44836 18806 139551 18808
rect 44836 18804 44842 18806
rect 139485 18803 139551 18806
rect 267733 18866 267799 18869
rect 558126 18866 558132 18868
rect 267733 18864 558132 18866
rect 267733 18808 267738 18864
rect 267794 18808 558132 18864
rect 267733 18806 558132 18808
rect 267733 18803 267799 18806
rect 558126 18804 558132 18806
rect 558196 18804 558202 18868
rect 278773 18730 278839 18733
rect 574134 18730 574140 18732
rect 278773 18728 574140 18730
rect 278773 18672 278778 18728
rect 278834 18672 574140 18728
rect 278773 18670 574140 18672
rect 278773 18667 278839 18670
rect 574134 18668 574140 18670
rect 574204 18668 574210 18732
rect 128353 18594 128419 18597
rect 553710 18594 553716 18596
rect 128353 18592 553716 18594
rect 128353 18536 128358 18592
rect 128414 18536 553716 18592
rect 128353 18534 553716 18536
rect 128353 18531 128419 18534
rect 553710 18532 553716 18534
rect 553780 18532 553786 18596
rect 178033 17778 178099 17781
rect 580942 17778 580948 17780
rect 178033 17776 580948 17778
rect 178033 17720 178038 17776
rect 178094 17720 580948 17776
rect 178033 17718 580948 17720
rect 178033 17715 178099 17718
rect 580942 17716 580948 17718
rect 581012 17716 581018 17780
rect 212625 17642 212691 17645
rect 542670 17642 542676 17644
rect 212625 17640 542676 17642
rect 212625 17584 212630 17640
rect 212686 17584 542676 17640
rect 212625 17582 542676 17584
rect 212625 17579 212691 17582
rect 542670 17580 542676 17582
rect 542740 17580 542746 17644
rect 560293 17642 560359 17645
rect 560702 17642 560708 17644
rect 560293 17640 560708 17642
rect 560293 17584 560298 17640
rect 560354 17584 560708 17640
rect 560293 17582 560708 17584
rect 560293 17579 560359 17582
rect 560702 17580 560708 17582
rect 560772 17580 560778 17644
rect 353293 17506 353359 17509
rect 575422 17506 575428 17508
rect 353293 17504 575428 17506
rect 353293 17448 353298 17504
rect 353354 17448 575428 17504
rect 353293 17446 575428 17448
rect 353293 17443 353359 17446
rect 575422 17444 575428 17446
rect 575492 17444 575498 17508
rect 335353 17370 335419 17373
rect 557574 17370 557580 17372
rect 335353 17368 557580 17370
rect 335353 17312 335358 17368
rect 335414 17312 557580 17368
rect 335353 17310 557580 17312
rect 335353 17307 335419 17310
rect 557574 17308 557580 17310
rect 557644 17308 557650 17372
rect 218053 17234 218119 17237
rect 556470 17234 556476 17236
rect 218053 17232 556476 17234
rect 218053 17176 218058 17232
rect 218114 17176 556476 17232
rect 218053 17174 556476 17176
rect 218053 17171 218119 17174
rect 556470 17172 556476 17174
rect 556540 17172 556546 17236
rect 402973 17098 403039 17101
rect 542854 17098 542860 17100
rect 402973 17096 542860 17098
rect 402973 17040 402978 17096
rect 403034 17040 542860 17096
rect 402973 17038 542860 17040
rect 402973 17035 403039 17038
rect 542854 17036 542860 17038
rect 542924 17036 542930 17100
rect 84193 16962 84259 16965
rect 563462 16962 563468 16964
rect 84193 16960 563468 16962
rect 84193 16904 84198 16960
rect 84254 16904 563468 16960
rect 84193 16902 563468 16904
rect 84193 16899 84259 16902
rect 563462 16900 563468 16902
rect 563532 16900 563538 16964
rect 39246 16492 39252 16556
rect 39316 16554 39322 16556
rect 150525 16554 150591 16557
rect 39316 16552 150591 16554
rect 39316 16496 150530 16552
rect 150586 16496 150591 16552
rect 39316 16494 150591 16496
rect 39316 16492 39322 16494
rect 150525 16491 150591 16494
rect 431953 16554 432019 16557
rect 547454 16554 547460 16556
rect 431953 16552 547460 16554
rect 431953 16496 431958 16552
rect 432014 16496 547460 16552
rect 431953 16494 547460 16496
rect 431953 16491 432019 16494
rect 547454 16492 547460 16494
rect 547524 16492 547530 16556
rect 440325 16418 440391 16421
rect 544142 16418 544148 16420
rect 440325 16416 544148 16418
rect 440325 16360 440330 16416
rect 440386 16360 544148 16416
rect 440325 16358 544148 16360
rect 440325 16355 440391 16358
rect 544142 16356 544148 16358
rect 544212 16356 544218 16420
rect 214465 16146 214531 16149
rect 580993 16146 581059 16149
rect 214465 16144 581059 16146
rect 214465 16088 214470 16144
rect 214526 16088 580998 16144
rect 581054 16088 581059 16144
rect 214465 16086 581059 16088
rect 214465 16083 214531 16086
rect 580993 16083 581059 16086
rect 143533 16010 143599 16013
rect 550582 16010 550588 16012
rect 143533 16008 550588 16010
rect 143533 15952 143538 16008
rect 143594 15952 550588 16008
rect 143533 15950 550588 15952
rect 143533 15947 143599 15950
rect 550582 15948 550588 15950
rect 550652 15948 550658 16012
rect 157793 15874 157859 15877
rect 582465 15874 582531 15877
rect 157793 15872 582531 15874
rect 157793 15816 157798 15872
rect 157854 15816 582470 15872
rect 582526 15816 582531 15872
rect 157793 15814 582531 15816
rect 157793 15811 157859 15814
rect 582465 15811 582531 15814
rect 220905 15194 220971 15197
rect 543038 15194 543044 15196
rect 220905 15192 543044 15194
rect 220905 15136 220910 15192
rect 220966 15136 543044 15192
rect 220905 15134 543044 15136
rect 220905 15131 220971 15134
rect 543038 15132 543044 15134
rect 543108 15132 543114 15196
rect 386413 15058 386479 15061
rect 541382 15058 541388 15060
rect 386413 15056 541388 15058
rect 386413 15000 386418 15056
rect 386474 15000 541388 15056
rect 386413 14998 541388 15000
rect 386413 14995 386479 14998
rect 541382 14996 541388 14998
rect 541452 14996 541458 15060
rect 438853 14922 438919 14925
rect 548006 14922 548012 14924
rect 438853 14920 548012 14922
rect 438853 14864 438858 14920
rect 438914 14864 548012 14920
rect 438853 14862 548012 14864
rect 438853 14859 438919 14862
rect 548006 14860 548012 14862
rect 548076 14860 548082 14924
rect 236545 14514 236611 14517
rect 549846 14514 549852 14516
rect 236545 14512 549852 14514
rect 236545 14456 236550 14512
rect 236606 14456 549852 14512
rect 236545 14454 549852 14456
rect 236545 14451 236611 14454
rect 549846 14452 549852 14454
rect 549916 14452 549922 14516
rect 339585 13698 339651 13701
rect 540094 13698 540100 13700
rect 339585 13696 540100 13698
rect 339585 13640 339590 13696
rect 339646 13640 540100 13696
rect 339585 13638 540100 13640
rect 339585 13635 339651 13638
rect 540094 13636 540100 13638
rect 540164 13636 540170 13700
rect 324405 13018 324471 13021
rect 545430 13018 545436 13020
rect 324405 13016 545436 13018
rect 324405 12960 324410 13016
rect 324466 12960 545436 13016
rect 324405 12958 545436 12960
rect 324405 12955 324471 12958
rect 545430 12956 545436 12958
rect 545500 12956 545506 13020
rect 484393 12338 484459 12341
rect 580165 12338 580231 12341
rect 484393 12336 580231 12338
rect 484393 12280 484398 12336
rect 484454 12280 580170 12336
rect 580226 12280 580231 12336
rect 484393 12278 580231 12280
rect 484393 12275 484459 12278
rect 580165 12275 580231 12278
rect 328729 11794 328795 11797
rect 557758 11794 557764 11796
rect 328729 11792 557764 11794
rect 328729 11736 328734 11792
rect 328790 11736 557764 11792
rect 328729 11734 557764 11736
rect 328729 11731 328795 11734
rect 557758 11732 557764 11734
rect 557828 11732 557834 11796
rect 46657 11658 46723 11661
rect 560886 11658 560892 11660
rect 46657 11656 560892 11658
rect 46657 11600 46662 11656
rect 46718 11600 560892 11656
rect 46657 11598 560892 11600
rect 46657 11595 46723 11598
rect 560886 11596 560892 11598
rect 560956 11596 560962 11660
rect 201493 10434 201559 10437
rect 556286 10434 556292 10436
rect 201493 10432 556292 10434
rect 201493 10376 201498 10432
rect 201554 10376 556292 10432
rect 201493 10374 556292 10376
rect 201493 10371 201559 10374
rect 556286 10372 556292 10374
rect 556356 10372 556362 10436
rect 35382 10236 35388 10300
rect 35452 10298 35458 10300
rect 132953 10298 133019 10301
rect 504357 10298 504423 10301
rect 35452 10296 504423 10298
rect 35452 10240 132958 10296
rect 133014 10240 504362 10296
rect 504418 10240 504423 10296
rect 35452 10238 504423 10240
rect 35452 10236 35458 10238
rect 132953 10235 133019 10238
rect 504357 10235 504423 10238
rect 276013 7714 276079 7717
rect 557942 7714 557948 7716
rect 276013 7712 557948 7714
rect 276013 7656 276018 7712
rect 276074 7656 557948 7712
rect 276013 7654 557948 7656
rect 276013 7651 276079 7654
rect 557942 7652 557948 7654
rect 558012 7652 558018 7716
rect 155401 7578 155467 7581
rect 556102 7578 556108 7580
rect 155401 7576 556108 7578
rect 155401 7520 155406 7576
rect 155462 7520 556108 7576
rect 155401 7518 556108 7520
rect 155401 7515 155467 7518
rect 556102 7516 556108 7518
rect 556172 7516 556178 7580
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 485221 6354 485287 6357
rect 562174 6354 562180 6356
rect 485221 6352 562180 6354
rect 485221 6296 485226 6352
rect 485282 6296 562180 6352
rect 485221 6294 562180 6296
rect 485221 6291 485287 6294
rect 562174 6292 562180 6294
rect 562244 6292 562250 6356
rect 179045 6218 179111 6221
rect 553526 6218 553532 6220
rect 179045 6216 553532 6218
rect 179045 6160 179050 6216
rect 179106 6160 553532 6216
rect 179045 6158 553532 6160
rect 179045 6155 179111 6158
rect 553526 6156 553532 6158
rect 553596 6156 553602 6220
rect 64321 4858 64387 4861
rect 559230 4858 559236 4860
rect 64321 4856 559236 4858
rect 64321 4800 64326 4856
rect 64382 4800 559236 4856
rect 64321 4798 559236 4800
rect 64321 4795 64387 4798
rect 559230 4796 559236 4798
rect 559300 4796 559306 4860
rect 531313 4042 531379 4045
rect 565854 4042 565860 4044
rect 531313 4040 565860 4042
rect 531313 3984 531318 4040
rect 531374 3984 565860 4040
rect 531313 3982 565860 3984
rect 531313 3979 531379 3982
rect 565854 3980 565860 3982
rect 565924 3980 565930 4044
rect 506473 3906 506539 3909
rect 563278 3906 563284 3908
rect 506473 3904 563284 3906
rect 506473 3848 506478 3904
rect 506534 3848 563284 3904
rect 506473 3846 563284 3848
rect 506473 3843 506539 3846
rect 563278 3844 563284 3846
rect 563348 3844 563354 3908
rect 242985 3770 243051 3773
rect 571558 3770 571564 3772
rect 242985 3768 571564 3770
rect 242985 3712 242990 3768
rect 243046 3712 571564 3768
rect 242985 3710 571564 3712
rect 242985 3707 243051 3710
rect 571558 3708 571564 3710
rect 571628 3708 571634 3772
rect 47894 3572 47900 3636
rect 47964 3634 47970 3636
rect 173157 3634 173223 3637
rect 47964 3632 173223 3634
rect 47964 3576 173162 3632
rect 173218 3576 173223 3632
rect 47964 3574 173223 3576
rect 47964 3572 47970 3574
rect 173157 3571 173223 3574
rect 203885 3634 203951 3637
rect 568614 3634 568620 3636
rect 203885 3632 568620 3634
rect 203885 3576 203890 3632
rect 203946 3576 568620 3632
rect 203885 3574 568620 3576
rect 203885 3571 203951 3574
rect 568614 3572 568620 3574
rect 568684 3572 568690 3636
rect 24209 3498 24275 3501
rect 25446 3498 25452 3500
rect 24209 3496 25452 3498
rect 24209 3440 24214 3496
rect 24270 3440 25452 3496
rect 24209 3438 25452 3440
rect 24209 3435 24275 3438
rect 25446 3436 25452 3438
rect 25516 3436 25522 3500
rect 35985 3498 36051 3501
rect 36670 3498 36676 3500
rect 35985 3496 36676 3498
rect 35985 3440 35990 3496
rect 36046 3440 36676 3496
rect 35985 3438 36676 3440
rect 35985 3435 36051 3438
rect 36670 3436 36676 3438
rect 36740 3436 36746 3500
rect 43069 3498 43135 3501
rect 43662 3498 43668 3500
rect 43069 3496 43668 3498
rect 43069 3440 43074 3496
rect 43130 3440 43668 3496
rect 43069 3438 43668 3440
rect 43069 3435 43135 3438
rect 43662 3436 43668 3438
rect 43732 3436 43738 3500
rect 50153 3498 50219 3501
rect 50838 3498 50844 3500
rect 50153 3496 50844 3498
rect 50153 3440 50158 3496
rect 50214 3440 50844 3496
rect 50153 3438 50844 3440
rect 50153 3435 50219 3438
rect 50838 3436 50844 3438
rect 50908 3436 50914 3500
rect 54886 3436 54892 3500
rect 54956 3498 54962 3500
rect 74993 3498 75059 3501
rect 54956 3496 75059 3498
rect 54956 3440 74998 3496
rect 75054 3440 75059 3496
rect 54956 3438 75059 3440
rect 54956 3436 54962 3438
rect 74993 3435 75059 3438
rect 169569 3498 169635 3501
rect 574318 3498 574324 3500
rect 169569 3496 574324 3498
rect 169569 3440 169574 3496
rect 169630 3440 574324 3496
rect 169569 3438 574324 3440
rect 169569 3435 169635 3438
rect 574318 3436 574324 3438
rect 574388 3436 574394 3500
rect 55070 3300 55076 3364
rect 55140 3362 55146 3364
rect 103329 3362 103395 3365
rect 55140 3360 103395 3362
rect 55140 3304 103334 3360
rect 103390 3304 103395 3360
rect 55140 3302 103395 3304
rect 55140 3300 55146 3302
rect 103329 3299 103395 3302
rect 126973 3362 127039 3365
rect 570086 3362 570092 3364
rect 126973 3360 570092 3362
rect 126973 3304 126978 3360
rect 127034 3304 570092 3360
rect 126973 3302 570092 3304
rect 126973 3299 127039 3302
rect 570086 3300 570092 3302
rect 570156 3300 570162 3364
rect 541566 3164 541572 3228
rect 541636 3226 541642 3228
rect 541985 3226 542051 3229
rect 541636 3224 542051 3226
rect 541636 3168 541990 3224
rect 542046 3168 542051 3224
rect 541636 3166 542051 3168
rect 541636 3164 541642 3166
rect 541985 3163 542051 3166
<< via3 >>
rect 551508 700300 551572 700364
rect 356652 686020 356716 686084
rect 28212 685884 28276 685948
rect 552244 685884 552308 685948
rect 407620 684660 407684 684724
rect 392532 683708 392596 683772
rect 393084 683572 393148 683636
rect 568620 683436 568684 683500
rect 409828 683300 409892 683364
rect 25452 683164 25516 683228
rect 403756 682620 403820 682684
rect 552060 682620 552124 682684
rect 403572 682484 403636 682548
rect 560524 682484 560588 682548
rect 395292 682348 395356 682412
rect 561628 682348 561692 682412
rect 358124 682212 358188 682276
rect 565124 682212 565188 682276
rect 399340 682076 399404 682140
rect 566964 682076 567028 682140
rect 397316 681940 397380 682004
rect 574140 681940 574204 682004
rect 356836 681804 356900 681868
rect 578556 681804 578620 681868
rect 405596 681124 405660 681188
rect 400076 680988 400140 681052
rect 575428 680988 575492 681052
rect 359412 680716 359476 680780
rect 565860 680716 565924 680780
rect 367692 680580 367756 680644
rect 409644 679764 409708 679828
rect 408356 678268 408420 678332
rect 409828 678268 409892 678332
rect 166764 676092 166828 676156
rect 155724 675004 155788 675068
rect 346900 675004 346964 675068
rect 154436 674928 154500 674932
rect 154436 674872 154486 674928
rect 154486 674872 154500 674928
rect 154436 674868 154500 674872
rect 328500 674928 328564 674932
rect 328500 674872 328550 674928
rect 328550 674872 328564 674928
rect 328500 674868 328564 674872
rect 329788 674928 329852 674932
rect 329788 674872 329802 674928
rect 329802 674872 329852 674928
rect 329788 674868 329852 674872
rect 340828 674928 340892 674932
rect 340828 674872 340878 674928
rect 340878 674872 340892 674928
rect 340828 674868 340892 674872
rect 552244 673916 552308 673980
rect 580948 669836 581012 669900
rect 557580 668476 557644 668540
rect 571380 666436 571444 666500
rect 566044 663716 566108 663780
rect 370452 657596 370516 657660
rect 402100 652156 402164 652220
rect 575612 650796 575676 650860
rect 556108 649436 556172 649500
rect 579660 646036 579724 646100
rect 401364 645356 401428 645420
rect 368980 635836 369044 635900
rect 557764 633796 557828 633860
rect 557948 630396 558012 630460
rect 404124 628356 404188 628420
rect 571564 628356 571628 628420
rect 406516 627676 406580 627740
rect 560708 626996 560772 627060
rect 405412 624276 405476 624340
rect 378732 622916 378796 622980
rect 561812 616116 561876 616180
rect 552244 614756 552308 614820
rect 556660 612036 556724 612100
rect 377260 611356 377324 611420
rect 556292 607956 556356 608020
rect 399524 607276 399588 607340
rect 387564 604420 387628 604484
rect 578740 602516 578804 602580
rect 570092 601836 570156 601900
rect 407804 601156 407868 601220
rect 556476 599116 556540 599180
rect 382780 598436 382844 598500
rect 551508 597484 551572 597548
rect 363460 593676 363524 593740
rect 550404 591568 550468 591632
rect 558868 590956 558932 591020
rect 550404 590684 550468 590748
rect 581132 590684 581196 590748
rect 84332 589520 84396 589524
rect 84332 589464 84382 589520
rect 84382 589464 84396 589520
rect 84332 589460 84396 589464
rect 407620 589052 407684 589116
rect 43852 588780 43916 588844
rect 44956 588644 45020 588708
rect 388300 588508 388364 588572
rect 53052 587828 53116 587892
rect 54156 587828 54220 587892
rect 56548 587888 56612 587892
rect 56548 587832 56598 587888
rect 56598 587832 56612 587888
rect 56548 587828 56612 587832
rect 57836 587888 57900 587892
rect 57836 587832 57886 587888
rect 57886 587832 57900 587888
rect 57836 587828 57900 587832
rect 59124 587828 59188 587892
rect 60228 587828 60292 587892
rect 62436 587828 62500 587892
rect 63540 587888 63604 587892
rect 63540 587832 63554 587888
rect 63554 587832 63604 587888
rect 63540 587828 63604 587832
rect 64276 587828 64340 587892
rect 66116 587828 66180 587892
rect 66668 587828 66732 587892
rect 68324 587828 68388 587892
rect 69612 587828 69676 587892
rect 70532 587828 70596 587892
rect 71820 587888 71884 587892
rect 71820 587832 71834 587888
rect 71834 587832 71884 587888
rect 71820 587828 71884 587832
rect 72924 587828 72988 587892
rect 74580 587888 74644 587892
rect 74580 587832 74630 587888
rect 74630 587832 74644 587888
rect 74580 587828 74644 587832
rect 77708 587828 77772 587892
rect 78812 587828 78876 587892
rect 79548 587828 79612 587892
rect 81204 587888 81268 587892
rect 81204 587832 81218 587888
rect 81218 587832 81268 587888
rect 81204 587828 81268 587832
rect 82308 587828 82372 587892
rect 83596 587828 83660 587892
rect 87092 587888 87156 587892
rect 87092 587832 87142 587888
rect 87142 587832 87156 587888
rect 87092 587828 87156 587832
rect 89484 587828 89548 587892
rect 91692 587828 91756 587892
rect 92980 587828 93044 587892
rect 94084 587828 94148 587892
rect 94452 587828 94516 587892
rect 99420 587888 99484 587892
rect 99420 587832 99470 587888
rect 99470 587832 99484 587888
rect 99420 587828 99484 587832
rect 101996 587888 102060 587892
rect 101996 587832 102010 587888
rect 102010 587832 102060 587888
rect 101996 587828 102060 587832
rect 106964 587888 107028 587892
rect 106964 587832 106978 587888
rect 106978 587832 107028 587888
rect 106964 587828 107028 587832
rect 109356 587828 109420 587892
rect 111932 587828 111996 587892
rect 114508 587828 114572 587892
rect 119476 587828 119540 587892
rect 124444 587888 124508 587892
rect 124444 587832 124458 587888
rect 124458 587832 124508 587888
rect 124444 587828 124508 587832
rect 129412 587828 129476 587892
rect 131804 587888 131868 587892
rect 131804 587832 131818 587888
rect 131818 587832 131868 587888
rect 131804 587828 131868 587832
rect 134380 587828 134444 587892
rect 136956 587828 137020 587892
rect 139348 587888 139412 587892
rect 139348 587832 139398 587888
rect 139398 587832 139412 587888
rect 139348 587828 139412 587832
rect 141924 587888 141988 587892
rect 141924 587832 141974 587888
rect 141974 587832 141988 587888
rect 141924 587828 141988 587832
rect 159404 587828 159468 587892
rect 226012 587828 226076 587892
rect 228220 587828 228284 587892
rect 230612 587828 230676 587892
rect 234292 587828 234356 587892
rect 236500 587828 236564 587892
rect 237604 587828 237668 587892
rect 238340 587828 238404 587892
rect 239996 587828 240060 587892
rect 241284 587828 241348 587892
rect 242388 587888 242452 587892
rect 242388 587832 242438 587888
rect 242438 587832 242452 587888
rect 242388 587828 242452 587832
rect 243308 587828 243372 587892
rect 244596 587828 244660 587892
rect 245884 587888 245948 587892
rect 245884 587832 245898 587888
rect 245898 587832 245948 587888
rect 245884 587828 245948 587832
rect 246988 587888 247052 587892
rect 246988 587832 247038 587888
rect 247038 587832 247052 587888
rect 246988 587828 247052 587832
rect 248092 587888 248156 587892
rect 248092 587832 248142 587888
rect 248142 587832 248156 587888
rect 248092 587828 248156 587832
rect 248460 587888 248524 587892
rect 248460 587832 248474 587888
rect 248474 587832 248524 587888
rect 248460 587828 248524 587832
rect 249564 587828 249628 587892
rect 252876 587828 252940 587892
rect 253980 587888 254044 587892
rect 253980 587832 253994 587888
rect 253994 587832 254044 587888
rect 253980 587828 254044 587832
rect 256004 587828 256068 587892
rect 256372 587828 256436 587892
rect 257660 587828 257724 587892
rect 259868 587828 259932 587892
rect 260972 587888 261036 587892
rect 260972 587832 261022 587888
rect 261022 587832 261036 587888
rect 260972 587828 261036 587832
rect 261156 587828 261220 587892
rect 262260 587888 262324 587892
rect 262260 587832 262274 587888
rect 262274 587832 262324 587888
rect 262260 587828 262324 587832
rect 263548 587828 263612 587892
rect 265756 587828 265820 587892
rect 268516 587828 268580 587892
rect 269252 587828 269316 587892
rect 270908 587828 270972 587892
rect 273484 587888 273548 587892
rect 273484 587832 273534 587888
rect 273534 587832 273548 587888
rect 273484 587828 273548 587832
rect 275876 587828 275940 587892
rect 281028 587888 281092 587892
rect 281028 587832 281078 587888
rect 281078 587832 281092 587888
rect 281028 587828 281092 587832
rect 283420 587828 283484 587892
rect 285996 587828 286060 587892
rect 288388 587888 288452 587892
rect 288388 587832 288438 587888
rect 288438 587832 288452 587888
rect 288388 587828 288452 587832
rect 290964 587888 291028 587892
rect 290964 587832 291014 587888
rect 291014 587832 291028 587888
rect 290964 587828 291028 587832
rect 298508 587828 298572 587892
rect 300900 587888 300964 587892
rect 300900 587832 300914 587888
rect 300914 587832 300964 587888
rect 300900 587828 300964 587832
rect 303476 587828 303540 587892
rect 305868 587828 305932 587892
rect 308444 587888 308508 587892
rect 308444 587832 308494 587888
rect 308494 587832 308508 587888
rect 308444 587828 308508 587832
rect 310836 587828 310900 587892
rect 313412 587828 313476 587892
rect 315988 587888 316052 587892
rect 315988 587832 316038 587888
rect 316038 587832 316052 587888
rect 315988 587828 316052 587832
rect 333468 587828 333532 587892
rect 55628 587692 55692 587756
rect 61516 587692 61580 587756
rect 64644 587692 64708 587756
rect 69428 587692 69492 587756
rect 72188 587692 72252 587756
rect 75500 587692 75564 587756
rect 77156 587752 77220 587756
rect 77156 587696 77206 587752
rect 77206 587696 77220 587752
rect 77156 587692 77220 587696
rect 79916 587692 79980 587756
rect 81940 587752 82004 587756
rect 81940 587696 81954 587752
rect 81954 587696 82004 587752
rect 81940 587692 82004 587696
rect 88196 587692 88260 587756
rect 95188 587752 95252 587756
rect 95188 587696 95238 587752
rect 95238 587696 95252 587752
rect 95188 587692 95252 587696
rect 127020 587692 127084 587756
rect 235396 587692 235460 587756
rect 240732 587752 240796 587756
rect 240732 587696 240782 587752
rect 240782 587696 240796 587752
rect 240732 587692 240796 587696
rect 246068 587692 246132 587756
rect 251036 587692 251100 587756
rect 253428 587692 253492 587756
rect 264468 587752 264532 587756
rect 264468 587696 264482 587752
rect 264482 587696 264532 587752
rect 264468 587692 264532 587696
rect 265940 587692 266004 587756
rect 74028 587556 74092 587620
rect 227116 587420 227180 587484
rect 229508 587284 229572 587348
rect 250668 587284 250732 587348
rect 348372 587284 348436 587348
rect 255268 587148 255332 587212
rect 238524 586740 238588 586804
rect 257844 586740 257908 586804
rect 48452 586332 48516 586396
rect 51948 586604 52012 586668
rect 67220 586604 67284 586668
rect 76604 586604 76668 586668
rect 86908 586604 86972 586668
rect 84148 586468 84212 586532
rect 85620 586468 85684 586532
rect 89300 586604 89364 586668
rect 90404 586604 90468 586668
rect 92060 586604 92124 586668
rect 96844 586604 96908 586668
rect 103468 586468 103532 586532
rect 116900 586604 116964 586668
rect 121868 586604 121932 586668
rect 159220 586604 159284 586668
rect 231716 586604 231780 586668
rect 233188 586604 233252 586668
rect 243676 586604 243740 586668
rect 251772 586604 251836 586668
rect 258580 586468 258644 586532
rect 263364 586604 263428 586668
rect 267044 586604 267108 586668
rect 267964 586468 268028 586532
rect 277348 586468 277412 586532
rect 293540 586604 293604 586668
rect 295932 586604 295996 586668
rect 333100 586604 333164 586668
rect 407804 584292 407868 584356
rect 46980 583068 47044 583132
rect 346348 582932 346412 582996
rect 570092 582116 570156 582180
rect 351132 581572 351196 581636
rect 391244 581436 391308 581500
rect 387012 580756 387076 580820
rect 567332 580756 567396 580820
rect 563100 579396 563164 579460
rect 349108 578852 349172 578916
rect 371740 578716 371804 578780
rect 46796 577492 46860 577556
rect 561996 576676 562060 576740
rect 347820 575996 347884 576060
rect 46612 574636 46676 574700
rect 559052 574092 559116 574156
rect 350948 571916 351012 571980
rect 47348 570692 47412 570756
rect 348004 570556 348068 570620
rect 47164 569196 47228 569260
rect 353524 568788 353588 568852
rect 396580 568652 396644 568716
rect 46244 567836 46308 567900
rect 347636 567428 347700 567492
rect 391060 567292 391124 567356
rect 398604 567156 398668 567220
rect 553348 566476 553412 566540
rect 363644 566340 363708 566404
rect 389772 566204 389836 566268
rect 359596 566068 359660 566132
rect 351868 565932 351932 565996
rect 352052 565796 352116 565860
rect 373212 565796 373276 565860
rect 563284 565116 563348 565180
rect 356100 564844 356164 564908
rect 46428 563620 46492 563684
rect 349292 563484 349356 563548
rect 381492 563348 381556 563412
rect 391428 563076 391492 563140
rect 39620 562668 39684 562732
rect 48452 562532 48516 562596
rect 48636 562396 48700 562460
rect 44772 562260 44836 562324
rect 364380 562124 364444 562188
rect 27476 561852 27540 561916
rect 360148 561852 360212 561916
rect 360332 561716 360396 561780
rect 41276 561172 41340 561236
rect 395476 560900 395540 560964
rect 400812 560492 400876 560556
rect 347636 560356 347700 560420
rect 346348 560084 346412 560148
rect 347268 560084 347332 560148
rect 48084 558724 48148 558788
rect 347636 558180 347700 558244
rect 39252 558044 39316 558108
rect 48268 558044 48332 558108
rect 389956 557636 390020 557700
rect 347636 557364 347700 557428
rect 348556 557364 348620 557428
rect 347636 557228 347700 557292
rect 558132 556276 558196 556340
rect 48268 556140 48332 556204
rect 347636 556140 347700 556204
rect 349476 556140 349540 556204
rect 566228 552196 566292 552260
rect 566412 551516 566476 551580
rect 352052 548932 352116 548996
rect 45324 548252 45388 548316
rect 574324 544716 574388 544780
rect 38516 534108 38580 534172
rect 41828 533292 41892 533356
rect 407620 533836 407684 533900
rect 560892 531796 560956 531860
rect 44036 530708 44100 530772
rect 37044 527308 37108 527372
rect 36860 527172 36924 527236
rect 378916 527036 378980 527100
rect 348004 523500 348068 523564
rect 348924 522956 348988 523020
rect 35756 520372 35820 520436
rect 350580 520236 350644 520300
rect 367140 518876 367204 518940
rect 42012 515068 42076 515132
rect 30972 514796 31036 514860
rect 34284 514796 34348 514860
rect 395660 510716 395724 510780
rect 41276 510444 41340 510508
rect 350764 507860 350828 507924
rect 374500 502420 374564 502484
rect 32996 499700 33060 499764
rect 41276 498748 41340 498812
rect 385540 497116 385604 497180
rect 550772 497116 550836 497180
rect 554820 494396 554884 494460
rect 553532 491676 553596 491740
rect 41092 490588 41156 490652
rect 352052 490588 352116 490652
rect 407804 488956 407868 489020
rect 45140 486508 45204 486572
rect 37596 482972 37660 483036
rect 349108 482972 349172 483036
rect 392716 480116 392780 480180
rect 39804 476308 39868 476372
rect 43852 476172 43916 476236
rect 408540 476172 408604 476236
rect 565308 472636 565372 472700
rect 353708 472228 353772 472292
rect 35572 470868 35636 470932
rect 41644 466516 41708 466580
rect 408356 466516 408420 466580
rect 40908 465156 40972 465220
rect 349108 463932 349172 463996
rect 355180 461756 355244 461820
rect 36676 458220 36740 458284
rect 43852 456860 43916 456924
rect 364564 456996 364628 457060
rect 348372 456860 348436 456924
rect 348372 456724 348436 456788
rect 377444 453596 377508 453660
rect 39436 450468 39500 450532
rect 561076 450196 561140 450260
rect 43668 449108 43732 449172
rect 551508 441356 551572 441420
rect 550220 440676 550284 440740
rect 40724 438908 40788 438972
rect 349660 434828 349724 434892
rect 349292 433196 349356 433260
rect 47532 428504 47596 428568
rect 46244 412932 46308 412996
rect 347820 411164 347884 411228
rect 567516 410756 567580 410820
rect 555004 404636 555068 404700
rect 46244 402052 46308 402116
rect 32812 400828 32876 400892
rect 565492 400284 565556 400348
rect 349476 385732 349540 385796
rect 44956 383012 45020 383076
rect 407988 378116 408052 378180
rect 349476 358804 349540 358868
rect 348740 341396 348804 341460
rect 559236 336636 559300 336700
rect 360700 325756 360764 325820
rect 44956 317324 45020 317388
rect 409460 316916 409524 316980
rect 553716 315556 553780 315620
rect 43484 313244 43548 313308
rect 44772 313244 44836 313308
rect 387748 311884 387812 311948
rect 406148 306036 406212 306100
rect 354444 304948 354508 305012
rect 372660 302228 372724 302292
rect 348556 299372 348620 299436
rect 44956 285228 45020 285292
rect 351132 278292 351196 278356
rect 409644 277476 409708 277540
rect 44772 275980 44836 276044
rect 31524 273668 31588 273732
rect 350948 268092 351012 268156
rect 35388 267956 35452 268020
rect 44588 264828 44652 264892
rect 43484 264556 43548 264620
rect 409092 262924 409156 262988
rect 36492 262244 36556 262308
rect 406332 262108 406396 262172
rect 44772 259524 44836 259588
rect 44956 258164 45020 258228
rect 46060 252452 46124 252516
rect 46428 251772 46492 251836
rect 404860 251772 404924 251836
rect 46428 247556 46492 247620
rect 46612 247012 46676 247076
rect 563468 246876 563532 246940
rect 350948 245516 351012 245580
rect 44588 245380 44652 245444
rect 44772 244292 44836 244356
rect 46612 244352 46676 244356
rect 46612 244296 46662 244352
rect 46662 244296 46676 244352
rect 46612 244292 46676 244296
rect 46796 244292 46860 244356
rect 396212 243476 396276 243540
rect 409828 242796 409892 242860
rect 410012 242524 410076 242588
rect 47716 241436 47780 241500
rect 47348 240892 47412 240956
rect 391428 240484 391492 240548
rect 388300 238308 388364 238372
rect 393084 236676 393148 236740
rect 547092 236676 547156 236740
rect 405596 235724 405660 235788
rect 548012 235724 548076 235788
rect 400076 235588 400140 235652
rect 544332 235588 544396 235652
rect 387564 235452 387628 235516
rect 540284 235452 540348 235516
rect 541572 235316 541636 235380
rect 556844 235316 556908 235380
rect 406148 235180 406212 235244
rect 556660 234636 556724 234700
rect 538812 234228 538876 234292
rect 405412 234092 405476 234156
rect 404124 233956 404188 234020
rect 549484 233956 549548 234020
rect 348924 233820 348988 233884
rect 538996 232460 539060 232524
rect 539180 231644 539244 231708
rect 402100 231508 402164 231572
rect 397316 231236 397380 231300
rect 401364 231100 401428 231164
rect 47716 226400 47780 226404
rect 47716 226344 47766 226400
rect 47766 226344 47780 226400
rect 47716 226340 47780 226344
rect 47716 222124 47780 222188
rect 39252 220764 39316 220828
rect 44772 220764 44836 220828
rect 47164 220492 47228 220556
rect 48084 220220 48148 220284
rect 44588 220084 44652 220148
rect 39252 218044 39316 218108
rect 46980 210292 47044 210356
rect 542676 210292 542740 210356
rect 406516 206212 406580 206276
rect 39068 205668 39132 205732
rect 39252 205668 39316 205732
rect 39620 204852 39684 204916
rect 47532 204444 47596 204508
rect 47900 204444 47964 204508
rect 47532 204308 47596 204372
rect 39252 203492 39316 203556
rect 44588 201588 44652 201652
rect 48268 201588 48332 201652
rect 44772 201452 44836 201516
rect 347820 201044 347884 201108
rect 48268 200500 48332 200564
rect 347636 200500 347700 200564
rect 41828 200016 41892 200020
rect 41828 199960 41878 200016
rect 41878 199960 41892 200016
rect 41828 199956 41892 199960
rect 49004 199548 49068 199612
rect 347452 199548 347516 199612
rect 350948 198868 351012 198932
rect 368980 198324 369044 198388
rect 356836 198188 356900 198252
rect 359412 198052 359476 198116
rect 47532 197916 47596 197980
rect 367692 196692 367756 196756
rect 47900 196556 47964 196620
rect 36676 195876 36740 195940
rect 403756 195740 403820 195804
rect 349108 195468 349172 195532
rect 46244 195196 46308 195260
rect 30972 194516 31036 194580
rect 395660 194380 395724 194444
rect 48268 193972 48332 194036
rect 53052 193836 53116 193900
rect 49004 192884 49068 192948
rect 356100 192884 356164 192948
rect 374500 192748 374564 192812
rect 45140 192612 45204 192676
rect 555004 192476 555068 192540
rect 347452 191660 347516 191724
rect 347084 191524 347148 191588
rect 55076 191252 55140 191316
rect 57836 191116 57900 191180
rect 550220 191116 550284 191180
rect 551508 190980 551572 191044
rect 350580 190300 350644 190364
rect 61332 190164 61396 190228
rect 50476 190028 50540 190092
rect 377260 189892 377324 189956
rect 53604 189756 53668 189820
rect 399524 189756 399588 189820
rect 55444 189620 55508 189684
rect 407620 189620 407684 189684
rect 378916 188804 378980 188868
rect 47900 188668 47964 188732
rect 385540 188668 385604 188732
rect 43668 188532 43732 188596
rect 55628 188396 55692 188460
rect 552244 188396 552308 188460
rect 36676 188260 36740 188324
rect 61516 187580 61580 187644
rect 58572 187444 58636 187508
rect 59124 187308 59188 187372
rect 54708 187172 54772 187236
rect 396212 187036 396276 187100
rect 539548 186900 539612 186964
rect 49556 185812 49620 185876
rect 360332 185812 360396 185876
rect 50660 185676 50724 185740
rect 36860 185540 36924 185604
rect 60596 184588 60660 184652
rect 353524 184588 353588 184652
rect 353708 184452 353772 184516
rect 407988 184316 408052 184380
rect 37044 184180 37108 184244
rect 54892 182820 54956 182884
rect 387012 182820 387076 182884
rect 348372 181596 348436 181660
rect 348740 181460 348804 181524
rect 50292 181324 50356 181388
rect 367140 181324 367204 181388
rect 395292 180644 395356 180708
rect 41092 180508 41156 180572
rect 49372 180372 49436 180436
rect 382780 180372 382844 180436
rect 391244 180236 391308 180300
rect 34284 180100 34348 180164
rect 539732 179964 539796 180028
rect 350764 179828 350828 179892
rect 364564 178740 364628 178804
rect 45876 178604 45940 178668
rect 61700 177788 61764 177852
rect 349660 177652 349724 177716
rect 378732 177516 378796 177580
rect 49188 177380 49252 177444
rect 392532 177380 392596 177444
rect 541020 177244 541084 177308
rect 60412 174932 60476 174996
rect 52316 174796 52380 174860
rect 46612 174660 46676 174724
rect 542676 174660 542740 174724
rect 41092 174524 41156 174588
rect 41276 173300 41340 173364
rect 50844 173164 50908 173228
rect 346900 172348 346964 172412
rect 53420 172212 53484 172276
rect 377444 172212 377508 172276
rect 41276 172076 41340 172140
rect 373212 172076 373276 172140
rect 46244 171940 46308 172004
rect 387748 171940 387812 172004
rect 389956 171804 390020 171868
rect 46060 171668 46124 171732
rect 543964 171668 544028 171732
rect 43668 170444 43732 170508
rect 392716 170444 392780 170508
rect 563284 170308 563348 170372
rect 41644 168948 41708 169012
rect 39436 167724 39500 167788
rect 559052 167588 559116 167652
rect 54524 166500 54588 166564
rect 363460 166500 363524 166564
rect 545436 166500 545500 166564
rect 53236 166364 53300 166428
rect 562180 166364 562244 166428
rect 40724 166228 40788 166292
rect 563284 166228 563348 166292
rect 399340 163644 399404 163708
rect 389772 163508 389836 163572
rect 358124 163372 358188 163436
rect 541204 163372 541268 163436
rect 403572 162012 403636 162076
rect 549852 161196 549916 161260
rect 548196 161060 548260 161124
rect 57652 160924 57716 160988
rect 371740 160924 371804 160988
rect 391060 160924 391124 160988
rect 552244 160924 552308 160988
rect 547460 160788 547524 160852
rect 552428 160652 552492 160716
rect 355180 159564 355244 159628
rect 543780 159564 543844 159628
rect 57468 159428 57532 159492
rect 545804 159428 545868 159492
rect 563100 159292 563164 159356
rect 539364 158612 539428 158676
rect 352052 158476 352116 158540
rect 549668 158476 549732 158540
rect 58940 158340 59004 158404
rect 46428 158204 46492 158268
rect 544148 158204 544212 158268
rect 398604 157252 398668 157316
rect 552612 157252 552676 157316
rect 409092 157116 409156 157180
rect 40908 156980 40972 157044
rect 409460 156980 409524 157044
rect 35572 156844 35636 156908
rect 539916 156708 539980 156772
rect 563100 156572 563164 156636
rect 46428 155952 46492 155956
rect 46428 155896 46442 155952
rect 46442 155896 46492 155952
rect 46428 155892 46492 155896
rect 351868 155756 351932 155820
rect 60044 155620 60108 155684
rect 543412 155620 543476 155684
rect 364380 155484 364444 155548
rect 360148 155348 360212 155412
rect 545252 155348 545316 155412
rect 58756 155212 58820 155276
rect 407804 155212 407868 155276
rect 406332 154260 406396 154324
rect 547828 154260 547892 154324
rect 542860 154124 542924 154188
rect 360700 153988 360764 154052
rect 363644 153988 363708 154052
rect 549300 153988 549364 154052
rect 545068 153852 545132 153916
rect 551508 153716 551572 153780
rect 396580 153036 396644 153100
rect 48820 152900 48884 152964
rect 356652 152900 356716 152964
rect 400812 152900 400876 152964
rect 47716 152764 47780 152828
rect 395476 152764 395540 152828
rect 408540 152628 408604 152692
rect 409828 152628 409892 152692
rect 354444 152492 354508 152556
rect 381492 152492 381556 152556
rect 553900 152492 553964 152556
rect 370452 152356 370516 152420
rect 541388 151676 541452 151740
rect 410196 151404 410260 151468
rect 559052 151268 559116 151332
rect 349476 151132 349540 151196
rect 359596 151132 359660 151196
rect 555004 151132 555068 151196
rect 57284 150996 57348 151060
rect 372660 150996 372724 151060
rect 404860 150996 404924 151060
rect 539180 150452 539244 150516
rect 540100 150452 540164 150516
rect 60228 150044 60292 150108
rect 61332 150044 61396 150108
rect 61516 149908 61580 149972
rect 547276 149908 547340 149972
rect 49004 149092 49068 149156
rect 563652 149092 563716 149156
rect 51028 148684 51092 148748
rect 60228 148684 60292 148748
rect 540100 148548 540164 148612
rect 47716 147732 47780 147796
rect 51028 147460 51092 147524
rect 52132 147460 52196 147524
rect 539364 147324 539428 147388
rect 540284 146916 540348 146980
rect 539364 146780 539428 146844
rect 60044 146508 60108 146572
rect 539364 146508 539428 146572
rect 544148 146236 544212 146300
rect 542860 146100 542924 146164
rect 544700 146100 544764 146164
rect 539364 145420 539428 145484
rect 59308 144876 59372 144940
rect 540836 144740 540900 144804
rect 58020 143516 58084 143580
rect 58756 143516 58820 143580
rect 52316 142292 52380 142356
rect 52316 142020 52380 142084
rect 59124 142020 59188 142084
rect 59492 142020 59556 142084
rect 539364 141748 539428 141812
rect 544332 139572 544396 139636
rect 545620 139572 545684 139636
rect 544516 139436 544580 139500
rect 545436 139436 545500 139500
rect 60596 139164 60660 139228
rect 547276 138620 547340 138684
rect 51028 138076 51092 138140
rect 52132 138076 52196 138140
rect 544700 138076 544764 138140
rect 547276 138076 547340 138140
rect 544700 137940 544764 138004
rect 59308 137260 59372 137324
rect 563652 137260 563716 137324
rect 59124 136580 59188 136644
rect 544332 136580 544396 136644
rect 544516 136640 544580 136644
rect 544516 136584 544566 136640
rect 544566 136584 544580 136640
rect 544516 136580 544580 136584
rect 564020 136580 564084 136644
rect 58572 135900 58636 135964
rect 41092 135220 41156 135284
rect 541388 133180 541452 133244
rect 547276 132772 547340 132836
rect 547644 132772 547708 132836
rect 541940 131276 542004 131340
rect 544700 131276 544764 131340
rect 544516 131200 544580 131204
rect 544516 131144 544566 131200
rect 544566 131144 544580 131200
rect 544516 131140 544580 131144
rect 541572 130460 541636 130524
rect 542124 130324 542188 130388
rect 548012 130324 548076 130388
rect 540652 129644 540716 129708
rect 548380 129508 548444 129572
rect 543044 128420 543108 128484
rect 544148 127604 544212 127668
rect 544332 127604 544396 127668
rect 545436 127604 545500 127668
rect 545620 127060 545684 127124
rect 545620 126924 545684 126988
rect 547644 126924 547708 126988
rect 545804 126788 545868 126852
rect 547276 126788 547340 126852
rect 540836 126244 540900 126308
rect 59492 125428 59556 125492
rect 58572 124748 58636 124812
rect 51028 124068 51092 124132
rect 52132 124068 52196 124132
rect 58940 124204 59004 124268
rect 544516 124128 544580 124132
rect 544516 124072 544566 124128
rect 544566 124072 544580 124128
rect 544516 124068 544580 124072
rect 544332 123932 544396 123996
rect 46428 123524 46492 123588
rect 58756 123524 58820 123588
rect 46244 123388 46308 123452
rect 59860 123388 59924 123452
rect 59676 122028 59740 122092
rect 59308 120184 59372 120188
rect 59308 120128 59322 120184
rect 59322 120128 59372 120184
rect 59308 120124 59372 120128
rect 58020 117948 58084 118012
rect 544148 117948 544212 118012
rect 544516 117328 544580 117332
rect 544516 117272 544566 117328
rect 544566 117272 544580 117328
rect 544516 117268 544580 117272
rect 541204 115908 541268 115972
rect 541756 115968 541820 115972
rect 541756 115912 541806 115968
rect 541806 115912 541820 115968
rect 541756 115908 541820 115912
rect 544516 114412 544580 114476
rect 547460 114276 547524 114340
rect 549484 113188 549548 113252
rect 542492 113052 542556 113116
rect 59308 111828 59372 111892
rect 542860 110876 542924 110940
rect 541940 110604 542004 110668
rect 547460 110604 547524 110668
rect 544148 110468 544212 110532
rect 540652 110196 540716 110260
rect 541204 110196 541268 110260
rect 541756 107476 541820 107540
rect 542492 107476 542556 107540
rect 541572 105436 541636 105500
rect 543412 104212 543476 104276
rect 541388 102308 541452 102372
rect 543044 102308 543108 102372
rect 542124 102172 542188 102236
rect 59308 99996 59372 100060
rect 541204 99452 541268 99516
rect 564020 99452 564084 99516
rect 540100 95100 540164 95164
rect 543228 88980 543292 89044
rect 553900 88980 553964 89044
rect 542308 87892 542372 87956
rect 543044 86124 543108 86188
rect 548380 85580 548444 85644
rect 548196 84628 548260 84692
rect 549852 83268 549916 83332
rect 541204 82860 541268 82924
rect 549852 81500 549916 81564
rect 57284 74972 57348 75036
rect 549668 72252 549732 72316
rect 541020 70892 541084 70956
rect 543964 68852 544028 68916
rect 57836 64772 57900 64836
rect 57468 59332 57532 59396
rect 55444 57972 55508 58036
rect 563100 55252 563164 55316
rect 552612 51036 552676 51100
rect 41276 48588 41340 48652
rect 539732 46820 539796 46884
rect 53052 44236 53116 44300
rect 551508 41652 551572 41716
rect 539916 38524 539980 38588
rect 552428 37300 552492 37364
rect 55628 35532 55692 35596
rect 539548 35260 539612 35324
rect 57652 34852 57716 34916
rect 45876 30908 45940 30972
rect 539364 31044 539428 31108
rect 540284 30908 540348 30972
rect 555004 30908 555068 30972
rect 59124 30772 59188 30836
rect 552244 30364 552308 30428
rect 59308 29820 59372 29884
rect 50292 29548 50356 29612
rect 545252 29548 545316 29612
rect 52132 29412 52196 29476
rect 547644 29412 547708 29476
rect 561812 29276 561876 29340
rect 561996 29140 562060 29204
rect 575612 29140 575676 29204
rect 543780 29004 543844 29068
rect 59860 28868 59924 28932
rect 39804 28732 39868 28796
rect 541204 28732 541268 28796
rect 44036 28460 44100 28524
rect 560524 28460 560588 28524
rect 50476 28324 50540 28388
rect 58756 28188 58820 28252
rect 552060 28188 552124 28252
rect 45324 28052 45388 28116
rect 49004 27508 49068 27572
rect 549300 27508 549364 27572
rect 561076 27372 561140 27436
rect 44956 27236 45020 27300
rect 566044 27236 566108 27300
rect 578556 27100 578620 27164
rect 43852 26964 43916 27028
rect 545068 26964 545132 27028
rect 561628 26828 561692 26892
rect 42012 26692 42076 26756
rect 545620 26692 545684 26756
rect 36492 26556 36556 26620
rect 567148 26148 567212 26212
rect 32996 26012 33060 26076
rect 38516 25876 38580 25940
rect 37596 25740 37660 25804
rect 60044 25604 60108 25668
rect 566412 25604 566476 25668
rect 53236 25468 53300 25532
rect 54524 25468 54588 25532
rect 53420 25332 53484 25396
rect 538812 25332 538876 25396
rect 32812 25196 32876 25260
rect 547276 24788 547340 24852
rect 54708 24516 54772 24580
rect 556660 24516 556724 24580
rect 52316 24380 52380 24444
rect 565308 24380 565372 24444
rect 567332 24244 567396 24308
rect 553348 24108 553412 24172
rect 39068 23972 39132 24036
rect 566228 23972 566292 24036
rect 53604 23020 53668 23084
rect 581132 23020 581196 23084
rect 548380 22884 548444 22948
rect 579660 22748 579724 22812
rect 48084 22612 48148 22676
rect 547092 22612 547156 22676
rect 578740 22476 578804 22540
rect 35756 21932 35820 21996
rect 540284 21932 540348 21996
rect 49556 21796 49620 21860
rect 565492 21796 565556 21860
rect 571380 21660 571444 21724
rect 565124 21524 565188 21588
rect 50660 21388 50724 21452
rect 567516 21388 567580 21452
rect 49188 21252 49252 21316
rect 570092 21252 570156 21316
rect 558868 21116 558932 21180
rect 31524 20572 31588 20636
rect 27476 20164 27540 20228
rect 543228 20164 543292 20228
rect 49372 19892 49436 19956
rect 554820 19892 554884 19956
rect 28212 19348 28276 19412
rect 47716 19076 47780 19140
rect 544332 19076 544396 19140
rect 58572 18940 58636 19004
rect 559052 18940 559116 19004
rect 44772 18804 44836 18868
rect 558132 18804 558196 18868
rect 574140 18668 574204 18732
rect 553716 18532 553780 18596
rect 580948 17716 581012 17780
rect 542676 17580 542740 17644
rect 560708 17580 560772 17644
rect 575428 17444 575492 17508
rect 557580 17308 557644 17372
rect 556476 17172 556540 17236
rect 542860 17036 542924 17100
rect 563468 16900 563532 16964
rect 39252 16492 39316 16556
rect 547460 16492 547524 16556
rect 544148 16356 544212 16420
rect 550588 15948 550652 16012
rect 543044 15132 543108 15196
rect 541388 14996 541452 15060
rect 548012 14860 548076 14924
rect 549852 14452 549916 14516
rect 540100 13636 540164 13700
rect 545436 12956 545500 13020
rect 557764 11732 557828 11796
rect 560892 11596 560956 11660
rect 556292 10372 556356 10436
rect 35388 10236 35452 10300
rect 557948 7652 558012 7716
rect 556108 7516 556172 7580
rect 562180 6292 562244 6356
rect 553532 6156 553596 6220
rect 559236 4796 559300 4860
rect 565860 3980 565924 4044
rect 563284 3844 563348 3908
rect 571564 3708 571628 3772
rect 47900 3572 47964 3636
rect 568620 3572 568684 3636
rect 25452 3436 25516 3500
rect 36676 3436 36740 3500
rect 43668 3436 43732 3500
rect 50844 3436 50908 3500
rect 54892 3436 54956 3500
rect 574324 3436 574388 3500
rect 55076 3300 55140 3364
rect 570092 3300 570156 3364
rect 541572 3164 541636 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28211 685948 28277 685949
rect 28211 685884 28212 685948
rect 28276 685884 28277 685948
rect 28211 685883 28277 685884
rect 25451 683228 25517 683229
rect 25451 683164 25452 683228
rect 25516 683164 25517 683228
rect 25451 683163 25517 683164
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 25454 3501 25514 683163
rect 27475 561916 27541 561917
rect 27475 561852 27476 561916
rect 27540 561852 27541 561916
rect 27475 561851 27541 561852
rect 27478 20229 27538 561851
rect 27475 20228 27541 20229
rect 27475 20164 27476 20228
rect 27540 20164 27541 20228
rect 27475 20163 27541 20164
rect 28214 19413 28274 685883
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 675308 38414 686898
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 675308 42914 691398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 675308 47414 695898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 675308 51914 700398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 675308 65414 677898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 675308 69914 682398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 675308 74414 686898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 675308 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 675308 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 675308 87914 700398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 675308 101414 677898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 675308 105914 682398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 675308 110414 686898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 675308 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 675308 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 675308 123914 700398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 675308 137414 677898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 675308 141914 682398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 675308 146414 686898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 675308 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 675308 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 675308 159914 700398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 166763 676156 166829 676157
rect 166763 676092 166764 676156
rect 166828 676092 166829 676156
rect 166763 676091 166829 676092
rect 155723 675068 155789 675069
rect 155723 675004 155724 675068
rect 155788 675004 155789 675068
rect 155723 675003 155789 675004
rect 154435 674932 154501 674933
rect 154435 674868 154436 674932
rect 154500 674868 154501 674932
rect 154435 674867 154501 674868
rect 154438 673470 154498 674867
rect 155726 673470 155786 675003
rect 154438 673410 154524 673470
rect 154464 673202 154524 673410
rect 155688 673410 155786 673470
rect 166766 673470 166826 676091
rect 172794 675308 173414 677898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 166766 673410 166900 673470
rect 155688 673202 155748 673410
rect 166840 673202 166900 673410
rect 36272 655954 36620 655986
rect 36272 655718 36328 655954
rect 36564 655718 36620 655954
rect 36272 655634 36620 655718
rect 36272 655398 36328 655634
rect 36564 655398 36620 655634
rect 36272 655366 36620 655398
rect 172000 655954 172348 655986
rect 172000 655718 172056 655954
rect 172292 655718 172348 655954
rect 172000 655634 172348 655718
rect 172000 655398 172056 655634
rect 172292 655398 172348 655634
rect 172000 655366 172348 655398
rect 36952 651454 37300 651486
rect 36952 651218 37008 651454
rect 37244 651218 37300 651454
rect 36952 651134 37300 651218
rect 36952 650898 37008 651134
rect 37244 650898 37300 651134
rect 36952 650866 37300 650898
rect 171320 651454 171668 651486
rect 171320 651218 171376 651454
rect 171612 651218 171668 651454
rect 171320 651134 171668 651218
rect 171320 650898 171376 651134
rect 171612 650898 171668 651134
rect 171320 650866 171668 650898
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 36272 619954 36620 619986
rect 36272 619718 36328 619954
rect 36564 619718 36620 619954
rect 36272 619634 36620 619718
rect 36272 619398 36328 619634
rect 36564 619398 36620 619634
rect 36272 619366 36620 619398
rect 172000 619954 172348 619986
rect 172000 619718 172056 619954
rect 172292 619718 172348 619954
rect 172000 619634 172348 619718
rect 172000 619398 172056 619634
rect 172292 619398 172348 619634
rect 172000 619366 172348 619398
rect 36952 615454 37300 615486
rect 36952 615218 37008 615454
rect 37244 615218 37300 615454
rect 36952 615134 37300 615218
rect 36952 614898 37008 615134
rect 37244 614898 37300 615134
rect 36952 614866 37300 614898
rect 171320 615454 171668 615486
rect 171320 615218 171376 615454
rect 171612 615218 171668 615454
rect 171320 615134 171668 615218
rect 171320 614898 171376 615134
rect 171612 614898 171668 615134
rect 171320 614866 171668 614898
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 52056 589930 52116 590106
rect 53144 589930 53204 590106
rect 54232 589930 54292 590106
rect 51950 589870 52116 589930
rect 53054 589870 53204 589930
rect 54158 589870 54292 589930
rect 55592 589930 55652 590106
rect 56544 589930 56604 590106
rect 57768 589930 57828 590106
rect 59128 589930 59188 590106
rect 55592 589870 55690 589930
rect 56544 589870 56610 589930
rect 57768 589870 57898 589930
rect 43851 588844 43917 588845
rect 43851 588780 43852 588844
rect 43916 588780 43917 588844
rect 43851 588779 43917 588780
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 30971 514860 31037 514861
rect 30971 514796 30972 514860
rect 31036 514796 31037 514860
rect 30971 514795 31037 514796
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 30974 194581 31034 514795
rect 33294 502954 33914 538398
rect 37794 579454 38414 588000
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 42294 583954 42914 588000
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 39619 562732 39685 562733
rect 39619 562668 39620 562732
rect 39684 562668 39685 562732
rect 39619 562667 39685 562668
rect 39251 558108 39317 558109
rect 39251 558044 39252 558108
rect 39316 558044 39317 558108
rect 39251 558043 39317 558044
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37043 527372 37109 527373
rect 37043 527308 37044 527372
rect 37108 527308 37109 527372
rect 37043 527307 37109 527308
rect 36859 527236 36925 527237
rect 36859 527172 36860 527236
rect 36924 527172 36925 527236
rect 36859 527171 36925 527172
rect 35755 520436 35821 520437
rect 35755 520372 35756 520436
rect 35820 520372 35821 520436
rect 35755 520371 35821 520372
rect 34283 514860 34349 514861
rect 34283 514796 34284 514860
rect 34348 514796 34349 514860
rect 34283 514795 34349 514796
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 32995 499764 33061 499765
rect 32995 499700 32996 499764
rect 33060 499700 33061 499764
rect 32995 499699 33061 499700
rect 32811 400892 32877 400893
rect 32811 400828 32812 400892
rect 32876 400828 32877 400892
rect 32811 400827 32877 400828
rect 31523 273732 31589 273733
rect 31523 273668 31524 273732
rect 31588 273668 31589 273732
rect 31523 273667 31589 273668
rect 30971 194580 31037 194581
rect 30971 194516 30972 194580
rect 31036 194516 31037 194580
rect 30971 194515 31037 194516
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28211 19412 28277 19413
rect 28211 19348 28212 19412
rect 28276 19348 28277 19412
rect 28211 19347 28277 19348
rect 25451 3500 25517 3501
rect 25451 3436 25452 3500
rect 25516 3436 25517 3500
rect 25451 3435 25517 3436
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 -6106 29414 29898
rect 31526 20637 31586 273667
rect 32814 25261 32874 400827
rect 32998 26077 33058 499699
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 34286 180165 34346 514795
rect 35571 470932 35637 470933
rect 35571 470868 35572 470932
rect 35636 470868 35637 470932
rect 35571 470867 35637 470868
rect 35387 268020 35453 268021
rect 35387 267956 35388 268020
rect 35452 267956 35453 268020
rect 35387 267955 35453 267956
rect 34283 180164 34349 180165
rect 34283 180100 34284 180164
rect 34348 180100 34349 180164
rect 34283 180099 34349 180100
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 32995 26076 33061 26077
rect 32995 26012 32996 26076
rect 33060 26012 33061 26076
rect 32995 26011 33061 26012
rect 32811 25260 32877 25261
rect 32811 25196 32812 25260
rect 32876 25196 32877 25260
rect 32811 25195 32877 25196
rect 31523 20636 31589 20637
rect 31523 20572 31524 20636
rect 31588 20572 31589 20636
rect 31523 20571 31589 20572
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 -7066 33914 34398
rect 35390 10301 35450 267955
rect 35574 156909 35634 470867
rect 35571 156908 35637 156909
rect 35571 156844 35572 156908
rect 35636 156844 35637 156908
rect 35571 156843 35637 156844
rect 35758 21997 35818 520371
rect 36675 458284 36741 458285
rect 36675 458220 36676 458284
rect 36740 458220 36741 458284
rect 36675 458219 36741 458220
rect 36491 262308 36557 262309
rect 36491 262244 36492 262308
rect 36556 262244 36557 262308
rect 36491 262243 36557 262244
rect 36494 26621 36554 262243
rect 36678 195941 36738 458219
rect 36675 195940 36741 195941
rect 36675 195876 36676 195940
rect 36740 195876 36741 195940
rect 36675 195875 36741 195876
rect 36675 188324 36741 188325
rect 36675 188260 36676 188324
rect 36740 188260 36741 188324
rect 36675 188259 36741 188260
rect 36491 26620 36557 26621
rect 36491 26556 36492 26620
rect 36556 26556 36557 26620
rect 36491 26555 36557 26556
rect 35755 21996 35821 21997
rect 35755 21932 35756 21996
rect 35820 21932 35821 21996
rect 35755 21931 35821 21932
rect 35387 10300 35453 10301
rect 35387 10236 35388 10300
rect 35452 10236 35453 10300
rect 35387 10235 35453 10236
rect 36678 3501 36738 188259
rect 36862 185605 36922 527171
rect 36859 185604 36925 185605
rect 36859 185540 36860 185604
rect 36924 185540 36925 185604
rect 36859 185539 36925 185540
rect 37046 184245 37106 527307
rect 37794 507454 38414 542898
rect 38515 534172 38581 534173
rect 38515 534108 38516 534172
rect 38580 534108 38581 534172
rect 38515 534107 38581 534108
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37595 483036 37661 483037
rect 37595 482972 37596 483036
rect 37660 482972 37661 483036
rect 37595 482971 37661 482972
rect 37043 184244 37109 184245
rect 37043 184180 37044 184244
rect 37108 184180 37109 184244
rect 37043 184179 37109 184180
rect 37598 25805 37658 482971
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37595 25804 37661 25805
rect 37595 25740 37596 25804
rect 37660 25740 37661 25804
rect 37595 25739 37661 25740
rect 36675 3500 36741 3501
rect 36675 3436 36676 3500
rect 36740 3436 36741 3500
rect 36675 3435 36741 3436
rect 37794 3454 38414 38898
rect 38518 25941 38578 534107
rect 39254 220829 39314 558043
rect 39435 450532 39501 450533
rect 39435 450468 39436 450532
rect 39500 450468 39501 450532
rect 39435 450467 39501 450468
rect 39251 220828 39317 220829
rect 39251 220764 39252 220828
rect 39316 220764 39317 220828
rect 39251 220763 39317 220764
rect 39251 218108 39317 218109
rect 39251 218044 39252 218108
rect 39316 218044 39317 218108
rect 39251 218043 39317 218044
rect 39254 205733 39314 218043
rect 39067 205732 39133 205733
rect 39067 205668 39068 205732
rect 39132 205668 39133 205732
rect 39067 205667 39133 205668
rect 39251 205732 39317 205733
rect 39251 205668 39252 205732
rect 39316 205668 39317 205732
rect 39251 205667 39317 205668
rect 38515 25940 38581 25941
rect 38515 25876 38516 25940
rect 38580 25876 38581 25940
rect 38515 25875 38581 25876
rect 39070 24037 39130 205667
rect 39251 203556 39317 203557
rect 39251 203492 39252 203556
rect 39316 203492 39317 203556
rect 39251 203491 39317 203492
rect 39067 24036 39133 24037
rect 39067 23972 39068 24036
rect 39132 23972 39133 24036
rect 39067 23971 39133 23972
rect 39254 16557 39314 203491
rect 39438 167789 39498 450467
rect 39622 204917 39682 562667
rect 41275 561236 41341 561237
rect 41275 561172 41276 561236
rect 41340 561172 41341 561236
rect 41275 561171 41341 561172
rect 41278 510509 41338 561171
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 41827 533356 41893 533357
rect 41827 533292 41828 533356
rect 41892 533292 41893 533356
rect 41827 533291 41893 533292
rect 41275 510508 41341 510509
rect 41275 510444 41276 510508
rect 41340 510444 41341 510508
rect 41275 510443 41341 510444
rect 41275 498812 41341 498813
rect 41275 498748 41276 498812
rect 41340 498748 41341 498812
rect 41275 498747 41341 498748
rect 41091 490652 41157 490653
rect 41091 490588 41092 490652
rect 41156 490588 41157 490652
rect 41091 490587 41157 490588
rect 39803 476372 39869 476373
rect 39803 476308 39804 476372
rect 39868 476308 39869 476372
rect 39803 476307 39869 476308
rect 39619 204916 39685 204917
rect 39619 204852 39620 204916
rect 39684 204852 39685 204916
rect 39619 204851 39685 204852
rect 39435 167788 39501 167789
rect 39435 167724 39436 167788
rect 39500 167724 39501 167788
rect 39435 167723 39501 167724
rect 39806 28797 39866 476307
rect 40907 465220 40973 465221
rect 40907 465156 40908 465220
rect 40972 465156 40973 465220
rect 40907 465155 40973 465156
rect 40723 438972 40789 438973
rect 40723 438908 40724 438972
rect 40788 438908 40789 438972
rect 40723 438907 40789 438908
rect 40726 166293 40786 438907
rect 40723 166292 40789 166293
rect 40723 166228 40724 166292
rect 40788 166228 40789 166292
rect 40723 166227 40789 166228
rect 40910 157045 40970 465155
rect 41094 180573 41154 490587
rect 41091 180572 41157 180573
rect 41091 180508 41092 180572
rect 41156 180508 41157 180572
rect 41091 180507 41157 180508
rect 41091 174588 41157 174589
rect 41091 174524 41092 174588
rect 41156 174524 41157 174588
rect 41091 174523 41157 174524
rect 40907 157044 40973 157045
rect 40907 156980 40908 157044
rect 40972 156980 40973 157044
rect 40907 156979 40973 156980
rect 41094 135285 41154 174523
rect 41278 173365 41338 498747
rect 41643 466580 41709 466581
rect 41643 466516 41644 466580
rect 41708 466516 41709 466580
rect 41643 466515 41709 466516
rect 41275 173364 41341 173365
rect 41275 173300 41276 173364
rect 41340 173300 41341 173364
rect 41275 173299 41341 173300
rect 41275 172140 41341 172141
rect 41275 172076 41276 172140
rect 41340 172076 41341 172140
rect 41275 172075 41341 172076
rect 41091 135284 41157 135285
rect 41091 135220 41092 135284
rect 41156 135220 41157 135284
rect 41091 135219 41157 135220
rect 41278 48653 41338 172075
rect 41646 169013 41706 466515
rect 41830 200021 41890 533291
rect 42011 515132 42077 515133
rect 42011 515068 42012 515132
rect 42076 515068 42077 515132
rect 42011 515067 42077 515068
rect 41827 200020 41893 200021
rect 41827 199956 41828 200020
rect 41892 199956 41893 200020
rect 41827 199955 41893 199956
rect 41643 169012 41709 169013
rect 41643 168948 41644 169012
rect 41708 168948 41709 169012
rect 41643 168947 41709 168948
rect 41275 48652 41341 48653
rect 41275 48588 41276 48652
rect 41340 48588 41341 48652
rect 41275 48587 41341 48588
rect 39803 28796 39869 28797
rect 39803 28732 39804 28796
rect 39868 28732 39869 28796
rect 39803 28731 39869 28732
rect 42014 26757 42074 515067
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 43854 476237 43914 588779
rect 44955 588708 45021 588709
rect 44955 588644 44956 588708
rect 45020 588644 45021 588708
rect 44955 588643 45021 588644
rect 44771 562324 44837 562325
rect 44771 562260 44772 562324
rect 44836 562260 44837 562324
rect 44771 562259 44837 562260
rect 44035 530772 44101 530773
rect 44035 530708 44036 530772
rect 44100 530708 44101 530772
rect 44035 530707 44101 530708
rect 43851 476236 43917 476237
rect 43851 476172 43852 476236
rect 43916 476172 43917 476236
rect 43851 476171 43917 476172
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 43851 456924 43917 456925
rect 43851 456860 43852 456924
rect 43916 456860 43917 456924
rect 43851 456859 43917 456860
rect 43667 449172 43733 449173
rect 43667 449108 43668 449172
rect 43732 449108 43733 449172
rect 43667 449107 43733 449108
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 43483 313308 43549 313309
rect 43483 313244 43484 313308
rect 43548 313244 43549 313308
rect 43483 313243 43549 313244
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 43486 264621 43546 313243
rect 43483 264620 43549 264621
rect 43483 264556 43484 264620
rect 43548 264556 43549 264620
rect 43483 264555 43549 264556
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 43670 188597 43730 449107
rect 43667 188596 43733 188597
rect 43667 188532 43668 188596
rect 43732 188532 43733 188596
rect 43667 188531 43733 188532
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 43667 170508 43733 170509
rect 43667 170444 43668 170508
rect 43732 170444 43733 170508
rect 43667 170443 43733 170444
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42011 26756 42077 26757
rect 42011 26692 42012 26756
rect 42076 26692 42077 26756
rect 42011 26691 42077 26692
rect 39251 16556 39317 16557
rect 39251 16492 39252 16556
rect 39316 16492 39317 16556
rect 39251 16491 39317 16492
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 43670 3501 43730 170443
rect 43854 27029 43914 456859
rect 44038 28525 44098 530707
rect 44774 313309 44834 562259
rect 44958 383077 45018 588643
rect 51950 586669 52010 589870
rect 53054 587893 53114 589870
rect 54158 587893 54218 589870
rect 53051 587892 53117 587893
rect 53051 587828 53052 587892
rect 53116 587828 53117 587892
rect 53051 587827 53117 587828
rect 54155 587892 54221 587893
rect 54155 587828 54156 587892
rect 54220 587828 54221 587892
rect 54155 587827 54221 587828
rect 55630 587757 55690 589870
rect 56550 587893 56610 589870
rect 57838 587893 57898 589870
rect 59126 589870 59188 589930
rect 60216 589930 60276 590106
rect 61440 589930 61500 590106
rect 62528 589930 62588 590106
rect 63616 589930 63676 590106
rect 64296 589930 64356 590106
rect 64704 589930 64764 590106
rect 60216 589870 60290 589930
rect 61440 589870 61578 589930
rect 59126 587893 59186 589870
rect 60230 587893 60290 589870
rect 56547 587892 56613 587893
rect 56547 587828 56548 587892
rect 56612 587828 56613 587892
rect 56547 587827 56613 587828
rect 57835 587892 57901 587893
rect 57835 587828 57836 587892
rect 57900 587828 57901 587892
rect 57835 587827 57901 587828
rect 59123 587892 59189 587893
rect 59123 587828 59124 587892
rect 59188 587828 59189 587892
rect 59123 587827 59189 587828
rect 60227 587892 60293 587893
rect 60227 587828 60228 587892
rect 60292 587828 60293 587892
rect 60227 587827 60293 587828
rect 61518 587757 61578 589870
rect 62438 589870 62588 589930
rect 63542 589870 63676 589930
rect 64278 589870 64356 589930
rect 64646 589870 64764 589930
rect 66064 589930 66124 590106
rect 66744 589930 66804 590106
rect 67288 589930 67348 590106
rect 68376 589930 68436 590106
rect 69464 589930 69524 590106
rect 66064 589870 66178 589930
rect 62438 587893 62498 589870
rect 63542 587893 63602 589870
rect 64278 587893 64338 589870
rect 62435 587892 62501 587893
rect 62435 587828 62436 587892
rect 62500 587828 62501 587892
rect 62435 587827 62501 587828
rect 63539 587892 63605 587893
rect 63539 587828 63540 587892
rect 63604 587828 63605 587892
rect 63539 587827 63605 587828
rect 64275 587892 64341 587893
rect 64275 587828 64276 587892
rect 64340 587828 64341 587892
rect 64275 587827 64341 587828
rect 64646 587757 64706 589870
rect 66118 587893 66178 589870
rect 66670 589870 66804 589930
rect 67222 589870 67348 589930
rect 68326 589870 68436 589930
rect 69430 589870 69524 589930
rect 69600 589930 69660 590106
rect 70552 589930 70612 590106
rect 71912 589930 71972 590106
rect 69600 589870 69674 589930
rect 66670 587893 66730 589870
rect 66115 587892 66181 587893
rect 66115 587828 66116 587892
rect 66180 587828 66181 587892
rect 66115 587827 66181 587828
rect 66667 587892 66733 587893
rect 66667 587828 66668 587892
rect 66732 587828 66733 587892
rect 66667 587827 66733 587828
rect 55627 587756 55693 587757
rect 55627 587692 55628 587756
rect 55692 587692 55693 587756
rect 55627 587691 55693 587692
rect 61515 587756 61581 587757
rect 61515 587692 61516 587756
rect 61580 587692 61581 587756
rect 61515 587691 61581 587692
rect 64643 587756 64709 587757
rect 64643 587692 64644 587756
rect 64708 587692 64709 587756
rect 64643 587691 64709 587692
rect 67222 586669 67282 589870
rect 68326 587893 68386 589870
rect 68323 587892 68389 587893
rect 68323 587828 68324 587892
rect 68388 587828 68389 587892
rect 68323 587827 68389 587828
rect 69430 587757 69490 589870
rect 69614 587893 69674 589870
rect 70534 589870 70612 589930
rect 71822 589870 71972 589930
rect 72048 589930 72108 590106
rect 73000 589930 73060 590106
rect 74088 589930 74148 590106
rect 72048 589870 72250 589930
rect 70534 587893 70594 589870
rect 71822 587893 71882 589870
rect 69611 587892 69677 587893
rect 69611 587828 69612 587892
rect 69676 587828 69677 587892
rect 69611 587827 69677 587828
rect 70531 587892 70597 587893
rect 70531 587828 70532 587892
rect 70596 587828 70597 587892
rect 70531 587827 70597 587828
rect 71819 587892 71885 587893
rect 71819 587828 71820 587892
rect 71884 587828 71885 587892
rect 71819 587827 71885 587828
rect 72190 587757 72250 589870
rect 72926 589870 73060 589930
rect 74030 589870 74148 589930
rect 74496 589930 74556 590106
rect 75448 589930 75508 590106
rect 76672 589930 76732 590106
rect 74496 589870 74642 589930
rect 75448 589870 75562 589930
rect 72926 587893 72986 589870
rect 72923 587892 72989 587893
rect 72923 587828 72924 587892
rect 72988 587828 72989 587892
rect 72923 587827 72989 587828
rect 69427 587756 69493 587757
rect 69427 587692 69428 587756
rect 69492 587692 69493 587756
rect 69427 587691 69493 587692
rect 72187 587756 72253 587757
rect 72187 587692 72188 587756
rect 72252 587692 72253 587756
rect 72187 587691 72253 587692
rect 74030 587621 74090 589870
rect 74582 587893 74642 589870
rect 74579 587892 74645 587893
rect 74579 587828 74580 587892
rect 74644 587828 74645 587892
rect 74579 587827 74645 587828
rect 75502 587757 75562 589870
rect 76606 589870 76732 589930
rect 77080 589930 77140 590106
rect 77760 589930 77820 590106
rect 78848 589930 78908 590106
rect 77080 589870 77218 589930
rect 75499 587756 75565 587757
rect 75499 587692 75500 587756
rect 75564 587692 75565 587756
rect 75499 587691 75565 587692
rect 74027 587620 74093 587621
rect 74027 587556 74028 587620
rect 74092 587556 74093 587620
rect 74027 587555 74093 587556
rect 76606 586669 76666 589870
rect 77158 587757 77218 589870
rect 77710 589870 77820 589930
rect 78814 589870 78908 589930
rect 79528 589930 79588 590106
rect 79936 589930 79996 590106
rect 81296 589930 81356 590106
rect 81976 589930 82036 590106
rect 82384 589930 82444 590106
rect 83608 589930 83668 590106
rect 79528 589870 79610 589930
rect 77710 587893 77770 589870
rect 78814 587893 78874 589870
rect 79550 587893 79610 589870
rect 79918 589870 79996 589930
rect 81206 589870 81356 589930
rect 81942 589870 82036 589930
rect 82310 589870 82444 589930
rect 83598 589870 83668 589930
rect 84288 589930 84348 590106
rect 84696 589930 84756 590106
rect 85784 589930 85844 590106
rect 87008 589930 87068 590106
rect 84288 589870 84394 589930
rect 77707 587892 77773 587893
rect 77707 587828 77708 587892
rect 77772 587828 77773 587892
rect 77707 587827 77773 587828
rect 78811 587892 78877 587893
rect 78811 587828 78812 587892
rect 78876 587828 78877 587892
rect 78811 587827 78877 587828
rect 79547 587892 79613 587893
rect 79547 587828 79548 587892
rect 79612 587828 79613 587892
rect 79547 587827 79613 587828
rect 79918 587757 79978 589870
rect 81206 587893 81266 589870
rect 81203 587892 81269 587893
rect 81203 587828 81204 587892
rect 81268 587828 81269 587892
rect 81203 587827 81269 587828
rect 81942 587757 82002 589870
rect 82310 587893 82370 589870
rect 83598 587893 83658 589870
rect 84334 589525 84394 589870
rect 84518 589870 84756 589930
rect 85622 589870 85844 589930
rect 86910 589870 87068 589930
rect 84331 589524 84397 589525
rect 84331 589460 84332 589524
rect 84396 589460 84397 589524
rect 84331 589459 84397 589460
rect 84518 589290 84578 589870
rect 83966 589230 84578 589290
rect 82307 587892 82373 587893
rect 82307 587828 82308 587892
rect 82372 587828 82373 587892
rect 82307 587827 82373 587828
rect 83595 587892 83661 587893
rect 83595 587828 83596 587892
rect 83660 587828 83661 587892
rect 83595 587827 83661 587828
rect 77155 587756 77221 587757
rect 77155 587692 77156 587756
rect 77220 587692 77221 587756
rect 77155 587691 77221 587692
rect 79915 587756 79981 587757
rect 79915 587692 79916 587756
rect 79980 587692 79981 587756
rect 79915 587691 79981 587692
rect 81939 587756 82005 587757
rect 81939 587692 81940 587756
rect 82004 587692 82005 587756
rect 81939 587691 82005 587692
rect 51947 586668 52013 586669
rect 51947 586604 51948 586668
rect 52012 586604 52013 586668
rect 51947 586603 52013 586604
rect 67219 586668 67285 586669
rect 67219 586604 67220 586668
rect 67284 586604 67285 586668
rect 67219 586603 67285 586604
rect 76603 586668 76669 586669
rect 76603 586604 76604 586668
rect 76668 586604 76669 586668
rect 76603 586603 76669 586604
rect 83966 586530 84026 589230
rect 85622 586533 85682 589870
rect 86910 586669 86970 589870
rect 87144 589290 87204 590106
rect 88232 589930 88292 590106
rect 89320 589930 89380 590106
rect 89592 589930 89652 590106
rect 90408 589930 90468 590106
rect 91768 589930 91828 590106
rect 87094 589230 87204 589290
rect 88198 589870 88292 589930
rect 89302 589870 89380 589930
rect 89486 589870 89652 589930
rect 90406 589870 90468 589930
rect 91694 589870 91828 589930
rect 92040 589930 92100 590106
rect 92992 589930 93052 590106
rect 92040 589870 92122 589930
rect 87094 587893 87154 589230
rect 87091 587892 87157 587893
rect 87091 587828 87092 587892
rect 87156 587828 87157 587892
rect 87091 587827 87157 587828
rect 88198 587757 88258 589870
rect 88195 587756 88261 587757
rect 88195 587692 88196 587756
rect 88260 587692 88261 587756
rect 88195 587691 88261 587692
rect 89302 586669 89362 589870
rect 89486 587893 89546 589870
rect 89483 587892 89549 587893
rect 89483 587828 89484 587892
rect 89548 587828 89549 587892
rect 89483 587827 89549 587828
rect 90406 586669 90466 589870
rect 91694 587893 91754 589870
rect 91691 587892 91757 587893
rect 91691 587828 91692 587892
rect 91756 587828 91757 587892
rect 91691 587827 91757 587828
rect 92062 586669 92122 589870
rect 92982 589870 93052 589930
rect 94080 589930 94140 590106
rect 94488 589930 94548 590106
rect 94080 589870 94146 589930
rect 92982 587893 93042 589870
rect 94086 587893 94146 589870
rect 94454 589870 94548 589930
rect 95168 589930 95228 590106
rect 96936 589930 96996 590106
rect 99520 589930 99580 590106
rect 95168 589870 95250 589930
rect 94454 587893 94514 589870
rect 92979 587892 93045 587893
rect 92979 587828 92980 587892
rect 93044 587828 93045 587892
rect 92979 587827 93045 587828
rect 94083 587892 94149 587893
rect 94083 587828 94084 587892
rect 94148 587828 94149 587892
rect 94083 587827 94149 587828
rect 94451 587892 94517 587893
rect 94451 587828 94452 587892
rect 94516 587828 94517 587892
rect 94451 587827 94517 587828
rect 95190 587757 95250 589870
rect 96846 589870 96996 589930
rect 99422 589870 99580 589930
rect 101968 589930 102028 590106
rect 104280 589930 104340 590106
rect 107000 589930 107060 590106
rect 109448 589930 109508 590106
rect 101968 589870 102058 589930
rect 95187 587756 95253 587757
rect 95187 587692 95188 587756
rect 95252 587692 95253 587756
rect 95187 587691 95253 587692
rect 96846 586669 96906 589870
rect 99422 587893 99482 589870
rect 101998 587893 102058 589870
rect 104206 589870 104340 589930
rect 106966 589870 107060 589930
rect 109358 589870 109508 589930
rect 111896 589930 111956 590106
rect 114480 589930 114540 590106
rect 116928 589930 116988 590106
rect 119512 589930 119572 590106
rect 121960 589930 122020 590106
rect 124544 589930 124604 590106
rect 111896 589870 111994 589930
rect 114480 589870 114570 589930
rect 104206 589290 104266 589870
rect 103286 589230 104266 589290
rect 99419 587892 99485 587893
rect 99419 587828 99420 587892
rect 99484 587828 99485 587892
rect 99419 587827 99485 587828
rect 101995 587892 102061 587893
rect 101995 587828 101996 587892
rect 102060 587828 102061 587892
rect 101995 587827 102061 587828
rect 86907 586668 86973 586669
rect 86907 586604 86908 586668
rect 86972 586604 86973 586668
rect 86907 586603 86973 586604
rect 89299 586668 89365 586669
rect 89299 586604 89300 586668
rect 89364 586604 89365 586668
rect 89299 586603 89365 586604
rect 90403 586668 90469 586669
rect 90403 586604 90404 586668
rect 90468 586604 90469 586668
rect 90403 586603 90469 586604
rect 92059 586668 92125 586669
rect 92059 586604 92060 586668
rect 92124 586604 92125 586668
rect 92059 586603 92125 586604
rect 96843 586668 96909 586669
rect 96843 586604 96844 586668
rect 96908 586604 96909 586668
rect 96843 586603 96909 586604
rect 84147 586532 84213 586533
rect 84147 586530 84148 586532
rect 83966 586470 84148 586530
rect 84147 586468 84148 586470
rect 84212 586468 84213 586532
rect 84147 586467 84213 586468
rect 85619 586532 85685 586533
rect 85619 586468 85620 586532
rect 85684 586468 85685 586532
rect 103286 586530 103346 589230
rect 106966 587893 107026 589870
rect 109358 587893 109418 589870
rect 111934 587893 111994 589870
rect 114510 587893 114570 589870
rect 116902 589870 116988 589930
rect 119478 589870 119572 589930
rect 121870 589870 122020 589930
rect 124446 589870 124604 589930
rect 126992 589930 127052 590106
rect 129440 589930 129500 590106
rect 131888 589930 131948 590106
rect 134472 589930 134532 590106
rect 126992 589870 127082 589930
rect 106963 587892 107029 587893
rect 106963 587828 106964 587892
rect 107028 587828 107029 587892
rect 106963 587827 107029 587828
rect 109355 587892 109421 587893
rect 109355 587828 109356 587892
rect 109420 587828 109421 587892
rect 109355 587827 109421 587828
rect 111931 587892 111997 587893
rect 111931 587828 111932 587892
rect 111996 587828 111997 587892
rect 111931 587827 111997 587828
rect 114507 587892 114573 587893
rect 114507 587828 114508 587892
rect 114572 587828 114573 587892
rect 114507 587827 114573 587828
rect 116902 586669 116962 589870
rect 119478 587893 119538 589870
rect 119475 587892 119541 587893
rect 119475 587828 119476 587892
rect 119540 587828 119541 587892
rect 119475 587827 119541 587828
rect 121870 586669 121930 589870
rect 124446 587893 124506 589870
rect 124443 587892 124509 587893
rect 124443 587828 124444 587892
rect 124508 587828 124509 587892
rect 124443 587827 124509 587828
rect 127022 587757 127082 589870
rect 129414 589870 129500 589930
rect 131806 589870 131948 589930
rect 134382 589870 134532 589930
rect 136920 589930 136980 590106
rect 139368 589930 139428 590106
rect 141952 589930 142012 590106
rect 159224 589930 159284 590106
rect 136920 589870 137018 589930
rect 129414 587893 129474 589870
rect 131806 587893 131866 589870
rect 134382 587893 134442 589870
rect 136958 587893 137018 589870
rect 139350 589870 139428 589930
rect 141926 589870 142012 589930
rect 159222 589870 159284 589930
rect 159360 589930 159420 590106
rect 159360 589870 159466 589930
rect 139350 587893 139410 589870
rect 141926 587893 141986 589870
rect 129411 587892 129477 587893
rect 129411 587828 129412 587892
rect 129476 587828 129477 587892
rect 129411 587827 129477 587828
rect 131803 587892 131869 587893
rect 131803 587828 131804 587892
rect 131868 587828 131869 587892
rect 131803 587827 131869 587828
rect 134379 587892 134445 587893
rect 134379 587828 134380 587892
rect 134444 587828 134445 587892
rect 134379 587827 134445 587828
rect 136955 587892 137021 587893
rect 136955 587828 136956 587892
rect 137020 587828 137021 587892
rect 136955 587827 137021 587828
rect 139347 587892 139413 587893
rect 139347 587828 139348 587892
rect 139412 587828 139413 587892
rect 139347 587827 139413 587828
rect 141923 587892 141989 587893
rect 141923 587828 141924 587892
rect 141988 587828 141989 587892
rect 141923 587827 141989 587828
rect 127019 587756 127085 587757
rect 127019 587692 127020 587756
rect 127084 587692 127085 587756
rect 127019 587691 127085 587692
rect 159222 586669 159282 589870
rect 159406 587893 159466 589870
rect 159403 587892 159469 587893
rect 159403 587828 159404 587892
rect 159468 587828 159469 587892
rect 159403 587827 159469 587828
rect 116899 586668 116965 586669
rect 116899 586604 116900 586668
rect 116964 586604 116965 586668
rect 116899 586603 116965 586604
rect 121867 586668 121933 586669
rect 121867 586604 121868 586668
rect 121932 586604 121933 586668
rect 121867 586603 121933 586604
rect 159219 586668 159285 586669
rect 159219 586604 159220 586668
rect 159284 586604 159285 586668
rect 159219 586603 159285 586604
rect 103467 586532 103533 586533
rect 103467 586530 103468 586532
rect 103286 586470 103468 586530
rect 85619 586467 85685 586468
rect 103467 586468 103468 586470
rect 103532 586468 103533 586532
rect 103467 586467 103533 586468
rect 48451 586396 48517 586397
rect 48451 586332 48452 586396
rect 48516 586332 48517 586396
rect 48451 586331 48517 586332
rect 46979 583132 47045 583133
rect 46979 583068 46980 583132
rect 47044 583068 47045 583132
rect 46979 583067 47045 583068
rect 46795 577556 46861 577557
rect 46795 577492 46796 577556
rect 46860 577492 46861 577556
rect 46795 577491 46861 577492
rect 46611 574700 46677 574701
rect 46611 574636 46612 574700
rect 46676 574636 46677 574700
rect 46611 574635 46677 574636
rect 46243 567900 46309 567901
rect 46243 567836 46244 567900
rect 46308 567836 46309 567900
rect 46243 567835 46309 567836
rect 45323 548316 45389 548317
rect 45323 548252 45324 548316
rect 45388 548252 45389 548316
rect 45323 548251 45389 548252
rect 45139 486572 45205 486573
rect 45139 486508 45140 486572
rect 45204 486508 45205 486572
rect 45139 486507 45205 486508
rect 44955 383076 45021 383077
rect 44955 383012 44956 383076
rect 45020 383012 45021 383076
rect 44955 383011 45021 383012
rect 44955 317388 45021 317389
rect 44955 317324 44956 317388
rect 45020 317324 45021 317388
rect 44955 317323 45021 317324
rect 44771 313308 44837 313309
rect 44771 313244 44772 313308
rect 44836 313244 44837 313308
rect 44771 313243 44837 313244
rect 44958 285293 45018 317323
rect 44955 285292 45021 285293
rect 44955 285228 44956 285292
rect 45020 285228 45021 285292
rect 44955 285227 45021 285228
rect 44771 276044 44837 276045
rect 44771 275980 44772 276044
rect 44836 275980 44837 276044
rect 44771 275979 44837 275980
rect 44587 264892 44653 264893
rect 44587 264828 44588 264892
rect 44652 264828 44653 264892
rect 44587 264827 44653 264828
rect 44590 245445 44650 264827
rect 44774 259589 44834 275979
rect 44771 259588 44837 259589
rect 44771 259524 44772 259588
rect 44836 259524 44837 259588
rect 44771 259523 44837 259524
rect 44955 258228 45021 258229
rect 44955 258164 44956 258228
rect 45020 258164 45021 258228
rect 44955 258163 45021 258164
rect 44587 245444 44653 245445
rect 44587 245380 44588 245444
rect 44652 245380 44653 245444
rect 44587 245379 44653 245380
rect 44771 244356 44837 244357
rect 44771 244292 44772 244356
rect 44836 244292 44837 244356
rect 44771 244291 44837 244292
rect 44774 220829 44834 244291
rect 44771 220828 44837 220829
rect 44771 220764 44772 220828
rect 44836 220764 44837 220828
rect 44771 220763 44837 220764
rect 44587 220148 44653 220149
rect 44587 220084 44588 220148
rect 44652 220084 44653 220148
rect 44587 220083 44653 220084
rect 44590 201653 44650 220083
rect 44587 201652 44653 201653
rect 44587 201588 44588 201652
rect 44652 201588 44653 201652
rect 44587 201587 44653 201588
rect 44771 201516 44837 201517
rect 44771 201452 44772 201516
rect 44836 201452 44837 201516
rect 44771 201451 44837 201452
rect 44035 28524 44101 28525
rect 44035 28460 44036 28524
rect 44100 28460 44101 28524
rect 44035 28459 44101 28460
rect 43851 27028 43917 27029
rect 43851 26964 43852 27028
rect 43916 26964 43917 27028
rect 43851 26963 43917 26964
rect 44774 18869 44834 201451
rect 44958 27301 45018 258163
rect 45142 192677 45202 486507
rect 45139 192676 45205 192677
rect 45139 192612 45140 192676
rect 45204 192612 45205 192676
rect 45139 192611 45205 192612
rect 45326 28117 45386 548251
rect 46246 412997 46306 567835
rect 46427 563684 46493 563685
rect 46427 563620 46428 563684
rect 46492 563620 46493 563684
rect 46427 563619 46493 563620
rect 46243 412996 46309 412997
rect 46243 412932 46244 412996
rect 46308 412932 46309 412996
rect 46243 412931 46309 412932
rect 46243 402116 46309 402117
rect 46243 402052 46244 402116
rect 46308 402052 46309 402116
rect 46243 402051 46309 402052
rect 46059 252516 46125 252517
rect 46059 252452 46060 252516
rect 46124 252452 46125 252516
rect 46059 252451 46125 252452
rect 45875 178668 45941 178669
rect 45875 178604 45876 178668
rect 45940 178604 45941 178668
rect 45875 178603 45941 178604
rect 45878 30973 45938 178603
rect 46062 171733 46122 252451
rect 46246 195261 46306 402051
rect 46430 251837 46490 563619
rect 46427 251836 46493 251837
rect 46427 251772 46428 251836
rect 46492 251772 46493 251836
rect 46427 251771 46493 251772
rect 46427 247620 46493 247621
rect 46427 247556 46428 247620
rect 46492 247556 46493 247620
rect 46427 247555 46493 247556
rect 46243 195260 46309 195261
rect 46243 195196 46244 195260
rect 46308 195196 46309 195260
rect 46243 195195 46309 195196
rect 46243 172004 46309 172005
rect 46243 171940 46244 172004
rect 46308 171940 46309 172004
rect 46243 171939 46309 171940
rect 46059 171732 46125 171733
rect 46059 171668 46060 171732
rect 46124 171668 46125 171732
rect 46059 171667 46125 171668
rect 46246 123453 46306 171939
rect 46430 158269 46490 247555
rect 46614 247077 46674 574635
rect 46611 247076 46677 247077
rect 46611 247012 46612 247076
rect 46676 247012 46677 247076
rect 46611 247011 46677 247012
rect 46798 244357 46858 577491
rect 46611 244356 46677 244357
rect 46611 244292 46612 244356
rect 46676 244292 46677 244356
rect 46611 244291 46677 244292
rect 46795 244356 46861 244357
rect 46795 244292 46796 244356
rect 46860 244292 46861 244356
rect 46795 244291 46861 244292
rect 46614 174725 46674 244291
rect 46982 210357 47042 583067
rect 48454 576870 48514 586331
rect 48454 576810 48882 576870
rect 47347 570756 47413 570757
rect 47347 570692 47348 570756
rect 47412 570692 47413 570756
rect 47347 570691 47413 570692
rect 47163 569260 47229 569261
rect 47163 569196 47164 569260
rect 47228 569196 47229 569260
rect 47163 569195 47229 569196
rect 47166 220557 47226 569195
rect 47350 240957 47410 570691
rect 48451 562596 48517 562597
rect 48451 562532 48452 562596
rect 48516 562532 48517 562596
rect 48451 562531 48517 562532
rect 48083 558788 48149 558789
rect 48083 558724 48084 558788
rect 48148 558724 48149 558788
rect 48083 558723 48149 558724
rect 48086 558650 48146 558723
rect 48454 558650 48514 562531
rect 48635 562460 48701 562461
rect 48635 562396 48636 562460
rect 48700 562396 48701 562460
rect 48635 562395 48701 562396
rect 48086 558590 48514 558650
rect 48267 558108 48333 558109
rect 48267 558044 48268 558108
rect 48332 558044 48333 558108
rect 48267 558043 48333 558044
rect 48270 557970 48330 558043
rect 48638 557970 48698 562395
rect 48270 557910 48698 557970
rect 48822 557550 48882 576810
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 562000 177914 574398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 562000 182414 578898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 562000 186914 583398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 562000 191414 587898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 562000 195914 592398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 562000 200414 596898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 675308 209414 677898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 675308 213914 682398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 675308 218414 686898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 675308 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 675308 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 675308 231914 700398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 675308 245414 677898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 675308 249914 682398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 675308 254414 686898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 675308 258914 691398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 675308 263414 695898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 675308 267914 700398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 675308 281414 677898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 675308 285914 682398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 675308 290414 686898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 675308 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 675308 299414 695898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 675308 303914 700398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 675308 317414 677898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 675308 321914 682398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 675308 326414 686898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 675308 330914 691398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 675308 335414 695898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 675308 339914 700398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 356651 686084 356717 686085
rect 356651 686020 356652 686084
rect 356716 686020 356717 686084
rect 356651 686019 356717 686020
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 346899 675068 346965 675069
rect 346899 675004 346900 675068
rect 346964 675004 346965 675068
rect 346899 675003 346965 675004
rect 328499 674932 328565 674933
rect 328499 674868 328500 674932
rect 328564 674868 328565 674932
rect 328499 674867 328565 674868
rect 329787 674932 329853 674933
rect 329787 674868 329788 674932
rect 329852 674868 329853 674932
rect 329787 674867 329853 674868
rect 340827 674932 340893 674933
rect 340827 674868 340828 674932
rect 340892 674868 340893 674932
rect 340827 674867 340893 674868
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 328502 673470 328562 674867
rect 329790 673470 329850 674867
rect 204294 637954 204914 673398
rect 328464 673410 328562 673470
rect 329688 673410 329850 673470
rect 340830 673470 340890 674867
rect 340830 673410 340900 673470
rect 328464 673202 328524 673410
rect 329688 673202 329748 673410
rect 340840 673202 340900 673410
rect 210272 655954 210620 655986
rect 210272 655718 210328 655954
rect 210564 655718 210620 655954
rect 210272 655634 210620 655718
rect 210272 655398 210328 655634
rect 210564 655398 210620 655634
rect 210272 655366 210620 655398
rect 346000 655954 346348 655986
rect 346000 655718 346056 655954
rect 346292 655718 346348 655954
rect 346000 655634 346348 655718
rect 346000 655398 346056 655634
rect 346292 655398 346348 655634
rect 346000 655366 346348 655398
rect 210952 651454 211300 651486
rect 210952 651218 211008 651454
rect 211244 651218 211300 651454
rect 210952 651134 211300 651218
rect 210952 650898 211008 651134
rect 211244 650898 211300 651134
rect 210952 650866 211300 650898
rect 345320 651454 345668 651486
rect 345320 651218 345376 651454
rect 345612 651218 345668 651454
rect 345320 651134 345668 651218
rect 345320 650898 345376 651134
rect 345612 650898 345668 651134
rect 345320 650866 345668 650898
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 210272 619954 210620 619986
rect 210272 619718 210328 619954
rect 210564 619718 210620 619954
rect 210272 619634 210620 619718
rect 210272 619398 210328 619634
rect 210564 619398 210620 619634
rect 210272 619366 210620 619398
rect 346000 619954 346348 619986
rect 346000 619718 346056 619954
rect 346292 619718 346348 619954
rect 346000 619634 346348 619718
rect 346000 619398 346056 619634
rect 346292 619398 346348 619634
rect 346000 619366 346348 619398
rect 210952 615454 211300 615486
rect 210952 615218 211008 615454
rect 211244 615218 211300 615454
rect 210952 615134 211300 615218
rect 210952 614898 211008 615134
rect 211244 614898 211300 615134
rect 210952 614866 211300 614898
rect 345320 615454 345668 615486
rect 345320 615218 345376 615454
rect 345612 615218 345668 615454
rect 345320 615134 345668 615218
rect 345320 614898 345376 615134
rect 345612 614898 345668 615134
rect 345320 614866 345668 614898
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 226056 589930 226116 590106
rect 227144 589930 227204 590106
rect 228232 589930 228292 590106
rect 229592 589930 229652 590106
rect 226014 589870 226116 589930
rect 227118 589870 227204 589930
rect 228222 589870 228292 589930
rect 229510 589870 229652 589930
rect 230544 589930 230604 590106
rect 231768 589930 231828 590106
rect 230544 589870 230674 589930
rect 226014 587893 226074 589870
rect 226011 587892 226077 587893
rect 226011 587828 226012 587892
rect 226076 587828 226077 587892
rect 226011 587827 226077 587828
rect 227118 587485 227178 589870
rect 228222 587893 228282 589870
rect 228219 587892 228285 587893
rect 228219 587828 228220 587892
rect 228284 587828 228285 587892
rect 228219 587827 228285 587828
rect 227115 587484 227181 587485
rect 227115 587420 227116 587484
rect 227180 587420 227181 587484
rect 227115 587419 227181 587420
rect 229510 587349 229570 589870
rect 230614 587893 230674 589870
rect 231718 589870 231828 589930
rect 233128 589930 233188 590106
rect 234216 589930 234276 590106
rect 235440 589930 235500 590106
rect 236528 589930 236588 590106
rect 237616 589930 237676 590106
rect 233128 589870 233250 589930
rect 234216 589870 234354 589930
rect 230611 587892 230677 587893
rect 230611 587828 230612 587892
rect 230676 587828 230677 587892
rect 230611 587827 230677 587828
rect 229507 587348 229573 587349
rect 229507 587284 229508 587348
rect 229572 587284 229573 587348
rect 229507 587283 229573 587284
rect 231718 586669 231778 589870
rect 233190 586669 233250 589870
rect 234294 587893 234354 589870
rect 235398 589870 235500 589930
rect 236502 589870 236588 589930
rect 237606 589870 237676 589930
rect 238296 589930 238356 590106
rect 238704 589930 238764 590106
rect 240064 589930 240124 590106
rect 240744 589930 240804 590106
rect 241288 589930 241348 590106
rect 238296 589870 238402 589930
rect 234291 587892 234357 587893
rect 234291 587828 234292 587892
rect 234356 587828 234357 587892
rect 234291 587827 234357 587828
rect 235398 587757 235458 589870
rect 236502 587893 236562 589870
rect 237606 587893 237666 589870
rect 238342 587893 238402 589870
rect 238526 589870 238764 589930
rect 239998 589870 240124 589930
rect 240734 589870 240804 589930
rect 241286 589870 241348 589930
rect 242376 589930 242436 590106
rect 243464 589930 243524 590106
rect 242376 589870 242450 589930
rect 236499 587892 236565 587893
rect 236499 587828 236500 587892
rect 236564 587828 236565 587892
rect 236499 587827 236565 587828
rect 237603 587892 237669 587893
rect 237603 587828 237604 587892
rect 237668 587828 237669 587892
rect 237603 587827 237669 587828
rect 238339 587892 238405 587893
rect 238339 587828 238340 587892
rect 238404 587828 238405 587892
rect 238339 587827 238405 587828
rect 235395 587756 235461 587757
rect 235395 587692 235396 587756
rect 235460 587692 235461 587756
rect 235395 587691 235461 587692
rect 238526 586805 238586 589870
rect 239998 587893 240058 589870
rect 239995 587892 240061 587893
rect 239995 587828 239996 587892
rect 240060 587828 240061 587892
rect 239995 587827 240061 587828
rect 240734 587757 240794 589870
rect 241286 587893 241346 589870
rect 242390 587893 242450 589870
rect 243310 589870 243524 589930
rect 243600 589930 243660 590106
rect 244552 589930 244612 590106
rect 245912 589930 245972 590106
rect 243600 589870 243738 589930
rect 244552 589870 244658 589930
rect 243310 587893 243370 589870
rect 241283 587892 241349 587893
rect 241283 587828 241284 587892
rect 241348 587828 241349 587892
rect 241283 587827 241349 587828
rect 242387 587892 242453 587893
rect 242387 587828 242388 587892
rect 242452 587828 242453 587892
rect 242387 587827 242453 587828
rect 243307 587892 243373 587893
rect 243307 587828 243308 587892
rect 243372 587828 243373 587892
rect 243307 587827 243373 587828
rect 240731 587756 240797 587757
rect 240731 587692 240732 587756
rect 240796 587692 240797 587756
rect 240731 587691 240797 587692
rect 238523 586804 238589 586805
rect 238523 586740 238524 586804
rect 238588 586740 238589 586804
rect 238523 586739 238589 586740
rect 243678 586669 243738 589870
rect 244598 587893 244658 589870
rect 245886 589870 245972 589930
rect 246048 589930 246108 590106
rect 247000 589930 247060 590106
rect 246048 589870 246130 589930
rect 245886 587893 245946 589870
rect 244595 587892 244661 587893
rect 244595 587828 244596 587892
rect 244660 587828 244661 587892
rect 244595 587827 244661 587828
rect 245883 587892 245949 587893
rect 245883 587828 245884 587892
rect 245948 587828 245949 587892
rect 245883 587827 245949 587828
rect 246070 587757 246130 589870
rect 246990 589870 247060 589930
rect 248088 589930 248148 590106
rect 248496 589930 248556 590106
rect 248088 589870 248154 589930
rect 246990 587893 247050 589870
rect 248094 587893 248154 589870
rect 248462 589870 248556 589930
rect 249448 589930 249508 590106
rect 250672 589930 250732 590106
rect 251080 589930 251140 590106
rect 249448 589870 249626 589930
rect 248462 587893 248522 589870
rect 249566 587893 249626 589870
rect 250670 589870 250732 589930
rect 251038 589870 251140 589930
rect 251760 589930 251820 590106
rect 252848 589930 252908 590106
rect 253528 589930 253588 590106
rect 251760 589870 251834 589930
rect 252848 589870 252938 589930
rect 246987 587892 247053 587893
rect 246987 587828 246988 587892
rect 247052 587828 247053 587892
rect 246987 587827 247053 587828
rect 248091 587892 248157 587893
rect 248091 587828 248092 587892
rect 248156 587828 248157 587892
rect 248091 587827 248157 587828
rect 248459 587892 248525 587893
rect 248459 587828 248460 587892
rect 248524 587828 248525 587892
rect 248459 587827 248525 587828
rect 249563 587892 249629 587893
rect 249563 587828 249564 587892
rect 249628 587828 249629 587892
rect 249563 587827 249629 587828
rect 246067 587756 246133 587757
rect 246067 587692 246068 587756
rect 246132 587692 246133 587756
rect 246067 587691 246133 587692
rect 250670 587349 250730 589870
rect 251038 587757 251098 589870
rect 251035 587756 251101 587757
rect 251035 587692 251036 587756
rect 251100 587692 251101 587756
rect 251035 587691 251101 587692
rect 250667 587348 250733 587349
rect 250667 587284 250668 587348
rect 250732 587284 250733 587348
rect 250667 587283 250733 587284
rect 251774 586669 251834 589870
rect 252878 587893 252938 589870
rect 253430 589870 253588 589930
rect 253936 589930 253996 590106
rect 255296 589930 255356 590106
rect 253936 589870 254042 589930
rect 252875 587892 252941 587893
rect 252875 587828 252876 587892
rect 252940 587828 252941 587892
rect 252875 587827 252941 587828
rect 253430 587757 253490 589870
rect 253982 587893 254042 589870
rect 255270 589870 255356 589930
rect 255976 589930 256036 590106
rect 256384 589930 256444 590106
rect 255976 589870 256066 589930
rect 253979 587892 254045 587893
rect 253979 587828 253980 587892
rect 254044 587828 254045 587892
rect 253979 587827 254045 587828
rect 253427 587756 253493 587757
rect 253427 587692 253428 587756
rect 253492 587692 253493 587756
rect 253427 587691 253493 587692
rect 255270 587213 255330 589870
rect 256006 587893 256066 589870
rect 256374 589870 256444 589930
rect 257608 589930 257668 590106
rect 258288 589930 258348 590106
rect 258696 589930 258756 590106
rect 257608 589870 257722 589930
rect 256374 587893 256434 589870
rect 257662 587893 257722 589870
rect 258214 589870 258348 589930
rect 258582 589870 258756 589930
rect 259784 589930 259844 590106
rect 261008 589930 261068 590106
rect 259784 589870 259930 589930
rect 258214 589290 258274 589870
rect 257846 589230 258274 589290
rect 256003 587892 256069 587893
rect 256003 587828 256004 587892
rect 256068 587828 256069 587892
rect 256003 587827 256069 587828
rect 256371 587892 256437 587893
rect 256371 587828 256372 587892
rect 256436 587828 256437 587892
rect 256371 587827 256437 587828
rect 257659 587892 257725 587893
rect 257659 587828 257660 587892
rect 257724 587828 257725 587892
rect 257659 587827 257725 587828
rect 255267 587212 255333 587213
rect 255267 587148 255268 587212
rect 255332 587148 255333 587212
rect 255267 587147 255333 587148
rect 257846 586805 257906 589230
rect 257843 586804 257909 586805
rect 257843 586740 257844 586804
rect 257908 586740 257909 586804
rect 257843 586739 257909 586740
rect 231715 586668 231781 586669
rect 231715 586604 231716 586668
rect 231780 586604 231781 586668
rect 231715 586603 231781 586604
rect 233187 586668 233253 586669
rect 233187 586604 233188 586668
rect 233252 586604 233253 586668
rect 233187 586603 233253 586604
rect 243675 586668 243741 586669
rect 243675 586604 243676 586668
rect 243740 586604 243741 586668
rect 243675 586603 243741 586604
rect 251771 586668 251837 586669
rect 251771 586604 251772 586668
rect 251836 586604 251837 586668
rect 251771 586603 251837 586604
rect 258582 586533 258642 589870
rect 259870 587893 259930 589870
rect 260974 589870 261068 589930
rect 261144 589930 261204 590106
rect 262232 589930 262292 590106
rect 263320 589930 263380 590106
rect 263592 589930 263652 590106
rect 261144 589870 261218 589930
rect 262232 589870 262322 589930
rect 263320 589870 263426 589930
rect 260974 587893 261034 589870
rect 261158 587893 261218 589870
rect 262262 587893 262322 589870
rect 259867 587892 259933 587893
rect 259867 587828 259868 587892
rect 259932 587828 259933 587892
rect 259867 587827 259933 587828
rect 260971 587892 261037 587893
rect 260971 587828 260972 587892
rect 261036 587828 261037 587892
rect 260971 587827 261037 587828
rect 261155 587892 261221 587893
rect 261155 587828 261156 587892
rect 261220 587828 261221 587892
rect 261155 587827 261221 587828
rect 262259 587892 262325 587893
rect 262259 587828 262260 587892
rect 262324 587828 262325 587892
rect 262259 587827 262325 587828
rect 263366 586669 263426 589870
rect 263550 589870 263652 589930
rect 264408 589930 264468 590106
rect 265768 589930 265828 590106
rect 266040 589930 266100 590106
rect 264408 589870 264530 589930
rect 263550 587893 263610 589870
rect 263547 587892 263613 587893
rect 263547 587828 263548 587892
rect 263612 587828 263613 587892
rect 263547 587827 263613 587828
rect 264470 587757 264530 589870
rect 265758 589870 265828 589930
rect 265942 589870 266100 589930
rect 266992 589930 267052 590106
rect 268080 589930 268140 590106
rect 266992 589870 267106 589930
rect 265758 587893 265818 589870
rect 265755 587892 265821 587893
rect 265755 587828 265756 587892
rect 265820 587828 265821 587892
rect 265755 587827 265821 587828
rect 265942 587757 266002 589870
rect 264467 587756 264533 587757
rect 264467 587692 264468 587756
rect 264532 587692 264533 587756
rect 264467 587691 264533 587692
rect 265939 587756 266005 587757
rect 265939 587692 265940 587756
rect 266004 587692 266005 587756
rect 265939 587691 266005 587692
rect 267046 586669 267106 589870
rect 267966 589870 268140 589930
rect 268488 589930 268548 590106
rect 269168 589930 269228 590106
rect 270936 589930 270996 590106
rect 273520 589930 273580 590106
rect 275968 589930 276028 590106
rect 278280 589930 278340 590106
rect 268488 589870 268578 589930
rect 269168 589870 269314 589930
rect 263363 586668 263429 586669
rect 263363 586604 263364 586668
rect 263428 586604 263429 586668
rect 263363 586603 263429 586604
rect 267043 586668 267109 586669
rect 267043 586604 267044 586668
rect 267108 586604 267109 586668
rect 267043 586603 267109 586604
rect 267966 586533 268026 589870
rect 268518 587893 268578 589870
rect 269254 587893 269314 589870
rect 270910 589870 270996 589930
rect 273486 589870 273580 589930
rect 275878 589870 276028 589930
rect 278270 589870 278340 589930
rect 281000 589930 281060 590106
rect 283448 589930 283508 590106
rect 281000 589870 281090 589930
rect 270910 587893 270970 589870
rect 273486 587893 273546 589870
rect 275878 587893 275938 589870
rect 278270 589290 278330 589870
rect 277166 589230 278330 589290
rect 268515 587892 268581 587893
rect 268515 587828 268516 587892
rect 268580 587828 268581 587892
rect 268515 587827 268581 587828
rect 269251 587892 269317 587893
rect 269251 587828 269252 587892
rect 269316 587828 269317 587892
rect 269251 587827 269317 587828
rect 270907 587892 270973 587893
rect 270907 587828 270908 587892
rect 270972 587828 270973 587892
rect 270907 587827 270973 587828
rect 273483 587892 273549 587893
rect 273483 587828 273484 587892
rect 273548 587828 273549 587892
rect 273483 587827 273549 587828
rect 275875 587892 275941 587893
rect 275875 587828 275876 587892
rect 275940 587828 275941 587892
rect 275875 587827 275941 587828
rect 258579 586532 258645 586533
rect 258579 586468 258580 586532
rect 258644 586468 258645 586532
rect 258579 586467 258645 586468
rect 267963 586532 268029 586533
rect 267963 586468 267964 586532
rect 268028 586468 268029 586532
rect 277166 586530 277226 589230
rect 281030 587893 281090 589870
rect 283422 589870 283508 589930
rect 285896 589930 285956 590106
rect 288480 589930 288540 590106
rect 285896 589870 286058 589930
rect 283422 587893 283482 589870
rect 285998 587893 286058 589870
rect 288390 589870 288540 589930
rect 290928 589930 290988 590106
rect 293512 589930 293572 590106
rect 295960 589930 296020 590106
rect 298544 589930 298604 590106
rect 300992 589930 301052 590106
rect 290928 589870 291026 589930
rect 293512 589870 293602 589930
rect 288390 587893 288450 589870
rect 290966 587893 291026 589870
rect 281027 587892 281093 587893
rect 281027 587828 281028 587892
rect 281092 587828 281093 587892
rect 281027 587827 281093 587828
rect 283419 587892 283485 587893
rect 283419 587828 283420 587892
rect 283484 587828 283485 587892
rect 283419 587827 283485 587828
rect 285995 587892 286061 587893
rect 285995 587828 285996 587892
rect 286060 587828 286061 587892
rect 285995 587827 286061 587828
rect 288387 587892 288453 587893
rect 288387 587828 288388 587892
rect 288452 587828 288453 587892
rect 288387 587827 288453 587828
rect 290963 587892 291029 587893
rect 290963 587828 290964 587892
rect 291028 587828 291029 587892
rect 290963 587827 291029 587828
rect 293542 586669 293602 589870
rect 295934 589870 296020 589930
rect 298510 589870 298604 589930
rect 300902 589870 301052 589930
rect 303440 589930 303500 590106
rect 305888 589930 305948 590106
rect 308472 589930 308532 590106
rect 310920 589930 310980 590106
rect 303440 589870 303538 589930
rect 295934 586669 295994 589870
rect 298510 587893 298570 589870
rect 300902 587893 300962 589870
rect 303478 587893 303538 589870
rect 305870 589870 305948 589930
rect 308446 589870 308532 589930
rect 310838 589870 310980 589930
rect 313368 589930 313428 590106
rect 315952 589930 316012 590106
rect 333224 589930 333284 590106
rect 313368 589870 313474 589930
rect 305870 587893 305930 589870
rect 308446 587893 308506 589870
rect 310838 587893 310898 589870
rect 313414 587893 313474 589870
rect 315806 589870 316012 589930
rect 333102 589870 333284 589930
rect 333360 589930 333420 590106
rect 333360 589870 333530 589930
rect 298507 587892 298573 587893
rect 298507 587828 298508 587892
rect 298572 587828 298573 587892
rect 298507 587827 298573 587828
rect 300899 587892 300965 587893
rect 300899 587828 300900 587892
rect 300964 587828 300965 587892
rect 300899 587827 300965 587828
rect 303475 587892 303541 587893
rect 303475 587828 303476 587892
rect 303540 587828 303541 587892
rect 303475 587827 303541 587828
rect 305867 587892 305933 587893
rect 305867 587828 305868 587892
rect 305932 587828 305933 587892
rect 305867 587827 305933 587828
rect 308443 587892 308509 587893
rect 308443 587828 308444 587892
rect 308508 587828 308509 587892
rect 308443 587827 308509 587828
rect 310835 587892 310901 587893
rect 310835 587828 310836 587892
rect 310900 587828 310901 587892
rect 310835 587827 310901 587828
rect 313411 587892 313477 587893
rect 313411 587828 313412 587892
rect 313476 587828 313477 587892
rect 315806 587890 315866 589870
rect 315987 587892 316053 587893
rect 315987 587890 315988 587892
rect 315806 587830 315988 587890
rect 313411 587827 313477 587828
rect 315987 587828 315988 587830
rect 316052 587828 316053 587892
rect 315987 587827 316053 587828
rect 333102 586669 333162 589870
rect 333470 587893 333530 589870
rect 333467 587892 333533 587893
rect 333467 587828 333468 587892
rect 333532 587828 333533 587892
rect 333467 587827 333533 587828
rect 293539 586668 293605 586669
rect 293539 586604 293540 586668
rect 293604 586604 293605 586668
rect 293539 586603 293605 586604
rect 295931 586668 295997 586669
rect 295931 586604 295932 586668
rect 295996 586604 295997 586668
rect 295931 586603 295997 586604
rect 333099 586668 333165 586669
rect 333099 586604 333100 586668
rect 333164 586604 333165 586668
rect 333099 586603 333165 586604
rect 277347 586532 277413 586533
rect 277347 586530 277348 586532
rect 277166 586470 277348 586530
rect 267963 586467 268029 586468
rect 277347 586468 277348 586470
rect 277412 586468 277413 586532
rect 277347 586467 277413 586468
rect 346347 582996 346413 582997
rect 346347 582932 346348 582996
rect 346412 582932 346413 582996
rect 346347 582931 346413 582932
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 562000 204914 565398
rect 346350 560149 346410 582931
rect 346347 560148 346413 560149
rect 346347 560084 346348 560148
rect 346412 560084 346413 560148
rect 346347 560083 346413 560084
rect 48270 557490 48882 557550
rect 48270 556205 48330 557490
rect 346902 556610 346962 675003
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 348371 587348 348437 587349
rect 348371 587284 348372 587348
rect 348436 587284 348437 587348
rect 348371 587283 348437 587284
rect 347819 576060 347885 576061
rect 347819 575996 347820 576060
rect 347884 575996 347885 576060
rect 347819 575995 347885 575996
rect 347635 567492 347701 567493
rect 347635 567428 347636 567492
rect 347700 567428 347701 567492
rect 347635 567427 347701 567428
rect 347638 563070 347698 567427
rect 347454 563010 347698 563070
rect 347267 560148 347333 560149
rect 347267 560084 347268 560148
rect 347332 560084 347333 560148
rect 347267 560083 347333 560084
rect 347270 557290 347330 560083
rect 347454 557970 347514 563010
rect 347635 560420 347701 560421
rect 347635 560356 347636 560420
rect 347700 560356 347701 560420
rect 347635 560355 347701 560356
rect 347638 558245 347698 560355
rect 347635 558244 347701 558245
rect 347635 558180 347636 558244
rect 347700 558180 347701 558244
rect 347635 558179 347701 558180
rect 347454 557910 347698 557970
rect 347638 557429 347698 557910
rect 347635 557428 347701 557429
rect 347635 557364 347636 557428
rect 347700 557364 347701 557428
rect 347635 557363 347701 557364
rect 347635 557292 347701 557293
rect 347635 557290 347636 557292
rect 347270 557230 347636 557290
rect 347635 557228 347636 557230
rect 347700 557228 347701 557292
rect 347635 557227 347701 557228
rect 346902 556550 347698 556610
rect 347638 556205 347698 556550
rect 48267 556204 48333 556205
rect 48267 556140 48268 556204
rect 48332 556140 48333 556204
rect 48267 556139 48333 556140
rect 347635 556204 347701 556205
rect 347635 556140 347636 556204
rect 347700 556140 347701 556204
rect 347635 556139 347701 556140
rect 67568 547954 67888 547986
rect 67568 547718 67610 547954
rect 67846 547718 67888 547954
rect 67568 547634 67888 547718
rect 67568 547398 67610 547634
rect 67846 547398 67888 547634
rect 67568 547366 67888 547398
rect 98288 547954 98608 547986
rect 98288 547718 98330 547954
rect 98566 547718 98608 547954
rect 98288 547634 98608 547718
rect 98288 547398 98330 547634
rect 98566 547398 98608 547634
rect 98288 547366 98608 547398
rect 129008 547954 129328 547986
rect 129008 547718 129050 547954
rect 129286 547718 129328 547954
rect 129008 547634 129328 547718
rect 129008 547398 129050 547634
rect 129286 547398 129328 547634
rect 129008 547366 129328 547398
rect 159728 547954 160048 547986
rect 159728 547718 159770 547954
rect 160006 547718 160048 547954
rect 159728 547634 160048 547718
rect 159728 547398 159770 547634
rect 160006 547398 160048 547634
rect 159728 547366 160048 547398
rect 190448 547954 190768 547986
rect 190448 547718 190490 547954
rect 190726 547718 190768 547954
rect 190448 547634 190768 547718
rect 190448 547398 190490 547634
rect 190726 547398 190768 547634
rect 190448 547366 190768 547398
rect 221168 547954 221488 547986
rect 221168 547718 221210 547954
rect 221446 547718 221488 547954
rect 221168 547634 221488 547718
rect 221168 547398 221210 547634
rect 221446 547398 221488 547634
rect 221168 547366 221488 547398
rect 251888 547954 252208 547986
rect 251888 547718 251930 547954
rect 252166 547718 252208 547954
rect 251888 547634 252208 547718
rect 251888 547398 251930 547634
rect 252166 547398 252208 547634
rect 251888 547366 252208 547398
rect 282608 547954 282928 547986
rect 282608 547718 282650 547954
rect 282886 547718 282928 547954
rect 282608 547634 282928 547718
rect 282608 547398 282650 547634
rect 282886 547398 282928 547634
rect 282608 547366 282928 547398
rect 313328 547954 313648 547986
rect 313328 547718 313370 547954
rect 313606 547718 313648 547954
rect 313328 547634 313648 547718
rect 313328 547398 313370 547634
rect 313606 547398 313648 547634
rect 313328 547366 313648 547398
rect 344048 547954 344368 547986
rect 344048 547718 344090 547954
rect 344326 547718 344368 547954
rect 344048 547634 344368 547718
rect 344048 547398 344090 547634
rect 344326 547398 344368 547634
rect 344048 547366 344368 547398
rect 52208 543454 52528 543486
rect 52208 543218 52250 543454
rect 52486 543218 52528 543454
rect 52208 543134 52528 543218
rect 52208 542898 52250 543134
rect 52486 542898 52528 543134
rect 52208 542866 52528 542898
rect 82928 543454 83248 543486
rect 82928 543218 82970 543454
rect 83206 543218 83248 543454
rect 82928 543134 83248 543218
rect 82928 542898 82970 543134
rect 83206 542898 83248 543134
rect 82928 542866 83248 542898
rect 113648 543454 113968 543486
rect 113648 543218 113690 543454
rect 113926 543218 113968 543454
rect 113648 543134 113968 543218
rect 113648 542898 113690 543134
rect 113926 542898 113968 543134
rect 113648 542866 113968 542898
rect 144368 543454 144688 543486
rect 144368 543218 144410 543454
rect 144646 543218 144688 543454
rect 144368 543134 144688 543218
rect 144368 542898 144410 543134
rect 144646 542898 144688 543134
rect 144368 542866 144688 542898
rect 175088 543454 175408 543486
rect 175088 543218 175130 543454
rect 175366 543218 175408 543454
rect 175088 543134 175408 543218
rect 175088 542898 175130 543134
rect 175366 542898 175408 543134
rect 175088 542866 175408 542898
rect 205808 543454 206128 543486
rect 205808 543218 205850 543454
rect 206086 543218 206128 543454
rect 205808 543134 206128 543218
rect 205808 542898 205850 543134
rect 206086 542898 206128 543134
rect 205808 542866 206128 542898
rect 236528 543454 236848 543486
rect 236528 543218 236570 543454
rect 236806 543218 236848 543454
rect 236528 543134 236848 543218
rect 236528 542898 236570 543134
rect 236806 542898 236848 543134
rect 236528 542866 236848 542898
rect 267248 543454 267568 543486
rect 267248 543218 267290 543454
rect 267526 543218 267568 543454
rect 267248 543134 267568 543218
rect 267248 542898 267290 543134
rect 267526 542898 267568 543134
rect 267248 542866 267568 542898
rect 297968 543454 298288 543486
rect 297968 543218 298010 543454
rect 298246 543218 298288 543454
rect 297968 543134 298288 543218
rect 297968 542898 298010 543134
rect 298246 542898 298288 543134
rect 297968 542866 298288 542898
rect 328688 543454 329008 543486
rect 328688 543218 328730 543454
rect 328966 543218 329008 543454
rect 328688 543134 329008 543218
rect 328688 542898 328730 543134
rect 328966 542898 329008 543134
rect 328688 542866 329008 542898
rect 67568 511954 67888 511986
rect 67568 511718 67610 511954
rect 67846 511718 67888 511954
rect 67568 511634 67888 511718
rect 67568 511398 67610 511634
rect 67846 511398 67888 511634
rect 67568 511366 67888 511398
rect 98288 511954 98608 511986
rect 98288 511718 98330 511954
rect 98566 511718 98608 511954
rect 98288 511634 98608 511718
rect 98288 511398 98330 511634
rect 98566 511398 98608 511634
rect 98288 511366 98608 511398
rect 129008 511954 129328 511986
rect 129008 511718 129050 511954
rect 129286 511718 129328 511954
rect 129008 511634 129328 511718
rect 129008 511398 129050 511634
rect 129286 511398 129328 511634
rect 129008 511366 129328 511398
rect 159728 511954 160048 511986
rect 159728 511718 159770 511954
rect 160006 511718 160048 511954
rect 159728 511634 160048 511718
rect 159728 511398 159770 511634
rect 160006 511398 160048 511634
rect 159728 511366 160048 511398
rect 190448 511954 190768 511986
rect 190448 511718 190490 511954
rect 190726 511718 190768 511954
rect 190448 511634 190768 511718
rect 190448 511398 190490 511634
rect 190726 511398 190768 511634
rect 190448 511366 190768 511398
rect 221168 511954 221488 511986
rect 221168 511718 221210 511954
rect 221446 511718 221488 511954
rect 221168 511634 221488 511718
rect 221168 511398 221210 511634
rect 221446 511398 221488 511634
rect 221168 511366 221488 511398
rect 251888 511954 252208 511986
rect 251888 511718 251930 511954
rect 252166 511718 252208 511954
rect 251888 511634 252208 511718
rect 251888 511398 251930 511634
rect 252166 511398 252208 511634
rect 251888 511366 252208 511398
rect 282608 511954 282928 511986
rect 282608 511718 282650 511954
rect 282886 511718 282928 511954
rect 282608 511634 282928 511718
rect 282608 511398 282650 511634
rect 282886 511398 282928 511634
rect 282608 511366 282928 511398
rect 313328 511954 313648 511986
rect 313328 511718 313370 511954
rect 313606 511718 313648 511954
rect 313328 511634 313648 511718
rect 313328 511398 313370 511634
rect 313606 511398 313648 511634
rect 313328 511366 313648 511398
rect 344048 511954 344368 511986
rect 344048 511718 344090 511954
rect 344326 511718 344368 511954
rect 344048 511634 344368 511718
rect 344048 511398 344090 511634
rect 344326 511398 344368 511634
rect 344048 511366 344368 511398
rect 52208 507454 52528 507486
rect 52208 507218 52250 507454
rect 52486 507218 52528 507454
rect 52208 507134 52528 507218
rect 52208 506898 52250 507134
rect 52486 506898 52528 507134
rect 52208 506866 52528 506898
rect 82928 507454 83248 507486
rect 82928 507218 82970 507454
rect 83206 507218 83248 507454
rect 82928 507134 83248 507218
rect 82928 506898 82970 507134
rect 83206 506898 83248 507134
rect 82928 506866 83248 506898
rect 113648 507454 113968 507486
rect 113648 507218 113690 507454
rect 113926 507218 113968 507454
rect 113648 507134 113968 507218
rect 113648 506898 113690 507134
rect 113926 506898 113968 507134
rect 113648 506866 113968 506898
rect 144368 507454 144688 507486
rect 144368 507218 144410 507454
rect 144646 507218 144688 507454
rect 144368 507134 144688 507218
rect 144368 506898 144410 507134
rect 144646 506898 144688 507134
rect 144368 506866 144688 506898
rect 175088 507454 175408 507486
rect 175088 507218 175130 507454
rect 175366 507218 175408 507454
rect 175088 507134 175408 507218
rect 175088 506898 175130 507134
rect 175366 506898 175408 507134
rect 175088 506866 175408 506898
rect 205808 507454 206128 507486
rect 205808 507218 205850 507454
rect 206086 507218 206128 507454
rect 205808 507134 206128 507218
rect 205808 506898 205850 507134
rect 206086 506898 206128 507134
rect 205808 506866 206128 506898
rect 236528 507454 236848 507486
rect 236528 507218 236570 507454
rect 236806 507218 236848 507454
rect 236528 507134 236848 507218
rect 236528 506898 236570 507134
rect 236806 506898 236848 507134
rect 236528 506866 236848 506898
rect 267248 507454 267568 507486
rect 267248 507218 267290 507454
rect 267526 507218 267568 507454
rect 267248 507134 267568 507218
rect 267248 506898 267290 507134
rect 267526 506898 267568 507134
rect 267248 506866 267568 506898
rect 297968 507454 298288 507486
rect 297968 507218 298010 507454
rect 298246 507218 298288 507454
rect 297968 507134 298288 507218
rect 297968 506898 298010 507134
rect 298246 506898 298288 507134
rect 297968 506866 298288 506898
rect 328688 507454 329008 507486
rect 328688 507218 328730 507454
rect 328966 507218 329008 507454
rect 328688 507134 329008 507218
rect 328688 506898 328730 507134
rect 328966 506898 329008 507134
rect 328688 506866 329008 506898
rect 67568 475954 67888 475986
rect 67568 475718 67610 475954
rect 67846 475718 67888 475954
rect 67568 475634 67888 475718
rect 67568 475398 67610 475634
rect 67846 475398 67888 475634
rect 67568 475366 67888 475398
rect 98288 475954 98608 475986
rect 98288 475718 98330 475954
rect 98566 475718 98608 475954
rect 98288 475634 98608 475718
rect 98288 475398 98330 475634
rect 98566 475398 98608 475634
rect 98288 475366 98608 475398
rect 129008 475954 129328 475986
rect 129008 475718 129050 475954
rect 129286 475718 129328 475954
rect 129008 475634 129328 475718
rect 129008 475398 129050 475634
rect 129286 475398 129328 475634
rect 129008 475366 129328 475398
rect 159728 475954 160048 475986
rect 159728 475718 159770 475954
rect 160006 475718 160048 475954
rect 159728 475634 160048 475718
rect 159728 475398 159770 475634
rect 160006 475398 160048 475634
rect 159728 475366 160048 475398
rect 190448 475954 190768 475986
rect 190448 475718 190490 475954
rect 190726 475718 190768 475954
rect 190448 475634 190768 475718
rect 190448 475398 190490 475634
rect 190726 475398 190768 475634
rect 190448 475366 190768 475398
rect 221168 475954 221488 475986
rect 221168 475718 221210 475954
rect 221446 475718 221488 475954
rect 221168 475634 221488 475718
rect 221168 475398 221210 475634
rect 221446 475398 221488 475634
rect 221168 475366 221488 475398
rect 251888 475954 252208 475986
rect 251888 475718 251930 475954
rect 252166 475718 252208 475954
rect 251888 475634 252208 475718
rect 251888 475398 251930 475634
rect 252166 475398 252208 475634
rect 251888 475366 252208 475398
rect 282608 475954 282928 475986
rect 282608 475718 282650 475954
rect 282886 475718 282928 475954
rect 282608 475634 282928 475718
rect 282608 475398 282650 475634
rect 282886 475398 282928 475634
rect 282608 475366 282928 475398
rect 313328 475954 313648 475986
rect 313328 475718 313370 475954
rect 313606 475718 313648 475954
rect 313328 475634 313648 475718
rect 313328 475398 313370 475634
rect 313606 475398 313648 475634
rect 313328 475366 313648 475398
rect 344048 475954 344368 475986
rect 344048 475718 344090 475954
rect 344326 475718 344368 475954
rect 344048 475634 344368 475718
rect 344048 475398 344090 475634
rect 344326 475398 344368 475634
rect 344048 475366 344368 475398
rect 52208 471454 52528 471486
rect 52208 471218 52250 471454
rect 52486 471218 52528 471454
rect 52208 471134 52528 471218
rect 52208 470898 52250 471134
rect 52486 470898 52528 471134
rect 52208 470866 52528 470898
rect 82928 471454 83248 471486
rect 82928 471218 82970 471454
rect 83206 471218 83248 471454
rect 82928 471134 83248 471218
rect 82928 470898 82970 471134
rect 83206 470898 83248 471134
rect 82928 470866 83248 470898
rect 113648 471454 113968 471486
rect 113648 471218 113690 471454
rect 113926 471218 113968 471454
rect 113648 471134 113968 471218
rect 113648 470898 113690 471134
rect 113926 470898 113968 471134
rect 113648 470866 113968 470898
rect 144368 471454 144688 471486
rect 144368 471218 144410 471454
rect 144646 471218 144688 471454
rect 144368 471134 144688 471218
rect 144368 470898 144410 471134
rect 144646 470898 144688 471134
rect 144368 470866 144688 470898
rect 175088 471454 175408 471486
rect 175088 471218 175130 471454
rect 175366 471218 175408 471454
rect 175088 471134 175408 471218
rect 175088 470898 175130 471134
rect 175366 470898 175408 471134
rect 175088 470866 175408 470898
rect 205808 471454 206128 471486
rect 205808 471218 205850 471454
rect 206086 471218 206128 471454
rect 205808 471134 206128 471218
rect 205808 470898 205850 471134
rect 206086 470898 206128 471134
rect 205808 470866 206128 470898
rect 236528 471454 236848 471486
rect 236528 471218 236570 471454
rect 236806 471218 236848 471454
rect 236528 471134 236848 471218
rect 236528 470898 236570 471134
rect 236806 470898 236848 471134
rect 236528 470866 236848 470898
rect 267248 471454 267568 471486
rect 267248 471218 267290 471454
rect 267526 471218 267568 471454
rect 267248 471134 267568 471218
rect 267248 470898 267290 471134
rect 267526 470898 267568 471134
rect 267248 470866 267568 470898
rect 297968 471454 298288 471486
rect 297968 471218 298010 471454
rect 298246 471218 298288 471454
rect 297968 471134 298288 471218
rect 297968 470898 298010 471134
rect 298246 470898 298288 471134
rect 297968 470866 298288 470898
rect 328688 471454 329008 471486
rect 328688 471218 328730 471454
rect 328966 471218 329008 471454
rect 328688 471134 329008 471218
rect 328688 470898 328730 471134
rect 328966 470898 329008 471134
rect 328688 470866 329008 470898
rect 67568 439954 67888 439986
rect 67568 439718 67610 439954
rect 67846 439718 67888 439954
rect 67568 439634 67888 439718
rect 67568 439398 67610 439634
rect 67846 439398 67888 439634
rect 67568 439366 67888 439398
rect 98288 439954 98608 439986
rect 98288 439718 98330 439954
rect 98566 439718 98608 439954
rect 98288 439634 98608 439718
rect 98288 439398 98330 439634
rect 98566 439398 98608 439634
rect 98288 439366 98608 439398
rect 129008 439954 129328 439986
rect 129008 439718 129050 439954
rect 129286 439718 129328 439954
rect 129008 439634 129328 439718
rect 129008 439398 129050 439634
rect 129286 439398 129328 439634
rect 129008 439366 129328 439398
rect 159728 439954 160048 439986
rect 159728 439718 159770 439954
rect 160006 439718 160048 439954
rect 159728 439634 160048 439718
rect 159728 439398 159770 439634
rect 160006 439398 160048 439634
rect 159728 439366 160048 439398
rect 190448 439954 190768 439986
rect 190448 439718 190490 439954
rect 190726 439718 190768 439954
rect 190448 439634 190768 439718
rect 190448 439398 190490 439634
rect 190726 439398 190768 439634
rect 190448 439366 190768 439398
rect 221168 439954 221488 439986
rect 221168 439718 221210 439954
rect 221446 439718 221488 439954
rect 221168 439634 221488 439718
rect 221168 439398 221210 439634
rect 221446 439398 221488 439634
rect 221168 439366 221488 439398
rect 251888 439954 252208 439986
rect 251888 439718 251930 439954
rect 252166 439718 252208 439954
rect 251888 439634 252208 439718
rect 251888 439398 251930 439634
rect 252166 439398 252208 439634
rect 251888 439366 252208 439398
rect 282608 439954 282928 439986
rect 282608 439718 282650 439954
rect 282886 439718 282928 439954
rect 282608 439634 282928 439718
rect 282608 439398 282650 439634
rect 282886 439398 282928 439634
rect 282608 439366 282928 439398
rect 313328 439954 313648 439986
rect 313328 439718 313370 439954
rect 313606 439718 313648 439954
rect 313328 439634 313648 439718
rect 313328 439398 313370 439634
rect 313606 439398 313648 439634
rect 313328 439366 313648 439398
rect 344048 439954 344368 439986
rect 344048 439718 344090 439954
rect 344326 439718 344368 439954
rect 344048 439634 344368 439718
rect 344048 439398 344090 439634
rect 344326 439398 344368 439634
rect 344048 439366 344368 439398
rect 52208 435454 52528 435486
rect 52208 435218 52250 435454
rect 52486 435218 52528 435454
rect 52208 435134 52528 435218
rect 52208 434898 52250 435134
rect 52486 434898 52528 435134
rect 52208 434866 52528 434898
rect 82928 435454 83248 435486
rect 82928 435218 82970 435454
rect 83206 435218 83248 435454
rect 82928 435134 83248 435218
rect 82928 434898 82970 435134
rect 83206 434898 83248 435134
rect 82928 434866 83248 434898
rect 113648 435454 113968 435486
rect 113648 435218 113690 435454
rect 113926 435218 113968 435454
rect 113648 435134 113968 435218
rect 113648 434898 113690 435134
rect 113926 434898 113968 435134
rect 113648 434866 113968 434898
rect 144368 435454 144688 435486
rect 144368 435218 144410 435454
rect 144646 435218 144688 435454
rect 144368 435134 144688 435218
rect 144368 434898 144410 435134
rect 144646 434898 144688 435134
rect 144368 434866 144688 434898
rect 175088 435454 175408 435486
rect 175088 435218 175130 435454
rect 175366 435218 175408 435454
rect 175088 435134 175408 435218
rect 175088 434898 175130 435134
rect 175366 434898 175408 435134
rect 175088 434866 175408 434898
rect 205808 435454 206128 435486
rect 205808 435218 205850 435454
rect 206086 435218 206128 435454
rect 205808 435134 206128 435218
rect 205808 434898 205850 435134
rect 206086 434898 206128 435134
rect 205808 434866 206128 434898
rect 236528 435454 236848 435486
rect 236528 435218 236570 435454
rect 236806 435218 236848 435454
rect 236528 435134 236848 435218
rect 236528 434898 236570 435134
rect 236806 434898 236848 435134
rect 236528 434866 236848 434898
rect 267248 435454 267568 435486
rect 267248 435218 267290 435454
rect 267526 435218 267568 435454
rect 267248 435134 267568 435218
rect 267248 434898 267290 435134
rect 267526 434898 267568 435134
rect 267248 434866 267568 434898
rect 297968 435454 298288 435486
rect 297968 435218 298010 435454
rect 298246 435218 298288 435454
rect 297968 435134 298288 435218
rect 297968 434898 298010 435134
rect 298246 434898 298288 435134
rect 297968 434866 298288 434898
rect 328688 435454 329008 435486
rect 328688 435218 328730 435454
rect 328966 435218 329008 435454
rect 328688 435134 329008 435218
rect 328688 434898 328730 435134
rect 328966 434898 329008 435134
rect 328688 434866 329008 434898
rect 47531 428568 47597 428569
rect 47531 428504 47532 428568
rect 47596 428504 47597 428568
rect 47531 428503 47597 428504
rect 47347 240956 47413 240957
rect 47347 240892 47348 240956
rect 47412 240892 47413 240956
rect 47347 240891 47413 240892
rect 47163 220556 47229 220557
rect 47163 220492 47164 220556
rect 47228 220492 47229 220556
rect 47163 220491 47229 220492
rect 46979 210356 47045 210357
rect 46979 210292 46980 210356
rect 47044 210292 47045 210356
rect 46979 210291 47045 210292
rect 47534 204509 47594 428503
rect 347822 411229 347882 575995
rect 348003 570620 348069 570621
rect 348003 570556 348004 570620
rect 348068 570556 348069 570620
rect 348003 570555 348069 570556
rect 348006 523565 348066 570555
rect 348003 523564 348069 523565
rect 348003 523500 348004 523564
rect 348068 523500 348069 523564
rect 348003 523499 348069 523500
rect 348374 456925 348434 587283
rect 351131 581636 351197 581637
rect 351131 581572 351132 581636
rect 351196 581572 351197 581636
rect 351131 581571 351197 581572
rect 349107 578916 349173 578917
rect 349107 578852 349108 578916
rect 349172 578852 349173 578916
rect 349107 578851 349173 578852
rect 348555 557428 348621 557429
rect 348555 557364 348556 557428
rect 348620 557364 348621 557428
rect 348555 557363 348621 557364
rect 348371 456924 348437 456925
rect 348371 456860 348372 456924
rect 348436 456860 348437 456924
rect 348371 456859 348437 456860
rect 348371 456788 348437 456789
rect 348371 456724 348372 456788
rect 348436 456724 348437 456788
rect 348371 456723 348437 456724
rect 347819 411228 347885 411229
rect 347819 411164 347820 411228
rect 347884 411164 347885 411228
rect 347819 411163 347885 411164
rect 67568 403954 67888 403986
rect 67568 403718 67610 403954
rect 67846 403718 67888 403954
rect 67568 403634 67888 403718
rect 67568 403398 67610 403634
rect 67846 403398 67888 403634
rect 67568 403366 67888 403398
rect 98288 403954 98608 403986
rect 98288 403718 98330 403954
rect 98566 403718 98608 403954
rect 98288 403634 98608 403718
rect 98288 403398 98330 403634
rect 98566 403398 98608 403634
rect 98288 403366 98608 403398
rect 129008 403954 129328 403986
rect 129008 403718 129050 403954
rect 129286 403718 129328 403954
rect 129008 403634 129328 403718
rect 129008 403398 129050 403634
rect 129286 403398 129328 403634
rect 129008 403366 129328 403398
rect 159728 403954 160048 403986
rect 159728 403718 159770 403954
rect 160006 403718 160048 403954
rect 159728 403634 160048 403718
rect 159728 403398 159770 403634
rect 160006 403398 160048 403634
rect 159728 403366 160048 403398
rect 190448 403954 190768 403986
rect 190448 403718 190490 403954
rect 190726 403718 190768 403954
rect 190448 403634 190768 403718
rect 190448 403398 190490 403634
rect 190726 403398 190768 403634
rect 190448 403366 190768 403398
rect 221168 403954 221488 403986
rect 221168 403718 221210 403954
rect 221446 403718 221488 403954
rect 221168 403634 221488 403718
rect 221168 403398 221210 403634
rect 221446 403398 221488 403634
rect 221168 403366 221488 403398
rect 251888 403954 252208 403986
rect 251888 403718 251930 403954
rect 252166 403718 252208 403954
rect 251888 403634 252208 403718
rect 251888 403398 251930 403634
rect 252166 403398 252208 403634
rect 251888 403366 252208 403398
rect 282608 403954 282928 403986
rect 282608 403718 282650 403954
rect 282886 403718 282928 403954
rect 282608 403634 282928 403718
rect 282608 403398 282650 403634
rect 282886 403398 282928 403634
rect 282608 403366 282928 403398
rect 313328 403954 313648 403986
rect 313328 403718 313370 403954
rect 313606 403718 313648 403954
rect 313328 403634 313648 403718
rect 313328 403398 313370 403634
rect 313606 403398 313648 403634
rect 313328 403366 313648 403398
rect 344048 403954 344368 403986
rect 344048 403718 344090 403954
rect 344326 403718 344368 403954
rect 344048 403634 344368 403718
rect 344048 403398 344090 403634
rect 344326 403398 344368 403634
rect 344048 403366 344368 403398
rect 52208 399454 52528 399486
rect 52208 399218 52250 399454
rect 52486 399218 52528 399454
rect 52208 399134 52528 399218
rect 52208 398898 52250 399134
rect 52486 398898 52528 399134
rect 52208 398866 52528 398898
rect 82928 399454 83248 399486
rect 82928 399218 82970 399454
rect 83206 399218 83248 399454
rect 82928 399134 83248 399218
rect 82928 398898 82970 399134
rect 83206 398898 83248 399134
rect 82928 398866 83248 398898
rect 113648 399454 113968 399486
rect 113648 399218 113690 399454
rect 113926 399218 113968 399454
rect 113648 399134 113968 399218
rect 113648 398898 113690 399134
rect 113926 398898 113968 399134
rect 113648 398866 113968 398898
rect 144368 399454 144688 399486
rect 144368 399218 144410 399454
rect 144646 399218 144688 399454
rect 144368 399134 144688 399218
rect 144368 398898 144410 399134
rect 144646 398898 144688 399134
rect 144368 398866 144688 398898
rect 175088 399454 175408 399486
rect 175088 399218 175130 399454
rect 175366 399218 175408 399454
rect 175088 399134 175408 399218
rect 175088 398898 175130 399134
rect 175366 398898 175408 399134
rect 175088 398866 175408 398898
rect 205808 399454 206128 399486
rect 205808 399218 205850 399454
rect 206086 399218 206128 399454
rect 205808 399134 206128 399218
rect 205808 398898 205850 399134
rect 206086 398898 206128 399134
rect 205808 398866 206128 398898
rect 236528 399454 236848 399486
rect 236528 399218 236570 399454
rect 236806 399218 236848 399454
rect 236528 399134 236848 399218
rect 236528 398898 236570 399134
rect 236806 398898 236848 399134
rect 236528 398866 236848 398898
rect 267248 399454 267568 399486
rect 267248 399218 267290 399454
rect 267526 399218 267568 399454
rect 267248 399134 267568 399218
rect 267248 398898 267290 399134
rect 267526 398898 267568 399134
rect 267248 398866 267568 398898
rect 297968 399454 298288 399486
rect 297968 399218 298010 399454
rect 298246 399218 298288 399454
rect 297968 399134 298288 399218
rect 297968 398898 298010 399134
rect 298246 398898 298288 399134
rect 297968 398866 298288 398898
rect 328688 399454 329008 399486
rect 328688 399218 328730 399454
rect 328966 399218 329008 399454
rect 328688 399134 329008 399218
rect 328688 398898 328730 399134
rect 328966 398898 329008 399134
rect 328688 398866 329008 398898
rect 67568 367954 67888 367986
rect 67568 367718 67610 367954
rect 67846 367718 67888 367954
rect 67568 367634 67888 367718
rect 67568 367398 67610 367634
rect 67846 367398 67888 367634
rect 67568 367366 67888 367398
rect 98288 367954 98608 367986
rect 98288 367718 98330 367954
rect 98566 367718 98608 367954
rect 98288 367634 98608 367718
rect 98288 367398 98330 367634
rect 98566 367398 98608 367634
rect 98288 367366 98608 367398
rect 129008 367954 129328 367986
rect 129008 367718 129050 367954
rect 129286 367718 129328 367954
rect 129008 367634 129328 367718
rect 129008 367398 129050 367634
rect 129286 367398 129328 367634
rect 129008 367366 129328 367398
rect 159728 367954 160048 367986
rect 159728 367718 159770 367954
rect 160006 367718 160048 367954
rect 159728 367634 160048 367718
rect 159728 367398 159770 367634
rect 160006 367398 160048 367634
rect 159728 367366 160048 367398
rect 190448 367954 190768 367986
rect 190448 367718 190490 367954
rect 190726 367718 190768 367954
rect 190448 367634 190768 367718
rect 190448 367398 190490 367634
rect 190726 367398 190768 367634
rect 190448 367366 190768 367398
rect 221168 367954 221488 367986
rect 221168 367718 221210 367954
rect 221446 367718 221488 367954
rect 221168 367634 221488 367718
rect 221168 367398 221210 367634
rect 221446 367398 221488 367634
rect 221168 367366 221488 367398
rect 251888 367954 252208 367986
rect 251888 367718 251930 367954
rect 252166 367718 252208 367954
rect 251888 367634 252208 367718
rect 251888 367398 251930 367634
rect 252166 367398 252208 367634
rect 251888 367366 252208 367398
rect 282608 367954 282928 367986
rect 282608 367718 282650 367954
rect 282886 367718 282928 367954
rect 282608 367634 282928 367718
rect 282608 367398 282650 367634
rect 282886 367398 282928 367634
rect 282608 367366 282928 367398
rect 313328 367954 313648 367986
rect 313328 367718 313370 367954
rect 313606 367718 313648 367954
rect 313328 367634 313648 367718
rect 313328 367398 313370 367634
rect 313606 367398 313648 367634
rect 313328 367366 313648 367398
rect 344048 367954 344368 367986
rect 344048 367718 344090 367954
rect 344326 367718 344368 367954
rect 344048 367634 344368 367718
rect 344048 367398 344090 367634
rect 344326 367398 344368 367634
rect 344048 367366 344368 367398
rect 52208 363454 52528 363486
rect 52208 363218 52250 363454
rect 52486 363218 52528 363454
rect 52208 363134 52528 363218
rect 52208 362898 52250 363134
rect 52486 362898 52528 363134
rect 52208 362866 52528 362898
rect 82928 363454 83248 363486
rect 82928 363218 82970 363454
rect 83206 363218 83248 363454
rect 82928 363134 83248 363218
rect 82928 362898 82970 363134
rect 83206 362898 83248 363134
rect 82928 362866 83248 362898
rect 113648 363454 113968 363486
rect 113648 363218 113690 363454
rect 113926 363218 113968 363454
rect 113648 363134 113968 363218
rect 113648 362898 113690 363134
rect 113926 362898 113968 363134
rect 113648 362866 113968 362898
rect 144368 363454 144688 363486
rect 144368 363218 144410 363454
rect 144646 363218 144688 363454
rect 144368 363134 144688 363218
rect 144368 362898 144410 363134
rect 144646 362898 144688 363134
rect 144368 362866 144688 362898
rect 175088 363454 175408 363486
rect 175088 363218 175130 363454
rect 175366 363218 175408 363454
rect 175088 363134 175408 363218
rect 175088 362898 175130 363134
rect 175366 362898 175408 363134
rect 175088 362866 175408 362898
rect 205808 363454 206128 363486
rect 205808 363218 205850 363454
rect 206086 363218 206128 363454
rect 205808 363134 206128 363218
rect 205808 362898 205850 363134
rect 206086 362898 206128 363134
rect 205808 362866 206128 362898
rect 236528 363454 236848 363486
rect 236528 363218 236570 363454
rect 236806 363218 236848 363454
rect 236528 363134 236848 363218
rect 236528 362898 236570 363134
rect 236806 362898 236848 363134
rect 236528 362866 236848 362898
rect 267248 363454 267568 363486
rect 267248 363218 267290 363454
rect 267526 363218 267568 363454
rect 267248 363134 267568 363218
rect 267248 362898 267290 363134
rect 267526 362898 267568 363134
rect 267248 362866 267568 362898
rect 297968 363454 298288 363486
rect 297968 363218 298010 363454
rect 298246 363218 298288 363454
rect 297968 363134 298288 363218
rect 297968 362898 298010 363134
rect 298246 362898 298288 363134
rect 297968 362866 298288 362898
rect 328688 363454 329008 363486
rect 328688 363218 328730 363454
rect 328966 363218 329008 363454
rect 328688 363134 329008 363218
rect 328688 362898 328730 363134
rect 328966 362898 329008 363134
rect 328688 362866 329008 362898
rect 67568 331954 67888 331986
rect 67568 331718 67610 331954
rect 67846 331718 67888 331954
rect 67568 331634 67888 331718
rect 67568 331398 67610 331634
rect 67846 331398 67888 331634
rect 67568 331366 67888 331398
rect 98288 331954 98608 331986
rect 98288 331718 98330 331954
rect 98566 331718 98608 331954
rect 98288 331634 98608 331718
rect 98288 331398 98330 331634
rect 98566 331398 98608 331634
rect 98288 331366 98608 331398
rect 129008 331954 129328 331986
rect 129008 331718 129050 331954
rect 129286 331718 129328 331954
rect 129008 331634 129328 331718
rect 129008 331398 129050 331634
rect 129286 331398 129328 331634
rect 129008 331366 129328 331398
rect 159728 331954 160048 331986
rect 159728 331718 159770 331954
rect 160006 331718 160048 331954
rect 159728 331634 160048 331718
rect 159728 331398 159770 331634
rect 160006 331398 160048 331634
rect 159728 331366 160048 331398
rect 190448 331954 190768 331986
rect 190448 331718 190490 331954
rect 190726 331718 190768 331954
rect 190448 331634 190768 331718
rect 190448 331398 190490 331634
rect 190726 331398 190768 331634
rect 190448 331366 190768 331398
rect 221168 331954 221488 331986
rect 221168 331718 221210 331954
rect 221446 331718 221488 331954
rect 221168 331634 221488 331718
rect 221168 331398 221210 331634
rect 221446 331398 221488 331634
rect 221168 331366 221488 331398
rect 251888 331954 252208 331986
rect 251888 331718 251930 331954
rect 252166 331718 252208 331954
rect 251888 331634 252208 331718
rect 251888 331398 251930 331634
rect 252166 331398 252208 331634
rect 251888 331366 252208 331398
rect 282608 331954 282928 331986
rect 282608 331718 282650 331954
rect 282886 331718 282928 331954
rect 282608 331634 282928 331718
rect 282608 331398 282650 331634
rect 282886 331398 282928 331634
rect 282608 331366 282928 331398
rect 313328 331954 313648 331986
rect 313328 331718 313370 331954
rect 313606 331718 313648 331954
rect 313328 331634 313648 331718
rect 313328 331398 313370 331634
rect 313606 331398 313648 331634
rect 313328 331366 313648 331398
rect 344048 331954 344368 331986
rect 344048 331718 344090 331954
rect 344326 331718 344368 331954
rect 344048 331634 344368 331718
rect 344048 331398 344090 331634
rect 344326 331398 344368 331634
rect 344048 331366 344368 331398
rect 52208 327454 52528 327486
rect 52208 327218 52250 327454
rect 52486 327218 52528 327454
rect 52208 327134 52528 327218
rect 52208 326898 52250 327134
rect 52486 326898 52528 327134
rect 52208 326866 52528 326898
rect 82928 327454 83248 327486
rect 82928 327218 82970 327454
rect 83206 327218 83248 327454
rect 82928 327134 83248 327218
rect 82928 326898 82970 327134
rect 83206 326898 83248 327134
rect 82928 326866 83248 326898
rect 113648 327454 113968 327486
rect 113648 327218 113690 327454
rect 113926 327218 113968 327454
rect 113648 327134 113968 327218
rect 113648 326898 113690 327134
rect 113926 326898 113968 327134
rect 113648 326866 113968 326898
rect 144368 327454 144688 327486
rect 144368 327218 144410 327454
rect 144646 327218 144688 327454
rect 144368 327134 144688 327218
rect 144368 326898 144410 327134
rect 144646 326898 144688 327134
rect 144368 326866 144688 326898
rect 175088 327454 175408 327486
rect 175088 327218 175130 327454
rect 175366 327218 175408 327454
rect 175088 327134 175408 327218
rect 175088 326898 175130 327134
rect 175366 326898 175408 327134
rect 175088 326866 175408 326898
rect 205808 327454 206128 327486
rect 205808 327218 205850 327454
rect 206086 327218 206128 327454
rect 205808 327134 206128 327218
rect 205808 326898 205850 327134
rect 206086 326898 206128 327134
rect 205808 326866 206128 326898
rect 236528 327454 236848 327486
rect 236528 327218 236570 327454
rect 236806 327218 236848 327454
rect 236528 327134 236848 327218
rect 236528 326898 236570 327134
rect 236806 326898 236848 327134
rect 236528 326866 236848 326898
rect 267248 327454 267568 327486
rect 267248 327218 267290 327454
rect 267526 327218 267568 327454
rect 267248 327134 267568 327218
rect 267248 326898 267290 327134
rect 267526 326898 267568 327134
rect 267248 326866 267568 326898
rect 297968 327454 298288 327486
rect 297968 327218 298010 327454
rect 298246 327218 298288 327454
rect 297968 327134 298288 327218
rect 297968 326898 298010 327134
rect 298246 326898 298288 327134
rect 297968 326866 298288 326898
rect 328688 327454 329008 327486
rect 328688 327218 328730 327454
rect 328966 327218 329008 327454
rect 328688 327134 329008 327218
rect 328688 326898 328730 327134
rect 328966 326898 329008 327134
rect 328688 326866 329008 326898
rect 67568 295954 67888 295986
rect 67568 295718 67610 295954
rect 67846 295718 67888 295954
rect 67568 295634 67888 295718
rect 67568 295398 67610 295634
rect 67846 295398 67888 295634
rect 67568 295366 67888 295398
rect 98288 295954 98608 295986
rect 98288 295718 98330 295954
rect 98566 295718 98608 295954
rect 98288 295634 98608 295718
rect 98288 295398 98330 295634
rect 98566 295398 98608 295634
rect 98288 295366 98608 295398
rect 129008 295954 129328 295986
rect 129008 295718 129050 295954
rect 129286 295718 129328 295954
rect 129008 295634 129328 295718
rect 129008 295398 129050 295634
rect 129286 295398 129328 295634
rect 129008 295366 129328 295398
rect 159728 295954 160048 295986
rect 159728 295718 159770 295954
rect 160006 295718 160048 295954
rect 159728 295634 160048 295718
rect 159728 295398 159770 295634
rect 160006 295398 160048 295634
rect 159728 295366 160048 295398
rect 190448 295954 190768 295986
rect 190448 295718 190490 295954
rect 190726 295718 190768 295954
rect 190448 295634 190768 295718
rect 190448 295398 190490 295634
rect 190726 295398 190768 295634
rect 190448 295366 190768 295398
rect 221168 295954 221488 295986
rect 221168 295718 221210 295954
rect 221446 295718 221488 295954
rect 221168 295634 221488 295718
rect 221168 295398 221210 295634
rect 221446 295398 221488 295634
rect 221168 295366 221488 295398
rect 251888 295954 252208 295986
rect 251888 295718 251930 295954
rect 252166 295718 252208 295954
rect 251888 295634 252208 295718
rect 251888 295398 251930 295634
rect 252166 295398 252208 295634
rect 251888 295366 252208 295398
rect 282608 295954 282928 295986
rect 282608 295718 282650 295954
rect 282886 295718 282928 295954
rect 282608 295634 282928 295718
rect 282608 295398 282650 295634
rect 282886 295398 282928 295634
rect 282608 295366 282928 295398
rect 313328 295954 313648 295986
rect 313328 295718 313370 295954
rect 313606 295718 313648 295954
rect 313328 295634 313648 295718
rect 313328 295398 313370 295634
rect 313606 295398 313648 295634
rect 313328 295366 313648 295398
rect 344048 295954 344368 295986
rect 344048 295718 344090 295954
rect 344326 295718 344368 295954
rect 344048 295634 344368 295718
rect 344048 295398 344090 295634
rect 344326 295398 344368 295634
rect 344048 295366 344368 295398
rect 52208 291454 52528 291486
rect 52208 291218 52250 291454
rect 52486 291218 52528 291454
rect 52208 291134 52528 291218
rect 52208 290898 52250 291134
rect 52486 290898 52528 291134
rect 52208 290866 52528 290898
rect 82928 291454 83248 291486
rect 82928 291218 82970 291454
rect 83206 291218 83248 291454
rect 82928 291134 83248 291218
rect 82928 290898 82970 291134
rect 83206 290898 83248 291134
rect 82928 290866 83248 290898
rect 113648 291454 113968 291486
rect 113648 291218 113690 291454
rect 113926 291218 113968 291454
rect 113648 291134 113968 291218
rect 113648 290898 113690 291134
rect 113926 290898 113968 291134
rect 113648 290866 113968 290898
rect 144368 291454 144688 291486
rect 144368 291218 144410 291454
rect 144646 291218 144688 291454
rect 144368 291134 144688 291218
rect 144368 290898 144410 291134
rect 144646 290898 144688 291134
rect 144368 290866 144688 290898
rect 175088 291454 175408 291486
rect 175088 291218 175130 291454
rect 175366 291218 175408 291454
rect 175088 291134 175408 291218
rect 175088 290898 175130 291134
rect 175366 290898 175408 291134
rect 175088 290866 175408 290898
rect 205808 291454 206128 291486
rect 205808 291218 205850 291454
rect 206086 291218 206128 291454
rect 205808 291134 206128 291218
rect 205808 290898 205850 291134
rect 206086 290898 206128 291134
rect 205808 290866 206128 290898
rect 236528 291454 236848 291486
rect 236528 291218 236570 291454
rect 236806 291218 236848 291454
rect 236528 291134 236848 291218
rect 236528 290898 236570 291134
rect 236806 290898 236848 291134
rect 236528 290866 236848 290898
rect 267248 291454 267568 291486
rect 267248 291218 267290 291454
rect 267526 291218 267568 291454
rect 267248 291134 267568 291218
rect 267248 290898 267290 291134
rect 267526 290898 267568 291134
rect 267248 290866 267568 290898
rect 297968 291454 298288 291486
rect 297968 291218 298010 291454
rect 298246 291218 298288 291454
rect 297968 291134 298288 291218
rect 297968 290898 298010 291134
rect 298246 290898 298288 291134
rect 297968 290866 298288 290898
rect 328688 291454 329008 291486
rect 328688 291218 328730 291454
rect 328966 291218 329008 291454
rect 328688 291134 329008 291218
rect 328688 290898 328730 291134
rect 328966 290898 329008 291134
rect 328688 290866 329008 290898
rect 67568 259954 67888 259986
rect 67568 259718 67610 259954
rect 67846 259718 67888 259954
rect 67568 259634 67888 259718
rect 67568 259398 67610 259634
rect 67846 259398 67888 259634
rect 67568 259366 67888 259398
rect 98288 259954 98608 259986
rect 98288 259718 98330 259954
rect 98566 259718 98608 259954
rect 98288 259634 98608 259718
rect 98288 259398 98330 259634
rect 98566 259398 98608 259634
rect 98288 259366 98608 259398
rect 129008 259954 129328 259986
rect 129008 259718 129050 259954
rect 129286 259718 129328 259954
rect 129008 259634 129328 259718
rect 129008 259398 129050 259634
rect 129286 259398 129328 259634
rect 129008 259366 129328 259398
rect 159728 259954 160048 259986
rect 159728 259718 159770 259954
rect 160006 259718 160048 259954
rect 159728 259634 160048 259718
rect 159728 259398 159770 259634
rect 160006 259398 160048 259634
rect 159728 259366 160048 259398
rect 190448 259954 190768 259986
rect 190448 259718 190490 259954
rect 190726 259718 190768 259954
rect 190448 259634 190768 259718
rect 190448 259398 190490 259634
rect 190726 259398 190768 259634
rect 190448 259366 190768 259398
rect 221168 259954 221488 259986
rect 221168 259718 221210 259954
rect 221446 259718 221488 259954
rect 221168 259634 221488 259718
rect 221168 259398 221210 259634
rect 221446 259398 221488 259634
rect 221168 259366 221488 259398
rect 251888 259954 252208 259986
rect 251888 259718 251930 259954
rect 252166 259718 252208 259954
rect 251888 259634 252208 259718
rect 251888 259398 251930 259634
rect 252166 259398 252208 259634
rect 251888 259366 252208 259398
rect 282608 259954 282928 259986
rect 282608 259718 282650 259954
rect 282886 259718 282928 259954
rect 282608 259634 282928 259718
rect 282608 259398 282650 259634
rect 282886 259398 282928 259634
rect 282608 259366 282928 259398
rect 313328 259954 313648 259986
rect 313328 259718 313370 259954
rect 313606 259718 313648 259954
rect 313328 259634 313648 259718
rect 313328 259398 313370 259634
rect 313606 259398 313648 259634
rect 313328 259366 313648 259398
rect 344048 259954 344368 259986
rect 344048 259718 344090 259954
rect 344326 259718 344368 259954
rect 344048 259634 344368 259718
rect 344048 259398 344090 259634
rect 344326 259398 344368 259634
rect 344048 259366 344368 259398
rect 52208 255454 52528 255486
rect 52208 255218 52250 255454
rect 52486 255218 52528 255454
rect 52208 255134 52528 255218
rect 52208 254898 52250 255134
rect 52486 254898 52528 255134
rect 52208 254866 52528 254898
rect 82928 255454 83248 255486
rect 82928 255218 82970 255454
rect 83206 255218 83248 255454
rect 82928 255134 83248 255218
rect 82928 254898 82970 255134
rect 83206 254898 83248 255134
rect 82928 254866 83248 254898
rect 113648 255454 113968 255486
rect 113648 255218 113690 255454
rect 113926 255218 113968 255454
rect 113648 255134 113968 255218
rect 113648 254898 113690 255134
rect 113926 254898 113968 255134
rect 113648 254866 113968 254898
rect 144368 255454 144688 255486
rect 144368 255218 144410 255454
rect 144646 255218 144688 255454
rect 144368 255134 144688 255218
rect 144368 254898 144410 255134
rect 144646 254898 144688 255134
rect 144368 254866 144688 254898
rect 175088 255454 175408 255486
rect 175088 255218 175130 255454
rect 175366 255218 175408 255454
rect 175088 255134 175408 255218
rect 175088 254898 175130 255134
rect 175366 254898 175408 255134
rect 175088 254866 175408 254898
rect 205808 255454 206128 255486
rect 205808 255218 205850 255454
rect 206086 255218 206128 255454
rect 205808 255134 206128 255218
rect 205808 254898 205850 255134
rect 206086 254898 206128 255134
rect 205808 254866 206128 254898
rect 236528 255454 236848 255486
rect 236528 255218 236570 255454
rect 236806 255218 236848 255454
rect 236528 255134 236848 255218
rect 236528 254898 236570 255134
rect 236806 254898 236848 255134
rect 236528 254866 236848 254898
rect 267248 255454 267568 255486
rect 267248 255218 267290 255454
rect 267526 255218 267568 255454
rect 267248 255134 267568 255218
rect 267248 254898 267290 255134
rect 267526 254898 267568 255134
rect 267248 254866 267568 254898
rect 297968 255454 298288 255486
rect 297968 255218 298010 255454
rect 298246 255218 298288 255454
rect 297968 255134 298288 255218
rect 297968 254898 298010 255134
rect 298246 254898 298288 255134
rect 297968 254866 298288 254898
rect 328688 255454 329008 255486
rect 328688 255218 328730 255454
rect 328966 255218 329008 255454
rect 328688 255134 329008 255218
rect 328688 254898 328730 255134
rect 328966 254898 329008 255134
rect 328688 254866 329008 254898
rect 47715 241500 47781 241501
rect 47715 241436 47716 241500
rect 47780 241436 47781 241500
rect 47715 241435 47781 241436
rect 47718 226405 47778 241435
rect 47715 226404 47781 226405
rect 47715 226340 47716 226404
rect 47780 226340 47781 226404
rect 47715 226339 47781 226340
rect 67568 223954 67888 223986
rect 67568 223718 67610 223954
rect 67846 223718 67888 223954
rect 67568 223634 67888 223718
rect 67568 223398 67610 223634
rect 67846 223398 67888 223634
rect 67568 223366 67888 223398
rect 98288 223954 98608 223986
rect 98288 223718 98330 223954
rect 98566 223718 98608 223954
rect 98288 223634 98608 223718
rect 98288 223398 98330 223634
rect 98566 223398 98608 223634
rect 98288 223366 98608 223398
rect 129008 223954 129328 223986
rect 129008 223718 129050 223954
rect 129286 223718 129328 223954
rect 129008 223634 129328 223718
rect 129008 223398 129050 223634
rect 129286 223398 129328 223634
rect 129008 223366 129328 223398
rect 159728 223954 160048 223986
rect 159728 223718 159770 223954
rect 160006 223718 160048 223954
rect 159728 223634 160048 223718
rect 159728 223398 159770 223634
rect 160006 223398 160048 223634
rect 159728 223366 160048 223398
rect 190448 223954 190768 223986
rect 190448 223718 190490 223954
rect 190726 223718 190768 223954
rect 190448 223634 190768 223718
rect 190448 223398 190490 223634
rect 190726 223398 190768 223634
rect 190448 223366 190768 223398
rect 221168 223954 221488 223986
rect 221168 223718 221210 223954
rect 221446 223718 221488 223954
rect 221168 223634 221488 223718
rect 221168 223398 221210 223634
rect 221446 223398 221488 223634
rect 221168 223366 221488 223398
rect 251888 223954 252208 223986
rect 251888 223718 251930 223954
rect 252166 223718 252208 223954
rect 251888 223634 252208 223718
rect 251888 223398 251930 223634
rect 252166 223398 252208 223634
rect 251888 223366 252208 223398
rect 282608 223954 282928 223986
rect 282608 223718 282650 223954
rect 282886 223718 282928 223954
rect 282608 223634 282928 223718
rect 282608 223398 282650 223634
rect 282886 223398 282928 223634
rect 282608 223366 282928 223398
rect 313328 223954 313648 223986
rect 313328 223718 313370 223954
rect 313606 223718 313648 223954
rect 313328 223634 313648 223718
rect 313328 223398 313370 223634
rect 313606 223398 313648 223634
rect 313328 223366 313648 223398
rect 344048 223954 344368 223986
rect 344048 223718 344090 223954
rect 344326 223718 344368 223954
rect 344048 223634 344368 223718
rect 344048 223398 344090 223634
rect 344326 223398 344368 223634
rect 344048 223366 344368 223398
rect 47715 222188 47781 222189
rect 47715 222124 47716 222188
rect 47780 222124 47781 222188
rect 47715 222123 47781 222124
rect 47531 204508 47597 204509
rect 47531 204444 47532 204508
rect 47596 204444 47597 204508
rect 47531 204443 47597 204444
rect 47531 204372 47597 204373
rect 47531 204308 47532 204372
rect 47596 204308 47597 204372
rect 47531 204307 47597 204308
rect 46794 192454 47414 198000
rect 47534 197981 47594 204307
rect 47531 197980 47597 197981
rect 47531 197916 47532 197980
rect 47596 197916 47597 197980
rect 47531 197915 47597 197916
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46611 174724 46677 174725
rect 46611 174660 46612 174724
rect 46676 174660 46677 174724
rect 46611 174659 46677 174660
rect 46427 158268 46493 158269
rect 46427 158204 46428 158268
rect 46492 158204 46493 158268
rect 46427 158203 46493 158204
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46427 155956 46493 155957
rect 46427 155892 46428 155956
rect 46492 155892 46493 155956
rect 46427 155891 46493 155892
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46430 123589 46490 155891
rect 46427 123588 46493 123589
rect 46427 123524 46428 123588
rect 46492 123524 46493 123588
rect 46427 123523 46493 123524
rect 46243 123452 46309 123453
rect 46243 123388 46244 123452
rect 46308 123388 46309 123452
rect 46243 123387 46309 123388
rect 46794 120454 47414 155898
rect 47718 152829 47778 222123
rect 48083 220284 48149 220285
rect 48083 220220 48084 220284
rect 48148 220220 48149 220284
rect 48083 220219 48149 220220
rect 47899 204508 47965 204509
rect 47899 204444 47900 204508
rect 47964 204444 47965 204508
rect 47899 204443 47965 204444
rect 47902 196621 47962 204443
rect 47899 196620 47965 196621
rect 47899 196556 47900 196620
rect 47964 196556 47965 196620
rect 47899 196555 47965 196556
rect 47899 188732 47965 188733
rect 47899 188668 47900 188732
rect 47964 188668 47965 188732
rect 47899 188667 47965 188668
rect 47715 152828 47781 152829
rect 47715 152764 47716 152828
rect 47780 152764 47781 152828
rect 47715 152763 47781 152764
rect 47715 147796 47781 147797
rect 47715 147732 47716 147796
rect 47780 147732 47781 147796
rect 47715 147731 47781 147732
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 45875 30972 45941 30973
rect 45875 30908 45876 30972
rect 45940 30908 45941 30972
rect 45875 30907 45941 30908
rect 45323 28116 45389 28117
rect 45323 28052 45324 28116
rect 45388 28052 45389 28116
rect 45323 28051 45389 28052
rect 44955 27300 45021 27301
rect 44955 27236 44956 27300
rect 45020 27236 45021 27300
rect 44955 27235 45021 27236
rect 44771 18868 44837 18869
rect 44771 18804 44772 18868
rect 44836 18804 44837 18868
rect 44771 18803 44837 18804
rect 46794 12454 47414 47898
rect 47718 19141 47778 147731
rect 47715 19140 47781 19141
rect 47715 19076 47716 19140
rect 47780 19076 47781 19140
rect 47715 19075 47781 19076
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 43667 3500 43733 3501
rect 43667 3436 43668 3500
rect 43732 3436 43733 3500
rect 43667 3435 43733 3436
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 -2266 47414 11898
rect 47902 3637 47962 188667
rect 48086 22677 48146 220219
rect 52208 219454 52528 219486
rect 52208 219218 52250 219454
rect 52486 219218 52528 219454
rect 52208 219134 52528 219218
rect 52208 218898 52250 219134
rect 52486 218898 52528 219134
rect 52208 218866 52528 218898
rect 82928 219454 83248 219486
rect 82928 219218 82970 219454
rect 83206 219218 83248 219454
rect 82928 219134 83248 219218
rect 82928 218898 82970 219134
rect 83206 218898 83248 219134
rect 82928 218866 83248 218898
rect 113648 219454 113968 219486
rect 113648 219218 113690 219454
rect 113926 219218 113968 219454
rect 113648 219134 113968 219218
rect 113648 218898 113690 219134
rect 113926 218898 113968 219134
rect 113648 218866 113968 218898
rect 144368 219454 144688 219486
rect 144368 219218 144410 219454
rect 144646 219218 144688 219454
rect 144368 219134 144688 219218
rect 144368 218898 144410 219134
rect 144646 218898 144688 219134
rect 144368 218866 144688 218898
rect 175088 219454 175408 219486
rect 175088 219218 175130 219454
rect 175366 219218 175408 219454
rect 175088 219134 175408 219218
rect 175088 218898 175130 219134
rect 175366 218898 175408 219134
rect 175088 218866 175408 218898
rect 205808 219454 206128 219486
rect 205808 219218 205850 219454
rect 206086 219218 206128 219454
rect 205808 219134 206128 219218
rect 205808 218898 205850 219134
rect 206086 218898 206128 219134
rect 205808 218866 206128 218898
rect 236528 219454 236848 219486
rect 236528 219218 236570 219454
rect 236806 219218 236848 219454
rect 236528 219134 236848 219218
rect 236528 218898 236570 219134
rect 236806 218898 236848 219134
rect 236528 218866 236848 218898
rect 267248 219454 267568 219486
rect 267248 219218 267290 219454
rect 267526 219218 267568 219454
rect 267248 219134 267568 219218
rect 267248 218898 267290 219134
rect 267526 218898 267568 219134
rect 267248 218866 267568 218898
rect 297968 219454 298288 219486
rect 297968 219218 298010 219454
rect 298246 219218 298288 219454
rect 297968 219134 298288 219218
rect 297968 218898 298010 219134
rect 298246 218898 298288 219134
rect 297968 218866 298288 218898
rect 328688 219454 329008 219486
rect 328688 219218 328730 219454
rect 328966 219218 329008 219454
rect 328688 219134 329008 219218
rect 328688 218898 328730 219134
rect 328966 218898 329008 219134
rect 328688 218866 329008 218898
rect 48267 201652 48333 201653
rect 48267 201588 48268 201652
rect 48332 201588 48333 201652
rect 48267 201587 48333 201588
rect 48270 200970 48330 201587
rect 347819 201108 347885 201109
rect 347819 201044 347820 201108
rect 347884 201044 347885 201108
rect 347819 201043 347885 201044
rect 347822 200970 347882 201043
rect 48270 200910 48514 200970
rect 48267 200564 48333 200565
rect 48267 200500 48268 200564
rect 48332 200500 48333 200564
rect 48267 200499 48333 200500
rect 48270 194037 48330 200499
rect 48454 195990 48514 200910
rect 346902 200910 347882 200970
rect 49003 199612 49069 199613
rect 49003 199548 49004 199612
rect 49068 199548 49069 199612
rect 49003 199547 49069 199548
rect 48454 195930 48882 195990
rect 48267 194036 48333 194037
rect 48267 193972 48268 194036
rect 48332 193972 48333 194036
rect 48267 193971 48333 193972
rect 48822 152965 48882 195930
rect 49006 192949 49066 199547
rect 51294 196954 51914 198000
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 49003 192948 49069 192949
rect 49003 192884 49004 192948
rect 49068 192884 49069 192948
rect 49003 192883 49069 192884
rect 50475 190092 50541 190093
rect 50475 190028 50476 190092
rect 50540 190028 50541 190092
rect 50475 190027 50541 190028
rect 49555 185876 49621 185877
rect 49555 185812 49556 185876
rect 49620 185812 49621 185876
rect 49555 185811 49621 185812
rect 49371 180436 49437 180437
rect 49371 180372 49372 180436
rect 49436 180372 49437 180436
rect 49371 180371 49437 180372
rect 49187 177444 49253 177445
rect 49187 177380 49188 177444
rect 49252 177380 49253 177444
rect 49187 177379 49253 177380
rect 48819 152964 48885 152965
rect 48819 152900 48820 152964
rect 48884 152900 48885 152964
rect 48819 152899 48885 152900
rect 49003 149156 49069 149157
rect 49003 149092 49004 149156
rect 49068 149092 49069 149156
rect 49003 149091 49069 149092
rect 49006 27573 49066 149091
rect 49003 27572 49069 27573
rect 49003 27508 49004 27572
rect 49068 27508 49069 27572
rect 49003 27507 49069 27508
rect 48083 22676 48149 22677
rect 48083 22612 48084 22676
rect 48148 22612 48149 22676
rect 48083 22611 48149 22612
rect 49190 21317 49250 177379
rect 49187 21316 49253 21317
rect 49187 21252 49188 21316
rect 49252 21252 49253 21316
rect 49187 21251 49253 21252
rect 49374 19957 49434 180371
rect 49558 21861 49618 185811
rect 50291 181388 50357 181389
rect 50291 181324 50292 181388
rect 50356 181324 50357 181388
rect 50291 181323 50357 181324
rect 50294 29613 50354 181323
rect 50291 29612 50357 29613
rect 50291 29548 50292 29612
rect 50356 29548 50357 29612
rect 50291 29547 50357 29548
rect 50478 28389 50538 190027
rect 50659 185740 50725 185741
rect 50659 185676 50660 185740
rect 50724 185676 50725 185740
rect 50659 185675 50725 185676
rect 50475 28388 50541 28389
rect 50475 28324 50476 28388
rect 50540 28324 50541 28388
rect 50475 28323 50541 28324
rect 49555 21860 49621 21861
rect 49555 21796 49556 21860
rect 49620 21796 49621 21860
rect 49555 21795 49621 21796
rect 50662 21453 50722 185675
rect 50843 173228 50909 173229
rect 50843 173164 50844 173228
rect 50908 173164 50909 173228
rect 50843 173163 50909 173164
rect 50659 21452 50725 21453
rect 50659 21388 50660 21452
rect 50724 21388 50725 21452
rect 50659 21387 50725 21388
rect 49371 19956 49437 19957
rect 49371 19892 49372 19956
rect 49436 19892 49437 19956
rect 49371 19891 49437 19892
rect 47899 3636 47965 3637
rect 47899 3572 47900 3636
rect 47964 3572 47965 3636
rect 47899 3571 47965 3572
rect 50846 3501 50906 173163
rect 51294 160954 51914 196398
rect 53051 193900 53117 193901
rect 53051 193836 53052 193900
rect 53116 193836 53117 193900
rect 53051 193835 53117 193836
rect 52315 174860 52381 174861
rect 52315 174796 52316 174860
rect 52380 174796 52381 174860
rect 52315 174795 52381 174796
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51027 148748 51093 148749
rect 51027 148684 51028 148748
rect 51092 148684 51093 148748
rect 51027 148683 51093 148684
rect 51030 147525 51090 148683
rect 51027 147524 51093 147525
rect 51027 147460 51028 147524
rect 51092 147460 51093 147524
rect 51027 147459 51093 147460
rect 51027 138140 51093 138141
rect 51027 138076 51028 138140
rect 51092 138076 51093 138140
rect 51027 138075 51093 138076
rect 51030 124133 51090 138075
rect 51294 124954 51914 160398
rect 52318 151830 52378 174795
rect 52134 151770 52378 151830
rect 52134 147690 52194 151770
rect 52134 147630 52378 147690
rect 52131 147524 52197 147525
rect 52131 147460 52132 147524
rect 52196 147460 52197 147524
rect 52131 147459 52197 147460
rect 52134 138141 52194 147459
rect 52318 142357 52378 147630
rect 52315 142356 52381 142357
rect 52315 142292 52316 142356
rect 52380 142292 52381 142356
rect 52315 142291 52381 142292
rect 52315 142084 52381 142085
rect 52315 142020 52316 142084
rect 52380 142020 52381 142084
rect 52315 142019 52381 142020
rect 52131 138140 52197 138141
rect 52131 138076 52132 138140
rect 52196 138076 52197 138140
rect 52131 138075 52197 138076
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51027 124132 51093 124133
rect 51027 124068 51028 124132
rect 51092 124068 51093 124132
rect 51027 124067 51093 124068
rect 51294 88954 51914 124398
rect 52131 124132 52197 124133
rect 52131 124068 52132 124132
rect 52196 124068 52197 124132
rect 52131 124067 52197 124068
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 52134 29477 52194 124067
rect 52131 29476 52197 29477
rect 52131 29412 52132 29476
rect 52196 29412 52197 29476
rect 52131 29411 52197 29412
rect 52318 24445 52378 142019
rect 53054 44301 53114 193835
rect 55075 191316 55141 191317
rect 55075 191252 55076 191316
rect 55140 191252 55141 191316
rect 55075 191251 55141 191252
rect 53603 189820 53669 189821
rect 53603 189756 53604 189820
rect 53668 189756 53669 189820
rect 53603 189755 53669 189756
rect 53419 172276 53485 172277
rect 53419 172212 53420 172276
rect 53484 172212 53485 172276
rect 53419 172211 53485 172212
rect 53235 166428 53301 166429
rect 53235 166364 53236 166428
rect 53300 166364 53301 166428
rect 53235 166363 53301 166364
rect 53051 44300 53117 44301
rect 53051 44236 53052 44300
rect 53116 44236 53117 44300
rect 53051 44235 53117 44236
rect 53238 25533 53298 166363
rect 53235 25532 53301 25533
rect 53235 25468 53236 25532
rect 53300 25468 53301 25532
rect 53235 25467 53301 25468
rect 53422 25397 53482 172211
rect 53419 25396 53485 25397
rect 53419 25332 53420 25396
rect 53484 25332 53485 25396
rect 53419 25331 53485 25332
rect 52315 24444 52381 24445
rect 52315 24380 52316 24444
rect 52380 24380 52381 24444
rect 52315 24379 52381 24380
rect 53606 23085 53666 189755
rect 54707 187236 54773 187237
rect 54707 187172 54708 187236
rect 54772 187172 54773 187236
rect 54707 187171 54773 187172
rect 54523 166564 54589 166565
rect 54523 166500 54524 166564
rect 54588 166500 54589 166564
rect 54523 166499 54589 166500
rect 54526 25533 54586 166499
rect 54523 25532 54589 25533
rect 54523 25468 54524 25532
rect 54588 25468 54589 25532
rect 54523 25467 54589 25468
rect 54710 24581 54770 187171
rect 54891 182884 54957 182885
rect 54891 182820 54892 182884
rect 54956 182820 54957 182884
rect 54891 182819 54957 182820
rect 54707 24580 54773 24581
rect 54707 24516 54708 24580
rect 54772 24516 54773 24580
rect 54707 24515 54773 24516
rect 53603 23084 53669 23085
rect 53603 23020 53604 23084
rect 53668 23020 53669 23084
rect 53603 23019 53669 23020
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 50843 3500 50909 3501
rect 50843 3436 50844 3500
rect 50908 3436 50909 3500
rect 50843 3435 50909 3436
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 -3226 51914 16398
rect 54894 3501 54954 182819
rect 54891 3500 54957 3501
rect 54891 3436 54892 3500
rect 54956 3436 54957 3500
rect 54891 3435 54957 3436
rect 55078 3365 55138 191251
rect 55443 189684 55509 189685
rect 55443 189620 55444 189684
rect 55508 189620 55509 189684
rect 55443 189619 55509 189620
rect 55446 58037 55506 189619
rect 55627 188460 55693 188461
rect 55627 188396 55628 188460
rect 55692 188396 55693 188460
rect 55627 188395 55693 188396
rect 55443 58036 55509 58037
rect 55443 57972 55444 58036
rect 55508 57972 55509 58036
rect 55443 57971 55509 57972
rect 55630 35597 55690 188395
rect 55794 165454 56414 198000
rect 82794 192454 83414 198000
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 57835 191180 57901 191181
rect 57835 191116 57836 191180
rect 57900 191116 57901 191180
rect 57835 191115 57901 191116
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57651 160988 57717 160989
rect 57651 160924 57652 160988
rect 57716 160924 57717 160988
rect 57651 160923 57717 160924
rect 57467 159492 57533 159493
rect 57467 159428 57468 159492
rect 57532 159428 57533 159492
rect 57467 159427 57533 159428
rect 57283 151060 57349 151061
rect 57283 150996 57284 151060
rect 57348 150996 57349 151060
rect 57283 150995 57349 150996
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 57286 75037 57346 150995
rect 57283 75036 57349 75037
rect 57283 74972 57284 75036
rect 57348 74972 57349 75036
rect 57283 74971 57349 74972
rect 57470 59397 57530 159427
rect 57467 59396 57533 59397
rect 57467 59332 57468 59396
rect 57532 59332 57533 59396
rect 57467 59331 57533 59332
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55627 35596 55693 35597
rect 55627 35532 55628 35596
rect 55692 35532 55693 35596
rect 55627 35531 55693 35532
rect 55794 21454 56414 56898
rect 57654 34917 57714 160923
rect 57838 64837 57898 191115
rect 61331 190228 61397 190229
rect 61331 190164 61332 190228
rect 61396 190164 61397 190228
rect 61331 190163 61397 190164
rect 58571 187508 58637 187509
rect 58571 187444 58572 187508
rect 58636 187444 58637 187508
rect 58571 187443 58637 187444
rect 58019 143580 58085 143581
rect 58019 143516 58020 143580
rect 58084 143516 58085 143580
rect 58019 143515 58085 143516
rect 58022 118013 58082 143515
rect 58574 135965 58634 187443
rect 59123 187372 59189 187373
rect 59123 187308 59124 187372
rect 59188 187308 59189 187372
rect 59123 187307 59189 187308
rect 58939 158404 59005 158405
rect 58939 158340 58940 158404
rect 59004 158340 59005 158404
rect 58939 158339 59005 158340
rect 58755 155276 58821 155277
rect 58755 155212 58756 155276
rect 58820 155212 58821 155276
rect 58755 155211 58821 155212
rect 58758 143581 58818 155211
rect 58755 143580 58821 143581
rect 58755 143516 58756 143580
rect 58820 143516 58821 143580
rect 58755 143515 58821 143516
rect 58571 135964 58637 135965
rect 58571 135900 58572 135964
rect 58636 135900 58637 135964
rect 58571 135899 58637 135900
rect 58571 124812 58637 124813
rect 58571 124748 58572 124812
rect 58636 124748 58637 124812
rect 58571 124747 58637 124748
rect 58019 118012 58085 118013
rect 58019 117948 58020 118012
rect 58084 117948 58085 118012
rect 58019 117947 58085 117948
rect 57835 64836 57901 64837
rect 57835 64772 57836 64836
rect 57900 64772 57901 64836
rect 57835 64771 57901 64772
rect 57651 34916 57717 34917
rect 57651 34852 57652 34916
rect 57716 34852 57717 34916
rect 57651 34851 57717 34852
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55075 3364 55141 3365
rect 55075 3300 55076 3364
rect 55140 3300 55141 3364
rect 55075 3299 55141 3300
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 -4186 56414 20898
rect 58574 19005 58634 124747
rect 58942 124269 59002 158339
rect 59126 142085 59186 187307
rect 60595 184652 60661 184653
rect 60595 184588 60596 184652
rect 60660 184588 60661 184652
rect 60595 184587 60661 184588
rect 60411 174996 60477 174997
rect 60411 174932 60412 174996
rect 60476 174932 60477 174996
rect 60411 174931 60477 174932
rect 60043 155684 60109 155685
rect 60043 155620 60044 155684
rect 60108 155620 60109 155684
rect 60043 155619 60109 155620
rect 60046 146573 60106 155619
rect 60227 150108 60293 150109
rect 60227 150044 60228 150108
rect 60292 150044 60293 150108
rect 60227 150043 60293 150044
rect 60230 148749 60290 150043
rect 60227 148748 60293 148749
rect 60227 148684 60228 148748
rect 60292 148684 60293 148748
rect 60227 148683 60293 148684
rect 60414 147930 60474 174931
rect 60230 147870 60474 147930
rect 60043 146572 60109 146573
rect 60043 146508 60044 146572
rect 60108 146508 60109 146572
rect 60043 146507 60109 146508
rect 59307 144940 59373 144941
rect 59307 144876 59308 144940
rect 59372 144876 59373 144940
rect 59307 144875 59373 144876
rect 59123 142084 59189 142085
rect 59123 142020 59124 142084
rect 59188 142020 59189 142084
rect 59123 142019 59189 142020
rect 59310 137325 59370 144875
rect 59491 142084 59557 142085
rect 59491 142020 59492 142084
rect 59556 142020 59557 142084
rect 59491 142019 59557 142020
rect 59307 137324 59373 137325
rect 59307 137260 59308 137324
rect 59372 137260 59373 137324
rect 59307 137259 59373 137260
rect 59123 136644 59189 136645
rect 59123 136580 59124 136644
rect 59188 136580 59189 136644
rect 59123 136579 59189 136580
rect 58939 124268 59005 124269
rect 58939 124204 58940 124268
rect 59004 124204 59005 124268
rect 58939 124203 59005 124204
rect 58755 123588 58821 123589
rect 58755 123524 58756 123588
rect 58820 123524 58821 123588
rect 58755 123523 58821 123524
rect 58758 28253 58818 123523
rect 59126 30837 59186 136579
rect 59494 125493 59554 142019
rect 60230 138030 60290 147870
rect 60598 147690 60658 184587
rect 61334 150109 61394 190163
rect 61515 187644 61581 187645
rect 61515 187580 61516 187644
rect 61580 187580 61581 187644
rect 61515 187579 61581 187580
rect 61331 150108 61397 150109
rect 61331 150044 61332 150108
rect 61396 150044 61397 150108
rect 61331 150043 61397 150044
rect 61518 149973 61578 187579
rect 61699 177852 61765 177853
rect 61699 177788 61700 177852
rect 61764 177788 61765 177852
rect 61699 177787 61765 177788
rect 61515 149972 61581 149973
rect 61515 149908 61516 149972
rect 61580 149908 61581 149972
rect 61515 149907 61581 149908
rect 59678 137970 60290 138030
rect 60414 147630 60658 147690
rect 60414 138030 60474 147630
rect 61702 146570 61762 177787
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 152000 83414 155898
rect 87294 196954 87914 198000
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 152000 87914 160398
rect 118794 192454 119414 198000
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 152000 119414 155898
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 152000 123914 160398
rect 154794 192454 155414 198000
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 152000 155414 155898
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 152000 159914 160398
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 152000 191414 155898
rect 195294 196954 195914 198000
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 152000 195914 160398
rect 226794 192454 227414 198000
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 152000 227414 155898
rect 231294 196954 231914 198000
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 152000 231914 160398
rect 262794 192454 263414 198000
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 152000 263414 155898
rect 267294 196954 267914 198000
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 152000 267914 160398
rect 298794 192454 299414 198000
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 152000 299414 155898
rect 303294 196954 303914 198000
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 152000 303914 160398
rect 334794 192454 335414 198000
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 152000 335414 155898
rect 339294 196954 339914 198000
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 346902 172413 346962 200910
rect 347635 200564 347701 200565
rect 347635 200500 347636 200564
rect 347700 200500 347701 200564
rect 347635 200499 347701 200500
rect 347638 200130 347698 200499
rect 347086 200070 347698 200130
rect 347086 191589 347146 200070
rect 347451 199612 347517 199613
rect 347451 199548 347452 199612
rect 347516 199548 347517 199612
rect 347451 199547 347517 199548
rect 347454 191725 347514 199547
rect 347451 191724 347517 191725
rect 347451 191660 347452 191724
rect 347516 191660 347517 191724
rect 347451 191659 347517 191660
rect 347083 191588 347149 191589
rect 347083 191524 347084 191588
rect 347148 191524 347149 191588
rect 347083 191523 347149 191524
rect 348374 181661 348434 456723
rect 348558 299437 348618 557363
rect 348923 523020 348989 523021
rect 348923 522956 348924 523020
rect 348988 522956 348989 523020
rect 348923 522955 348989 522956
rect 348739 341460 348805 341461
rect 348739 341396 348740 341460
rect 348804 341396 348805 341460
rect 348739 341395 348805 341396
rect 348555 299436 348621 299437
rect 348555 299372 348556 299436
rect 348620 299372 348621 299436
rect 348555 299371 348621 299372
rect 348371 181660 348437 181661
rect 348371 181596 348372 181660
rect 348436 181596 348437 181660
rect 348371 181595 348437 181596
rect 348742 181525 348802 341395
rect 348926 233885 348986 522955
rect 349110 483037 349170 578851
rect 350947 571980 351013 571981
rect 350947 571916 350948 571980
rect 351012 571916 351013 571980
rect 350947 571915 351013 571916
rect 349291 563548 349357 563549
rect 349291 563484 349292 563548
rect 349356 563484 349357 563548
rect 349291 563483 349357 563484
rect 349107 483036 349173 483037
rect 349107 482972 349108 483036
rect 349172 482972 349173 483036
rect 349107 482971 349173 482972
rect 349107 463996 349173 463997
rect 349107 463932 349108 463996
rect 349172 463932 349173 463996
rect 349107 463931 349173 463932
rect 348923 233884 348989 233885
rect 348923 233820 348924 233884
rect 348988 233820 348989 233884
rect 348923 233819 348989 233820
rect 349110 195533 349170 463931
rect 349294 433261 349354 563483
rect 349475 556204 349541 556205
rect 349475 556140 349476 556204
rect 349540 556140 349541 556204
rect 349475 556139 349541 556140
rect 349291 433260 349357 433261
rect 349291 433196 349292 433260
rect 349356 433196 349357 433260
rect 349291 433195 349357 433196
rect 349478 385797 349538 556139
rect 350579 520300 350645 520301
rect 350579 520236 350580 520300
rect 350644 520236 350645 520300
rect 350579 520235 350645 520236
rect 349659 434892 349725 434893
rect 349659 434828 349660 434892
rect 349724 434828 349725 434892
rect 349659 434827 349725 434828
rect 349475 385796 349541 385797
rect 349475 385732 349476 385796
rect 349540 385732 349541 385796
rect 349475 385731 349541 385732
rect 349475 358868 349541 358869
rect 349475 358804 349476 358868
rect 349540 358804 349541 358868
rect 349475 358803 349541 358804
rect 349107 195532 349173 195533
rect 349107 195468 349108 195532
rect 349172 195468 349173 195532
rect 349107 195467 349173 195468
rect 348739 181524 348805 181525
rect 348739 181460 348740 181524
rect 348804 181460 348805 181524
rect 348739 181459 348805 181460
rect 346899 172412 346965 172413
rect 346899 172348 346900 172412
rect 346964 172348 346965 172412
rect 346899 172347 346965 172348
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 152000 339914 160398
rect 349478 151197 349538 358803
rect 349662 177717 349722 434827
rect 350582 190365 350642 520235
rect 350763 507924 350829 507925
rect 350763 507860 350764 507924
rect 350828 507860 350829 507924
rect 350763 507859 350829 507860
rect 350579 190364 350645 190365
rect 350579 190300 350580 190364
rect 350644 190300 350645 190364
rect 350579 190299 350645 190300
rect 350766 179893 350826 507859
rect 350950 268157 351010 571915
rect 351134 278357 351194 581571
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 351867 565996 351933 565997
rect 351867 565932 351868 565996
rect 351932 565932 351933 565996
rect 351867 565931 351933 565932
rect 351131 278356 351197 278357
rect 351131 278292 351132 278356
rect 351196 278292 351197 278356
rect 351131 278291 351197 278292
rect 350947 268156 351013 268157
rect 350947 268092 350948 268156
rect 351012 268092 351013 268156
rect 350947 268091 351013 268092
rect 350947 245580 351013 245581
rect 350947 245516 350948 245580
rect 351012 245516 351013 245580
rect 350947 245515 351013 245516
rect 350950 198933 351010 245515
rect 350947 198932 351013 198933
rect 350947 198868 350948 198932
rect 351012 198868 351013 198932
rect 350947 198867 351013 198868
rect 350763 179892 350829 179893
rect 350763 179828 350764 179892
rect 350828 179828 350829 179892
rect 350763 179827 350829 179828
rect 349659 177716 349725 177717
rect 349659 177652 349660 177716
rect 349724 177652 349725 177716
rect 349659 177651 349725 177652
rect 351870 155821 351930 565931
rect 352051 565860 352117 565861
rect 352051 565796 352052 565860
rect 352116 565796 352117 565860
rect 352051 565795 352117 565796
rect 352054 548997 352114 565795
rect 352051 548996 352117 548997
rect 352051 548932 352052 548996
rect 352116 548932 352117 548996
rect 352051 548931 352117 548932
rect 352794 534454 353414 569898
rect 353523 568852 353589 568853
rect 353523 568788 353524 568852
rect 353588 568788 353589 568852
rect 353523 568787 353589 568788
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352051 490652 352117 490653
rect 352051 490588 352052 490652
rect 352116 490588 352117 490652
rect 352051 490587 352117 490588
rect 352054 158541 352114 490587
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 353526 184653 353586 568787
rect 356099 564908 356165 564909
rect 356099 564844 356100 564908
rect 356164 564844 356165 564908
rect 356099 564843 356165 564844
rect 353707 472292 353773 472293
rect 353707 472228 353708 472292
rect 353772 472228 353773 472292
rect 353707 472227 353773 472228
rect 353523 184652 353589 184653
rect 353523 184588 353524 184652
rect 353588 184588 353589 184652
rect 353523 184587 353589 184588
rect 353710 184517 353770 472227
rect 355179 461820 355245 461821
rect 355179 461756 355180 461820
rect 355244 461756 355245 461820
rect 355179 461755 355245 461756
rect 354443 305012 354509 305013
rect 354443 304948 354444 305012
rect 354508 304948 354509 305012
rect 354443 304947 354509 304948
rect 354446 292590 354506 304947
rect 354446 292530 354690 292590
rect 354630 282930 354690 292530
rect 354446 282870 354690 282930
rect 353707 184516 353773 184517
rect 353707 184452 353708 184516
rect 353772 184452 353773 184516
rect 353707 184451 353773 184452
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352051 158540 352117 158541
rect 352051 158476 352052 158540
rect 352116 158476 352117 158540
rect 352051 158475 352117 158476
rect 351867 155820 351933 155821
rect 351867 155756 351868 155820
rect 351932 155756 351933 155820
rect 351867 155755 351933 155756
rect 352794 152000 353414 173898
rect 354446 152557 354506 282870
rect 355182 159629 355242 461755
rect 356102 192949 356162 564843
rect 356099 192948 356165 192949
rect 356099 192884 356100 192948
rect 356164 192884 356165 192948
rect 356099 192883 356165 192884
rect 355179 159628 355245 159629
rect 355179 159564 355180 159628
rect 355244 159564 355245 159628
rect 355179 159563 355245 159564
rect 356654 152965 356714 686019
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 356835 681868 356901 681869
rect 356835 681804 356836 681868
rect 356900 681804 356901 681868
rect 356835 681803 356901 681804
rect 356838 198253 356898 681803
rect 357294 646954 357914 682398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 358123 682276 358189 682277
rect 358123 682212 358124 682276
rect 358188 682212 358189 682276
rect 358123 682211 358189 682212
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 356835 198252 356901 198253
rect 356835 198188 356836 198252
rect 356900 198188 356901 198252
rect 356835 198187 356901 198188
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 356651 152964 356717 152965
rect 356651 152900 356652 152964
rect 356716 152900 356717 152964
rect 356651 152899 356717 152900
rect 354443 152556 354509 152557
rect 354443 152492 354444 152556
rect 354508 152492 354509 152556
rect 354443 152491 354509 152492
rect 357294 152000 357914 178398
rect 358126 163437 358186 682211
rect 359411 680780 359477 680781
rect 359411 680716 359412 680780
rect 359476 680716 359477 680780
rect 359411 680715 359477 680716
rect 359414 198117 359474 680715
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 367691 680644 367757 680645
rect 367691 680580 367692 680644
rect 367756 680580 367757 680644
rect 367691 680579 367757 680580
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 363459 593740 363525 593741
rect 363459 593676 363460 593740
rect 363524 593676 363525 593740
rect 363459 593675 363525 593676
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 359595 566132 359661 566133
rect 359595 566068 359596 566132
rect 359660 566068 359661 566132
rect 359595 566067 359661 566068
rect 359411 198116 359477 198117
rect 359411 198052 359412 198116
rect 359476 198052 359477 198116
rect 359411 198051 359477 198052
rect 358123 163436 358189 163437
rect 358123 163372 358124 163436
rect 358188 163372 358189 163436
rect 358123 163371 358189 163372
rect 359598 151197 359658 566067
rect 360147 561916 360213 561917
rect 360147 561852 360148 561916
rect 360212 561852 360213 561916
rect 360147 561851 360213 561852
rect 360150 292590 360210 561851
rect 360331 561780 360397 561781
rect 360331 561716 360332 561780
rect 360396 561716 360397 561780
rect 360331 561715 360397 561716
rect 359966 292530 360210 292590
rect 359966 282930 360026 292530
rect 359966 282870 360210 282930
rect 360150 155413 360210 282870
rect 360334 185877 360394 561715
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 360699 325820 360765 325821
rect 360699 325756 360700 325820
rect 360764 325756 360765 325820
rect 360699 325755 360765 325756
rect 360331 185876 360397 185877
rect 360331 185812 360332 185876
rect 360396 185812 360397 185876
rect 360331 185811 360397 185812
rect 360147 155412 360213 155413
rect 360147 155348 360148 155412
rect 360212 155348 360213 155412
rect 360147 155347 360213 155348
rect 360702 154053 360762 325755
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360699 154052 360765 154053
rect 360699 153988 360700 154052
rect 360764 153988 360765 154052
rect 360699 153987 360765 153988
rect 361794 152000 362414 182898
rect 363462 166565 363522 593675
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 363643 566404 363709 566405
rect 363643 566340 363644 566404
rect 363708 566340 363709 566404
rect 363643 566339 363709 566340
rect 363459 166564 363525 166565
rect 363459 166500 363460 166564
rect 363524 166500 363525 166564
rect 363459 166499 363525 166500
rect 363646 154053 363706 566339
rect 364379 562188 364445 562189
rect 364379 562124 364380 562188
rect 364444 562124 364445 562188
rect 364379 562123 364445 562124
rect 364382 155549 364442 562123
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 367139 518940 367205 518941
rect 367139 518876 367140 518940
rect 367204 518876 367205 518940
rect 367139 518875 367205 518876
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 364563 457060 364629 457061
rect 364563 456996 364564 457060
rect 364628 456996 364629 457060
rect 364563 456995 364629 456996
rect 364566 178805 364626 456995
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 364563 178804 364629 178805
rect 364563 178740 364564 178804
rect 364628 178740 364629 178804
rect 364563 178739 364629 178740
rect 364379 155548 364445 155549
rect 364379 155484 364380 155548
rect 364444 155484 364445 155548
rect 364379 155483 364445 155484
rect 363643 154052 363709 154053
rect 363643 153988 363644 154052
rect 363708 153988 363709 154052
rect 363643 153987 363709 153988
rect 366294 152000 366914 187398
rect 367142 181389 367202 518875
rect 367694 196757 367754 680579
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370451 657660 370517 657661
rect 370451 657596 370452 657660
rect 370516 657596 370517 657660
rect 370451 657595 370517 657596
rect 368979 635900 369045 635901
rect 368979 635836 368980 635900
rect 369044 635836 369045 635900
rect 368979 635835 369045 635836
rect 368982 198389 369042 635835
rect 368979 198388 369045 198389
rect 368979 198324 368980 198388
rect 369044 198324 369045 198388
rect 368979 198323 369045 198324
rect 367691 196756 367757 196757
rect 367691 196692 367692 196756
rect 367756 196692 367757 196756
rect 367691 196691 367757 196692
rect 367139 181388 367205 181389
rect 367139 181324 367140 181388
rect 367204 181324 367205 181388
rect 367139 181323 367205 181324
rect 370454 152421 370514 657595
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 378731 622980 378797 622981
rect 378731 622916 378732 622980
rect 378796 622916 378797 622980
rect 378731 622915 378797 622916
rect 377259 611420 377325 611421
rect 377259 611356 377260 611420
rect 377324 611356 377325 611420
rect 377259 611355 377325 611356
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 371739 578780 371805 578781
rect 371739 578716 371740 578780
rect 371804 578716 371805 578780
rect 371739 578715 371805 578716
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 371742 160989 371802 578715
rect 373211 565860 373277 565861
rect 373211 565796 373212 565860
rect 373276 565796 373277 565860
rect 373211 565795 373277 565796
rect 372659 302292 372725 302293
rect 372659 302228 372660 302292
rect 372724 302228 372725 302292
rect 372659 302227 372725 302228
rect 371739 160988 371805 160989
rect 371739 160924 371740 160988
rect 371804 160924 371805 160988
rect 371739 160923 371805 160924
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370451 152420 370517 152421
rect 370451 152356 370452 152420
rect 370516 152356 370517 152420
rect 370451 152355 370517 152356
rect 370794 152000 371414 155898
rect 349475 151196 349541 151197
rect 349475 151132 349476 151196
rect 349540 151132 349541 151196
rect 349475 151131 349541 151132
rect 359595 151196 359661 151197
rect 359595 151132 359596 151196
rect 359660 151132 359661 151196
rect 359595 151131 359661 151132
rect 372662 151061 372722 302227
rect 373214 172141 373274 565795
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 374499 502484 374565 502485
rect 374499 502420 374500 502484
rect 374564 502420 374565 502484
rect 374499 502419 374565 502420
rect 374502 192813 374562 502419
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 374499 192812 374565 192813
rect 374499 192748 374500 192812
rect 374564 192748 374565 192812
rect 374499 192747 374565 192748
rect 373211 172140 373277 172141
rect 373211 172076 373212 172140
rect 373276 172076 373277 172140
rect 373211 172075 373277 172076
rect 375294 160954 375914 196398
rect 377262 189957 377322 611355
rect 377443 453660 377509 453661
rect 377443 453596 377444 453660
rect 377508 453596 377509 453660
rect 377443 453595 377509 453596
rect 377259 189956 377325 189957
rect 377259 189892 377260 189956
rect 377324 189892 377325 189956
rect 377259 189891 377325 189892
rect 377446 172277 377506 453595
rect 378734 177581 378794 622915
rect 379794 597454 380414 632898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 392531 683772 392597 683773
rect 392531 683708 392532 683772
rect 392596 683708 392597 683772
rect 392531 683707 392597 683708
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 387563 604484 387629 604485
rect 387563 604420 387564 604484
rect 387628 604420 387629 604484
rect 387563 604419 387629 604420
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 382779 598500 382845 598501
rect 382779 598436 382780 598500
rect 382844 598436 382845 598500
rect 382779 598435 382845 598436
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 381491 563412 381557 563413
rect 381491 563348 381492 563412
rect 381556 563348 381557 563412
rect 381491 563347 381557 563348
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 378915 527100 378981 527101
rect 378915 527036 378916 527100
rect 378980 527036 378981 527100
rect 378915 527035 378981 527036
rect 378918 188869 378978 527035
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 378915 188868 378981 188869
rect 378915 188804 378916 188868
rect 378980 188804 378981 188868
rect 378915 188803 378981 188804
rect 378731 177580 378797 177581
rect 378731 177516 378732 177580
rect 378796 177516 378797 177580
rect 378731 177515 378797 177516
rect 377443 172276 377509 172277
rect 377443 172212 377444 172276
rect 377508 172212 377509 172276
rect 377443 172211 377509 172212
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 152000 375914 160398
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 152000 380414 164898
rect 381494 152557 381554 563347
rect 382782 180437 382842 598435
rect 384294 565954 384914 601398
rect 387011 580820 387077 580821
rect 387011 580756 387012 580820
rect 387076 580756 387077 580820
rect 387011 580755 387077 580756
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 385539 497180 385605 497181
rect 385539 497116 385540 497180
rect 385604 497116 385605 497180
rect 385539 497115 385605 497116
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 382779 180436 382845 180437
rect 382779 180372 382780 180436
rect 382844 180372 382845 180436
rect 382779 180371 382845 180372
rect 384294 169954 384914 205398
rect 385542 188733 385602 497115
rect 385539 188732 385605 188733
rect 385539 188668 385540 188732
rect 385604 188668 385605 188732
rect 385539 188667 385605 188668
rect 387014 182885 387074 580755
rect 387566 235517 387626 604419
rect 388299 588572 388365 588573
rect 388299 588508 388300 588572
rect 388364 588508 388365 588572
rect 388299 588507 388365 588508
rect 387747 311948 387813 311949
rect 387747 311884 387748 311948
rect 387812 311884 387813 311948
rect 387747 311883 387813 311884
rect 387563 235516 387629 235517
rect 387563 235452 387564 235516
rect 387628 235452 387629 235516
rect 387563 235451 387629 235452
rect 387011 182884 387077 182885
rect 387011 182820 387012 182884
rect 387076 182820 387077 182884
rect 387011 182819 387077 182820
rect 387750 172005 387810 311883
rect 388302 238373 388362 588507
rect 388794 570454 389414 605898
rect 391243 581500 391309 581501
rect 391243 581436 391244 581500
rect 391308 581436 391309 581500
rect 391243 581435 391309 581436
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 391059 567356 391125 567357
rect 391059 567292 391060 567356
rect 391124 567292 391125 567356
rect 391059 567291 391125 567292
rect 389771 566268 389837 566269
rect 389771 566204 389772 566268
rect 389836 566204 389837 566268
rect 389771 566203 389837 566204
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388299 238372 388365 238373
rect 388299 238308 388300 238372
rect 388364 238308 388365 238372
rect 388299 238307 388365 238308
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 387747 172004 387813 172005
rect 387747 171940 387748 172004
rect 387812 171940 387813 172004
rect 387747 171939 387813 171940
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 381491 152556 381557 152557
rect 381491 152492 381492 152556
rect 381556 152492 381557 152556
rect 381491 152491 381557 152492
rect 384294 152000 384914 169398
rect 388794 152000 389414 173898
rect 389774 163573 389834 566203
rect 389955 557700 390021 557701
rect 389955 557636 389956 557700
rect 390020 557636 390021 557700
rect 389955 557635 390021 557636
rect 389958 171869 390018 557635
rect 389955 171868 390021 171869
rect 389955 171804 389956 171868
rect 390020 171804 390021 171868
rect 389955 171803 390021 171804
rect 389771 163572 389837 163573
rect 389771 163508 389772 163572
rect 389836 163508 389837 163572
rect 389771 163507 389837 163508
rect 391062 160989 391122 567291
rect 391246 180301 391306 581435
rect 391427 563140 391493 563141
rect 391427 563076 391428 563140
rect 391492 563076 391493 563140
rect 391427 563075 391493 563076
rect 391430 240549 391490 563075
rect 391427 240548 391493 240549
rect 391427 240484 391428 240548
rect 391492 240484 391493 240548
rect 391427 240483 391493 240484
rect 391243 180300 391309 180301
rect 391243 180236 391244 180300
rect 391308 180236 391309 180300
rect 391243 180235 391309 180236
rect 392534 177445 392594 683707
rect 393083 683636 393149 683637
rect 393083 683572 393084 683636
rect 393148 683572 393149 683636
rect 393083 683571 393149 683572
rect 392715 480180 392781 480181
rect 392715 480116 392716 480180
rect 392780 480116 392781 480180
rect 392715 480115 392781 480116
rect 392531 177444 392597 177445
rect 392531 177380 392532 177444
rect 392596 177380 392597 177444
rect 392531 177379 392597 177380
rect 392718 170509 392778 480115
rect 393086 236741 393146 683571
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 393294 646954 393914 682398
rect 395291 682412 395357 682413
rect 395291 682348 395292 682412
rect 395356 682348 395357 682412
rect 395291 682347 395357 682348
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393083 236740 393149 236741
rect 393083 236676 393084 236740
rect 393148 236676 393149 236740
rect 393083 236675 393149 236676
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 395294 180709 395354 682347
rect 397315 682004 397381 682005
rect 397315 681940 397316 682004
rect 397380 681940 397381 682004
rect 397315 681939 397381 681940
rect 396579 568716 396645 568717
rect 396579 568652 396580 568716
rect 396644 568652 396645 568716
rect 396579 568651 396645 568652
rect 395475 560964 395541 560965
rect 395475 560900 395476 560964
rect 395540 560900 395541 560964
rect 395475 560899 395541 560900
rect 395291 180708 395357 180709
rect 395291 180644 395292 180708
rect 395356 180644 395357 180708
rect 395291 180643 395357 180644
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 392715 170508 392781 170509
rect 392715 170444 392716 170508
rect 392780 170444 392781 170508
rect 392715 170443 392781 170444
rect 391059 160988 391125 160989
rect 391059 160924 391060 160988
rect 391124 160924 391125 160988
rect 391059 160923 391125 160924
rect 393294 152000 393914 178398
rect 395478 152829 395538 560899
rect 395659 510780 395725 510781
rect 395659 510716 395660 510780
rect 395724 510716 395725 510780
rect 395659 510715 395725 510716
rect 395662 194445 395722 510715
rect 396211 243540 396277 243541
rect 396211 243476 396212 243540
rect 396276 243476 396277 243540
rect 396211 243475 396277 243476
rect 395659 194444 395725 194445
rect 395659 194380 395660 194444
rect 395724 194380 395725 194444
rect 395659 194379 395725 194380
rect 396214 187101 396274 243475
rect 396211 187100 396277 187101
rect 396211 187036 396212 187100
rect 396276 187036 396277 187100
rect 396211 187035 396277 187036
rect 396582 153101 396642 568651
rect 397318 231301 397378 681939
rect 397794 651454 398414 686898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 399339 682140 399405 682141
rect 399339 682076 399340 682140
rect 399404 682076 399405 682140
rect 399339 682075 399405 682076
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 398603 567220 398669 567221
rect 398603 567156 398604 567220
rect 398668 567156 398669 567220
rect 398603 567155 398669 567156
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397315 231300 397381 231301
rect 397315 231236 397316 231300
rect 397380 231236 397381 231300
rect 397315 231235 397381 231236
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 396579 153100 396645 153101
rect 396579 153036 396580 153100
rect 396644 153036 396645 153100
rect 396579 153035 396645 153036
rect 395475 152828 395541 152829
rect 395475 152764 395476 152828
rect 395540 152764 395541 152828
rect 395475 152763 395541 152764
rect 397794 152000 398414 182898
rect 398606 157317 398666 567155
rect 399342 163709 399402 682075
rect 400075 681052 400141 681053
rect 400075 680988 400076 681052
rect 400140 680988 400141 681052
rect 400075 680987 400141 680988
rect 399523 607340 399589 607341
rect 399523 607276 399524 607340
rect 399588 607276 399589 607340
rect 399523 607275 399589 607276
rect 399526 189821 399586 607275
rect 400078 235653 400138 680987
rect 402294 655954 402914 691398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 403755 682684 403821 682685
rect 403755 682620 403756 682684
rect 403820 682620 403821 682684
rect 403755 682619 403821 682620
rect 403571 682548 403637 682549
rect 403571 682484 403572 682548
rect 403636 682484 403637 682548
rect 403571 682483 403637 682484
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402099 652220 402165 652221
rect 402099 652156 402100 652220
rect 402164 652156 402165 652220
rect 402099 652155 402165 652156
rect 401363 645420 401429 645421
rect 401363 645356 401364 645420
rect 401428 645356 401429 645420
rect 401363 645355 401429 645356
rect 400811 560556 400877 560557
rect 400811 560492 400812 560556
rect 400876 560492 400877 560556
rect 400811 560491 400877 560492
rect 400075 235652 400141 235653
rect 400075 235588 400076 235652
rect 400140 235588 400141 235652
rect 400075 235587 400141 235588
rect 399523 189820 399589 189821
rect 399523 189756 399524 189820
rect 399588 189756 399589 189820
rect 399523 189755 399589 189756
rect 399339 163708 399405 163709
rect 399339 163644 399340 163708
rect 399404 163644 399405 163708
rect 399339 163643 399405 163644
rect 398603 157316 398669 157317
rect 398603 157252 398604 157316
rect 398668 157252 398669 157316
rect 398603 157251 398669 157252
rect 400814 152965 400874 560491
rect 401366 231165 401426 645355
rect 402102 231573 402162 652155
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402099 231572 402165 231573
rect 402099 231508 402100 231572
rect 402164 231508 402165 231572
rect 402099 231507 402165 231508
rect 401363 231164 401429 231165
rect 401363 231100 401364 231164
rect 401428 231100 401429 231164
rect 401363 231099 401429 231100
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 400811 152964 400877 152965
rect 400811 152900 400812 152964
rect 400876 152900 400877 152964
rect 400811 152899 400877 152900
rect 402294 152000 402914 187398
rect 403574 162077 403634 682483
rect 403758 195805 403818 682619
rect 405595 681188 405661 681189
rect 405595 681124 405596 681188
rect 405660 681124 405661 681188
rect 405595 681123 405661 681124
rect 404123 628420 404189 628421
rect 404123 628356 404124 628420
rect 404188 628356 404189 628420
rect 404123 628355 404189 628356
rect 404126 234021 404186 628355
rect 405411 624340 405477 624341
rect 405411 624276 405412 624340
rect 405476 624276 405477 624340
rect 405411 624275 405477 624276
rect 404859 251836 404925 251837
rect 404859 251772 404860 251836
rect 404924 251772 404925 251836
rect 404859 251771 404925 251772
rect 404123 234020 404189 234021
rect 404123 233956 404124 234020
rect 404188 233956 404189 234020
rect 404123 233955 404189 233956
rect 403755 195804 403821 195805
rect 403755 195740 403756 195804
rect 403820 195740 403821 195804
rect 403755 195739 403821 195740
rect 403571 162076 403637 162077
rect 403571 162012 403572 162076
rect 403636 162012 403637 162076
rect 403571 162011 403637 162012
rect 404862 151061 404922 251771
rect 405414 234157 405474 624275
rect 405598 235789 405658 681123
rect 406794 660454 407414 695898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 407619 684724 407685 684725
rect 407619 684660 407620 684724
rect 407684 684660 407685 684724
rect 407619 684659 407685 684660
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406515 627740 406581 627741
rect 406515 627676 406516 627740
rect 406580 627676 406581 627740
rect 406515 627675 406581 627676
rect 406147 306100 406213 306101
rect 406147 306036 406148 306100
rect 406212 306036 406213 306100
rect 406147 306035 406213 306036
rect 405595 235788 405661 235789
rect 405595 235724 405596 235788
rect 405660 235724 405661 235788
rect 405595 235723 405661 235724
rect 406150 235245 406210 306035
rect 406331 262172 406397 262173
rect 406331 262108 406332 262172
rect 406396 262108 406397 262172
rect 406331 262107 406397 262108
rect 406147 235244 406213 235245
rect 406147 235180 406148 235244
rect 406212 235180 406213 235244
rect 406147 235179 406213 235180
rect 405411 234156 405477 234157
rect 405411 234092 405412 234156
rect 405476 234092 405477 234156
rect 405411 234091 405477 234092
rect 406334 154325 406394 262107
rect 406518 206277 406578 627675
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 407622 589117 407682 684659
rect 409827 683364 409893 683365
rect 409827 683300 409828 683364
rect 409892 683300 409893 683364
rect 409827 683299 409893 683300
rect 409643 679828 409709 679829
rect 409643 679764 409644 679828
rect 409708 679764 409709 679828
rect 409643 679763 409709 679764
rect 408355 678332 408421 678333
rect 408355 678268 408356 678332
rect 408420 678268 408421 678332
rect 408355 678267 408421 678268
rect 407803 601220 407869 601221
rect 407803 601156 407804 601220
rect 407868 601156 407869 601220
rect 407803 601155 407869 601156
rect 407619 589116 407685 589117
rect 407619 589052 407620 589116
rect 407684 589052 407685 589116
rect 407619 589051 407685 589052
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 407806 584357 407866 601155
rect 407803 584356 407869 584357
rect 407803 584292 407804 584356
rect 407868 584292 407869 584356
rect 407803 584291 407869 584292
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 407619 533900 407685 533901
rect 407619 533836 407620 533900
rect 407684 533836 407685 533900
rect 407619 533835 407685 533836
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406515 206276 406581 206277
rect 406515 206212 406516 206276
rect 406580 206212 406581 206276
rect 406515 206211 406581 206212
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 407622 189685 407682 533835
rect 407803 489020 407869 489021
rect 407803 488956 407804 489020
rect 407868 488956 407869 489020
rect 407803 488955 407869 488956
rect 407619 189684 407685 189685
rect 407619 189620 407620 189684
rect 407684 189620 407685 189684
rect 407619 189619 407685 189620
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406331 154324 406397 154325
rect 406331 154260 406332 154324
rect 406396 154260 406397 154324
rect 406331 154259 406397 154260
rect 406794 152000 407414 155898
rect 407806 155277 407866 488955
rect 408358 466581 408418 678267
rect 408539 476236 408605 476237
rect 408539 476172 408540 476236
rect 408604 476172 408605 476236
rect 408539 476171 408605 476172
rect 408355 466580 408421 466581
rect 408355 466516 408356 466580
rect 408420 466516 408421 466580
rect 408355 466515 408421 466516
rect 407987 378180 408053 378181
rect 407987 378116 407988 378180
rect 408052 378116 408053 378180
rect 407987 378115 408053 378116
rect 407990 184381 408050 378115
rect 407987 184380 408053 184381
rect 407987 184316 407988 184380
rect 408052 184316 408053 184380
rect 407987 184315 408053 184316
rect 407803 155276 407869 155277
rect 407803 155212 407804 155276
rect 407868 155212 407869 155276
rect 407803 155211 407869 155212
rect 408542 152693 408602 476171
rect 409459 316980 409525 316981
rect 409459 316916 409460 316980
rect 409524 316916 409525 316980
rect 409459 316915 409525 316916
rect 409091 262988 409157 262989
rect 409091 262924 409092 262988
rect 409156 262924 409157 262988
rect 409091 262923 409157 262924
rect 409094 157181 409154 262923
rect 409091 157180 409157 157181
rect 409091 157116 409092 157180
rect 409156 157116 409157 157180
rect 409091 157115 409157 157116
rect 409462 157045 409522 316915
rect 409646 277541 409706 679763
rect 409830 678333 409890 683299
rect 411294 682000 411914 700398
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 682000 429914 682398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 682000 434414 686898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 682000 438914 691398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 682000 443414 695898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 682000 447914 700398
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 682000 465914 682398
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 682000 470414 686898
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 682000 474914 691398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 682000 479414 695898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 682000 483914 700398
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 682000 501914 682398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 682000 506414 686898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 682000 510914 691398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 682000 515414 695898
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 682000 519914 700398
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 682000 537914 682398
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 682000 542414 686898
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 682000 546914 691398
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 551507 700364 551573 700365
rect 551507 700300 551508 700364
rect 551572 700300 551573 700364
rect 551507 700299 551573 700300
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 682000 551414 695898
rect 409827 678332 409893 678333
rect 409827 678268 409828 678332
rect 409892 678268 409893 678332
rect 409827 678267 409893 678268
rect 429568 655954 429888 655986
rect 429568 655718 429610 655954
rect 429846 655718 429888 655954
rect 429568 655634 429888 655718
rect 429568 655398 429610 655634
rect 429846 655398 429888 655634
rect 429568 655366 429888 655398
rect 460288 655954 460608 655986
rect 460288 655718 460330 655954
rect 460566 655718 460608 655954
rect 460288 655634 460608 655718
rect 460288 655398 460330 655634
rect 460566 655398 460608 655634
rect 460288 655366 460608 655398
rect 491008 655954 491328 655986
rect 491008 655718 491050 655954
rect 491286 655718 491328 655954
rect 491008 655634 491328 655718
rect 491008 655398 491050 655634
rect 491286 655398 491328 655634
rect 491008 655366 491328 655398
rect 521728 655954 522048 655986
rect 521728 655718 521770 655954
rect 522006 655718 522048 655954
rect 521728 655634 522048 655718
rect 521728 655398 521770 655634
rect 522006 655398 522048 655634
rect 521728 655366 522048 655398
rect 414208 651454 414528 651486
rect 414208 651218 414250 651454
rect 414486 651218 414528 651454
rect 414208 651134 414528 651218
rect 414208 650898 414250 651134
rect 414486 650898 414528 651134
rect 414208 650866 414528 650898
rect 444928 651454 445248 651486
rect 444928 651218 444970 651454
rect 445206 651218 445248 651454
rect 444928 651134 445248 651218
rect 444928 650898 444970 651134
rect 445206 650898 445248 651134
rect 444928 650866 445248 650898
rect 475648 651454 475968 651486
rect 475648 651218 475690 651454
rect 475926 651218 475968 651454
rect 475648 651134 475968 651218
rect 475648 650898 475690 651134
rect 475926 650898 475968 651134
rect 475648 650866 475968 650898
rect 506368 651454 506688 651486
rect 506368 651218 506410 651454
rect 506646 651218 506688 651454
rect 506368 651134 506688 651218
rect 506368 650898 506410 651134
rect 506646 650898 506688 651134
rect 506368 650866 506688 650898
rect 537088 651454 537408 651486
rect 537088 651218 537130 651454
rect 537366 651218 537408 651454
rect 537088 651134 537408 651218
rect 537088 650898 537130 651134
rect 537366 650898 537408 651134
rect 537088 650866 537408 650898
rect 429568 619954 429888 619986
rect 429568 619718 429610 619954
rect 429846 619718 429888 619954
rect 429568 619634 429888 619718
rect 429568 619398 429610 619634
rect 429846 619398 429888 619634
rect 429568 619366 429888 619398
rect 460288 619954 460608 619986
rect 460288 619718 460330 619954
rect 460566 619718 460608 619954
rect 460288 619634 460608 619718
rect 460288 619398 460330 619634
rect 460566 619398 460608 619634
rect 460288 619366 460608 619398
rect 491008 619954 491328 619986
rect 491008 619718 491050 619954
rect 491286 619718 491328 619954
rect 491008 619634 491328 619718
rect 491008 619398 491050 619634
rect 491286 619398 491328 619634
rect 491008 619366 491328 619398
rect 521728 619954 522048 619986
rect 521728 619718 521770 619954
rect 522006 619718 522048 619954
rect 521728 619634 522048 619718
rect 521728 619398 521770 619634
rect 522006 619398 522048 619634
rect 521728 619366 522048 619398
rect 414208 615454 414528 615486
rect 414208 615218 414250 615454
rect 414486 615218 414528 615454
rect 414208 615134 414528 615218
rect 414208 614898 414250 615134
rect 414486 614898 414528 615134
rect 414208 614866 414528 614898
rect 444928 615454 445248 615486
rect 444928 615218 444970 615454
rect 445206 615218 445248 615454
rect 444928 615134 445248 615218
rect 444928 614898 444970 615134
rect 445206 614898 445248 615134
rect 444928 614866 445248 614898
rect 475648 615454 475968 615486
rect 475648 615218 475690 615454
rect 475926 615218 475968 615454
rect 475648 615134 475968 615218
rect 475648 614898 475690 615134
rect 475926 614898 475968 615134
rect 475648 614866 475968 614898
rect 506368 615454 506688 615486
rect 506368 615218 506410 615454
rect 506646 615218 506688 615454
rect 506368 615134 506688 615218
rect 506368 614898 506410 615134
rect 506646 614898 506688 615134
rect 506368 614866 506688 614898
rect 537088 615454 537408 615486
rect 537088 615218 537130 615454
rect 537366 615218 537408 615454
rect 537088 615134 537408 615218
rect 537088 614898 537130 615134
rect 537366 614898 537408 615134
rect 537088 614866 537408 614898
rect 551510 597549 551570 700299
rect 552243 685948 552309 685949
rect 552243 685884 552244 685948
rect 552308 685884 552309 685948
rect 552243 685883 552309 685884
rect 552059 682684 552125 682685
rect 552059 682620 552060 682684
rect 552124 682620 552125 682684
rect 552059 682619 552125 682620
rect 551507 597548 551573 597549
rect 551507 597484 551508 597548
rect 551572 597484 551573 597548
rect 551507 597483 551573 597484
rect 550403 591632 550469 591633
rect 550403 591568 550404 591632
rect 550468 591568 550469 591632
rect 550403 591567 550469 591568
rect 550406 590749 550466 591567
rect 550403 590748 550469 590749
rect 550403 590684 550404 590748
rect 550468 590684 550469 590748
rect 550403 590683 550469 590684
rect 429568 583954 429888 583986
rect 429568 583718 429610 583954
rect 429846 583718 429888 583954
rect 429568 583634 429888 583718
rect 429568 583398 429610 583634
rect 429846 583398 429888 583634
rect 429568 583366 429888 583398
rect 460288 583954 460608 583986
rect 460288 583718 460330 583954
rect 460566 583718 460608 583954
rect 460288 583634 460608 583718
rect 460288 583398 460330 583634
rect 460566 583398 460608 583634
rect 460288 583366 460608 583398
rect 491008 583954 491328 583986
rect 491008 583718 491050 583954
rect 491286 583718 491328 583954
rect 491008 583634 491328 583718
rect 491008 583398 491050 583634
rect 491286 583398 491328 583634
rect 491008 583366 491328 583398
rect 521728 583954 522048 583986
rect 521728 583718 521770 583954
rect 522006 583718 522048 583954
rect 521728 583634 522048 583718
rect 521728 583398 521770 583634
rect 522006 583398 522048 583634
rect 521728 583366 522048 583398
rect 414208 579454 414528 579486
rect 414208 579218 414250 579454
rect 414486 579218 414528 579454
rect 414208 579134 414528 579218
rect 414208 578898 414250 579134
rect 414486 578898 414528 579134
rect 414208 578866 414528 578898
rect 444928 579454 445248 579486
rect 444928 579218 444970 579454
rect 445206 579218 445248 579454
rect 444928 579134 445248 579218
rect 444928 578898 444970 579134
rect 445206 578898 445248 579134
rect 444928 578866 445248 578898
rect 475648 579454 475968 579486
rect 475648 579218 475690 579454
rect 475926 579218 475968 579454
rect 475648 579134 475968 579218
rect 475648 578898 475690 579134
rect 475926 578898 475968 579134
rect 475648 578866 475968 578898
rect 506368 579454 506688 579486
rect 506368 579218 506410 579454
rect 506646 579218 506688 579454
rect 506368 579134 506688 579218
rect 506368 578898 506410 579134
rect 506646 578898 506688 579134
rect 506368 578866 506688 578898
rect 537088 579454 537408 579486
rect 537088 579218 537130 579454
rect 537366 579218 537408 579454
rect 537088 579134 537408 579218
rect 537088 578898 537130 579134
rect 537366 578898 537408 579134
rect 537088 578866 537408 578898
rect 429568 547954 429888 547986
rect 429568 547718 429610 547954
rect 429846 547718 429888 547954
rect 429568 547634 429888 547718
rect 429568 547398 429610 547634
rect 429846 547398 429888 547634
rect 429568 547366 429888 547398
rect 460288 547954 460608 547986
rect 460288 547718 460330 547954
rect 460566 547718 460608 547954
rect 460288 547634 460608 547718
rect 460288 547398 460330 547634
rect 460566 547398 460608 547634
rect 460288 547366 460608 547398
rect 491008 547954 491328 547986
rect 491008 547718 491050 547954
rect 491286 547718 491328 547954
rect 491008 547634 491328 547718
rect 491008 547398 491050 547634
rect 491286 547398 491328 547634
rect 491008 547366 491328 547398
rect 521728 547954 522048 547986
rect 521728 547718 521770 547954
rect 522006 547718 522048 547954
rect 521728 547634 522048 547718
rect 521728 547398 521770 547634
rect 522006 547398 522048 547634
rect 521728 547366 522048 547398
rect 414208 543454 414528 543486
rect 414208 543218 414250 543454
rect 414486 543218 414528 543454
rect 414208 543134 414528 543218
rect 414208 542898 414250 543134
rect 414486 542898 414528 543134
rect 414208 542866 414528 542898
rect 444928 543454 445248 543486
rect 444928 543218 444970 543454
rect 445206 543218 445248 543454
rect 444928 543134 445248 543218
rect 444928 542898 444970 543134
rect 445206 542898 445248 543134
rect 444928 542866 445248 542898
rect 475648 543454 475968 543486
rect 475648 543218 475690 543454
rect 475926 543218 475968 543454
rect 475648 543134 475968 543218
rect 475648 542898 475690 543134
rect 475926 542898 475968 543134
rect 475648 542866 475968 542898
rect 506368 543454 506688 543486
rect 506368 543218 506410 543454
rect 506646 543218 506688 543454
rect 506368 543134 506688 543218
rect 506368 542898 506410 543134
rect 506646 542898 506688 543134
rect 506368 542866 506688 542898
rect 537088 543454 537408 543486
rect 537088 543218 537130 543454
rect 537366 543218 537408 543454
rect 537088 543134 537408 543218
rect 537088 542898 537130 543134
rect 537366 542898 537408 543134
rect 537088 542866 537408 542898
rect 429568 511954 429888 511986
rect 429568 511718 429610 511954
rect 429846 511718 429888 511954
rect 429568 511634 429888 511718
rect 429568 511398 429610 511634
rect 429846 511398 429888 511634
rect 429568 511366 429888 511398
rect 460288 511954 460608 511986
rect 460288 511718 460330 511954
rect 460566 511718 460608 511954
rect 460288 511634 460608 511718
rect 460288 511398 460330 511634
rect 460566 511398 460608 511634
rect 460288 511366 460608 511398
rect 491008 511954 491328 511986
rect 491008 511718 491050 511954
rect 491286 511718 491328 511954
rect 491008 511634 491328 511718
rect 491008 511398 491050 511634
rect 491286 511398 491328 511634
rect 491008 511366 491328 511398
rect 521728 511954 522048 511986
rect 521728 511718 521770 511954
rect 522006 511718 522048 511954
rect 521728 511634 522048 511718
rect 521728 511398 521770 511634
rect 522006 511398 522048 511634
rect 521728 511366 522048 511398
rect 414208 507454 414528 507486
rect 414208 507218 414250 507454
rect 414486 507218 414528 507454
rect 414208 507134 414528 507218
rect 414208 506898 414250 507134
rect 414486 506898 414528 507134
rect 414208 506866 414528 506898
rect 444928 507454 445248 507486
rect 444928 507218 444970 507454
rect 445206 507218 445248 507454
rect 444928 507134 445248 507218
rect 444928 506898 444970 507134
rect 445206 506898 445248 507134
rect 444928 506866 445248 506898
rect 475648 507454 475968 507486
rect 475648 507218 475690 507454
rect 475926 507218 475968 507454
rect 475648 507134 475968 507218
rect 475648 506898 475690 507134
rect 475926 506898 475968 507134
rect 475648 506866 475968 506898
rect 506368 507454 506688 507486
rect 506368 507218 506410 507454
rect 506646 507218 506688 507454
rect 506368 507134 506688 507218
rect 506368 506898 506410 507134
rect 506646 506898 506688 507134
rect 506368 506866 506688 506898
rect 537088 507454 537408 507486
rect 537088 507218 537130 507454
rect 537366 507218 537408 507454
rect 537088 507134 537408 507218
rect 537088 506898 537130 507134
rect 537366 506898 537408 507134
rect 537088 506866 537408 506898
rect 550771 497180 550837 497181
rect 550771 497116 550772 497180
rect 550836 497116 550837 497180
rect 550771 497115 550837 497116
rect 429568 475954 429888 475986
rect 429568 475718 429610 475954
rect 429846 475718 429888 475954
rect 429568 475634 429888 475718
rect 429568 475398 429610 475634
rect 429846 475398 429888 475634
rect 429568 475366 429888 475398
rect 460288 475954 460608 475986
rect 460288 475718 460330 475954
rect 460566 475718 460608 475954
rect 460288 475634 460608 475718
rect 460288 475398 460330 475634
rect 460566 475398 460608 475634
rect 460288 475366 460608 475398
rect 491008 475954 491328 475986
rect 491008 475718 491050 475954
rect 491286 475718 491328 475954
rect 491008 475634 491328 475718
rect 491008 475398 491050 475634
rect 491286 475398 491328 475634
rect 491008 475366 491328 475398
rect 521728 475954 522048 475986
rect 521728 475718 521770 475954
rect 522006 475718 522048 475954
rect 521728 475634 522048 475718
rect 521728 475398 521770 475634
rect 522006 475398 522048 475634
rect 521728 475366 522048 475398
rect 414208 471454 414528 471486
rect 414208 471218 414250 471454
rect 414486 471218 414528 471454
rect 414208 471134 414528 471218
rect 414208 470898 414250 471134
rect 414486 470898 414528 471134
rect 414208 470866 414528 470898
rect 444928 471454 445248 471486
rect 444928 471218 444970 471454
rect 445206 471218 445248 471454
rect 444928 471134 445248 471218
rect 444928 470898 444970 471134
rect 445206 470898 445248 471134
rect 444928 470866 445248 470898
rect 475648 471454 475968 471486
rect 475648 471218 475690 471454
rect 475926 471218 475968 471454
rect 475648 471134 475968 471218
rect 475648 470898 475690 471134
rect 475926 470898 475968 471134
rect 475648 470866 475968 470898
rect 506368 471454 506688 471486
rect 506368 471218 506410 471454
rect 506646 471218 506688 471454
rect 506368 471134 506688 471218
rect 506368 470898 506410 471134
rect 506646 470898 506688 471134
rect 506368 470866 506688 470898
rect 537088 471454 537408 471486
rect 537088 471218 537130 471454
rect 537366 471218 537408 471454
rect 537088 471134 537408 471218
rect 537088 470898 537130 471134
rect 537366 470898 537408 471134
rect 537088 470866 537408 470898
rect 550219 440740 550285 440741
rect 550219 440676 550220 440740
rect 550284 440676 550285 440740
rect 550219 440675 550285 440676
rect 429568 439954 429888 439986
rect 429568 439718 429610 439954
rect 429846 439718 429888 439954
rect 429568 439634 429888 439718
rect 429568 439398 429610 439634
rect 429846 439398 429888 439634
rect 429568 439366 429888 439398
rect 460288 439954 460608 439986
rect 460288 439718 460330 439954
rect 460566 439718 460608 439954
rect 460288 439634 460608 439718
rect 460288 439398 460330 439634
rect 460566 439398 460608 439634
rect 460288 439366 460608 439398
rect 491008 439954 491328 439986
rect 491008 439718 491050 439954
rect 491286 439718 491328 439954
rect 491008 439634 491328 439718
rect 491008 439398 491050 439634
rect 491286 439398 491328 439634
rect 491008 439366 491328 439398
rect 521728 439954 522048 439986
rect 521728 439718 521770 439954
rect 522006 439718 522048 439954
rect 521728 439634 522048 439718
rect 521728 439398 521770 439634
rect 522006 439398 522048 439634
rect 521728 439366 522048 439398
rect 414208 435454 414528 435486
rect 414208 435218 414250 435454
rect 414486 435218 414528 435454
rect 414208 435134 414528 435218
rect 414208 434898 414250 435134
rect 414486 434898 414528 435134
rect 414208 434866 414528 434898
rect 444928 435454 445248 435486
rect 444928 435218 444970 435454
rect 445206 435218 445248 435454
rect 444928 435134 445248 435218
rect 444928 434898 444970 435134
rect 445206 434898 445248 435134
rect 444928 434866 445248 434898
rect 475648 435454 475968 435486
rect 475648 435218 475690 435454
rect 475926 435218 475968 435454
rect 475648 435134 475968 435218
rect 475648 434898 475690 435134
rect 475926 434898 475968 435134
rect 475648 434866 475968 434898
rect 506368 435454 506688 435486
rect 506368 435218 506410 435454
rect 506646 435218 506688 435454
rect 506368 435134 506688 435218
rect 506368 434898 506410 435134
rect 506646 434898 506688 435134
rect 506368 434866 506688 434898
rect 537088 435454 537408 435486
rect 537088 435218 537130 435454
rect 537366 435218 537408 435454
rect 537088 435134 537408 435218
rect 537088 434898 537130 435134
rect 537366 434898 537408 435134
rect 537088 434866 537408 434898
rect 429568 403954 429888 403986
rect 429568 403718 429610 403954
rect 429846 403718 429888 403954
rect 429568 403634 429888 403718
rect 429568 403398 429610 403634
rect 429846 403398 429888 403634
rect 429568 403366 429888 403398
rect 460288 403954 460608 403986
rect 460288 403718 460330 403954
rect 460566 403718 460608 403954
rect 460288 403634 460608 403718
rect 460288 403398 460330 403634
rect 460566 403398 460608 403634
rect 460288 403366 460608 403398
rect 491008 403954 491328 403986
rect 491008 403718 491050 403954
rect 491286 403718 491328 403954
rect 491008 403634 491328 403718
rect 491008 403398 491050 403634
rect 491286 403398 491328 403634
rect 491008 403366 491328 403398
rect 521728 403954 522048 403986
rect 521728 403718 521770 403954
rect 522006 403718 522048 403954
rect 521728 403634 522048 403718
rect 521728 403398 521770 403634
rect 522006 403398 522048 403634
rect 521728 403366 522048 403398
rect 414208 399454 414528 399486
rect 414208 399218 414250 399454
rect 414486 399218 414528 399454
rect 414208 399134 414528 399218
rect 414208 398898 414250 399134
rect 414486 398898 414528 399134
rect 414208 398866 414528 398898
rect 444928 399454 445248 399486
rect 444928 399218 444970 399454
rect 445206 399218 445248 399454
rect 444928 399134 445248 399218
rect 444928 398898 444970 399134
rect 445206 398898 445248 399134
rect 444928 398866 445248 398898
rect 475648 399454 475968 399486
rect 475648 399218 475690 399454
rect 475926 399218 475968 399454
rect 475648 399134 475968 399218
rect 475648 398898 475690 399134
rect 475926 398898 475968 399134
rect 475648 398866 475968 398898
rect 506368 399454 506688 399486
rect 506368 399218 506410 399454
rect 506646 399218 506688 399454
rect 506368 399134 506688 399218
rect 506368 398898 506410 399134
rect 506646 398898 506688 399134
rect 506368 398866 506688 398898
rect 537088 399454 537408 399486
rect 537088 399218 537130 399454
rect 537366 399218 537408 399454
rect 537088 399134 537408 399218
rect 537088 398898 537130 399134
rect 537366 398898 537408 399134
rect 537088 398866 537408 398898
rect 429568 367954 429888 367986
rect 429568 367718 429610 367954
rect 429846 367718 429888 367954
rect 429568 367634 429888 367718
rect 429568 367398 429610 367634
rect 429846 367398 429888 367634
rect 429568 367366 429888 367398
rect 460288 367954 460608 367986
rect 460288 367718 460330 367954
rect 460566 367718 460608 367954
rect 460288 367634 460608 367718
rect 460288 367398 460330 367634
rect 460566 367398 460608 367634
rect 460288 367366 460608 367398
rect 491008 367954 491328 367986
rect 491008 367718 491050 367954
rect 491286 367718 491328 367954
rect 491008 367634 491328 367718
rect 491008 367398 491050 367634
rect 491286 367398 491328 367634
rect 491008 367366 491328 367398
rect 521728 367954 522048 367986
rect 521728 367718 521770 367954
rect 522006 367718 522048 367954
rect 521728 367634 522048 367718
rect 521728 367398 521770 367634
rect 522006 367398 522048 367634
rect 521728 367366 522048 367398
rect 414208 363454 414528 363486
rect 414208 363218 414250 363454
rect 414486 363218 414528 363454
rect 414208 363134 414528 363218
rect 414208 362898 414250 363134
rect 414486 362898 414528 363134
rect 414208 362866 414528 362898
rect 444928 363454 445248 363486
rect 444928 363218 444970 363454
rect 445206 363218 445248 363454
rect 444928 363134 445248 363218
rect 444928 362898 444970 363134
rect 445206 362898 445248 363134
rect 444928 362866 445248 362898
rect 475648 363454 475968 363486
rect 475648 363218 475690 363454
rect 475926 363218 475968 363454
rect 475648 363134 475968 363218
rect 475648 362898 475690 363134
rect 475926 362898 475968 363134
rect 475648 362866 475968 362898
rect 506368 363454 506688 363486
rect 506368 363218 506410 363454
rect 506646 363218 506688 363454
rect 506368 363134 506688 363218
rect 506368 362898 506410 363134
rect 506646 362898 506688 363134
rect 506368 362866 506688 362898
rect 537088 363454 537408 363486
rect 537088 363218 537130 363454
rect 537366 363218 537408 363454
rect 537088 363134 537408 363218
rect 537088 362898 537130 363134
rect 537366 362898 537408 363134
rect 537088 362866 537408 362898
rect 429568 331954 429888 331986
rect 429568 331718 429610 331954
rect 429846 331718 429888 331954
rect 429568 331634 429888 331718
rect 429568 331398 429610 331634
rect 429846 331398 429888 331634
rect 429568 331366 429888 331398
rect 460288 331954 460608 331986
rect 460288 331718 460330 331954
rect 460566 331718 460608 331954
rect 460288 331634 460608 331718
rect 460288 331398 460330 331634
rect 460566 331398 460608 331634
rect 460288 331366 460608 331398
rect 491008 331954 491328 331986
rect 491008 331718 491050 331954
rect 491286 331718 491328 331954
rect 491008 331634 491328 331718
rect 491008 331398 491050 331634
rect 491286 331398 491328 331634
rect 491008 331366 491328 331398
rect 521728 331954 522048 331986
rect 521728 331718 521770 331954
rect 522006 331718 522048 331954
rect 521728 331634 522048 331718
rect 521728 331398 521770 331634
rect 522006 331398 522048 331634
rect 521728 331366 522048 331398
rect 414208 327454 414528 327486
rect 414208 327218 414250 327454
rect 414486 327218 414528 327454
rect 414208 327134 414528 327218
rect 414208 326898 414250 327134
rect 414486 326898 414528 327134
rect 414208 326866 414528 326898
rect 444928 327454 445248 327486
rect 444928 327218 444970 327454
rect 445206 327218 445248 327454
rect 444928 327134 445248 327218
rect 444928 326898 444970 327134
rect 445206 326898 445248 327134
rect 444928 326866 445248 326898
rect 475648 327454 475968 327486
rect 475648 327218 475690 327454
rect 475926 327218 475968 327454
rect 475648 327134 475968 327218
rect 475648 326898 475690 327134
rect 475926 326898 475968 327134
rect 475648 326866 475968 326898
rect 506368 327454 506688 327486
rect 506368 327218 506410 327454
rect 506646 327218 506688 327454
rect 506368 327134 506688 327218
rect 506368 326898 506410 327134
rect 506646 326898 506688 327134
rect 506368 326866 506688 326898
rect 537088 327454 537408 327486
rect 537088 327218 537130 327454
rect 537366 327218 537408 327454
rect 537088 327134 537408 327218
rect 537088 326898 537130 327134
rect 537366 326898 537408 327134
rect 537088 326866 537408 326898
rect 429568 295954 429888 295986
rect 429568 295718 429610 295954
rect 429846 295718 429888 295954
rect 429568 295634 429888 295718
rect 429568 295398 429610 295634
rect 429846 295398 429888 295634
rect 429568 295366 429888 295398
rect 460288 295954 460608 295986
rect 460288 295718 460330 295954
rect 460566 295718 460608 295954
rect 460288 295634 460608 295718
rect 460288 295398 460330 295634
rect 460566 295398 460608 295634
rect 460288 295366 460608 295398
rect 491008 295954 491328 295986
rect 491008 295718 491050 295954
rect 491286 295718 491328 295954
rect 491008 295634 491328 295718
rect 491008 295398 491050 295634
rect 491286 295398 491328 295634
rect 491008 295366 491328 295398
rect 521728 295954 522048 295986
rect 521728 295718 521770 295954
rect 522006 295718 522048 295954
rect 521728 295634 522048 295718
rect 521728 295398 521770 295634
rect 522006 295398 522048 295634
rect 521728 295366 522048 295398
rect 414208 291454 414528 291486
rect 414208 291218 414250 291454
rect 414486 291218 414528 291454
rect 414208 291134 414528 291218
rect 414208 290898 414250 291134
rect 414486 290898 414528 291134
rect 414208 290866 414528 290898
rect 444928 291454 445248 291486
rect 444928 291218 444970 291454
rect 445206 291218 445248 291454
rect 444928 291134 445248 291218
rect 444928 290898 444970 291134
rect 445206 290898 445248 291134
rect 444928 290866 445248 290898
rect 475648 291454 475968 291486
rect 475648 291218 475690 291454
rect 475926 291218 475968 291454
rect 475648 291134 475968 291218
rect 475648 290898 475690 291134
rect 475926 290898 475968 291134
rect 475648 290866 475968 290898
rect 506368 291454 506688 291486
rect 506368 291218 506410 291454
rect 506646 291218 506688 291454
rect 506368 291134 506688 291218
rect 506368 290898 506410 291134
rect 506646 290898 506688 291134
rect 506368 290866 506688 290898
rect 537088 291454 537408 291486
rect 537088 291218 537130 291454
rect 537366 291218 537408 291454
rect 537088 291134 537408 291218
rect 537088 290898 537130 291134
rect 537366 290898 537408 291134
rect 537088 290866 537408 290898
rect 409643 277540 409709 277541
rect 409643 277476 409644 277540
rect 409708 277476 409709 277540
rect 409643 277475 409709 277476
rect 429568 259954 429888 259986
rect 429568 259718 429610 259954
rect 429846 259718 429888 259954
rect 429568 259634 429888 259718
rect 429568 259398 429610 259634
rect 429846 259398 429888 259634
rect 429568 259366 429888 259398
rect 460288 259954 460608 259986
rect 460288 259718 460330 259954
rect 460566 259718 460608 259954
rect 460288 259634 460608 259718
rect 460288 259398 460330 259634
rect 460566 259398 460608 259634
rect 460288 259366 460608 259398
rect 491008 259954 491328 259986
rect 491008 259718 491050 259954
rect 491286 259718 491328 259954
rect 491008 259634 491328 259718
rect 491008 259398 491050 259634
rect 491286 259398 491328 259634
rect 491008 259366 491328 259398
rect 521728 259954 522048 259986
rect 521728 259718 521770 259954
rect 522006 259718 522048 259954
rect 521728 259634 522048 259718
rect 521728 259398 521770 259634
rect 522006 259398 522048 259634
rect 521728 259366 522048 259398
rect 414208 255454 414528 255486
rect 414208 255218 414250 255454
rect 414486 255218 414528 255454
rect 414208 255134 414528 255218
rect 414208 254898 414250 255134
rect 414486 254898 414528 255134
rect 414208 254866 414528 254898
rect 444928 255454 445248 255486
rect 444928 255218 444970 255454
rect 445206 255218 445248 255454
rect 444928 255134 445248 255218
rect 444928 254898 444970 255134
rect 445206 254898 445248 255134
rect 444928 254866 445248 254898
rect 475648 255454 475968 255486
rect 475648 255218 475690 255454
rect 475926 255218 475968 255454
rect 475648 255134 475968 255218
rect 475648 254898 475690 255134
rect 475926 254898 475968 255134
rect 475648 254866 475968 254898
rect 506368 255454 506688 255486
rect 506368 255218 506410 255454
rect 506646 255218 506688 255454
rect 506368 255134 506688 255218
rect 506368 254898 506410 255134
rect 506646 254898 506688 255134
rect 506368 254866 506688 254898
rect 537088 255454 537408 255486
rect 537088 255218 537130 255454
rect 537366 255218 537408 255454
rect 537088 255134 537408 255218
rect 537088 254898 537130 255134
rect 537366 254898 537408 255134
rect 537088 254866 537408 254898
rect 409827 242860 409893 242861
rect 409827 242796 409828 242860
rect 409892 242796 409893 242860
rect 409827 242795 409893 242796
rect 409459 157044 409525 157045
rect 409459 156980 409460 157044
rect 409524 156980 409525 157044
rect 409459 156979 409525 156980
rect 409830 152693 409890 242795
rect 410011 242588 410077 242589
rect 410011 242524 410012 242588
rect 410076 242524 410077 242588
rect 410011 242523 410077 242524
rect 410014 238770 410074 242523
rect 410014 238710 410258 238770
rect 408539 152692 408605 152693
rect 408539 152628 408540 152692
rect 408604 152628 408605 152692
rect 408539 152627 408605 152628
rect 409827 152692 409893 152693
rect 409827 152628 409828 152692
rect 409892 152628 409893 152692
rect 409827 152627 409893 152628
rect 410198 151469 410258 238710
rect 411294 232954 411914 238000
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 152000 411914 160398
rect 415794 237454 416414 238000
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 152000 416414 164898
rect 420294 205954 420914 238000
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 152000 420914 169398
rect 424794 210454 425414 238000
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 152000 425414 173898
rect 429294 214954 429914 238000
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 152000 429914 178398
rect 433794 219454 434414 238000
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 152000 434414 182898
rect 438294 223954 438914 238000
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 152000 438914 187398
rect 442794 228454 443414 238000
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 152000 443414 155898
rect 447294 232954 447914 238000
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 152000 447914 160398
rect 451794 237454 452414 238000
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 152000 452414 164898
rect 456294 205954 456914 238000
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 152000 456914 169398
rect 460794 210454 461414 238000
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 152000 461414 173898
rect 465294 214954 465914 238000
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 152000 465914 178398
rect 469794 219454 470414 238000
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 152000 470414 182898
rect 474294 223954 474914 238000
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 152000 474914 187398
rect 478794 228454 479414 238000
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 152000 479414 155898
rect 483294 232954 483914 238000
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 152000 483914 160398
rect 487794 237454 488414 238000
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 152000 488414 164898
rect 492294 205954 492914 238000
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 152000 492914 169398
rect 496794 210454 497414 238000
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 152000 497414 173898
rect 501294 214954 501914 238000
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 152000 501914 178398
rect 505794 219454 506414 238000
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 152000 506414 182898
rect 510294 223954 510914 238000
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 152000 510914 187398
rect 514794 228454 515414 238000
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 152000 515414 155898
rect 519294 232954 519914 238000
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 152000 519914 160398
rect 523794 237454 524414 238000
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 152000 524414 164898
rect 528294 205954 528914 238000
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 152000 528914 169398
rect 532794 210454 533414 238000
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 152000 533414 173898
rect 537294 214954 537914 238000
rect 540283 235516 540349 235517
rect 540283 235452 540284 235516
rect 540348 235452 540349 235516
rect 540283 235451 540349 235452
rect 538811 234292 538877 234293
rect 538811 234228 538812 234292
rect 538876 234228 538877 234292
rect 538811 234227 538877 234228
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 152000 537914 178398
rect 410195 151468 410261 151469
rect 410195 151404 410196 151468
rect 410260 151404 410261 151468
rect 410195 151403 410261 151404
rect 372659 151060 372725 151061
rect 372659 150996 372660 151060
rect 372724 150996 372725 151060
rect 372659 150995 372725 150996
rect 404859 151060 404925 151061
rect 404859 150996 404860 151060
rect 404924 150996 404925 151060
rect 404859 150995 404925 150996
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 248528 147454 248848 147486
rect 248528 147218 248570 147454
rect 248806 147218 248848 147454
rect 248528 147134 248848 147218
rect 248528 146898 248570 147134
rect 248806 146898 248848 147134
rect 248528 146866 248848 146898
rect 279248 147454 279568 147486
rect 279248 147218 279290 147454
rect 279526 147218 279568 147454
rect 279248 147134 279568 147218
rect 279248 146898 279290 147134
rect 279526 146898 279568 147134
rect 279248 146866 279568 146898
rect 309968 147454 310288 147486
rect 309968 147218 310010 147454
rect 310246 147218 310288 147454
rect 309968 147134 310288 147218
rect 309968 146898 310010 147134
rect 310246 146898 310288 147134
rect 309968 146866 310288 146898
rect 340688 147454 341008 147486
rect 340688 147218 340730 147454
rect 340966 147218 341008 147454
rect 340688 147134 341008 147218
rect 340688 146898 340730 147134
rect 340966 146898 341008 147134
rect 340688 146866 341008 146898
rect 371408 147454 371728 147486
rect 371408 147218 371450 147454
rect 371686 147218 371728 147454
rect 371408 147134 371728 147218
rect 371408 146898 371450 147134
rect 371686 146898 371728 147134
rect 371408 146866 371728 146898
rect 402128 147454 402448 147486
rect 402128 147218 402170 147454
rect 402406 147218 402448 147454
rect 402128 147134 402448 147218
rect 402128 146898 402170 147134
rect 402406 146898 402448 147134
rect 402128 146866 402448 146898
rect 432848 147454 433168 147486
rect 432848 147218 432890 147454
rect 433126 147218 433168 147454
rect 432848 147134 433168 147218
rect 432848 146898 432890 147134
rect 433126 146898 433168 147134
rect 432848 146866 433168 146898
rect 463568 147454 463888 147486
rect 463568 147218 463610 147454
rect 463846 147218 463888 147454
rect 463568 147134 463888 147218
rect 463568 146898 463610 147134
rect 463846 146898 463888 147134
rect 463568 146866 463888 146898
rect 494288 147454 494608 147486
rect 494288 147218 494330 147454
rect 494566 147218 494608 147454
rect 494288 147134 494608 147218
rect 494288 146898 494330 147134
rect 494566 146898 494608 147134
rect 494288 146866 494608 146898
rect 525008 147454 525328 147486
rect 525008 147218 525050 147454
rect 525286 147218 525328 147454
rect 525008 147134 525328 147218
rect 525008 146898 525050 147134
rect 525286 146898 525328 147134
rect 525008 146866 525328 146898
rect 60782 146510 61762 146570
rect 538814 146570 538874 234227
rect 538995 232524 539061 232525
rect 538995 232460 538996 232524
rect 539060 232460 539061 232524
rect 538995 232459 539061 232460
rect 538998 147250 539058 232459
rect 539179 231708 539245 231709
rect 539179 231644 539180 231708
rect 539244 231644 539245 231708
rect 539179 231643 539245 231644
rect 539182 150517 539242 231643
rect 539547 186964 539613 186965
rect 539547 186900 539548 186964
rect 539612 186900 539613 186964
rect 539547 186899 539613 186900
rect 539363 158676 539429 158677
rect 539363 158612 539364 158676
rect 539428 158612 539429 158676
rect 539363 158611 539429 158612
rect 539179 150516 539245 150517
rect 539179 150452 539180 150516
rect 539244 150452 539245 150516
rect 539179 150451 539245 150452
rect 539366 147389 539426 158611
rect 539363 147388 539429 147389
rect 539363 147324 539364 147388
rect 539428 147324 539429 147388
rect 539363 147323 539429 147324
rect 538998 147190 539426 147250
rect 539366 146845 539426 147190
rect 539363 146844 539429 146845
rect 539363 146780 539364 146844
rect 539428 146780 539429 146844
rect 539363 146779 539429 146780
rect 539363 146572 539429 146573
rect 539363 146570 539364 146572
rect 538814 146510 539364 146570
rect 60782 145890 60842 146510
rect 539363 146508 539364 146510
rect 539428 146508 539429 146572
rect 539363 146507 539429 146508
rect 60598 145830 60842 145890
rect 60598 139229 60658 145830
rect 539363 145484 539429 145485
rect 539363 145420 539364 145484
rect 539428 145420 539429 145484
rect 539363 145419 539429 145420
rect 539366 141813 539426 145419
rect 539363 141812 539429 141813
rect 539363 141748 539364 141812
rect 539428 141748 539429 141812
rect 539363 141747 539429 141748
rect 60595 139228 60661 139229
rect 60595 139164 60596 139228
rect 60660 139164 60661 139228
rect 60595 139163 60661 139164
rect 60414 137970 60658 138030
rect 59491 125492 59557 125493
rect 59491 125428 59492 125492
rect 59556 125428 59557 125492
rect 59491 125427 59557 125428
rect 59678 122093 59738 137970
rect 59859 123452 59925 123453
rect 59859 123388 59860 123452
rect 59924 123388 59925 123452
rect 59859 123387 59925 123388
rect 59675 122092 59741 122093
rect 59675 122028 59676 122092
rect 59740 122028 59741 122092
rect 59675 122027 59741 122028
rect 59307 120188 59373 120189
rect 59307 120124 59308 120188
rect 59372 120124 59373 120188
rect 59307 120123 59373 120124
rect 59310 111893 59370 120123
rect 59307 111892 59373 111893
rect 59307 111828 59308 111892
rect 59372 111828 59373 111892
rect 59307 111827 59373 111828
rect 59307 100060 59373 100061
rect 59307 99996 59308 100060
rect 59372 99996 59373 100060
rect 59307 99995 59373 99996
rect 59123 30836 59189 30837
rect 59123 30772 59124 30836
rect 59188 30772 59189 30836
rect 59123 30771 59189 30772
rect 59310 29885 59370 99995
rect 59307 29884 59373 29885
rect 59307 29820 59308 29884
rect 59372 29820 59373 29884
rect 59307 29819 59373 29820
rect 59862 28933 59922 123387
rect 60598 122850 60658 137970
rect 60046 122790 60658 122850
rect 59859 28932 59925 28933
rect 59859 28868 59860 28932
rect 59924 28868 59925 28932
rect 59859 28867 59925 28868
rect 58755 28252 58821 28253
rect 58755 28188 58756 28252
rect 58820 28188 58821 28252
rect 58755 28187 58821 28188
rect 60046 25669 60106 122790
rect 79568 115954 79888 115986
rect 79568 115718 79610 115954
rect 79846 115718 79888 115954
rect 79568 115634 79888 115718
rect 79568 115398 79610 115634
rect 79846 115398 79888 115634
rect 79568 115366 79888 115398
rect 110288 115954 110608 115986
rect 110288 115718 110330 115954
rect 110566 115718 110608 115954
rect 110288 115634 110608 115718
rect 110288 115398 110330 115634
rect 110566 115398 110608 115634
rect 110288 115366 110608 115398
rect 141008 115954 141328 115986
rect 141008 115718 141050 115954
rect 141286 115718 141328 115954
rect 141008 115634 141328 115718
rect 141008 115398 141050 115634
rect 141286 115398 141328 115634
rect 141008 115366 141328 115398
rect 171728 115954 172048 115986
rect 171728 115718 171770 115954
rect 172006 115718 172048 115954
rect 171728 115634 172048 115718
rect 171728 115398 171770 115634
rect 172006 115398 172048 115634
rect 171728 115366 172048 115398
rect 202448 115954 202768 115986
rect 202448 115718 202490 115954
rect 202726 115718 202768 115954
rect 202448 115634 202768 115718
rect 202448 115398 202490 115634
rect 202726 115398 202768 115634
rect 202448 115366 202768 115398
rect 233168 115954 233488 115986
rect 233168 115718 233210 115954
rect 233446 115718 233488 115954
rect 233168 115634 233488 115718
rect 233168 115398 233210 115634
rect 233446 115398 233488 115634
rect 233168 115366 233488 115398
rect 263888 115954 264208 115986
rect 263888 115718 263930 115954
rect 264166 115718 264208 115954
rect 263888 115634 264208 115718
rect 263888 115398 263930 115634
rect 264166 115398 264208 115634
rect 263888 115366 264208 115398
rect 294608 115954 294928 115986
rect 294608 115718 294650 115954
rect 294886 115718 294928 115954
rect 294608 115634 294928 115718
rect 294608 115398 294650 115634
rect 294886 115398 294928 115634
rect 294608 115366 294928 115398
rect 325328 115954 325648 115986
rect 325328 115718 325370 115954
rect 325606 115718 325648 115954
rect 325328 115634 325648 115718
rect 325328 115398 325370 115634
rect 325606 115398 325648 115634
rect 325328 115366 325648 115398
rect 356048 115954 356368 115986
rect 356048 115718 356090 115954
rect 356326 115718 356368 115954
rect 356048 115634 356368 115718
rect 356048 115398 356090 115634
rect 356326 115398 356368 115634
rect 356048 115366 356368 115398
rect 386768 115954 387088 115986
rect 386768 115718 386810 115954
rect 387046 115718 387088 115954
rect 386768 115634 387088 115718
rect 386768 115398 386810 115634
rect 387046 115398 387088 115634
rect 386768 115366 387088 115398
rect 417488 115954 417808 115986
rect 417488 115718 417530 115954
rect 417766 115718 417808 115954
rect 417488 115634 417808 115718
rect 417488 115398 417530 115634
rect 417766 115398 417808 115634
rect 417488 115366 417808 115398
rect 448208 115954 448528 115986
rect 448208 115718 448250 115954
rect 448486 115718 448528 115954
rect 448208 115634 448528 115718
rect 448208 115398 448250 115634
rect 448486 115398 448528 115634
rect 448208 115366 448528 115398
rect 478928 115954 479248 115986
rect 478928 115718 478970 115954
rect 479206 115718 479248 115954
rect 478928 115634 479248 115718
rect 478928 115398 478970 115634
rect 479206 115398 479248 115634
rect 478928 115366 479248 115398
rect 509648 115954 509968 115986
rect 509648 115718 509690 115954
rect 509926 115718 509968 115954
rect 509648 115634 509968 115718
rect 509648 115398 509690 115634
rect 509926 115398 509968 115634
rect 509648 115366 509968 115398
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 248528 111454 248848 111486
rect 248528 111218 248570 111454
rect 248806 111218 248848 111454
rect 248528 111134 248848 111218
rect 248528 110898 248570 111134
rect 248806 110898 248848 111134
rect 248528 110866 248848 110898
rect 279248 111454 279568 111486
rect 279248 111218 279290 111454
rect 279526 111218 279568 111454
rect 279248 111134 279568 111218
rect 279248 110898 279290 111134
rect 279526 110898 279568 111134
rect 279248 110866 279568 110898
rect 309968 111454 310288 111486
rect 309968 111218 310010 111454
rect 310246 111218 310288 111454
rect 309968 111134 310288 111218
rect 309968 110898 310010 111134
rect 310246 110898 310288 111134
rect 309968 110866 310288 110898
rect 340688 111454 341008 111486
rect 340688 111218 340730 111454
rect 340966 111218 341008 111454
rect 340688 111134 341008 111218
rect 340688 110898 340730 111134
rect 340966 110898 341008 111134
rect 340688 110866 341008 110898
rect 371408 111454 371728 111486
rect 371408 111218 371450 111454
rect 371686 111218 371728 111454
rect 371408 111134 371728 111218
rect 371408 110898 371450 111134
rect 371686 110898 371728 111134
rect 371408 110866 371728 110898
rect 402128 111454 402448 111486
rect 402128 111218 402170 111454
rect 402406 111218 402448 111454
rect 402128 111134 402448 111218
rect 402128 110898 402170 111134
rect 402406 110898 402448 111134
rect 402128 110866 402448 110898
rect 432848 111454 433168 111486
rect 432848 111218 432890 111454
rect 433126 111218 433168 111454
rect 432848 111134 433168 111218
rect 432848 110898 432890 111134
rect 433126 110898 433168 111134
rect 432848 110866 433168 110898
rect 463568 111454 463888 111486
rect 463568 111218 463610 111454
rect 463846 111218 463888 111454
rect 463568 111134 463888 111218
rect 463568 110898 463610 111134
rect 463846 110898 463888 111134
rect 463568 110866 463888 110898
rect 494288 111454 494608 111486
rect 494288 111218 494330 111454
rect 494566 111218 494608 111454
rect 494288 111134 494608 111218
rect 494288 110898 494330 111134
rect 494566 110898 494608 111134
rect 494288 110866 494608 110898
rect 525008 111454 525328 111486
rect 525008 111218 525050 111454
rect 525286 111218 525328 111454
rect 525008 111134 525328 111218
rect 525008 110898 525050 111134
rect 525286 110898 525328 111134
rect 525008 110866 525328 110898
rect 79568 79954 79888 79986
rect 79568 79718 79610 79954
rect 79846 79718 79888 79954
rect 79568 79634 79888 79718
rect 79568 79398 79610 79634
rect 79846 79398 79888 79634
rect 79568 79366 79888 79398
rect 110288 79954 110608 79986
rect 110288 79718 110330 79954
rect 110566 79718 110608 79954
rect 110288 79634 110608 79718
rect 110288 79398 110330 79634
rect 110566 79398 110608 79634
rect 110288 79366 110608 79398
rect 141008 79954 141328 79986
rect 141008 79718 141050 79954
rect 141286 79718 141328 79954
rect 141008 79634 141328 79718
rect 141008 79398 141050 79634
rect 141286 79398 141328 79634
rect 141008 79366 141328 79398
rect 171728 79954 172048 79986
rect 171728 79718 171770 79954
rect 172006 79718 172048 79954
rect 171728 79634 172048 79718
rect 171728 79398 171770 79634
rect 172006 79398 172048 79634
rect 171728 79366 172048 79398
rect 202448 79954 202768 79986
rect 202448 79718 202490 79954
rect 202726 79718 202768 79954
rect 202448 79634 202768 79718
rect 202448 79398 202490 79634
rect 202726 79398 202768 79634
rect 202448 79366 202768 79398
rect 233168 79954 233488 79986
rect 233168 79718 233210 79954
rect 233446 79718 233488 79954
rect 233168 79634 233488 79718
rect 233168 79398 233210 79634
rect 233446 79398 233488 79634
rect 233168 79366 233488 79398
rect 263888 79954 264208 79986
rect 263888 79718 263930 79954
rect 264166 79718 264208 79954
rect 263888 79634 264208 79718
rect 263888 79398 263930 79634
rect 264166 79398 264208 79634
rect 263888 79366 264208 79398
rect 294608 79954 294928 79986
rect 294608 79718 294650 79954
rect 294886 79718 294928 79954
rect 294608 79634 294928 79718
rect 294608 79398 294650 79634
rect 294886 79398 294928 79634
rect 294608 79366 294928 79398
rect 325328 79954 325648 79986
rect 325328 79718 325370 79954
rect 325606 79718 325648 79954
rect 325328 79634 325648 79718
rect 325328 79398 325370 79634
rect 325606 79398 325648 79634
rect 325328 79366 325648 79398
rect 356048 79954 356368 79986
rect 356048 79718 356090 79954
rect 356326 79718 356368 79954
rect 356048 79634 356368 79718
rect 356048 79398 356090 79634
rect 356326 79398 356368 79634
rect 356048 79366 356368 79398
rect 386768 79954 387088 79986
rect 386768 79718 386810 79954
rect 387046 79718 387088 79954
rect 386768 79634 387088 79718
rect 386768 79398 386810 79634
rect 387046 79398 387088 79634
rect 386768 79366 387088 79398
rect 417488 79954 417808 79986
rect 417488 79718 417530 79954
rect 417766 79718 417808 79954
rect 417488 79634 417808 79718
rect 417488 79398 417530 79634
rect 417766 79398 417808 79634
rect 417488 79366 417808 79398
rect 448208 79954 448528 79986
rect 448208 79718 448250 79954
rect 448486 79718 448528 79954
rect 448208 79634 448528 79718
rect 448208 79398 448250 79634
rect 448486 79398 448528 79634
rect 448208 79366 448528 79398
rect 478928 79954 479248 79986
rect 478928 79718 478970 79954
rect 479206 79718 479248 79954
rect 478928 79634 479248 79718
rect 478928 79398 478970 79634
rect 479206 79398 479248 79634
rect 478928 79366 479248 79398
rect 509648 79954 509968 79986
rect 509648 79718 509690 79954
rect 509926 79718 509968 79954
rect 509648 79634 509968 79718
rect 509648 79398 509690 79634
rect 509926 79398 509968 79634
rect 509648 79366 509968 79398
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 248528 75454 248848 75486
rect 248528 75218 248570 75454
rect 248806 75218 248848 75454
rect 248528 75134 248848 75218
rect 248528 74898 248570 75134
rect 248806 74898 248848 75134
rect 248528 74866 248848 74898
rect 279248 75454 279568 75486
rect 279248 75218 279290 75454
rect 279526 75218 279568 75454
rect 279248 75134 279568 75218
rect 279248 74898 279290 75134
rect 279526 74898 279568 75134
rect 279248 74866 279568 74898
rect 309968 75454 310288 75486
rect 309968 75218 310010 75454
rect 310246 75218 310288 75454
rect 309968 75134 310288 75218
rect 309968 74898 310010 75134
rect 310246 74898 310288 75134
rect 309968 74866 310288 74898
rect 340688 75454 341008 75486
rect 340688 75218 340730 75454
rect 340966 75218 341008 75454
rect 340688 75134 341008 75218
rect 340688 74898 340730 75134
rect 340966 74898 341008 75134
rect 340688 74866 341008 74898
rect 371408 75454 371728 75486
rect 371408 75218 371450 75454
rect 371686 75218 371728 75454
rect 371408 75134 371728 75218
rect 371408 74898 371450 75134
rect 371686 74898 371728 75134
rect 371408 74866 371728 74898
rect 402128 75454 402448 75486
rect 402128 75218 402170 75454
rect 402406 75218 402448 75454
rect 402128 75134 402448 75218
rect 402128 74898 402170 75134
rect 402406 74898 402448 75134
rect 402128 74866 402448 74898
rect 432848 75454 433168 75486
rect 432848 75218 432890 75454
rect 433126 75218 433168 75454
rect 432848 75134 433168 75218
rect 432848 74898 432890 75134
rect 433126 74898 433168 75134
rect 432848 74866 433168 74898
rect 463568 75454 463888 75486
rect 463568 75218 463610 75454
rect 463846 75218 463888 75454
rect 463568 75134 463888 75218
rect 463568 74898 463610 75134
rect 463846 74898 463888 75134
rect 463568 74866 463888 74898
rect 494288 75454 494608 75486
rect 494288 75218 494330 75454
rect 494566 75218 494608 75454
rect 494288 75134 494608 75218
rect 494288 74898 494330 75134
rect 494566 74898 494608 75134
rect 494288 74866 494608 74898
rect 525008 75454 525328 75486
rect 525008 75218 525050 75454
rect 525286 75218 525328 75454
rect 525008 75134 525328 75218
rect 525008 74898 525050 75134
rect 525286 74898 525328 75134
rect 525008 74866 525328 74898
rect 79568 43954 79888 43986
rect 79568 43718 79610 43954
rect 79846 43718 79888 43954
rect 79568 43634 79888 43718
rect 79568 43398 79610 43634
rect 79846 43398 79888 43634
rect 79568 43366 79888 43398
rect 110288 43954 110608 43986
rect 110288 43718 110330 43954
rect 110566 43718 110608 43954
rect 110288 43634 110608 43718
rect 110288 43398 110330 43634
rect 110566 43398 110608 43634
rect 110288 43366 110608 43398
rect 141008 43954 141328 43986
rect 141008 43718 141050 43954
rect 141286 43718 141328 43954
rect 141008 43634 141328 43718
rect 141008 43398 141050 43634
rect 141286 43398 141328 43634
rect 141008 43366 141328 43398
rect 171728 43954 172048 43986
rect 171728 43718 171770 43954
rect 172006 43718 172048 43954
rect 171728 43634 172048 43718
rect 171728 43398 171770 43634
rect 172006 43398 172048 43634
rect 171728 43366 172048 43398
rect 202448 43954 202768 43986
rect 202448 43718 202490 43954
rect 202726 43718 202768 43954
rect 202448 43634 202768 43718
rect 202448 43398 202490 43634
rect 202726 43398 202768 43634
rect 202448 43366 202768 43398
rect 233168 43954 233488 43986
rect 233168 43718 233210 43954
rect 233446 43718 233488 43954
rect 233168 43634 233488 43718
rect 233168 43398 233210 43634
rect 233446 43398 233488 43634
rect 233168 43366 233488 43398
rect 263888 43954 264208 43986
rect 263888 43718 263930 43954
rect 264166 43718 264208 43954
rect 263888 43634 264208 43718
rect 263888 43398 263930 43634
rect 264166 43398 264208 43634
rect 263888 43366 264208 43398
rect 294608 43954 294928 43986
rect 294608 43718 294650 43954
rect 294886 43718 294928 43954
rect 294608 43634 294928 43718
rect 294608 43398 294650 43634
rect 294886 43398 294928 43634
rect 294608 43366 294928 43398
rect 325328 43954 325648 43986
rect 325328 43718 325370 43954
rect 325606 43718 325648 43954
rect 325328 43634 325648 43718
rect 325328 43398 325370 43634
rect 325606 43398 325648 43634
rect 325328 43366 325648 43398
rect 356048 43954 356368 43986
rect 356048 43718 356090 43954
rect 356326 43718 356368 43954
rect 356048 43634 356368 43718
rect 356048 43398 356090 43634
rect 356326 43398 356368 43634
rect 356048 43366 356368 43398
rect 386768 43954 387088 43986
rect 386768 43718 386810 43954
rect 387046 43718 387088 43954
rect 386768 43634 387088 43718
rect 386768 43398 386810 43634
rect 387046 43398 387088 43634
rect 386768 43366 387088 43398
rect 417488 43954 417808 43986
rect 417488 43718 417530 43954
rect 417766 43718 417808 43954
rect 417488 43634 417808 43718
rect 417488 43398 417530 43634
rect 417766 43398 417808 43634
rect 417488 43366 417808 43398
rect 448208 43954 448528 43986
rect 448208 43718 448250 43954
rect 448486 43718 448528 43954
rect 448208 43634 448528 43718
rect 448208 43398 448250 43634
rect 448486 43398 448528 43634
rect 448208 43366 448528 43398
rect 478928 43954 479248 43986
rect 478928 43718 478970 43954
rect 479206 43718 479248 43954
rect 478928 43634 479248 43718
rect 478928 43398 478970 43634
rect 479206 43398 479248 43634
rect 478928 43366 479248 43398
rect 509648 43954 509968 43986
rect 509648 43718 509690 43954
rect 509926 43718 509968 43954
rect 509648 43634 509968 43718
rect 509648 43398 509690 43634
rect 509926 43398 509968 43634
rect 509648 43366 509968 43398
rect 64208 39454 64528 39486
rect 64208 39218 64250 39454
rect 64486 39218 64528 39454
rect 64208 39134 64528 39218
rect 64208 38898 64250 39134
rect 64486 38898 64528 39134
rect 64208 38866 64528 38898
rect 94928 39454 95248 39486
rect 94928 39218 94970 39454
rect 95206 39218 95248 39454
rect 94928 39134 95248 39218
rect 94928 38898 94970 39134
rect 95206 38898 95248 39134
rect 94928 38866 95248 38898
rect 125648 39454 125968 39486
rect 125648 39218 125690 39454
rect 125926 39218 125968 39454
rect 125648 39134 125968 39218
rect 125648 38898 125690 39134
rect 125926 38898 125968 39134
rect 125648 38866 125968 38898
rect 156368 39454 156688 39486
rect 156368 39218 156410 39454
rect 156646 39218 156688 39454
rect 156368 39134 156688 39218
rect 156368 38898 156410 39134
rect 156646 38898 156688 39134
rect 156368 38866 156688 38898
rect 187088 39454 187408 39486
rect 187088 39218 187130 39454
rect 187366 39218 187408 39454
rect 187088 39134 187408 39218
rect 187088 38898 187130 39134
rect 187366 38898 187408 39134
rect 187088 38866 187408 38898
rect 217808 39454 218128 39486
rect 217808 39218 217850 39454
rect 218086 39218 218128 39454
rect 217808 39134 218128 39218
rect 217808 38898 217850 39134
rect 218086 38898 218128 39134
rect 217808 38866 218128 38898
rect 248528 39454 248848 39486
rect 248528 39218 248570 39454
rect 248806 39218 248848 39454
rect 248528 39134 248848 39218
rect 248528 38898 248570 39134
rect 248806 38898 248848 39134
rect 248528 38866 248848 38898
rect 279248 39454 279568 39486
rect 279248 39218 279290 39454
rect 279526 39218 279568 39454
rect 279248 39134 279568 39218
rect 279248 38898 279290 39134
rect 279526 38898 279568 39134
rect 279248 38866 279568 38898
rect 309968 39454 310288 39486
rect 309968 39218 310010 39454
rect 310246 39218 310288 39454
rect 309968 39134 310288 39218
rect 309968 38898 310010 39134
rect 310246 38898 310288 39134
rect 309968 38866 310288 38898
rect 340688 39454 341008 39486
rect 340688 39218 340730 39454
rect 340966 39218 341008 39454
rect 340688 39134 341008 39218
rect 340688 38898 340730 39134
rect 340966 38898 341008 39134
rect 340688 38866 341008 38898
rect 371408 39454 371728 39486
rect 371408 39218 371450 39454
rect 371686 39218 371728 39454
rect 371408 39134 371728 39218
rect 371408 38898 371450 39134
rect 371686 38898 371728 39134
rect 371408 38866 371728 38898
rect 402128 39454 402448 39486
rect 402128 39218 402170 39454
rect 402406 39218 402448 39454
rect 402128 39134 402448 39218
rect 402128 38898 402170 39134
rect 402406 38898 402448 39134
rect 402128 38866 402448 38898
rect 432848 39454 433168 39486
rect 432848 39218 432890 39454
rect 433126 39218 433168 39454
rect 432848 39134 433168 39218
rect 432848 38898 432890 39134
rect 433126 38898 433168 39134
rect 432848 38866 433168 38898
rect 463568 39454 463888 39486
rect 463568 39218 463610 39454
rect 463846 39218 463888 39454
rect 463568 39134 463888 39218
rect 463568 38898 463610 39134
rect 463846 38898 463888 39134
rect 463568 38866 463888 38898
rect 494288 39454 494608 39486
rect 494288 39218 494330 39454
rect 494566 39218 494608 39454
rect 494288 39134 494608 39218
rect 494288 38898 494330 39134
rect 494566 38898 494608 39134
rect 494288 38866 494608 38898
rect 525008 39454 525328 39486
rect 525008 39218 525050 39454
rect 525286 39218 525328 39454
rect 525008 39134 525328 39218
rect 525008 38898 525050 39134
rect 525286 38898 525328 39134
rect 525008 38866 525328 38898
rect 539550 35325 539610 186899
rect 539731 180028 539797 180029
rect 539731 179964 539732 180028
rect 539796 179964 539797 180028
rect 539731 179963 539797 179964
rect 539734 46885 539794 179963
rect 539915 156772 539981 156773
rect 539915 156708 539916 156772
rect 539980 156708 539981 156772
rect 539915 156707 539981 156708
rect 539731 46884 539797 46885
rect 539731 46820 539732 46884
rect 539796 46820 539797 46884
rect 539731 46819 539797 46820
rect 539918 38589 539978 156707
rect 540099 150516 540165 150517
rect 540099 150452 540100 150516
rect 540164 150452 540165 150516
rect 540099 150451 540165 150452
rect 540102 148613 540162 150451
rect 540099 148612 540165 148613
rect 540099 148548 540100 148612
rect 540164 148548 540165 148612
rect 540099 148547 540165 148548
rect 540286 146981 540346 235451
rect 541571 235380 541637 235381
rect 541571 235316 541572 235380
rect 541636 235316 541637 235380
rect 541571 235315 541637 235316
rect 541019 177308 541085 177309
rect 541019 177244 541020 177308
rect 541084 177244 541085 177308
rect 541019 177243 541085 177244
rect 540283 146980 540349 146981
rect 540283 146916 540284 146980
rect 540348 146916 540349 146980
rect 540283 146915 540349 146916
rect 540835 144804 540901 144805
rect 540835 144740 540836 144804
rect 540900 144740 540901 144804
rect 540835 144739 540901 144740
rect 540651 129708 540717 129709
rect 540651 129644 540652 129708
rect 540716 129644 540717 129708
rect 540651 129643 540717 129644
rect 540654 110261 540714 129643
rect 540838 126309 540898 144739
rect 540835 126308 540901 126309
rect 540835 126244 540836 126308
rect 540900 126244 540901 126308
rect 540835 126243 540901 126244
rect 540651 110260 540717 110261
rect 540651 110196 540652 110260
rect 540716 110196 540717 110260
rect 540651 110195 540717 110196
rect 540099 95164 540165 95165
rect 540099 95100 540100 95164
rect 540164 95100 540165 95164
rect 540099 95099 540165 95100
rect 539915 38588 539981 38589
rect 539915 38524 539916 38588
rect 539980 38524 539981 38588
rect 539915 38523 539981 38524
rect 539547 35324 539613 35325
rect 539547 35260 539548 35324
rect 539612 35260 539613 35324
rect 539547 35259 539613 35260
rect 539363 31108 539429 31109
rect 539363 31044 539364 31108
rect 539428 31044 539429 31108
rect 539363 31043 539429 31044
rect 60294 25954 60914 28000
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60043 25668 60109 25669
rect 60043 25604 60044 25668
rect 60108 25604 60109 25668
rect 60043 25603 60109 25604
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 58571 19004 58637 19005
rect 58571 18940 58572 19004
rect 58636 18940 58637 19004
rect 58571 18939 58637 18940
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 73794 3454 74414 28000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 7954 78914 28000
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 12454 83414 28000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 16954 87914 28000
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 21454 92414 28000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 25954 96914 28000
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 109794 3454 110414 28000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 7954 114914 28000
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 28000
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 16954 123914 28000
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 21454 128414 28000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 25954 132914 28000
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 145794 3454 146414 28000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 28000
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 28000
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 28000
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 28000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 28000
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 181794 3454 182414 28000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 7954 186914 28000
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 12454 191414 28000
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 28000
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 28000
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7954 222914 28000
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 12454 227414 28000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 16954 231914 28000
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 25954 240914 28000
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 7954 258914 28000
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 12454 263414 28000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 28000
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 25954 276914 28000
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 289794 3454 290414 28000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 28000
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 28000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 28000
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 28000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 25954 312914 28000
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 325794 3454 326414 28000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 7954 330914 28000
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 12454 335414 28000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 28000
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 28000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 25954 348914 28000
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 361794 3454 362414 28000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 7954 366914 28000
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 12454 371414 28000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 16954 375914 28000
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 21454 380414 28000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 25954 384914 28000
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 7954 402914 28000
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 12454 407414 28000
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 16954 411914 28000
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 21454 416414 28000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 25954 420914 28000
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 433794 3454 434414 28000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 7954 438914 28000
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 12454 443414 28000
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 16954 447914 28000
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 25954 456914 28000
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 7954 474914 28000
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 12454 479414 28000
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 16954 483914 28000
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 25954 492914 28000
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 7954 510914 28000
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 12454 515414 28000
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 16954 519914 28000
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 21454 524414 28000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 25954 528914 28000
rect 539366 26250 539426 31043
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 538814 26190 539426 26250
rect 538814 25397 538874 26190
rect 538811 25396 538877 25397
rect 538811 25332 538812 25396
rect 538876 25332 538877 25396
rect 538811 25331 538877 25332
rect 540102 13701 540162 95099
rect 541022 70957 541082 177243
rect 541203 163436 541269 163437
rect 541203 163372 541204 163436
rect 541268 163372 541269 163436
rect 541203 163371 541269 163372
rect 541206 115973 541266 163371
rect 541387 151740 541453 151741
rect 541387 151676 541388 151740
rect 541452 151676 541453 151740
rect 541387 151675 541453 151676
rect 541390 133245 541450 151675
rect 541387 133244 541453 133245
rect 541387 133180 541388 133244
rect 541452 133180 541453 133244
rect 541387 133179 541453 133180
rect 541574 130525 541634 235315
rect 541794 219454 542414 238000
rect 544331 235652 544397 235653
rect 544331 235588 544332 235652
rect 544396 235588 544397 235652
rect 544331 235587 544397 235588
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 542675 210356 542741 210357
rect 542675 210292 542676 210356
rect 542740 210292 542741 210356
rect 542675 210291 542741 210292
rect 542678 200130 542738 210291
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 152000 542414 182898
rect 542494 200070 542738 200130
rect 541939 131340 542005 131341
rect 541939 131276 541940 131340
rect 542004 131276 542005 131340
rect 541939 131275 542005 131276
rect 541571 130524 541637 130525
rect 541571 130460 541572 130524
rect 541636 130460 541637 130524
rect 541571 130459 541637 130460
rect 541203 115972 541269 115973
rect 541203 115908 541204 115972
rect 541268 115908 541269 115972
rect 541203 115907 541269 115908
rect 541755 115972 541821 115973
rect 541755 115908 541756 115972
rect 541820 115908 541821 115972
rect 541755 115907 541821 115908
rect 541203 110260 541269 110261
rect 541203 110196 541204 110260
rect 541268 110196 541269 110260
rect 541203 110195 541269 110196
rect 541206 99517 541266 110195
rect 541758 107541 541818 115907
rect 541942 110669 542002 131275
rect 542123 130388 542189 130389
rect 542123 130324 542124 130388
rect 542188 130324 542189 130388
rect 542123 130323 542189 130324
rect 541939 110668 542005 110669
rect 541939 110604 541940 110668
rect 542004 110604 542005 110668
rect 541939 110603 542005 110604
rect 541755 107540 541821 107541
rect 541755 107476 541756 107540
rect 541820 107476 541821 107540
rect 541755 107475 541821 107476
rect 541571 105500 541637 105501
rect 541571 105436 541572 105500
rect 541636 105436 541637 105500
rect 541571 105435 541637 105436
rect 541387 102372 541453 102373
rect 541387 102308 541388 102372
rect 541452 102308 541453 102372
rect 541387 102307 541453 102308
rect 541203 99516 541269 99517
rect 541203 99452 541204 99516
rect 541268 99452 541269 99516
rect 541203 99451 541269 99452
rect 541203 82924 541269 82925
rect 541203 82860 541204 82924
rect 541268 82860 541269 82924
rect 541203 82859 541269 82860
rect 541019 70956 541085 70957
rect 541019 70892 541020 70956
rect 541084 70892 541085 70956
rect 541019 70891 541085 70892
rect 540283 30972 540349 30973
rect 540283 30908 540284 30972
rect 540348 30908 540349 30972
rect 540283 30907 540349 30908
rect 540286 21997 540346 30907
rect 541206 28797 541266 82859
rect 541203 28796 541269 28797
rect 541203 28732 541204 28796
rect 541268 28732 541269 28796
rect 541203 28731 541269 28732
rect 540283 21996 540349 21997
rect 540283 21932 540284 21996
rect 540348 21932 540349 21996
rect 540283 21931 540349 21932
rect 541390 15061 541450 102307
rect 541387 15060 541453 15061
rect 541387 14996 541388 15060
rect 541452 14996 541453 15060
rect 541387 14995 541453 14996
rect 540099 13700 540165 13701
rect 540099 13636 540100 13700
rect 540164 13636 540165 13700
rect 540099 13635 540165 13636
rect 541574 3229 541634 105435
rect 542126 102237 542186 130323
rect 542494 113117 542554 200070
rect 542675 174724 542741 174725
rect 542675 174660 542676 174724
rect 542740 174660 542741 174724
rect 542675 174659 542741 174660
rect 542491 113116 542557 113117
rect 542491 113052 542492 113116
rect 542556 113052 542557 113116
rect 542491 113051 542557 113052
rect 542678 108490 542738 174659
rect 543963 171732 544029 171733
rect 543963 171668 543964 171732
rect 544028 171668 544029 171732
rect 543963 171667 544029 171668
rect 543779 159628 543845 159629
rect 543779 159564 543780 159628
rect 543844 159564 543845 159628
rect 543779 159563 543845 159564
rect 543411 155684 543477 155685
rect 543411 155620 543412 155684
rect 543476 155620 543477 155684
rect 543411 155619 543477 155620
rect 542859 154188 542925 154189
rect 542859 154124 542860 154188
rect 542924 154124 542925 154188
rect 542859 154123 542925 154124
rect 542862 146165 542922 154123
rect 542859 146164 542925 146165
rect 542859 146100 542860 146164
rect 542924 146100 542925 146164
rect 542859 146099 542925 146100
rect 543043 128484 543109 128485
rect 543043 128420 543044 128484
rect 543108 128420 543109 128484
rect 543043 128419 543109 128420
rect 542859 110940 542925 110941
rect 542859 110876 542860 110940
rect 542924 110876 542925 110940
rect 542859 110875 542925 110876
rect 542310 108430 542738 108490
rect 542123 102236 542189 102237
rect 542123 102172 542124 102236
rect 542188 102172 542189 102236
rect 542123 102171 542189 102172
rect 542310 87957 542370 108430
rect 542491 107540 542557 107541
rect 542491 107476 542492 107540
rect 542556 107476 542557 107540
rect 542491 107475 542557 107476
rect 542307 87956 542373 87957
rect 542307 87892 542308 87956
rect 542372 87892 542373 87956
rect 542307 87891 542373 87892
rect 542494 35910 542554 107475
rect 542494 35850 542738 35910
rect 541794 3454 542414 28000
rect 542678 17645 542738 35850
rect 542675 17644 542741 17645
rect 542675 17580 542676 17644
rect 542740 17580 542741 17644
rect 542675 17579 542741 17580
rect 542862 17101 542922 110875
rect 543046 102373 543106 128419
rect 543414 104277 543474 155619
rect 543411 104276 543477 104277
rect 543411 104212 543412 104276
rect 543476 104212 543477 104276
rect 543411 104211 543477 104212
rect 543043 102372 543109 102373
rect 543043 102308 543044 102372
rect 543108 102308 543109 102372
rect 543043 102307 543109 102308
rect 543227 89044 543293 89045
rect 543227 88980 543228 89044
rect 543292 88980 543293 89044
rect 543227 88979 543293 88980
rect 543043 86188 543109 86189
rect 543043 86124 543044 86188
rect 543108 86124 543109 86188
rect 543043 86123 543109 86124
rect 542859 17100 542925 17101
rect 542859 17036 542860 17100
rect 542924 17036 542925 17100
rect 542859 17035 542925 17036
rect 543046 15197 543106 86123
rect 543230 20229 543290 88979
rect 543782 29069 543842 159563
rect 543966 68917 544026 171667
rect 544147 158268 544213 158269
rect 544147 158204 544148 158268
rect 544212 158204 544213 158268
rect 544147 158203 544213 158204
rect 544150 146301 544210 158203
rect 544147 146300 544213 146301
rect 544147 146236 544148 146300
rect 544212 146236 544213 146300
rect 544147 146235 544213 146236
rect 544334 139637 544394 235587
rect 546294 223954 546914 238000
rect 547091 236740 547157 236741
rect 547091 236676 547092 236740
rect 547156 236676 547157 236740
rect 547091 236675 547157 236676
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 545435 166564 545501 166565
rect 545435 166500 545436 166564
rect 545500 166500 545501 166564
rect 545435 166499 545501 166500
rect 545251 155412 545317 155413
rect 545251 155348 545252 155412
rect 545316 155348 545317 155412
rect 545251 155347 545317 155348
rect 545067 153916 545133 153917
rect 545067 153852 545068 153916
rect 545132 153852 545133 153916
rect 545067 153851 545133 153852
rect 544699 146164 544765 146165
rect 544699 146100 544700 146164
rect 544764 146100 544765 146164
rect 544699 146099 544765 146100
rect 544331 139636 544397 139637
rect 544331 139572 544332 139636
rect 544396 139572 544397 139636
rect 544331 139571 544397 139572
rect 544515 139500 544581 139501
rect 544515 139436 544516 139500
rect 544580 139436 544581 139500
rect 544515 139435 544581 139436
rect 544518 136645 544578 139435
rect 544702 138141 544762 146099
rect 544699 138140 544765 138141
rect 544699 138076 544700 138140
rect 544764 138076 544765 138140
rect 544699 138075 544765 138076
rect 544699 138004 544765 138005
rect 544699 137940 544700 138004
rect 544764 137940 544765 138004
rect 544699 137939 544765 137940
rect 544331 136644 544397 136645
rect 544331 136580 544332 136644
rect 544396 136580 544397 136644
rect 544331 136579 544397 136580
rect 544515 136644 544581 136645
rect 544515 136580 544516 136644
rect 544580 136580 544581 136644
rect 544515 136579 544581 136580
rect 544334 127669 544394 136579
rect 544702 131341 544762 137939
rect 544699 131340 544765 131341
rect 544699 131276 544700 131340
rect 544764 131276 544765 131340
rect 544699 131275 544765 131276
rect 544515 131204 544581 131205
rect 544515 131140 544516 131204
rect 544580 131140 544581 131204
rect 544515 131139 544581 131140
rect 544147 127668 544213 127669
rect 544147 127604 544148 127668
rect 544212 127604 544213 127668
rect 544147 127603 544213 127604
rect 544331 127668 544397 127669
rect 544331 127604 544332 127668
rect 544396 127604 544397 127668
rect 544331 127603 544397 127604
rect 544150 118013 544210 127603
rect 544518 124133 544578 131139
rect 544515 124132 544581 124133
rect 544515 124068 544516 124132
rect 544580 124068 544581 124132
rect 544515 124067 544581 124068
rect 544331 123996 544397 123997
rect 544331 123932 544332 123996
rect 544396 123932 544397 123996
rect 544331 123931 544397 123932
rect 544147 118012 544213 118013
rect 544147 117948 544148 118012
rect 544212 117948 544213 118012
rect 544147 117947 544213 117948
rect 544147 110532 544213 110533
rect 544147 110468 544148 110532
rect 544212 110468 544213 110532
rect 544147 110467 544213 110468
rect 543963 68916 544029 68917
rect 543963 68852 543964 68916
rect 544028 68852 544029 68916
rect 543963 68851 544029 68852
rect 543779 29068 543845 29069
rect 543779 29004 543780 29068
rect 543844 29004 543845 29068
rect 543779 29003 543845 29004
rect 543227 20228 543293 20229
rect 543227 20164 543228 20228
rect 543292 20164 543293 20228
rect 543227 20163 543293 20164
rect 544150 16421 544210 110467
rect 544334 19141 544394 123931
rect 544515 117332 544581 117333
rect 544515 117268 544516 117332
rect 544580 117268 544581 117332
rect 544515 117267 544581 117268
rect 544518 114477 544578 117267
rect 544515 114476 544581 114477
rect 544515 114412 544516 114476
rect 544580 114412 544581 114476
rect 544515 114411 544581 114412
rect 545070 27029 545130 153851
rect 545254 29613 545314 155347
rect 545438 139501 545498 166499
rect 545803 159492 545869 159493
rect 545803 159428 545804 159492
rect 545868 159428 545869 159492
rect 545803 159427 545869 159428
rect 545619 139636 545685 139637
rect 545619 139572 545620 139636
rect 545684 139572 545685 139636
rect 545619 139571 545685 139572
rect 545435 139500 545501 139501
rect 545435 139436 545436 139500
rect 545500 139436 545501 139500
rect 545435 139435 545501 139436
rect 545435 127668 545501 127669
rect 545435 127604 545436 127668
rect 545500 127604 545501 127668
rect 545435 127603 545501 127604
rect 545251 29612 545317 29613
rect 545251 29548 545252 29612
rect 545316 29548 545317 29612
rect 545251 29547 545317 29548
rect 545067 27028 545133 27029
rect 545067 26964 545068 27028
rect 545132 26964 545133 27028
rect 545067 26963 545133 26964
rect 544331 19140 544397 19141
rect 544331 19076 544332 19140
rect 544396 19076 544397 19140
rect 544331 19075 544397 19076
rect 544147 16420 544213 16421
rect 544147 16356 544148 16420
rect 544212 16356 544213 16420
rect 544147 16355 544213 16356
rect 543043 15196 543109 15197
rect 543043 15132 543044 15196
rect 543108 15132 543109 15196
rect 543043 15131 543109 15132
rect 545438 13021 545498 127603
rect 545622 127125 545682 139571
rect 545619 127124 545685 127125
rect 545619 127060 545620 127124
rect 545684 127060 545685 127124
rect 545619 127059 545685 127060
rect 545619 126988 545685 126989
rect 545619 126924 545620 126988
rect 545684 126924 545685 126988
rect 545619 126923 545685 126924
rect 545622 26757 545682 126923
rect 545806 126853 545866 159427
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 545803 126852 545869 126853
rect 545803 126788 545804 126852
rect 545868 126788 545869 126852
rect 545803 126787 545869 126788
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 545619 26756 545685 26757
rect 545619 26692 545620 26756
rect 545684 26692 545685 26756
rect 545619 26691 545685 26692
rect 545435 13020 545501 13021
rect 545435 12956 545436 13020
rect 545500 12956 545501 13020
rect 545435 12955 545501 12956
rect 541571 3228 541637 3229
rect 541571 3164 541572 3228
rect 541636 3164 541637 3228
rect 541571 3163 541637 3164
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 7954 546914 43398
rect 547094 22677 547154 236675
rect 548011 235788 548077 235789
rect 548011 235724 548012 235788
rect 548076 235724 548077 235788
rect 548011 235723 548077 235724
rect 547459 160852 547525 160853
rect 547459 160788 547460 160852
rect 547524 160788 547525 160852
rect 547459 160787 547525 160788
rect 547275 149972 547341 149973
rect 547275 149908 547276 149972
rect 547340 149908 547341 149972
rect 547275 149907 547341 149908
rect 547278 138685 547338 149907
rect 547275 138684 547341 138685
rect 547275 138620 547276 138684
rect 547340 138620 547341 138684
rect 547275 138619 547341 138620
rect 547275 138140 547341 138141
rect 547275 138076 547276 138140
rect 547340 138076 547341 138140
rect 547275 138075 547341 138076
rect 547278 132837 547338 138075
rect 547275 132836 547341 132837
rect 547275 132772 547276 132836
rect 547340 132772 547341 132836
rect 547275 132771 547341 132772
rect 547275 126852 547341 126853
rect 547275 126788 547276 126852
rect 547340 126788 547341 126852
rect 547275 126787 547341 126788
rect 547278 24853 547338 126787
rect 547462 114341 547522 160787
rect 547827 154324 547893 154325
rect 547827 154260 547828 154324
rect 547892 154260 547893 154324
rect 547827 154259 547893 154260
rect 547830 147690 547890 154259
rect 547646 147630 547890 147690
rect 547646 132970 547706 147630
rect 547646 132910 547890 132970
rect 547643 132836 547709 132837
rect 547643 132772 547644 132836
rect 547708 132772 547709 132836
rect 547643 132771 547709 132772
rect 547646 126989 547706 132771
rect 547830 130250 547890 132910
rect 548014 130389 548074 235723
rect 549483 234020 549549 234021
rect 549483 233956 549484 234020
rect 549548 233956 549549 234020
rect 549483 233955 549549 233956
rect 548195 161124 548261 161125
rect 548195 161060 548196 161124
rect 548260 161060 548261 161124
rect 548195 161059 548261 161060
rect 548198 132510 548258 161059
rect 549299 154052 549365 154053
rect 549299 153988 549300 154052
rect 549364 153988 549365 154052
rect 549299 153987 549365 153988
rect 548198 132450 548626 132510
rect 548011 130388 548077 130389
rect 548011 130324 548012 130388
rect 548076 130324 548077 130388
rect 548011 130323 548077 130324
rect 547830 130190 548074 130250
rect 547643 126988 547709 126989
rect 547643 126924 547644 126988
rect 547708 126924 547709 126988
rect 547643 126923 547709 126924
rect 548014 126850 548074 130190
rect 548379 129572 548445 129573
rect 548379 129508 548380 129572
rect 548444 129508 548445 129572
rect 548379 129507 548445 129508
rect 547646 126790 548074 126850
rect 547459 114340 547525 114341
rect 547459 114276 547460 114340
rect 547524 114276 547525 114340
rect 547459 114275 547525 114276
rect 547459 110668 547525 110669
rect 547459 110604 547460 110668
rect 547524 110604 547525 110668
rect 547459 110603 547525 110604
rect 547275 24852 547341 24853
rect 547275 24788 547276 24852
rect 547340 24788 547341 24852
rect 547275 24787 547341 24788
rect 547091 22676 547157 22677
rect 547091 22612 547092 22676
rect 547156 22612 547157 22676
rect 547091 22611 547157 22612
rect 547462 16557 547522 110603
rect 547646 29477 547706 126790
rect 548382 125490 548442 129507
rect 548014 125430 548442 125490
rect 547643 29476 547709 29477
rect 547643 29412 547644 29476
rect 547708 29412 547709 29476
rect 547643 29411 547709 29412
rect 547459 16556 547525 16557
rect 547459 16492 547460 16556
rect 547524 16492 547525 16556
rect 547459 16491 547525 16492
rect 548014 14925 548074 125430
rect 548566 122850 548626 132450
rect 548198 122790 548626 122850
rect 548198 84693 548258 122790
rect 548379 85644 548445 85645
rect 548379 85580 548380 85644
rect 548444 85580 548445 85644
rect 548379 85579 548445 85580
rect 548195 84692 548261 84693
rect 548195 84628 548196 84692
rect 548260 84628 548261 84692
rect 548195 84627 548261 84628
rect 548382 22949 548442 85579
rect 549302 27573 549362 153987
rect 549486 113253 549546 233955
rect 550222 191181 550282 440675
rect 550774 238770 550834 497115
rect 551507 441420 551573 441421
rect 551507 441356 551508 441420
rect 551572 441356 551573 441420
rect 551507 441355 551573 441356
rect 550590 238710 550834 238770
rect 550219 191180 550285 191181
rect 550219 191116 550220 191180
rect 550284 191116 550285 191180
rect 550219 191115 550285 191116
rect 549851 161260 549917 161261
rect 549851 161196 549852 161260
rect 549916 161196 549917 161260
rect 549851 161195 549917 161196
rect 549667 158540 549733 158541
rect 549667 158476 549668 158540
rect 549732 158476 549733 158540
rect 549667 158475 549733 158476
rect 549483 113252 549549 113253
rect 549483 113188 549484 113252
rect 549548 113188 549549 113252
rect 549483 113187 549549 113188
rect 549670 72317 549730 158475
rect 549854 83333 549914 161195
rect 549851 83332 549917 83333
rect 549851 83268 549852 83332
rect 549916 83268 549917 83332
rect 549851 83267 549917 83268
rect 549851 81564 549917 81565
rect 549851 81500 549852 81564
rect 549916 81500 549917 81564
rect 549851 81499 549917 81500
rect 549667 72316 549733 72317
rect 549667 72252 549668 72316
rect 549732 72252 549733 72316
rect 549667 72251 549733 72252
rect 549299 27572 549365 27573
rect 549299 27508 549300 27572
rect 549364 27508 549365 27572
rect 549299 27507 549365 27508
rect 548379 22948 548445 22949
rect 548379 22884 548380 22948
rect 548444 22884 548445 22948
rect 548379 22883 548445 22884
rect 548011 14924 548077 14925
rect 548011 14860 548012 14924
rect 548076 14860 548077 14924
rect 548011 14859 548077 14860
rect 549854 14517 549914 81499
rect 550590 16013 550650 238710
rect 550794 228454 551414 238000
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 551510 191045 551570 441355
rect 551507 191044 551573 191045
rect 551507 190980 551508 191044
rect 551572 190980 551573 191044
rect 551507 190979 551573 190980
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 551507 153780 551573 153781
rect 551507 153716 551508 153780
rect 551572 153716 551573 153780
rect 551507 153715 551573 153716
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550587 16012 550653 16013
rect 550587 15948 550588 16012
rect 550652 15948 550653 16012
rect 550587 15947 550653 15948
rect 549851 14516 549917 14517
rect 549851 14452 549852 14516
rect 549916 14452 549917 14516
rect 549851 14451 549917 14452
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 12454 551414 47898
rect 551510 41717 551570 153715
rect 551507 41716 551573 41717
rect 551507 41652 551508 41716
rect 551572 41652 551573 41716
rect 551507 41651 551573 41652
rect 552062 28253 552122 682619
rect 552246 673981 552306 685883
rect 552243 673980 552309 673981
rect 552243 673916 552244 673980
rect 552308 673916 552309 673980
rect 552243 673915 552309 673916
rect 555294 664954 555914 700398
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 560523 682548 560589 682549
rect 560523 682484 560524 682548
rect 560588 682484 560589 682548
rect 560523 682483 560589 682484
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 557579 668540 557645 668541
rect 557579 668476 557580 668540
rect 557644 668476 557645 668540
rect 557579 668475 557645 668476
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 556107 649500 556173 649501
rect 556107 649436 556108 649500
rect 556172 649436 556173 649500
rect 556107 649435 556173 649436
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 552243 614820 552309 614821
rect 552243 614756 552244 614820
rect 552308 614756 552309 614820
rect 552243 614755 552309 614756
rect 552246 188461 552306 614755
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 553347 566540 553413 566541
rect 553347 566476 553348 566540
rect 553412 566476 553413 566540
rect 553347 566475 553413 566476
rect 553350 524430 553410 566475
rect 553166 524370 553410 524430
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 553166 514770 553226 524370
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 553166 514710 553410 514770
rect 553350 466470 553410 514710
rect 554819 494460 554885 494461
rect 554819 494396 554820 494460
rect 554884 494396 554885 494460
rect 554819 494395 554885 494396
rect 553531 491740 553597 491741
rect 553531 491676 553532 491740
rect 553596 491676 553597 491740
rect 553531 491675 553597 491676
rect 553166 466410 553410 466470
rect 553166 456810 553226 466410
rect 553166 456750 553410 456810
rect 553350 418170 553410 456750
rect 553166 418110 553410 418170
rect 553166 408510 553226 418110
rect 553166 408450 553410 408510
rect 552243 188460 552309 188461
rect 552243 188396 552244 188460
rect 552308 188396 552309 188460
rect 552243 188395 552309 188396
rect 552243 160988 552309 160989
rect 552243 160924 552244 160988
rect 552308 160924 552309 160988
rect 552243 160923 552309 160924
rect 552246 30429 552306 160923
rect 552427 160716 552493 160717
rect 552427 160652 552428 160716
rect 552492 160652 552493 160716
rect 552427 160651 552493 160652
rect 552430 37365 552490 160651
rect 553350 157350 553410 408450
rect 552611 157316 552677 157317
rect 552611 157252 552612 157316
rect 552676 157252 552677 157316
rect 552611 157251 552677 157252
rect 553166 157290 553410 157350
rect 552614 51101 552674 157251
rect 553166 147690 553226 157290
rect 553166 147630 553410 147690
rect 552611 51100 552677 51101
rect 552611 51036 552612 51100
rect 552676 51036 552677 51100
rect 552611 51035 552677 51036
rect 552427 37364 552493 37365
rect 552427 37300 552428 37364
rect 552492 37300 552493 37364
rect 552427 37299 552493 37300
rect 552243 30428 552309 30429
rect 552243 30364 552244 30428
rect 552308 30364 552309 30428
rect 552243 30363 552309 30364
rect 552059 28252 552125 28253
rect 552059 28188 552060 28252
rect 552124 28188 552125 28252
rect 552059 28187 552125 28188
rect 553350 24173 553410 147630
rect 553347 24172 553413 24173
rect 553347 24108 553348 24172
rect 553412 24108 553413 24172
rect 553347 24107 553413 24108
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 553534 6221 553594 491675
rect 553715 315620 553781 315621
rect 553715 315556 553716 315620
rect 553780 315556 553781 315620
rect 553715 315555 553781 315556
rect 553718 18597 553778 315555
rect 553899 152556 553965 152557
rect 553899 152492 553900 152556
rect 553964 152492 553965 152556
rect 553899 152491 553965 152492
rect 553902 89045 553962 152491
rect 553899 89044 553965 89045
rect 553899 88980 553900 89044
rect 553964 88980 553965 89044
rect 553899 88979 553965 88980
rect 554822 19957 554882 494395
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555003 404700 555069 404701
rect 555003 404636 555004 404700
rect 555068 404636 555069 404700
rect 555003 404635 555069 404636
rect 555006 192541 555066 404635
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555003 192540 555069 192541
rect 555003 192476 555004 192540
rect 555068 192476 555069 192540
rect 555003 192475 555069 192476
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555003 151196 555069 151197
rect 555003 151132 555004 151196
rect 555068 151132 555069 151196
rect 555003 151131 555069 151132
rect 555006 30973 555066 151131
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555003 30972 555069 30973
rect 555003 30908 555004 30972
rect 555068 30908 555069 30972
rect 555003 30907 555069 30908
rect 554819 19956 554885 19957
rect 554819 19892 554820 19956
rect 554884 19892 554885 19956
rect 554819 19891 554885 19892
rect 553715 18596 553781 18597
rect 553715 18532 553716 18596
rect 553780 18532 553781 18596
rect 553715 18531 553781 18532
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 553531 6220 553597 6221
rect 553531 6156 553532 6220
rect 553596 6156 553597 6220
rect 553531 6155 553597 6156
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 -3226 555914 16398
rect 556110 7581 556170 649435
rect 556659 612100 556725 612101
rect 556659 612036 556660 612100
rect 556724 612036 556725 612100
rect 556659 612035 556725 612036
rect 556291 608020 556357 608021
rect 556291 607956 556292 608020
rect 556356 607956 556357 608020
rect 556291 607955 556357 607956
rect 556294 10437 556354 607955
rect 556475 599180 556541 599181
rect 556475 599116 556476 599180
rect 556540 599116 556541 599180
rect 556475 599115 556541 599116
rect 556478 17237 556538 599115
rect 556662 234701 556722 612035
rect 556843 235380 556909 235381
rect 556843 235316 556844 235380
rect 556908 235316 556909 235380
rect 556843 235315 556909 235316
rect 556659 234700 556725 234701
rect 556659 234636 556660 234700
rect 556724 234636 556725 234700
rect 556659 234635 556725 234636
rect 556846 219450 556906 235315
rect 556662 219390 556906 219450
rect 556662 24581 556722 219390
rect 556659 24580 556725 24581
rect 556659 24516 556660 24580
rect 556724 24516 556725 24580
rect 556659 24515 556725 24516
rect 557582 17373 557642 668475
rect 557763 633860 557829 633861
rect 557763 633796 557764 633860
rect 557828 633796 557829 633860
rect 557763 633795 557829 633796
rect 557579 17372 557645 17373
rect 557579 17308 557580 17372
rect 557644 17308 557645 17372
rect 557579 17307 557645 17308
rect 556475 17236 556541 17237
rect 556475 17172 556476 17236
rect 556540 17172 556541 17236
rect 556475 17171 556541 17172
rect 557766 11797 557826 633795
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 557947 630460 558013 630461
rect 557947 630396 557948 630460
rect 558012 630396 558013 630460
rect 557947 630395 558013 630396
rect 557763 11796 557829 11797
rect 557763 11732 557764 11796
rect 557828 11732 557829 11796
rect 557763 11731 557829 11732
rect 556291 10436 556357 10437
rect 556291 10372 556292 10436
rect 556356 10372 556357 10436
rect 556291 10371 556357 10372
rect 557950 7717 558010 630395
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 558867 591020 558933 591021
rect 558867 590956 558868 591020
rect 558932 590956 558933 591020
rect 558867 590955 558933 590956
rect 558131 556340 558197 556341
rect 558131 556276 558132 556340
rect 558196 556276 558197 556340
rect 558131 556275 558197 556276
rect 558134 18869 558194 556275
rect 558870 21181 558930 590955
rect 559051 574156 559117 574157
rect 559051 574092 559052 574156
rect 559116 574092 559117 574156
rect 559051 574091 559117 574092
rect 559054 167653 559114 574091
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559235 336700 559301 336701
rect 559235 336636 559236 336700
rect 559300 336636 559301 336700
rect 559235 336635 559301 336636
rect 559051 167652 559117 167653
rect 559051 167588 559052 167652
rect 559116 167588 559117 167652
rect 559051 167587 559117 167588
rect 559051 151332 559117 151333
rect 559051 151268 559052 151332
rect 559116 151268 559117 151332
rect 559051 151267 559117 151268
rect 558867 21180 558933 21181
rect 558867 21116 558868 21180
rect 558932 21116 558933 21180
rect 558867 21115 558933 21116
rect 559054 19005 559114 151267
rect 559051 19004 559117 19005
rect 559051 18940 559052 19004
rect 559116 18940 559117 19004
rect 559051 18939 559117 18940
rect 558131 18868 558197 18869
rect 558131 18804 558132 18868
rect 558196 18804 558197 18868
rect 558131 18803 558197 18804
rect 557947 7716 558013 7717
rect 557947 7652 557948 7716
rect 558012 7652 558013 7716
rect 557947 7651 558013 7652
rect 556107 7580 556173 7581
rect 556107 7516 556108 7580
rect 556172 7516 556173 7580
rect 556107 7515 556173 7516
rect 559238 4861 559298 336635
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 560526 28525 560586 682483
rect 561627 682412 561693 682413
rect 561627 682348 561628 682412
rect 561692 682348 561693 682412
rect 561627 682347 561693 682348
rect 560707 627060 560773 627061
rect 560707 626996 560708 627060
rect 560772 626996 560773 627060
rect 560707 626995 560773 626996
rect 560523 28524 560589 28525
rect 560523 28460 560524 28524
rect 560588 28460 560589 28524
rect 560523 28459 560589 28460
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559235 4860 559301 4861
rect 559235 4796 559236 4860
rect 559300 4796 559301 4860
rect 559235 4795 559301 4796
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 -4186 560414 20898
rect 560710 17645 560770 626995
rect 560891 531860 560957 531861
rect 560891 531796 560892 531860
rect 560956 531796 560957 531860
rect 560891 531795 560957 531796
rect 560707 17644 560773 17645
rect 560707 17580 560708 17644
rect 560772 17580 560773 17644
rect 560707 17579 560773 17580
rect 560894 11661 560954 531795
rect 561075 450260 561141 450261
rect 561075 450196 561076 450260
rect 561140 450196 561141 450260
rect 561075 450195 561141 450196
rect 561078 27437 561138 450195
rect 561075 27436 561141 27437
rect 561075 27372 561076 27436
rect 561140 27372 561141 27436
rect 561075 27371 561141 27372
rect 561630 26893 561690 682347
rect 564294 673954 564914 709082
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568619 683500 568685 683501
rect 568619 683436 568620 683500
rect 568684 683436 568685 683500
rect 568619 683435 568685 683436
rect 565123 682276 565189 682277
rect 565123 682212 565124 682276
rect 565188 682212 565189 682276
rect 565123 682211 565189 682212
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 561811 616180 561877 616181
rect 561811 616116 561812 616180
rect 561876 616116 561877 616180
rect 561811 616115 561877 616116
rect 561814 29341 561874 616115
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 563099 579460 563165 579461
rect 563099 579396 563100 579460
rect 563164 579396 563165 579460
rect 563099 579395 563165 579396
rect 561995 576740 562061 576741
rect 561995 576676 561996 576740
rect 562060 576676 562061 576740
rect 561995 576675 562061 576676
rect 561811 29340 561877 29341
rect 561811 29276 561812 29340
rect 561876 29276 561877 29340
rect 561811 29275 561877 29276
rect 561998 29205 562058 576675
rect 562179 166428 562245 166429
rect 562179 166364 562180 166428
rect 562244 166364 562245 166428
rect 562179 166363 562245 166364
rect 561995 29204 562061 29205
rect 561995 29140 561996 29204
rect 562060 29140 562061 29204
rect 561995 29139 562061 29140
rect 561627 26892 561693 26893
rect 561627 26828 561628 26892
rect 561692 26828 561693 26892
rect 561627 26827 561693 26828
rect 560891 11660 560957 11661
rect 560891 11596 560892 11660
rect 560956 11596 560957 11660
rect 560891 11595 560957 11596
rect 562182 6357 562242 166363
rect 563102 159357 563162 579395
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 563283 565180 563349 565181
rect 563283 565116 563284 565180
rect 563348 565116 563349 565180
rect 563283 565115 563349 565116
rect 563286 170373 563346 565115
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 563467 246940 563533 246941
rect 563467 246876 563468 246940
rect 563532 246876 563533 246940
rect 563467 246875 563533 246876
rect 563283 170372 563349 170373
rect 563283 170308 563284 170372
rect 563348 170308 563349 170372
rect 563283 170307 563349 170308
rect 563283 166292 563349 166293
rect 563283 166228 563284 166292
rect 563348 166228 563349 166292
rect 563283 166227 563349 166228
rect 563099 159356 563165 159357
rect 563099 159292 563100 159356
rect 563164 159292 563165 159356
rect 563099 159291 563165 159292
rect 563099 156636 563165 156637
rect 563099 156572 563100 156636
rect 563164 156572 563165 156636
rect 563099 156571 563165 156572
rect 563102 55317 563162 156571
rect 563099 55316 563165 55317
rect 563099 55252 563100 55316
rect 563164 55252 563165 55316
rect 563099 55251 563165 55252
rect 562179 6356 562245 6357
rect 562179 6292 562180 6356
rect 562244 6292 562245 6356
rect 562179 6291 562245 6292
rect 563286 3909 563346 166227
rect 563470 16965 563530 246875
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 563651 149156 563717 149157
rect 563651 149092 563652 149156
rect 563716 149092 563717 149156
rect 563651 149091 563717 149092
rect 563654 137325 563714 149091
rect 563651 137324 563717 137325
rect 563651 137260 563652 137324
rect 563716 137260 563717 137324
rect 563651 137259 563717 137260
rect 564019 136644 564085 136645
rect 564019 136580 564020 136644
rect 564084 136580 564085 136644
rect 564019 136579 564085 136580
rect 564022 99517 564082 136579
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564019 99516 564085 99517
rect 564019 99452 564020 99516
rect 564084 99452 564085 99516
rect 564019 99451 564085 99452
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 563467 16964 563533 16965
rect 563467 16900 563468 16964
rect 563532 16900 563533 16964
rect 563467 16899 563533 16900
rect 563283 3908 563349 3909
rect 563283 3844 563284 3908
rect 563348 3844 563349 3908
rect 563283 3843 563349 3844
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 -5146 564914 25398
rect 565126 21589 565186 682211
rect 566963 682140 567029 682141
rect 566963 682076 566964 682140
rect 567028 682076 567029 682140
rect 566963 682075 567029 682076
rect 565859 680780 565925 680781
rect 565859 680716 565860 680780
rect 565924 680716 565925 680780
rect 565859 680715 565925 680716
rect 565307 472700 565373 472701
rect 565307 472636 565308 472700
rect 565372 472636 565373 472700
rect 565307 472635 565373 472636
rect 565310 24445 565370 472635
rect 565491 400348 565557 400349
rect 565491 400284 565492 400348
rect 565556 400284 565557 400348
rect 565491 400283 565557 400284
rect 565307 24444 565373 24445
rect 565307 24380 565308 24444
rect 565372 24380 565373 24444
rect 565307 24379 565373 24380
rect 565494 21861 565554 400283
rect 565491 21860 565557 21861
rect 565491 21796 565492 21860
rect 565556 21796 565557 21860
rect 565491 21795 565557 21796
rect 565123 21588 565189 21589
rect 565123 21524 565124 21588
rect 565188 21524 565189 21588
rect 565123 21523 565189 21524
rect 565862 4045 565922 680715
rect 566043 663780 566109 663781
rect 566043 663716 566044 663780
rect 566108 663716 566109 663780
rect 566043 663715 566109 663716
rect 566046 27301 566106 663715
rect 566227 552260 566293 552261
rect 566227 552196 566228 552260
rect 566292 552196 566293 552260
rect 566227 552195 566293 552196
rect 566043 27300 566109 27301
rect 566043 27236 566044 27300
rect 566108 27236 566109 27300
rect 566043 27235 566109 27236
rect 566230 24037 566290 552195
rect 566411 551580 566477 551581
rect 566411 551516 566412 551580
rect 566476 551516 566477 551580
rect 566411 551515 566477 551516
rect 566414 25669 566474 551515
rect 566966 26250 567026 682075
rect 567331 580820 567397 580821
rect 567331 580756 567332 580820
rect 567396 580756 567397 580820
rect 567331 580755 567397 580756
rect 566966 26213 567210 26250
rect 566966 26212 567213 26213
rect 566966 26190 567148 26212
rect 567147 26148 567148 26190
rect 567212 26148 567213 26212
rect 567147 26147 567213 26148
rect 566411 25668 566477 25669
rect 566411 25604 566412 25668
rect 566476 25604 566477 25668
rect 566411 25603 566477 25604
rect 567334 24309 567394 580755
rect 567515 410820 567581 410821
rect 567515 410756 567516 410820
rect 567580 410756 567581 410820
rect 567515 410755 567581 410756
rect 567331 24308 567397 24309
rect 567331 24244 567332 24308
rect 567396 24244 567397 24308
rect 567331 24243 567397 24244
rect 566227 24036 566293 24037
rect 566227 23972 566228 24036
rect 566292 23972 566293 24036
rect 566227 23971 566293 23972
rect 567518 21453 567578 410755
rect 567515 21452 567581 21453
rect 567515 21388 567516 21452
rect 567580 21388 567581 21452
rect 567515 21387 567581 21388
rect 565859 4044 565925 4045
rect 565859 3980 565860 4044
rect 565924 3980 565925 4044
rect 565859 3979 565925 3980
rect 568622 3637 568682 683435
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 571379 666500 571445 666501
rect 571379 666436 571380 666500
rect 571444 666436 571445 666500
rect 571379 666435 571445 666436
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 570091 601900 570157 601901
rect 570091 601836 570092 601900
rect 570156 601836 570157 601900
rect 570091 601835 570157 601836
rect 570094 586530 570154 601835
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568619 3636 568685 3637
rect 568619 3572 568620 3636
rect 568684 3572 568685 3636
rect 568619 3571 568685 3572
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 -6106 569414 29898
rect 569910 586470 570154 586530
rect 569910 16590 569970 586470
rect 570091 582180 570157 582181
rect 570091 582116 570092 582180
rect 570156 582116 570157 582180
rect 570091 582115 570157 582116
rect 570094 21317 570154 582115
rect 571382 21725 571442 666435
rect 573294 646954 573914 682398
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 574139 682004 574205 682005
rect 574139 681940 574140 682004
rect 574204 681940 574205 682004
rect 574139 681939 574205 681940
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 571563 628420 571629 628421
rect 571563 628356 571564 628420
rect 571628 628356 571629 628420
rect 571563 628355 571629 628356
rect 571379 21724 571445 21725
rect 571379 21660 571380 21724
rect 571444 21660 571445 21724
rect 571379 21659 571445 21660
rect 570091 21316 570157 21317
rect 570091 21252 570092 21316
rect 570156 21252 570157 21316
rect 570091 21251 570157 21252
rect 569910 16530 570154 16590
rect 570094 3365 570154 16530
rect 571566 3773 571626 628355
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 571563 3772 571629 3773
rect 571563 3708 571564 3772
rect 571628 3708 571629 3772
rect 571563 3707 571629 3708
rect 570091 3364 570157 3365
rect 570091 3300 570092 3364
rect 570156 3300 570157 3364
rect 570091 3299 570157 3300
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 -7066 573914 34398
rect 574142 18733 574202 681939
rect 575427 681052 575493 681053
rect 575427 680988 575428 681052
rect 575492 680988 575493 681052
rect 575427 680987 575493 680988
rect 574323 544780 574389 544781
rect 574323 544716 574324 544780
rect 574388 544716 574389 544780
rect 574323 544715 574389 544716
rect 574139 18732 574205 18733
rect 574139 18668 574140 18732
rect 574204 18668 574205 18732
rect 574139 18667 574205 18668
rect 574326 3501 574386 544715
rect 575430 17509 575490 680987
rect 577794 651454 578414 686898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 578555 681868 578621 681869
rect 578555 681804 578556 681868
rect 578620 681804 578621 681868
rect 578555 681803 578621 681804
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 575611 650860 575677 650861
rect 575611 650796 575612 650860
rect 575676 650796 575677 650860
rect 575611 650795 575677 650796
rect 575614 29205 575674 650795
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 575611 29204 575677 29205
rect 575611 29140 575612 29204
rect 575676 29140 575677 29204
rect 575611 29139 575677 29140
rect 575427 17508 575493 17509
rect 575427 17444 575428 17508
rect 575492 17444 575493 17508
rect 575427 17443 575493 17444
rect 574323 3500 574389 3501
rect 574323 3436 574324 3500
rect 574388 3436 574389 3500
rect 574323 3435 574389 3436
rect 577794 3454 578414 38898
rect 578558 27165 578618 681803
rect 580947 669900 581013 669901
rect 580947 669836 580948 669900
rect 581012 669836 581013 669900
rect 580947 669835 581013 669836
rect 579659 646100 579725 646101
rect 579659 646036 579660 646100
rect 579724 646036 579725 646100
rect 579659 646035 579725 646036
rect 578739 602580 578805 602581
rect 578739 602516 578740 602580
rect 578804 602516 578805 602580
rect 578739 602515 578805 602516
rect 578555 27164 578621 27165
rect 578555 27100 578556 27164
rect 578620 27100 578621 27164
rect 578555 27099 578621 27100
rect 578742 22541 578802 602515
rect 579662 22813 579722 646035
rect 579659 22812 579725 22813
rect 579659 22748 579660 22812
rect 579724 22748 579725 22812
rect 579659 22747 579725 22748
rect 578739 22540 578805 22541
rect 578739 22476 578740 22540
rect 578804 22476 578805 22540
rect 578739 22475 578805 22476
rect 580950 17781 581010 669835
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 581131 590748 581197 590749
rect 581131 590684 581132 590748
rect 581196 590684 581197 590748
rect 581131 590683 581197 590684
rect 581134 23085 581194 590683
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 581131 23084 581197 23085
rect 581131 23020 581132 23084
rect 581196 23020 581197 23084
rect 581131 23019 581197 23020
rect 580947 17780 581013 17781
rect 580947 17716 580948 17780
rect 581012 17716 581013 17780
rect 580947 17715 581013 17716
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 36328 655718 36564 655954
rect 36328 655398 36564 655634
rect 172056 655718 172292 655954
rect 172056 655398 172292 655634
rect 37008 651218 37244 651454
rect 37008 650898 37244 651134
rect 171376 651218 171612 651454
rect 171376 650898 171612 651134
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 36328 619718 36564 619954
rect 36328 619398 36564 619634
rect 172056 619718 172292 619954
rect 172056 619398 172292 619634
rect 37008 615218 37244 615454
rect 37008 614898 37244 615134
rect 171376 615218 171612 615454
rect 171376 614898 171612 615134
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 210328 655718 210564 655954
rect 210328 655398 210564 655634
rect 346056 655718 346292 655954
rect 346056 655398 346292 655634
rect 211008 651218 211244 651454
rect 211008 650898 211244 651134
rect 345376 651218 345612 651454
rect 345376 650898 345612 651134
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 210328 619718 210564 619954
rect 210328 619398 210564 619634
rect 346056 619718 346292 619954
rect 346056 619398 346292 619634
rect 211008 615218 211244 615454
rect 211008 614898 211244 615134
rect 345376 615218 345612 615454
rect 345376 614898 345612 615134
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 67610 547718 67846 547954
rect 67610 547398 67846 547634
rect 98330 547718 98566 547954
rect 98330 547398 98566 547634
rect 129050 547718 129286 547954
rect 129050 547398 129286 547634
rect 159770 547718 160006 547954
rect 159770 547398 160006 547634
rect 190490 547718 190726 547954
rect 190490 547398 190726 547634
rect 221210 547718 221446 547954
rect 221210 547398 221446 547634
rect 251930 547718 252166 547954
rect 251930 547398 252166 547634
rect 282650 547718 282886 547954
rect 282650 547398 282886 547634
rect 313370 547718 313606 547954
rect 313370 547398 313606 547634
rect 344090 547718 344326 547954
rect 344090 547398 344326 547634
rect 52250 543218 52486 543454
rect 52250 542898 52486 543134
rect 82970 543218 83206 543454
rect 82970 542898 83206 543134
rect 113690 543218 113926 543454
rect 113690 542898 113926 543134
rect 144410 543218 144646 543454
rect 144410 542898 144646 543134
rect 175130 543218 175366 543454
rect 175130 542898 175366 543134
rect 205850 543218 206086 543454
rect 205850 542898 206086 543134
rect 236570 543218 236806 543454
rect 236570 542898 236806 543134
rect 267290 543218 267526 543454
rect 267290 542898 267526 543134
rect 298010 543218 298246 543454
rect 298010 542898 298246 543134
rect 328730 543218 328966 543454
rect 328730 542898 328966 543134
rect 67610 511718 67846 511954
rect 67610 511398 67846 511634
rect 98330 511718 98566 511954
rect 98330 511398 98566 511634
rect 129050 511718 129286 511954
rect 129050 511398 129286 511634
rect 159770 511718 160006 511954
rect 159770 511398 160006 511634
rect 190490 511718 190726 511954
rect 190490 511398 190726 511634
rect 221210 511718 221446 511954
rect 221210 511398 221446 511634
rect 251930 511718 252166 511954
rect 251930 511398 252166 511634
rect 282650 511718 282886 511954
rect 282650 511398 282886 511634
rect 313370 511718 313606 511954
rect 313370 511398 313606 511634
rect 344090 511718 344326 511954
rect 344090 511398 344326 511634
rect 52250 507218 52486 507454
rect 52250 506898 52486 507134
rect 82970 507218 83206 507454
rect 82970 506898 83206 507134
rect 113690 507218 113926 507454
rect 113690 506898 113926 507134
rect 144410 507218 144646 507454
rect 144410 506898 144646 507134
rect 175130 507218 175366 507454
rect 175130 506898 175366 507134
rect 205850 507218 206086 507454
rect 205850 506898 206086 507134
rect 236570 507218 236806 507454
rect 236570 506898 236806 507134
rect 267290 507218 267526 507454
rect 267290 506898 267526 507134
rect 298010 507218 298246 507454
rect 298010 506898 298246 507134
rect 328730 507218 328966 507454
rect 328730 506898 328966 507134
rect 67610 475718 67846 475954
rect 67610 475398 67846 475634
rect 98330 475718 98566 475954
rect 98330 475398 98566 475634
rect 129050 475718 129286 475954
rect 129050 475398 129286 475634
rect 159770 475718 160006 475954
rect 159770 475398 160006 475634
rect 190490 475718 190726 475954
rect 190490 475398 190726 475634
rect 221210 475718 221446 475954
rect 221210 475398 221446 475634
rect 251930 475718 252166 475954
rect 251930 475398 252166 475634
rect 282650 475718 282886 475954
rect 282650 475398 282886 475634
rect 313370 475718 313606 475954
rect 313370 475398 313606 475634
rect 344090 475718 344326 475954
rect 344090 475398 344326 475634
rect 52250 471218 52486 471454
rect 52250 470898 52486 471134
rect 82970 471218 83206 471454
rect 82970 470898 83206 471134
rect 113690 471218 113926 471454
rect 113690 470898 113926 471134
rect 144410 471218 144646 471454
rect 144410 470898 144646 471134
rect 175130 471218 175366 471454
rect 175130 470898 175366 471134
rect 205850 471218 206086 471454
rect 205850 470898 206086 471134
rect 236570 471218 236806 471454
rect 236570 470898 236806 471134
rect 267290 471218 267526 471454
rect 267290 470898 267526 471134
rect 298010 471218 298246 471454
rect 298010 470898 298246 471134
rect 328730 471218 328966 471454
rect 328730 470898 328966 471134
rect 67610 439718 67846 439954
rect 67610 439398 67846 439634
rect 98330 439718 98566 439954
rect 98330 439398 98566 439634
rect 129050 439718 129286 439954
rect 129050 439398 129286 439634
rect 159770 439718 160006 439954
rect 159770 439398 160006 439634
rect 190490 439718 190726 439954
rect 190490 439398 190726 439634
rect 221210 439718 221446 439954
rect 221210 439398 221446 439634
rect 251930 439718 252166 439954
rect 251930 439398 252166 439634
rect 282650 439718 282886 439954
rect 282650 439398 282886 439634
rect 313370 439718 313606 439954
rect 313370 439398 313606 439634
rect 344090 439718 344326 439954
rect 344090 439398 344326 439634
rect 52250 435218 52486 435454
rect 52250 434898 52486 435134
rect 82970 435218 83206 435454
rect 82970 434898 83206 435134
rect 113690 435218 113926 435454
rect 113690 434898 113926 435134
rect 144410 435218 144646 435454
rect 144410 434898 144646 435134
rect 175130 435218 175366 435454
rect 175130 434898 175366 435134
rect 205850 435218 206086 435454
rect 205850 434898 206086 435134
rect 236570 435218 236806 435454
rect 236570 434898 236806 435134
rect 267290 435218 267526 435454
rect 267290 434898 267526 435134
rect 298010 435218 298246 435454
rect 298010 434898 298246 435134
rect 328730 435218 328966 435454
rect 328730 434898 328966 435134
rect 67610 403718 67846 403954
rect 67610 403398 67846 403634
rect 98330 403718 98566 403954
rect 98330 403398 98566 403634
rect 129050 403718 129286 403954
rect 129050 403398 129286 403634
rect 159770 403718 160006 403954
rect 159770 403398 160006 403634
rect 190490 403718 190726 403954
rect 190490 403398 190726 403634
rect 221210 403718 221446 403954
rect 221210 403398 221446 403634
rect 251930 403718 252166 403954
rect 251930 403398 252166 403634
rect 282650 403718 282886 403954
rect 282650 403398 282886 403634
rect 313370 403718 313606 403954
rect 313370 403398 313606 403634
rect 344090 403718 344326 403954
rect 344090 403398 344326 403634
rect 52250 399218 52486 399454
rect 52250 398898 52486 399134
rect 82970 399218 83206 399454
rect 82970 398898 83206 399134
rect 113690 399218 113926 399454
rect 113690 398898 113926 399134
rect 144410 399218 144646 399454
rect 144410 398898 144646 399134
rect 175130 399218 175366 399454
rect 175130 398898 175366 399134
rect 205850 399218 206086 399454
rect 205850 398898 206086 399134
rect 236570 399218 236806 399454
rect 236570 398898 236806 399134
rect 267290 399218 267526 399454
rect 267290 398898 267526 399134
rect 298010 399218 298246 399454
rect 298010 398898 298246 399134
rect 328730 399218 328966 399454
rect 328730 398898 328966 399134
rect 67610 367718 67846 367954
rect 67610 367398 67846 367634
rect 98330 367718 98566 367954
rect 98330 367398 98566 367634
rect 129050 367718 129286 367954
rect 129050 367398 129286 367634
rect 159770 367718 160006 367954
rect 159770 367398 160006 367634
rect 190490 367718 190726 367954
rect 190490 367398 190726 367634
rect 221210 367718 221446 367954
rect 221210 367398 221446 367634
rect 251930 367718 252166 367954
rect 251930 367398 252166 367634
rect 282650 367718 282886 367954
rect 282650 367398 282886 367634
rect 313370 367718 313606 367954
rect 313370 367398 313606 367634
rect 344090 367718 344326 367954
rect 344090 367398 344326 367634
rect 52250 363218 52486 363454
rect 52250 362898 52486 363134
rect 82970 363218 83206 363454
rect 82970 362898 83206 363134
rect 113690 363218 113926 363454
rect 113690 362898 113926 363134
rect 144410 363218 144646 363454
rect 144410 362898 144646 363134
rect 175130 363218 175366 363454
rect 175130 362898 175366 363134
rect 205850 363218 206086 363454
rect 205850 362898 206086 363134
rect 236570 363218 236806 363454
rect 236570 362898 236806 363134
rect 267290 363218 267526 363454
rect 267290 362898 267526 363134
rect 298010 363218 298246 363454
rect 298010 362898 298246 363134
rect 328730 363218 328966 363454
rect 328730 362898 328966 363134
rect 67610 331718 67846 331954
rect 67610 331398 67846 331634
rect 98330 331718 98566 331954
rect 98330 331398 98566 331634
rect 129050 331718 129286 331954
rect 129050 331398 129286 331634
rect 159770 331718 160006 331954
rect 159770 331398 160006 331634
rect 190490 331718 190726 331954
rect 190490 331398 190726 331634
rect 221210 331718 221446 331954
rect 221210 331398 221446 331634
rect 251930 331718 252166 331954
rect 251930 331398 252166 331634
rect 282650 331718 282886 331954
rect 282650 331398 282886 331634
rect 313370 331718 313606 331954
rect 313370 331398 313606 331634
rect 344090 331718 344326 331954
rect 344090 331398 344326 331634
rect 52250 327218 52486 327454
rect 52250 326898 52486 327134
rect 82970 327218 83206 327454
rect 82970 326898 83206 327134
rect 113690 327218 113926 327454
rect 113690 326898 113926 327134
rect 144410 327218 144646 327454
rect 144410 326898 144646 327134
rect 175130 327218 175366 327454
rect 175130 326898 175366 327134
rect 205850 327218 206086 327454
rect 205850 326898 206086 327134
rect 236570 327218 236806 327454
rect 236570 326898 236806 327134
rect 267290 327218 267526 327454
rect 267290 326898 267526 327134
rect 298010 327218 298246 327454
rect 298010 326898 298246 327134
rect 328730 327218 328966 327454
rect 328730 326898 328966 327134
rect 67610 295718 67846 295954
rect 67610 295398 67846 295634
rect 98330 295718 98566 295954
rect 98330 295398 98566 295634
rect 129050 295718 129286 295954
rect 129050 295398 129286 295634
rect 159770 295718 160006 295954
rect 159770 295398 160006 295634
rect 190490 295718 190726 295954
rect 190490 295398 190726 295634
rect 221210 295718 221446 295954
rect 221210 295398 221446 295634
rect 251930 295718 252166 295954
rect 251930 295398 252166 295634
rect 282650 295718 282886 295954
rect 282650 295398 282886 295634
rect 313370 295718 313606 295954
rect 313370 295398 313606 295634
rect 344090 295718 344326 295954
rect 344090 295398 344326 295634
rect 52250 291218 52486 291454
rect 52250 290898 52486 291134
rect 82970 291218 83206 291454
rect 82970 290898 83206 291134
rect 113690 291218 113926 291454
rect 113690 290898 113926 291134
rect 144410 291218 144646 291454
rect 144410 290898 144646 291134
rect 175130 291218 175366 291454
rect 175130 290898 175366 291134
rect 205850 291218 206086 291454
rect 205850 290898 206086 291134
rect 236570 291218 236806 291454
rect 236570 290898 236806 291134
rect 267290 291218 267526 291454
rect 267290 290898 267526 291134
rect 298010 291218 298246 291454
rect 298010 290898 298246 291134
rect 328730 291218 328966 291454
rect 328730 290898 328966 291134
rect 67610 259718 67846 259954
rect 67610 259398 67846 259634
rect 98330 259718 98566 259954
rect 98330 259398 98566 259634
rect 129050 259718 129286 259954
rect 129050 259398 129286 259634
rect 159770 259718 160006 259954
rect 159770 259398 160006 259634
rect 190490 259718 190726 259954
rect 190490 259398 190726 259634
rect 221210 259718 221446 259954
rect 221210 259398 221446 259634
rect 251930 259718 252166 259954
rect 251930 259398 252166 259634
rect 282650 259718 282886 259954
rect 282650 259398 282886 259634
rect 313370 259718 313606 259954
rect 313370 259398 313606 259634
rect 344090 259718 344326 259954
rect 344090 259398 344326 259634
rect 52250 255218 52486 255454
rect 52250 254898 52486 255134
rect 82970 255218 83206 255454
rect 82970 254898 83206 255134
rect 113690 255218 113926 255454
rect 113690 254898 113926 255134
rect 144410 255218 144646 255454
rect 144410 254898 144646 255134
rect 175130 255218 175366 255454
rect 175130 254898 175366 255134
rect 205850 255218 206086 255454
rect 205850 254898 206086 255134
rect 236570 255218 236806 255454
rect 236570 254898 236806 255134
rect 267290 255218 267526 255454
rect 267290 254898 267526 255134
rect 298010 255218 298246 255454
rect 298010 254898 298246 255134
rect 328730 255218 328966 255454
rect 328730 254898 328966 255134
rect 67610 223718 67846 223954
rect 67610 223398 67846 223634
rect 98330 223718 98566 223954
rect 98330 223398 98566 223634
rect 129050 223718 129286 223954
rect 129050 223398 129286 223634
rect 159770 223718 160006 223954
rect 159770 223398 160006 223634
rect 190490 223718 190726 223954
rect 190490 223398 190726 223634
rect 221210 223718 221446 223954
rect 221210 223398 221446 223634
rect 251930 223718 252166 223954
rect 251930 223398 252166 223634
rect 282650 223718 282886 223954
rect 282650 223398 282886 223634
rect 313370 223718 313606 223954
rect 313370 223398 313606 223634
rect 344090 223718 344326 223954
rect 344090 223398 344326 223634
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 52250 219218 52486 219454
rect 52250 218898 52486 219134
rect 82970 219218 83206 219454
rect 82970 218898 83206 219134
rect 113690 219218 113926 219454
rect 113690 218898 113926 219134
rect 144410 219218 144646 219454
rect 144410 218898 144646 219134
rect 175130 219218 175366 219454
rect 175130 218898 175366 219134
rect 205850 219218 206086 219454
rect 205850 218898 206086 219134
rect 236570 219218 236806 219454
rect 236570 218898 236806 219134
rect 267290 219218 267526 219454
rect 267290 218898 267526 219134
rect 298010 219218 298246 219454
rect 298010 218898 298246 219134
rect 328730 219218 328966 219454
rect 328730 218898 328966 219134
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 429610 655718 429846 655954
rect 429610 655398 429846 655634
rect 460330 655718 460566 655954
rect 460330 655398 460566 655634
rect 491050 655718 491286 655954
rect 491050 655398 491286 655634
rect 521770 655718 522006 655954
rect 521770 655398 522006 655634
rect 414250 651218 414486 651454
rect 414250 650898 414486 651134
rect 444970 651218 445206 651454
rect 444970 650898 445206 651134
rect 475690 651218 475926 651454
rect 475690 650898 475926 651134
rect 506410 651218 506646 651454
rect 506410 650898 506646 651134
rect 537130 651218 537366 651454
rect 537130 650898 537366 651134
rect 429610 619718 429846 619954
rect 429610 619398 429846 619634
rect 460330 619718 460566 619954
rect 460330 619398 460566 619634
rect 491050 619718 491286 619954
rect 491050 619398 491286 619634
rect 521770 619718 522006 619954
rect 521770 619398 522006 619634
rect 414250 615218 414486 615454
rect 414250 614898 414486 615134
rect 444970 615218 445206 615454
rect 444970 614898 445206 615134
rect 475690 615218 475926 615454
rect 475690 614898 475926 615134
rect 506410 615218 506646 615454
rect 506410 614898 506646 615134
rect 537130 615218 537366 615454
rect 537130 614898 537366 615134
rect 429610 583718 429846 583954
rect 429610 583398 429846 583634
rect 460330 583718 460566 583954
rect 460330 583398 460566 583634
rect 491050 583718 491286 583954
rect 491050 583398 491286 583634
rect 521770 583718 522006 583954
rect 521770 583398 522006 583634
rect 414250 579218 414486 579454
rect 414250 578898 414486 579134
rect 444970 579218 445206 579454
rect 444970 578898 445206 579134
rect 475690 579218 475926 579454
rect 475690 578898 475926 579134
rect 506410 579218 506646 579454
rect 506410 578898 506646 579134
rect 537130 579218 537366 579454
rect 537130 578898 537366 579134
rect 429610 547718 429846 547954
rect 429610 547398 429846 547634
rect 460330 547718 460566 547954
rect 460330 547398 460566 547634
rect 491050 547718 491286 547954
rect 491050 547398 491286 547634
rect 521770 547718 522006 547954
rect 521770 547398 522006 547634
rect 414250 543218 414486 543454
rect 414250 542898 414486 543134
rect 444970 543218 445206 543454
rect 444970 542898 445206 543134
rect 475690 543218 475926 543454
rect 475690 542898 475926 543134
rect 506410 543218 506646 543454
rect 506410 542898 506646 543134
rect 537130 543218 537366 543454
rect 537130 542898 537366 543134
rect 429610 511718 429846 511954
rect 429610 511398 429846 511634
rect 460330 511718 460566 511954
rect 460330 511398 460566 511634
rect 491050 511718 491286 511954
rect 491050 511398 491286 511634
rect 521770 511718 522006 511954
rect 521770 511398 522006 511634
rect 414250 507218 414486 507454
rect 414250 506898 414486 507134
rect 444970 507218 445206 507454
rect 444970 506898 445206 507134
rect 475690 507218 475926 507454
rect 475690 506898 475926 507134
rect 506410 507218 506646 507454
rect 506410 506898 506646 507134
rect 537130 507218 537366 507454
rect 537130 506898 537366 507134
rect 429610 475718 429846 475954
rect 429610 475398 429846 475634
rect 460330 475718 460566 475954
rect 460330 475398 460566 475634
rect 491050 475718 491286 475954
rect 491050 475398 491286 475634
rect 521770 475718 522006 475954
rect 521770 475398 522006 475634
rect 414250 471218 414486 471454
rect 414250 470898 414486 471134
rect 444970 471218 445206 471454
rect 444970 470898 445206 471134
rect 475690 471218 475926 471454
rect 475690 470898 475926 471134
rect 506410 471218 506646 471454
rect 506410 470898 506646 471134
rect 537130 471218 537366 471454
rect 537130 470898 537366 471134
rect 429610 439718 429846 439954
rect 429610 439398 429846 439634
rect 460330 439718 460566 439954
rect 460330 439398 460566 439634
rect 491050 439718 491286 439954
rect 491050 439398 491286 439634
rect 521770 439718 522006 439954
rect 521770 439398 522006 439634
rect 414250 435218 414486 435454
rect 414250 434898 414486 435134
rect 444970 435218 445206 435454
rect 444970 434898 445206 435134
rect 475690 435218 475926 435454
rect 475690 434898 475926 435134
rect 506410 435218 506646 435454
rect 506410 434898 506646 435134
rect 537130 435218 537366 435454
rect 537130 434898 537366 435134
rect 429610 403718 429846 403954
rect 429610 403398 429846 403634
rect 460330 403718 460566 403954
rect 460330 403398 460566 403634
rect 491050 403718 491286 403954
rect 491050 403398 491286 403634
rect 521770 403718 522006 403954
rect 521770 403398 522006 403634
rect 414250 399218 414486 399454
rect 414250 398898 414486 399134
rect 444970 399218 445206 399454
rect 444970 398898 445206 399134
rect 475690 399218 475926 399454
rect 475690 398898 475926 399134
rect 506410 399218 506646 399454
rect 506410 398898 506646 399134
rect 537130 399218 537366 399454
rect 537130 398898 537366 399134
rect 429610 367718 429846 367954
rect 429610 367398 429846 367634
rect 460330 367718 460566 367954
rect 460330 367398 460566 367634
rect 491050 367718 491286 367954
rect 491050 367398 491286 367634
rect 521770 367718 522006 367954
rect 521770 367398 522006 367634
rect 414250 363218 414486 363454
rect 414250 362898 414486 363134
rect 444970 363218 445206 363454
rect 444970 362898 445206 363134
rect 475690 363218 475926 363454
rect 475690 362898 475926 363134
rect 506410 363218 506646 363454
rect 506410 362898 506646 363134
rect 537130 363218 537366 363454
rect 537130 362898 537366 363134
rect 429610 331718 429846 331954
rect 429610 331398 429846 331634
rect 460330 331718 460566 331954
rect 460330 331398 460566 331634
rect 491050 331718 491286 331954
rect 491050 331398 491286 331634
rect 521770 331718 522006 331954
rect 521770 331398 522006 331634
rect 414250 327218 414486 327454
rect 414250 326898 414486 327134
rect 444970 327218 445206 327454
rect 444970 326898 445206 327134
rect 475690 327218 475926 327454
rect 475690 326898 475926 327134
rect 506410 327218 506646 327454
rect 506410 326898 506646 327134
rect 537130 327218 537366 327454
rect 537130 326898 537366 327134
rect 429610 295718 429846 295954
rect 429610 295398 429846 295634
rect 460330 295718 460566 295954
rect 460330 295398 460566 295634
rect 491050 295718 491286 295954
rect 491050 295398 491286 295634
rect 521770 295718 522006 295954
rect 521770 295398 522006 295634
rect 414250 291218 414486 291454
rect 414250 290898 414486 291134
rect 444970 291218 445206 291454
rect 444970 290898 445206 291134
rect 475690 291218 475926 291454
rect 475690 290898 475926 291134
rect 506410 291218 506646 291454
rect 506410 290898 506646 291134
rect 537130 291218 537366 291454
rect 537130 290898 537366 291134
rect 429610 259718 429846 259954
rect 429610 259398 429846 259634
rect 460330 259718 460566 259954
rect 460330 259398 460566 259634
rect 491050 259718 491286 259954
rect 491050 259398 491286 259634
rect 521770 259718 522006 259954
rect 521770 259398 522006 259634
rect 414250 255218 414486 255454
rect 414250 254898 414486 255134
rect 444970 255218 445206 255454
rect 444970 254898 445206 255134
rect 475690 255218 475926 255454
rect 475690 254898 475926 255134
rect 506410 255218 506646 255454
rect 506410 254898 506646 255134
rect 537130 255218 537366 255454
rect 537130 254898 537366 255134
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 248570 147218 248806 147454
rect 248570 146898 248806 147134
rect 279290 147218 279526 147454
rect 279290 146898 279526 147134
rect 310010 147218 310246 147454
rect 310010 146898 310246 147134
rect 340730 147218 340966 147454
rect 340730 146898 340966 147134
rect 371450 147218 371686 147454
rect 371450 146898 371686 147134
rect 402170 147218 402406 147454
rect 402170 146898 402406 147134
rect 432890 147218 433126 147454
rect 432890 146898 433126 147134
rect 463610 147218 463846 147454
rect 463610 146898 463846 147134
rect 494330 147218 494566 147454
rect 494330 146898 494566 147134
rect 525050 147218 525286 147454
rect 525050 146898 525286 147134
rect 79610 115718 79846 115954
rect 79610 115398 79846 115634
rect 110330 115718 110566 115954
rect 110330 115398 110566 115634
rect 141050 115718 141286 115954
rect 141050 115398 141286 115634
rect 171770 115718 172006 115954
rect 171770 115398 172006 115634
rect 202490 115718 202726 115954
rect 202490 115398 202726 115634
rect 233210 115718 233446 115954
rect 233210 115398 233446 115634
rect 263930 115718 264166 115954
rect 263930 115398 264166 115634
rect 294650 115718 294886 115954
rect 294650 115398 294886 115634
rect 325370 115718 325606 115954
rect 325370 115398 325606 115634
rect 356090 115718 356326 115954
rect 356090 115398 356326 115634
rect 386810 115718 387046 115954
rect 386810 115398 387046 115634
rect 417530 115718 417766 115954
rect 417530 115398 417766 115634
rect 448250 115718 448486 115954
rect 448250 115398 448486 115634
rect 478970 115718 479206 115954
rect 478970 115398 479206 115634
rect 509690 115718 509926 115954
rect 509690 115398 509926 115634
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 248570 111218 248806 111454
rect 248570 110898 248806 111134
rect 279290 111218 279526 111454
rect 279290 110898 279526 111134
rect 310010 111218 310246 111454
rect 310010 110898 310246 111134
rect 340730 111218 340966 111454
rect 340730 110898 340966 111134
rect 371450 111218 371686 111454
rect 371450 110898 371686 111134
rect 402170 111218 402406 111454
rect 402170 110898 402406 111134
rect 432890 111218 433126 111454
rect 432890 110898 433126 111134
rect 463610 111218 463846 111454
rect 463610 110898 463846 111134
rect 494330 111218 494566 111454
rect 494330 110898 494566 111134
rect 525050 111218 525286 111454
rect 525050 110898 525286 111134
rect 79610 79718 79846 79954
rect 79610 79398 79846 79634
rect 110330 79718 110566 79954
rect 110330 79398 110566 79634
rect 141050 79718 141286 79954
rect 141050 79398 141286 79634
rect 171770 79718 172006 79954
rect 171770 79398 172006 79634
rect 202490 79718 202726 79954
rect 202490 79398 202726 79634
rect 233210 79718 233446 79954
rect 233210 79398 233446 79634
rect 263930 79718 264166 79954
rect 263930 79398 264166 79634
rect 294650 79718 294886 79954
rect 294650 79398 294886 79634
rect 325370 79718 325606 79954
rect 325370 79398 325606 79634
rect 356090 79718 356326 79954
rect 356090 79398 356326 79634
rect 386810 79718 387046 79954
rect 386810 79398 387046 79634
rect 417530 79718 417766 79954
rect 417530 79398 417766 79634
rect 448250 79718 448486 79954
rect 448250 79398 448486 79634
rect 478970 79718 479206 79954
rect 478970 79398 479206 79634
rect 509690 79718 509926 79954
rect 509690 79398 509926 79634
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 248570 75218 248806 75454
rect 248570 74898 248806 75134
rect 279290 75218 279526 75454
rect 279290 74898 279526 75134
rect 310010 75218 310246 75454
rect 310010 74898 310246 75134
rect 340730 75218 340966 75454
rect 340730 74898 340966 75134
rect 371450 75218 371686 75454
rect 371450 74898 371686 75134
rect 402170 75218 402406 75454
rect 402170 74898 402406 75134
rect 432890 75218 433126 75454
rect 432890 74898 433126 75134
rect 463610 75218 463846 75454
rect 463610 74898 463846 75134
rect 494330 75218 494566 75454
rect 494330 74898 494566 75134
rect 525050 75218 525286 75454
rect 525050 74898 525286 75134
rect 79610 43718 79846 43954
rect 79610 43398 79846 43634
rect 110330 43718 110566 43954
rect 110330 43398 110566 43634
rect 141050 43718 141286 43954
rect 141050 43398 141286 43634
rect 171770 43718 172006 43954
rect 171770 43398 172006 43634
rect 202490 43718 202726 43954
rect 202490 43398 202726 43634
rect 233210 43718 233446 43954
rect 233210 43398 233446 43634
rect 263930 43718 264166 43954
rect 263930 43398 264166 43634
rect 294650 43718 294886 43954
rect 294650 43398 294886 43634
rect 325370 43718 325606 43954
rect 325370 43398 325606 43634
rect 356090 43718 356326 43954
rect 356090 43398 356326 43634
rect 386810 43718 387046 43954
rect 386810 43398 387046 43634
rect 417530 43718 417766 43954
rect 417530 43398 417766 43634
rect 448250 43718 448486 43954
rect 448250 43398 448486 43634
rect 478970 43718 479206 43954
rect 478970 43398 479206 43634
rect 509690 43718 509926 43954
rect 509690 43398 509926 43634
rect 64250 39218 64486 39454
rect 64250 38898 64486 39134
rect 94970 39218 95206 39454
rect 94970 38898 95206 39134
rect 125690 39218 125926 39454
rect 125690 38898 125926 39134
rect 156410 39218 156646 39454
rect 156410 38898 156646 39134
rect 187130 39218 187366 39454
rect 187130 38898 187366 39134
rect 217850 39218 218086 39454
rect 217850 38898 218086 39134
rect 248570 39218 248806 39454
rect 248570 38898 248806 39134
rect 279290 39218 279526 39454
rect 279290 38898 279526 39134
rect 310010 39218 310246 39454
rect 310010 38898 310246 39134
rect 340730 39218 340966 39454
rect 340730 38898 340966 39134
rect 371450 39218 371686 39454
rect 371450 38898 371686 39134
rect 402170 39218 402406 39454
rect 402170 38898 402406 39134
rect 432890 39218 433126 39454
rect 432890 38898 433126 39134
rect 463610 39218 463846 39454
rect 463610 38898 463846 39134
rect 494330 39218 494566 39454
rect 494330 38898 494566 39134
rect 525050 39218 525286 39454
rect 525050 38898 525286 39134
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 36328 655954
rect 36564 655718 172056 655954
rect 172292 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 210328 655954
rect 210564 655718 346056 655954
rect 346292 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 429610 655954
rect 429846 655718 460330 655954
rect 460566 655718 491050 655954
rect 491286 655718 521770 655954
rect 522006 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 36328 655634
rect 36564 655398 172056 655634
rect 172292 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 210328 655634
rect 210564 655398 346056 655634
rect 346292 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 429610 655634
rect 429846 655398 460330 655634
rect 460566 655398 491050 655634
rect 491286 655398 521770 655634
rect 522006 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37008 651454
rect 37244 651218 171376 651454
rect 171612 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 211008 651454
rect 211244 651218 345376 651454
rect 345612 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 414250 651454
rect 414486 651218 444970 651454
rect 445206 651218 475690 651454
rect 475926 651218 506410 651454
rect 506646 651218 537130 651454
rect 537366 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37008 651134
rect 37244 650898 171376 651134
rect 171612 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 211008 651134
rect 211244 650898 345376 651134
rect 345612 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 414250 651134
rect 414486 650898 444970 651134
rect 445206 650898 475690 651134
rect 475926 650898 506410 651134
rect 506646 650898 537130 651134
rect 537366 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 36328 619954
rect 36564 619718 172056 619954
rect 172292 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 210328 619954
rect 210564 619718 346056 619954
rect 346292 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 429610 619954
rect 429846 619718 460330 619954
rect 460566 619718 491050 619954
rect 491286 619718 521770 619954
rect 522006 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 36328 619634
rect 36564 619398 172056 619634
rect 172292 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 210328 619634
rect 210564 619398 346056 619634
rect 346292 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 429610 619634
rect 429846 619398 460330 619634
rect 460566 619398 491050 619634
rect 491286 619398 521770 619634
rect 522006 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37008 615454
rect 37244 615218 171376 615454
rect 171612 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 211008 615454
rect 211244 615218 345376 615454
rect 345612 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 414250 615454
rect 414486 615218 444970 615454
rect 445206 615218 475690 615454
rect 475926 615218 506410 615454
rect 506646 615218 537130 615454
rect 537366 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37008 615134
rect 37244 614898 171376 615134
rect 171612 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 211008 615134
rect 211244 614898 345376 615134
rect 345612 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 414250 615134
rect 414486 614898 444970 615134
rect 445206 614898 475690 615134
rect 475926 614898 506410 615134
rect 506646 614898 537130 615134
rect 537366 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 429610 583954
rect 429846 583718 460330 583954
rect 460566 583718 491050 583954
rect 491286 583718 521770 583954
rect 522006 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 429610 583634
rect 429846 583398 460330 583634
rect 460566 583398 491050 583634
rect 491286 583398 521770 583634
rect 522006 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 414250 579454
rect 414486 579218 444970 579454
rect 445206 579218 475690 579454
rect 475926 579218 506410 579454
rect 506646 579218 537130 579454
rect 537366 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 414250 579134
rect 414486 578898 444970 579134
rect 445206 578898 475690 579134
rect 475926 578898 506410 579134
rect 506646 578898 537130 579134
rect 537366 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 67610 547954
rect 67846 547718 98330 547954
rect 98566 547718 129050 547954
rect 129286 547718 159770 547954
rect 160006 547718 190490 547954
rect 190726 547718 221210 547954
rect 221446 547718 251930 547954
rect 252166 547718 282650 547954
rect 282886 547718 313370 547954
rect 313606 547718 344090 547954
rect 344326 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 429610 547954
rect 429846 547718 460330 547954
rect 460566 547718 491050 547954
rect 491286 547718 521770 547954
rect 522006 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 67610 547634
rect 67846 547398 98330 547634
rect 98566 547398 129050 547634
rect 129286 547398 159770 547634
rect 160006 547398 190490 547634
rect 190726 547398 221210 547634
rect 221446 547398 251930 547634
rect 252166 547398 282650 547634
rect 282886 547398 313370 547634
rect 313606 547398 344090 547634
rect 344326 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 429610 547634
rect 429846 547398 460330 547634
rect 460566 547398 491050 547634
rect 491286 547398 521770 547634
rect 522006 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 52250 543454
rect 52486 543218 82970 543454
rect 83206 543218 113690 543454
rect 113926 543218 144410 543454
rect 144646 543218 175130 543454
rect 175366 543218 205850 543454
rect 206086 543218 236570 543454
rect 236806 543218 267290 543454
rect 267526 543218 298010 543454
rect 298246 543218 328730 543454
rect 328966 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 414250 543454
rect 414486 543218 444970 543454
rect 445206 543218 475690 543454
rect 475926 543218 506410 543454
rect 506646 543218 537130 543454
rect 537366 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 52250 543134
rect 52486 542898 82970 543134
rect 83206 542898 113690 543134
rect 113926 542898 144410 543134
rect 144646 542898 175130 543134
rect 175366 542898 205850 543134
rect 206086 542898 236570 543134
rect 236806 542898 267290 543134
rect 267526 542898 298010 543134
rect 298246 542898 328730 543134
rect 328966 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 414250 543134
rect 414486 542898 444970 543134
rect 445206 542898 475690 543134
rect 475926 542898 506410 543134
rect 506646 542898 537130 543134
rect 537366 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 67610 511954
rect 67846 511718 98330 511954
rect 98566 511718 129050 511954
rect 129286 511718 159770 511954
rect 160006 511718 190490 511954
rect 190726 511718 221210 511954
rect 221446 511718 251930 511954
rect 252166 511718 282650 511954
rect 282886 511718 313370 511954
rect 313606 511718 344090 511954
rect 344326 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 429610 511954
rect 429846 511718 460330 511954
rect 460566 511718 491050 511954
rect 491286 511718 521770 511954
rect 522006 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 67610 511634
rect 67846 511398 98330 511634
rect 98566 511398 129050 511634
rect 129286 511398 159770 511634
rect 160006 511398 190490 511634
rect 190726 511398 221210 511634
rect 221446 511398 251930 511634
rect 252166 511398 282650 511634
rect 282886 511398 313370 511634
rect 313606 511398 344090 511634
rect 344326 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 429610 511634
rect 429846 511398 460330 511634
rect 460566 511398 491050 511634
rect 491286 511398 521770 511634
rect 522006 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 52250 507454
rect 52486 507218 82970 507454
rect 83206 507218 113690 507454
rect 113926 507218 144410 507454
rect 144646 507218 175130 507454
rect 175366 507218 205850 507454
rect 206086 507218 236570 507454
rect 236806 507218 267290 507454
rect 267526 507218 298010 507454
rect 298246 507218 328730 507454
rect 328966 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 414250 507454
rect 414486 507218 444970 507454
rect 445206 507218 475690 507454
rect 475926 507218 506410 507454
rect 506646 507218 537130 507454
rect 537366 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 52250 507134
rect 52486 506898 82970 507134
rect 83206 506898 113690 507134
rect 113926 506898 144410 507134
rect 144646 506898 175130 507134
rect 175366 506898 205850 507134
rect 206086 506898 236570 507134
rect 236806 506898 267290 507134
rect 267526 506898 298010 507134
rect 298246 506898 328730 507134
rect 328966 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 414250 507134
rect 414486 506898 444970 507134
rect 445206 506898 475690 507134
rect 475926 506898 506410 507134
rect 506646 506898 537130 507134
rect 537366 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 67610 475954
rect 67846 475718 98330 475954
rect 98566 475718 129050 475954
rect 129286 475718 159770 475954
rect 160006 475718 190490 475954
rect 190726 475718 221210 475954
rect 221446 475718 251930 475954
rect 252166 475718 282650 475954
rect 282886 475718 313370 475954
rect 313606 475718 344090 475954
rect 344326 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 429610 475954
rect 429846 475718 460330 475954
rect 460566 475718 491050 475954
rect 491286 475718 521770 475954
rect 522006 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 67610 475634
rect 67846 475398 98330 475634
rect 98566 475398 129050 475634
rect 129286 475398 159770 475634
rect 160006 475398 190490 475634
rect 190726 475398 221210 475634
rect 221446 475398 251930 475634
rect 252166 475398 282650 475634
rect 282886 475398 313370 475634
rect 313606 475398 344090 475634
rect 344326 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 429610 475634
rect 429846 475398 460330 475634
rect 460566 475398 491050 475634
rect 491286 475398 521770 475634
rect 522006 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 52250 471454
rect 52486 471218 82970 471454
rect 83206 471218 113690 471454
rect 113926 471218 144410 471454
rect 144646 471218 175130 471454
rect 175366 471218 205850 471454
rect 206086 471218 236570 471454
rect 236806 471218 267290 471454
rect 267526 471218 298010 471454
rect 298246 471218 328730 471454
rect 328966 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 414250 471454
rect 414486 471218 444970 471454
rect 445206 471218 475690 471454
rect 475926 471218 506410 471454
rect 506646 471218 537130 471454
rect 537366 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 52250 471134
rect 52486 470898 82970 471134
rect 83206 470898 113690 471134
rect 113926 470898 144410 471134
rect 144646 470898 175130 471134
rect 175366 470898 205850 471134
rect 206086 470898 236570 471134
rect 236806 470898 267290 471134
rect 267526 470898 298010 471134
rect 298246 470898 328730 471134
rect 328966 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 414250 471134
rect 414486 470898 444970 471134
rect 445206 470898 475690 471134
rect 475926 470898 506410 471134
rect 506646 470898 537130 471134
rect 537366 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 67610 439954
rect 67846 439718 98330 439954
rect 98566 439718 129050 439954
rect 129286 439718 159770 439954
rect 160006 439718 190490 439954
rect 190726 439718 221210 439954
rect 221446 439718 251930 439954
rect 252166 439718 282650 439954
rect 282886 439718 313370 439954
rect 313606 439718 344090 439954
rect 344326 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 429610 439954
rect 429846 439718 460330 439954
rect 460566 439718 491050 439954
rect 491286 439718 521770 439954
rect 522006 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 67610 439634
rect 67846 439398 98330 439634
rect 98566 439398 129050 439634
rect 129286 439398 159770 439634
rect 160006 439398 190490 439634
rect 190726 439398 221210 439634
rect 221446 439398 251930 439634
rect 252166 439398 282650 439634
rect 282886 439398 313370 439634
rect 313606 439398 344090 439634
rect 344326 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 429610 439634
rect 429846 439398 460330 439634
rect 460566 439398 491050 439634
rect 491286 439398 521770 439634
rect 522006 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 52250 435454
rect 52486 435218 82970 435454
rect 83206 435218 113690 435454
rect 113926 435218 144410 435454
rect 144646 435218 175130 435454
rect 175366 435218 205850 435454
rect 206086 435218 236570 435454
rect 236806 435218 267290 435454
rect 267526 435218 298010 435454
rect 298246 435218 328730 435454
rect 328966 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 414250 435454
rect 414486 435218 444970 435454
rect 445206 435218 475690 435454
rect 475926 435218 506410 435454
rect 506646 435218 537130 435454
rect 537366 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 52250 435134
rect 52486 434898 82970 435134
rect 83206 434898 113690 435134
rect 113926 434898 144410 435134
rect 144646 434898 175130 435134
rect 175366 434898 205850 435134
rect 206086 434898 236570 435134
rect 236806 434898 267290 435134
rect 267526 434898 298010 435134
rect 298246 434898 328730 435134
rect 328966 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 414250 435134
rect 414486 434898 444970 435134
rect 445206 434898 475690 435134
rect 475926 434898 506410 435134
rect 506646 434898 537130 435134
rect 537366 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 67610 403954
rect 67846 403718 98330 403954
rect 98566 403718 129050 403954
rect 129286 403718 159770 403954
rect 160006 403718 190490 403954
rect 190726 403718 221210 403954
rect 221446 403718 251930 403954
rect 252166 403718 282650 403954
rect 282886 403718 313370 403954
rect 313606 403718 344090 403954
rect 344326 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 429610 403954
rect 429846 403718 460330 403954
rect 460566 403718 491050 403954
rect 491286 403718 521770 403954
rect 522006 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 67610 403634
rect 67846 403398 98330 403634
rect 98566 403398 129050 403634
rect 129286 403398 159770 403634
rect 160006 403398 190490 403634
rect 190726 403398 221210 403634
rect 221446 403398 251930 403634
rect 252166 403398 282650 403634
rect 282886 403398 313370 403634
rect 313606 403398 344090 403634
rect 344326 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 429610 403634
rect 429846 403398 460330 403634
rect 460566 403398 491050 403634
rect 491286 403398 521770 403634
rect 522006 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 52250 399454
rect 52486 399218 82970 399454
rect 83206 399218 113690 399454
rect 113926 399218 144410 399454
rect 144646 399218 175130 399454
rect 175366 399218 205850 399454
rect 206086 399218 236570 399454
rect 236806 399218 267290 399454
rect 267526 399218 298010 399454
rect 298246 399218 328730 399454
rect 328966 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 414250 399454
rect 414486 399218 444970 399454
rect 445206 399218 475690 399454
rect 475926 399218 506410 399454
rect 506646 399218 537130 399454
rect 537366 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 52250 399134
rect 52486 398898 82970 399134
rect 83206 398898 113690 399134
rect 113926 398898 144410 399134
rect 144646 398898 175130 399134
rect 175366 398898 205850 399134
rect 206086 398898 236570 399134
rect 236806 398898 267290 399134
rect 267526 398898 298010 399134
rect 298246 398898 328730 399134
rect 328966 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 414250 399134
rect 414486 398898 444970 399134
rect 445206 398898 475690 399134
rect 475926 398898 506410 399134
rect 506646 398898 537130 399134
rect 537366 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 67610 367954
rect 67846 367718 98330 367954
rect 98566 367718 129050 367954
rect 129286 367718 159770 367954
rect 160006 367718 190490 367954
rect 190726 367718 221210 367954
rect 221446 367718 251930 367954
rect 252166 367718 282650 367954
rect 282886 367718 313370 367954
rect 313606 367718 344090 367954
rect 344326 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 429610 367954
rect 429846 367718 460330 367954
rect 460566 367718 491050 367954
rect 491286 367718 521770 367954
rect 522006 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 67610 367634
rect 67846 367398 98330 367634
rect 98566 367398 129050 367634
rect 129286 367398 159770 367634
rect 160006 367398 190490 367634
rect 190726 367398 221210 367634
rect 221446 367398 251930 367634
rect 252166 367398 282650 367634
rect 282886 367398 313370 367634
rect 313606 367398 344090 367634
rect 344326 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 429610 367634
rect 429846 367398 460330 367634
rect 460566 367398 491050 367634
rect 491286 367398 521770 367634
rect 522006 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 52250 363454
rect 52486 363218 82970 363454
rect 83206 363218 113690 363454
rect 113926 363218 144410 363454
rect 144646 363218 175130 363454
rect 175366 363218 205850 363454
rect 206086 363218 236570 363454
rect 236806 363218 267290 363454
rect 267526 363218 298010 363454
rect 298246 363218 328730 363454
rect 328966 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 414250 363454
rect 414486 363218 444970 363454
rect 445206 363218 475690 363454
rect 475926 363218 506410 363454
rect 506646 363218 537130 363454
rect 537366 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 52250 363134
rect 52486 362898 82970 363134
rect 83206 362898 113690 363134
rect 113926 362898 144410 363134
rect 144646 362898 175130 363134
rect 175366 362898 205850 363134
rect 206086 362898 236570 363134
rect 236806 362898 267290 363134
rect 267526 362898 298010 363134
rect 298246 362898 328730 363134
rect 328966 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 414250 363134
rect 414486 362898 444970 363134
rect 445206 362898 475690 363134
rect 475926 362898 506410 363134
rect 506646 362898 537130 363134
rect 537366 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 67610 331954
rect 67846 331718 98330 331954
rect 98566 331718 129050 331954
rect 129286 331718 159770 331954
rect 160006 331718 190490 331954
rect 190726 331718 221210 331954
rect 221446 331718 251930 331954
rect 252166 331718 282650 331954
rect 282886 331718 313370 331954
rect 313606 331718 344090 331954
rect 344326 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 429610 331954
rect 429846 331718 460330 331954
rect 460566 331718 491050 331954
rect 491286 331718 521770 331954
rect 522006 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 67610 331634
rect 67846 331398 98330 331634
rect 98566 331398 129050 331634
rect 129286 331398 159770 331634
rect 160006 331398 190490 331634
rect 190726 331398 221210 331634
rect 221446 331398 251930 331634
rect 252166 331398 282650 331634
rect 282886 331398 313370 331634
rect 313606 331398 344090 331634
rect 344326 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 429610 331634
rect 429846 331398 460330 331634
rect 460566 331398 491050 331634
rect 491286 331398 521770 331634
rect 522006 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 52250 327454
rect 52486 327218 82970 327454
rect 83206 327218 113690 327454
rect 113926 327218 144410 327454
rect 144646 327218 175130 327454
rect 175366 327218 205850 327454
rect 206086 327218 236570 327454
rect 236806 327218 267290 327454
rect 267526 327218 298010 327454
rect 298246 327218 328730 327454
rect 328966 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 414250 327454
rect 414486 327218 444970 327454
rect 445206 327218 475690 327454
rect 475926 327218 506410 327454
rect 506646 327218 537130 327454
rect 537366 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 52250 327134
rect 52486 326898 82970 327134
rect 83206 326898 113690 327134
rect 113926 326898 144410 327134
rect 144646 326898 175130 327134
rect 175366 326898 205850 327134
rect 206086 326898 236570 327134
rect 236806 326898 267290 327134
rect 267526 326898 298010 327134
rect 298246 326898 328730 327134
rect 328966 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 414250 327134
rect 414486 326898 444970 327134
rect 445206 326898 475690 327134
rect 475926 326898 506410 327134
rect 506646 326898 537130 327134
rect 537366 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 67610 295954
rect 67846 295718 98330 295954
rect 98566 295718 129050 295954
rect 129286 295718 159770 295954
rect 160006 295718 190490 295954
rect 190726 295718 221210 295954
rect 221446 295718 251930 295954
rect 252166 295718 282650 295954
rect 282886 295718 313370 295954
rect 313606 295718 344090 295954
rect 344326 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 429610 295954
rect 429846 295718 460330 295954
rect 460566 295718 491050 295954
rect 491286 295718 521770 295954
rect 522006 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 67610 295634
rect 67846 295398 98330 295634
rect 98566 295398 129050 295634
rect 129286 295398 159770 295634
rect 160006 295398 190490 295634
rect 190726 295398 221210 295634
rect 221446 295398 251930 295634
rect 252166 295398 282650 295634
rect 282886 295398 313370 295634
rect 313606 295398 344090 295634
rect 344326 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 429610 295634
rect 429846 295398 460330 295634
rect 460566 295398 491050 295634
rect 491286 295398 521770 295634
rect 522006 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 52250 291454
rect 52486 291218 82970 291454
rect 83206 291218 113690 291454
rect 113926 291218 144410 291454
rect 144646 291218 175130 291454
rect 175366 291218 205850 291454
rect 206086 291218 236570 291454
rect 236806 291218 267290 291454
rect 267526 291218 298010 291454
rect 298246 291218 328730 291454
rect 328966 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 414250 291454
rect 414486 291218 444970 291454
rect 445206 291218 475690 291454
rect 475926 291218 506410 291454
rect 506646 291218 537130 291454
rect 537366 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 52250 291134
rect 52486 290898 82970 291134
rect 83206 290898 113690 291134
rect 113926 290898 144410 291134
rect 144646 290898 175130 291134
rect 175366 290898 205850 291134
rect 206086 290898 236570 291134
rect 236806 290898 267290 291134
rect 267526 290898 298010 291134
rect 298246 290898 328730 291134
rect 328966 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 414250 291134
rect 414486 290898 444970 291134
rect 445206 290898 475690 291134
rect 475926 290898 506410 291134
rect 506646 290898 537130 291134
rect 537366 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 67610 259954
rect 67846 259718 98330 259954
rect 98566 259718 129050 259954
rect 129286 259718 159770 259954
rect 160006 259718 190490 259954
rect 190726 259718 221210 259954
rect 221446 259718 251930 259954
rect 252166 259718 282650 259954
rect 282886 259718 313370 259954
rect 313606 259718 344090 259954
rect 344326 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 429610 259954
rect 429846 259718 460330 259954
rect 460566 259718 491050 259954
rect 491286 259718 521770 259954
rect 522006 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 67610 259634
rect 67846 259398 98330 259634
rect 98566 259398 129050 259634
rect 129286 259398 159770 259634
rect 160006 259398 190490 259634
rect 190726 259398 221210 259634
rect 221446 259398 251930 259634
rect 252166 259398 282650 259634
rect 282886 259398 313370 259634
rect 313606 259398 344090 259634
rect 344326 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 429610 259634
rect 429846 259398 460330 259634
rect 460566 259398 491050 259634
rect 491286 259398 521770 259634
rect 522006 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 52250 255454
rect 52486 255218 82970 255454
rect 83206 255218 113690 255454
rect 113926 255218 144410 255454
rect 144646 255218 175130 255454
rect 175366 255218 205850 255454
rect 206086 255218 236570 255454
rect 236806 255218 267290 255454
rect 267526 255218 298010 255454
rect 298246 255218 328730 255454
rect 328966 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 414250 255454
rect 414486 255218 444970 255454
rect 445206 255218 475690 255454
rect 475926 255218 506410 255454
rect 506646 255218 537130 255454
rect 537366 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 52250 255134
rect 52486 254898 82970 255134
rect 83206 254898 113690 255134
rect 113926 254898 144410 255134
rect 144646 254898 175130 255134
rect 175366 254898 205850 255134
rect 206086 254898 236570 255134
rect 236806 254898 267290 255134
rect 267526 254898 298010 255134
rect 298246 254898 328730 255134
rect 328966 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 414250 255134
rect 414486 254898 444970 255134
rect 445206 254898 475690 255134
rect 475926 254898 506410 255134
rect 506646 254898 537130 255134
rect 537366 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 67610 223954
rect 67846 223718 98330 223954
rect 98566 223718 129050 223954
rect 129286 223718 159770 223954
rect 160006 223718 190490 223954
rect 190726 223718 221210 223954
rect 221446 223718 251930 223954
rect 252166 223718 282650 223954
rect 282886 223718 313370 223954
rect 313606 223718 344090 223954
rect 344326 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 67610 223634
rect 67846 223398 98330 223634
rect 98566 223398 129050 223634
rect 129286 223398 159770 223634
rect 160006 223398 190490 223634
rect 190726 223398 221210 223634
rect 221446 223398 251930 223634
rect 252166 223398 282650 223634
rect 282886 223398 313370 223634
rect 313606 223398 344090 223634
rect 344326 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 52250 219454
rect 52486 219218 82970 219454
rect 83206 219218 113690 219454
rect 113926 219218 144410 219454
rect 144646 219218 175130 219454
rect 175366 219218 205850 219454
rect 206086 219218 236570 219454
rect 236806 219218 267290 219454
rect 267526 219218 298010 219454
rect 298246 219218 328730 219454
rect 328966 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 52250 219134
rect 52486 218898 82970 219134
rect 83206 218898 113690 219134
rect 113926 218898 144410 219134
rect 144646 218898 175130 219134
rect 175366 218898 205850 219134
rect 206086 218898 236570 219134
rect 236806 218898 267290 219134
rect 267526 218898 298010 219134
rect 298246 218898 328730 219134
rect 328966 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 248570 147454
rect 248806 147218 279290 147454
rect 279526 147218 310010 147454
rect 310246 147218 340730 147454
rect 340966 147218 371450 147454
rect 371686 147218 402170 147454
rect 402406 147218 432890 147454
rect 433126 147218 463610 147454
rect 463846 147218 494330 147454
rect 494566 147218 525050 147454
rect 525286 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 248570 147134
rect 248806 146898 279290 147134
rect 279526 146898 310010 147134
rect 310246 146898 340730 147134
rect 340966 146898 371450 147134
rect 371686 146898 402170 147134
rect 402406 146898 432890 147134
rect 433126 146898 463610 147134
rect 463846 146898 494330 147134
rect 494566 146898 525050 147134
rect 525286 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 79610 115954
rect 79846 115718 110330 115954
rect 110566 115718 141050 115954
rect 141286 115718 171770 115954
rect 172006 115718 202490 115954
rect 202726 115718 233210 115954
rect 233446 115718 263930 115954
rect 264166 115718 294650 115954
rect 294886 115718 325370 115954
rect 325606 115718 356090 115954
rect 356326 115718 386810 115954
rect 387046 115718 417530 115954
rect 417766 115718 448250 115954
rect 448486 115718 478970 115954
rect 479206 115718 509690 115954
rect 509926 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 79610 115634
rect 79846 115398 110330 115634
rect 110566 115398 141050 115634
rect 141286 115398 171770 115634
rect 172006 115398 202490 115634
rect 202726 115398 233210 115634
rect 233446 115398 263930 115634
rect 264166 115398 294650 115634
rect 294886 115398 325370 115634
rect 325606 115398 356090 115634
rect 356326 115398 386810 115634
rect 387046 115398 417530 115634
rect 417766 115398 448250 115634
rect 448486 115398 478970 115634
rect 479206 115398 509690 115634
rect 509926 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 248570 111454
rect 248806 111218 279290 111454
rect 279526 111218 310010 111454
rect 310246 111218 340730 111454
rect 340966 111218 371450 111454
rect 371686 111218 402170 111454
rect 402406 111218 432890 111454
rect 433126 111218 463610 111454
rect 463846 111218 494330 111454
rect 494566 111218 525050 111454
rect 525286 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 248570 111134
rect 248806 110898 279290 111134
rect 279526 110898 310010 111134
rect 310246 110898 340730 111134
rect 340966 110898 371450 111134
rect 371686 110898 402170 111134
rect 402406 110898 432890 111134
rect 433126 110898 463610 111134
rect 463846 110898 494330 111134
rect 494566 110898 525050 111134
rect 525286 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 79610 79954
rect 79846 79718 110330 79954
rect 110566 79718 141050 79954
rect 141286 79718 171770 79954
rect 172006 79718 202490 79954
rect 202726 79718 233210 79954
rect 233446 79718 263930 79954
rect 264166 79718 294650 79954
rect 294886 79718 325370 79954
rect 325606 79718 356090 79954
rect 356326 79718 386810 79954
rect 387046 79718 417530 79954
rect 417766 79718 448250 79954
rect 448486 79718 478970 79954
rect 479206 79718 509690 79954
rect 509926 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 79610 79634
rect 79846 79398 110330 79634
rect 110566 79398 141050 79634
rect 141286 79398 171770 79634
rect 172006 79398 202490 79634
rect 202726 79398 233210 79634
rect 233446 79398 263930 79634
rect 264166 79398 294650 79634
rect 294886 79398 325370 79634
rect 325606 79398 356090 79634
rect 356326 79398 386810 79634
rect 387046 79398 417530 79634
rect 417766 79398 448250 79634
rect 448486 79398 478970 79634
rect 479206 79398 509690 79634
rect 509926 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 248570 75454
rect 248806 75218 279290 75454
rect 279526 75218 310010 75454
rect 310246 75218 340730 75454
rect 340966 75218 371450 75454
rect 371686 75218 402170 75454
rect 402406 75218 432890 75454
rect 433126 75218 463610 75454
rect 463846 75218 494330 75454
rect 494566 75218 525050 75454
rect 525286 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 248570 75134
rect 248806 74898 279290 75134
rect 279526 74898 310010 75134
rect 310246 74898 340730 75134
rect 340966 74898 371450 75134
rect 371686 74898 402170 75134
rect 402406 74898 432890 75134
rect 433126 74898 463610 75134
rect 463846 74898 494330 75134
rect 494566 74898 525050 75134
rect 525286 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 79610 43954
rect 79846 43718 110330 43954
rect 110566 43718 141050 43954
rect 141286 43718 171770 43954
rect 172006 43718 202490 43954
rect 202726 43718 233210 43954
rect 233446 43718 263930 43954
rect 264166 43718 294650 43954
rect 294886 43718 325370 43954
rect 325606 43718 356090 43954
rect 356326 43718 386810 43954
rect 387046 43718 417530 43954
rect 417766 43718 448250 43954
rect 448486 43718 478970 43954
rect 479206 43718 509690 43954
rect 509926 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 79610 43634
rect 79846 43398 110330 43634
rect 110566 43398 141050 43634
rect 141286 43398 171770 43634
rect 172006 43398 202490 43634
rect 202726 43398 233210 43634
rect 233446 43398 263930 43634
rect 264166 43398 294650 43634
rect 294886 43398 325370 43634
rect 325606 43398 356090 43634
rect 356326 43398 386810 43634
rect 387046 43398 417530 43634
rect 417766 43398 448250 43634
rect 448486 43398 478970 43634
rect 479206 43398 509690 43634
rect 509926 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 64250 39454
rect 64486 39218 94970 39454
rect 95206 39218 125690 39454
rect 125926 39218 156410 39454
rect 156646 39218 187130 39454
rect 187366 39218 217850 39454
rect 218086 39218 248570 39454
rect 248806 39218 279290 39454
rect 279526 39218 310010 39454
rect 310246 39218 340730 39454
rect 340966 39218 371450 39454
rect 371686 39218 402170 39454
rect 402406 39218 432890 39454
rect 433126 39218 463610 39454
rect 463846 39218 494330 39454
rect 494566 39218 525050 39454
rect 525286 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 64250 39134
rect 64486 38898 94970 39134
rect 95206 38898 125690 39134
rect 125926 38898 156410 39134
rect 156646 38898 187130 39134
rect 187366 38898 217850 39134
rect 218086 38898 248570 39134
rect 248806 38898 279290 39134
rect 279526 38898 310010 39134
rect 310246 38898 340730 39134
rect 340966 38898 371450 39134
rect 371686 38898 402170 39134
rect 402406 38898 432890 39134
rect 433126 38898 463610 39134
rect 463846 38898 494330 39134
rect 494566 38898 525050 39134
rect 525286 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use axi_node_intf_wrap  axi_interconnect_i
timestamp 0
transform 1 0 60000 0 1 30000
box 0 0 480000 120000
use mba_core_region  core_region_i
timestamp 0
transform 1 0 48000 0 1 200000
box 0 0 300000 360000
use sky130_sram_2kbyte_1rw1r_32x512_8  data_ram
timestamp 0
transform 1 0 210000 0 1 590000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_ram
timestamp 0
transform 1 0 36000 0 1 590000
box 0 0 136620 83308
use peripherals  peripherals_i
timestamp 0
transform 1 0 410000 0 1 240000
box 0 0 140000 440000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 588000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 675308 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 675308 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 675308 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 675308 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 562000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 675308 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 675308 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 675308 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 675308 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 152000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 152000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 152000 434414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 682000 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 152000 470414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 682000 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 152000 506414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 682000 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 152000 542414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 682000 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 675308 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 152000 83414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 675308 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 152000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 675308 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 152000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 675308 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 152000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 562000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 152000 227414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 675308 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 152000 263414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 675308 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 152000 299414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 675308 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 152000 335414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 675308 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 152000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 152000 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 152000 443414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 682000 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 152000 479414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 682000 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 152000 515414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 682000 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 682000 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 198000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 562000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 152000 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 152000 416414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 152000 452414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 152000 488414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 152000 524414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 675308 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 675308 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 675308 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 675308 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 675308 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 675308 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 675308 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 675308 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 152000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 152000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 152000 425414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 152000 461414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 152000 497414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 152000 533414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 562000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 152000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 152000 420914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 152000 456914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 152000 492914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 152000 528914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 675308 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 675308 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 675308 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 562000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 675308 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 675308 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 675308 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 675308 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 152000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 152000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 152000 429914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 682000 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 152000 465914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 682000 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 152000 501914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 682000 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 152000 537914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 682000 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 588000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 675308 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 675308 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 675308 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 675308 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 562000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 675308 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 675308 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 675308 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 675308 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 152000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 152000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 152000 438914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 682000 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 152000 474914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 682000 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 152000 510914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 682000 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 682000 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 675308 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 152000 87914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 675308 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 152000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 675308 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 152000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 675308 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 152000 195914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 562000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 152000 231914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 675308 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 152000 267914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 675308 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 152000 303914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 675308 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 152000 339914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 675308 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 152000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 152000 411914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 682000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 152000 447914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 682000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 152000 483914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 682000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 152000 519914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 682000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
