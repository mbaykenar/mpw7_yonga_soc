* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for axi_node_intf_wrap abstract view
.subckt axi_node_intf_wrap clk m00_ar_addr[0] m00_ar_addr[10] m00_ar_addr[11] m00_ar_addr[12]
+ m00_ar_addr[13] m00_ar_addr[14] m00_ar_addr[15] m00_ar_addr[16] m00_ar_addr[17]
+ m00_ar_addr[18] m00_ar_addr[19] m00_ar_addr[1] m00_ar_addr[20] m00_ar_addr[21] m00_ar_addr[22]
+ m00_ar_addr[23] m00_ar_addr[24] m00_ar_addr[25] m00_ar_addr[26] m00_ar_addr[27]
+ m00_ar_addr[28] m00_ar_addr[29] m00_ar_addr[2] m00_ar_addr[30] m00_ar_addr[31] m00_ar_addr[3]
+ m00_ar_addr[4] m00_ar_addr[5] m00_ar_addr[6] m00_ar_addr[7] m00_ar_addr[8] m00_ar_addr[9]
+ m00_ar_burst[0] m00_ar_burst[1] m00_ar_cache[0] m00_ar_cache[1] m00_ar_cache[2]
+ m00_ar_cache[3] m00_ar_id[0] m00_ar_id[10] m00_ar_id[11] m00_ar_id[1] m00_ar_id[2]
+ m00_ar_id[3] m00_ar_id[4] m00_ar_id[5] m00_ar_id[6] m00_ar_id[7] m00_ar_id[8] m00_ar_id[9]
+ m00_ar_len[0] m00_ar_len[1] m00_ar_len[2] m00_ar_len[3] m00_ar_len[4] m00_ar_len[5]
+ m00_ar_len[6] m00_ar_len[7] m00_ar_lock m00_ar_prot[0] m00_ar_prot[1] m00_ar_prot[2]
+ m00_ar_qos[0] m00_ar_qos[1] m00_ar_qos[2] m00_ar_qos[3] m00_ar_ready m00_ar_region[0]
+ m00_ar_region[1] m00_ar_region[2] m00_ar_region[3] m00_ar_size[0] m00_ar_size[1]
+ m00_ar_size[2] m00_ar_user[-1] m00_ar_user[0] m00_ar_valid m00_aw_addr[0] m00_aw_addr[10]
+ m00_aw_addr[11] m00_aw_addr[12] m00_aw_addr[13] m00_aw_addr[14] m00_aw_addr[15]
+ m00_aw_addr[16] m00_aw_addr[17] m00_aw_addr[18] m00_aw_addr[19] m00_aw_addr[1] m00_aw_addr[20]
+ m00_aw_addr[21] m00_aw_addr[22] m00_aw_addr[23] m00_aw_addr[24] m00_aw_addr[25]
+ m00_aw_addr[26] m00_aw_addr[27] m00_aw_addr[28] m00_aw_addr[29] m00_aw_addr[2] m00_aw_addr[30]
+ m00_aw_addr[31] m00_aw_addr[3] m00_aw_addr[4] m00_aw_addr[5] m00_aw_addr[6] m00_aw_addr[7]
+ m00_aw_addr[8] m00_aw_addr[9] m00_aw_burst[0] m00_aw_burst[1] m00_aw_cache[0] m00_aw_cache[1]
+ m00_aw_cache[2] m00_aw_cache[3] m00_aw_id[0] m00_aw_id[10] m00_aw_id[11] m00_aw_id[1]
+ m00_aw_id[2] m00_aw_id[3] m00_aw_id[4] m00_aw_id[5] m00_aw_id[6] m00_aw_id[7] m00_aw_id[8]
+ m00_aw_id[9] m00_aw_len[0] m00_aw_len[1] m00_aw_len[2] m00_aw_len[3] m00_aw_len[4]
+ m00_aw_len[5] m00_aw_len[6] m00_aw_len[7] m00_aw_lock m00_aw_prot[0] m00_aw_prot[1]
+ m00_aw_prot[2] m00_aw_qos[0] m00_aw_qos[1] m00_aw_qos[2] m00_aw_qos[3] m00_aw_ready
+ m00_aw_region[0] m00_aw_region[1] m00_aw_region[2] m00_aw_region[3] m00_aw_size[0]
+ m00_aw_size[1] m00_aw_size[2] m00_aw_user[-1] m00_aw_user[0] m00_aw_valid m00_b_id[0]
+ m00_b_id[10] m00_b_id[11] m00_b_id[1] m00_b_id[2] m00_b_id[3] m00_b_id[4] m00_b_id[5]
+ m00_b_id[6] m00_b_id[7] m00_b_id[8] m00_b_id[9] m00_b_ready m00_b_resp[0] m00_b_resp[1]
+ m00_b_user[-1] m00_b_user[0] m00_b_valid m00_r_data[0] m00_r_data[10] m00_r_data[11]
+ m00_r_data[12] m00_r_data[13] m00_r_data[14] m00_r_data[15] m00_r_data[16] m00_r_data[17]
+ m00_r_data[18] m00_r_data[19] m00_r_data[1] m00_r_data[20] m00_r_data[21] m00_r_data[22]
+ m00_r_data[23] m00_r_data[24] m00_r_data[25] m00_r_data[26] m00_r_data[27] m00_r_data[28]
+ m00_r_data[29] m00_r_data[2] m00_r_data[30] m00_r_data[31] m00_r_data[3] m00_r_data[4]
+ m00_r_data[5] m00_r_data[6] m00_r_data[7] m00_r_data[8] m00_r_data[9] m00_r_id[0]
+ m00_r_id[10] m00_r_id[11] m00_r_id[1] m00_r_id[2] m00_r_id[3] m00_r_id[4] m00_r_id[5]
+ m00_r_id[6] m00_r_id[7] m00_r_id[8] m00_r_id[9] m00_r_last m00_r_ready m00_r_resp[0]
+ m00_r_resp[1] m00_r_user[-1] m00_r_user[0] m00_r_valid m00_w_data[0] m00_w_data[10]
+ m00_w_data[11] m00_w_data[12] m00_w_data[13] m00_w_data[14] m00_w_data[15] m00_w_data[16]
+ m00_w_data[17] m00_w_data[18] m00_w_data[19] m00_w_data[1] m00_w_data[20] m00_w_data[21]
+ m00_w_data[22] m00_w_data[23] m00_w_data[24] m00_w_data[25] m00_w_data[26] m00_w_data[27]
+ m00_w_data[28] m00_w_data[29] m00_w_data[2] m00_w_data[30] m00_w_data[31] m00_w_data[3]
+ m00_w_data[4] m00_w_data[5] m00_w_data[6] m00_w_data[7] m00_w_data[8] m00_w_data[9]
+ m00_w_last m00_w_ready m00_w_strb[0] m00_w_strb[1] m00_w_strb[2] m00_w_strb[3] m00_w_user[-1]
+ m00_w_user[0] m00_w_valid m01_ar_addr[0] m01_ar_addr[10] m01_ar_addr[11] m01_ar_addr[12]
+ m01_ar_addr[13] m01_ar_addr[14] m01_ar_addr[15] m01_ar_addr[16] m01_ar_addr[17]
+ m01_ar_addr[18] m01_ar_addr[19] m01_ar_addr[1] m01_ar_addr[20] m01_ar_addr[21] m01_ar_addr[22]
+ m01_ar_addr[23] m01_ar_addr[24] m01_ar_addr[25] m01_ar_addr[26] m01_ar_addr[27]
+ m01_ar_addr[28] m01_ar_addr[29] m01_ar_addr[2] m01_ar_addr[30] m01_ar_addr[31] m01_ar_addr[3]
+ m01_ar_addr[4] m01_ar_addr[5] m01_ar_addr[6] m01_ar_addr[7] m01_ar_addr[8] m01_ar_addr[9]
+ m01_ar_burst[0] m01_ar_burst[1] m01_ar_cache[0] m01_ar_cache[1] m01_ar_cache[2]
+ m01_ar_cache[3] m01_ar_id[0] m01_ar_id[10] m01_ar_id[11] m01_ar_id[1] m01_ar_id[2]
+ m01_ar_id[3] m01_ar_id[4] m01_ar_id[5] m01_ar_id[6] m01_ar_id[7] m01_ar_id[8] m01_ar_id[9]
+ m01_ar_len[0] m01_ar_len[1] m01_ar_len[2] m01_ar_len[3] m01_ar_len[4] m01_ar_len[5]
+ m01_ar_len[6] m01_ar_len[7] m01_ar_lock m01_ar_prot[0] m01_ar_prot[1] m01_ar_prot[2]
+ m01_ar_qos[0] m01_ar_qos[1] m01_ar_qos[2] m01_ar_qos[3] m01_ar_ready m01_ar_region[0]
+ m01_ar_region[1] m01_ar_region[2] m01_ar_region[3] m01_ar_size[0] m01_ar_size[1]
+ m01_ar_size[2] m01_ar_user[-1] m01_ar_user[0] m01_ar_valid m01_aw_addr[0] m01_aw_addr[10]
+ m01_aw_addr[11] m01_aw_addr[12] m01_aw_addr[13] m01_aw_addr[14] m01_aw_addr[15]
+ m01_aw_addr[16] m01_aw_addr[17] m01_aw_addr[18] m01_aw_addr[19] m01_aw_addr[1] m01_aw_addr[20]
+ m01_aw_addr[21] m01_aw_addr[22] m01_aw_addr[23] m01_aw_addr[24] m01_aw_addr[25]
+ m01_aw_addr[26] m01_aw_addr[27] m01_aw_addr[28] m01_aw_addr[29] m01_aw_addr[2] m01_aw_addr[30]
+ m01_aw_addr[31] m01_aw_addr[3] m01_aw_addr[4] m01_aw_addr[5] m01_aw_addr[6] m01_aw_addr[7]
+ m01_aw_addr[8] m01_aw_addr[9] m01_aw_burst[0] m01_aw_burst[1] m01_aw_cache[0] m01_aw_cache[1]
+ m01_aw_cache[2] m01_aw_cache[3] m01_aw_id[0] m01_aw_id[10] m01_aw_id[11] m01_aw_id[1]
+ m01_aw_id[2] m01_aw_id[3] m01_aw_id[4] m01_aw_id[5] m01_aw_id[6] m01_aw_id[7] m01_aw_id[8]
+ m01_aw_id[9] m01_aw_len[0] m01_aw_len[1] m01_aw_len[2] m01_aw_len[3] m01_aw_len[4]
+ m01_aw_len[5] m01_aw_len[6] m01_aw_len[7] m01_aw_lock m01_aw_prot[0] m01_aw_prot[1]
+ m01_aw_prot[2] m01_aw_qos[0] m01_aw_qos[1] m01_aw_qos[2] m01_aw_qos[3] m01_aw_ready
+ m01_aw_region[0] m01_aw_region[1] m01_aw_region[2] m01_aw_region[3] m01_aw_size[0]
+ m01_aw_size[1] m01_aw_size[2] m01_aw_user[-1] m01_aw_user[0] m01_aw_valid m01_b_id[0]
+ m01_b_id[10] m01_b_id[11] m01_b_id[1] m01_b_id[2] m01_b_id[3] m01_b_id[4] m01_b_id[5]
+ m01_b_id[6] m01_b_id[7] m01_b_id[8] m01_b_id[9] m01_b_ready m01_b_resp[0] m01_b_resp[1]
+ m01_b_user[-1] m01_b_user[0] m01_b_valid m01_r_data[0] m01_r_data[10] m01_r_data[11]
+ m01_r_data[12] m01_r_data[13] m01_r_data[14] m01_r_data[15] m01_r_data[16] m01_r_data[17]
+ m01_r_data[18] m01_r_data[19] m01_r_data[1] m01_r_data[20] m01_r_data[21] m01_r_data[22]
+ m01_r_data[23] m01_r_data[24] m01_r_data[25] m01_r_data[26] m01_r_data[27] m01_r_data[28]
+ m01_r_data[29] m01_r_data[2] m01_r_data[30] m01_r_data[31] m01_r_data[3] m01_r_data[4]
+ m01_r_data[5] m01_r_data[6] m01_r_data[7] m01_r_data[8] m01_r_data[9] m01_r_id[0]
+ m01_r_id[10] m01_r_id[11] m01_r_id[1] m01_r_id[2] m01_r_id[3] m01_r_id[4] m01_r_id[5]
+ m01_r_id[6] m01_r_id[7] m01_r_id[8] m01_r_id[9] m01_r_last m01_r_ready m01_r_resp[0]
+ m01_r_resp[1] m01_r_user[-1] m01_r_user[0] m01_r_valid m01_w_data[0] m01_w_data[10]
+ m01_w_data[11] m01_w_data[12] m01_w_data[13] m01_w_data[14] m01_w_data[15] m01_w_data[16]
+ m01_w_data[17] m01_w_data[18] m01_w_data[19] m01_w_data[1] m01_w_data[20] m01_w_data[21]
+ m01_w_data[22] m01_w_data[23] m01_w_data[24] m01_w_data[25] m01_w_data[26] m01_w_data[27]
+ m01_w_data[28] m01_w_data[29] m01_w_data[2] m01_w_data[30] m01_w_data[31] m01_w_data[3]
+ m01_w_data[4] m01_w_data[5] m01_w_data[6] m01_w_data[7] m01_w_data[8] m01_w_data[9]
+ m01_w_last m01_w_ready m01_w_strb[0] m01_w_strb[1] m01_w_strb[2] m01_w_strb[3] m01_w_user[-1]
+ m01_w_user[0] m01_w_valid m02_ar_addr[0] m02_ar_addr[10] m02_ar_addr[11] m02_ar_addr[12]
+ m02_ar_addr[13] m02_ar_addr[14] m02_ar_addr[15] m02_ar_addr[16] m02_ar_addr[17]
+ m02_ar_addr[18] m02_ar_addr[19] m02_ar_addr[1] m02_ar_addr[20] m02_ar_addr[21] m02_ar_addr[22]
+ m02_ar_addr[23] m02_ar_addr[24] m02_ar_addr[25] m02_ar_addr[26] m02_ar_addr[27]
+ m02_ar_addr[28] m02_ar_addr[29] m02_ar_addr[2] m02_ar_addr[30] m02_ar_addr[31] m02_ar_addr[3]
+ m02_ar_addr[4] m02_ar_addr[5] m02_ar_addr[6] m02_ar_addr[7] m02_ar_addr[8] m02_ar_addr[9]
+ m02_ar_burst[0] m02_ar_burst[1] m02_ar_cache[0] m02_ar_cache[1] m02_ar_cache[2]
+ m02_ar_cache[3] m02_ar_id[0] m02_ar_id[10] m02_ar_id[11] m02_ar_id[1] m02_ar_id[2]
+ m02_ar_id[3] m02_ar_id[4] m02_ar_id[5] m02_ar_id[6] m02_ar_id[7] m02_ar_id[8] m02_ar_id[9]
+ m02_ar_len[0] m02_ar_len[1] m02_ar_len[2] m02_ar_len[3] m02_ar_len[4] m02_ar_len[5]
+ m02_ar_len[6] m02_ar_len[7] m02_ar_lock m02_ar_prot[0] m02_ar_prot[1] m02_ar_prot[2]
+ m02_ar_qos[0] m02_ar_qos[1] m02_ar_qos[2] m02_ar_qos[3] m02_ar_ready m02_ar_region[0]
+ m02_ar_region[1] m02_ar_region[2] m02_ar_region[3] m02_ar_size[0] m02_ar_size[1]
+ m02_ar_size[2] m02_ar_user[-1] m02_ar_user[0] m02_ar_valid m02_aw_addr[0] m02_aw_addr[10]
+ m02_aw_addr[11] m02_aw_addr[12] m02_aw_addr[13] m02_aw_addr[14] m02_aw_addr[15]
+ m02_aw_addr[16] m02_aw_addr[17] m02_aw_addr[18] m02_aw_addr[19] m02_aw_addr[1] m02_aw_addr[20]
+ m02_aw_addr[21] m02_aw_addr[22] m02_aw_addr[23] m02_aw_addr[24] m02_aw_addr[25]
+ m02_aw_addr[26] m02_aw_addr[27] m02_aw_addr[28] m02_aw_addr[29] m02_aw_addr[2] m02_aw_addr[30]
+ m02_aw_addr[31] m02_aw_addr[3] m02_aw_addr[4] m02_aw_addr[5] m02_aw_addr[6] m02_aw_addr[7]
+ m02_aw_addr[8] m02_aw_addr[9] m02_aw_burst[0] m02_aw_burst[1] m02_aw_cache[0] m02_aw_cache[1]
+ m02_aw_cache[2] m02_aw_cache[3] m02_aw_id[0] m02_aw_id[10] m02_aw_id[11] m02_aw_id[1]
+ m02_aw_id[2] m02_aw_id[3] m02_aw_id[4] m02_aw_id[5] m02_aw_id[6] m02_aw_id[7] m02_aw_id[8]
+ m02_aw_id[9] m02_aw_len[0] m02_aw_len[1] m02_aw_len[2] m02_aw_len[3] m02_aw_len[4]
+ m02_aw_len[5] m02_aw_len[6] m02_aw_len[7] m02_aw_lock m02_aw_prot[0] m02_aw_prot[1]
+ m02_aw_prot[2] m02_aw_qos[0] m02_aw_qos[1] m02_aw_qos[2] m02_aw_qos[3] m02_aw_ready
+ m02_aw_region[0] m02_aw_region[1] m02_aw_region[2] m02_aw_region[3] m02_aw_size[0]
+ m02_aw_size[1] m02_aw_size[2] m02_aw_user[-1] m02_aw_user[0] m02_aw_valid m02_b_id[0]
+ m02_b_id[10] m02_b_id[11] m02_b_id[1] m02_b_id[2] m02_b_id[3] m02_b_id[4] m02_b_id[5]
+ m02_b_id[6] m02_b_id[7] m02_b_id[8] m02_b_id[9] m02_b_ready m02_b_resp[0] m02_b_resp[1]
+ m02_b_user[-1] m02_b_user[0] m02_b_valid m02_r_data[0] m02_r_data[10] m02_r_data[11]
+ m02_r_data[12] m02_r_data[13] m02_r_data[14] m02_r_data[15] m02_r_data[16] m02_r_data[17]
+ m02_r_data[18] m02_r_data[19] m02_r_data[1] m02_r_data[20] m02_r_data[21] m02_r_data[22]
+ m02_r_data[23] m02_r_data[24] m02_r_data[25] m02_r_data[26] m02_r_data[27] m02_r_data[28]
+ m02_r_data[29] m02_r_data[2] m02_r_data[30] m02_r_data[31] m02_r_data[3] m02_r_data[4]
+ m02_r_data[5] m02_r_data[6] m02_r_data[7] m02_r_data[8] m02_r_data[9] m02_r_id[0]
+ m02_r_id[10] m02_r_id[11] m02_r_id[1] m02_r_id[2] m02_r_id[3] m02_r_id[4] m02_r_id[5]
+ m02_r_id[6] m02_r_id[7] m02_r_id[8] m02_r_id[9] m02_r_last m02_r_ready m02_r_resp[0]
+ m02_r_resp[1] m02_r_user[-1] m02_r_user[0] m02_r_valid m02_w_data[0] m02_w_data[10]
+ m02_w_data[11] m02_w_data[12] m02_w_data[13] m02_w_data[14] m02_w_data[15] m02_w_data[16]
+ m02_w_data[17] m02_w_data[18] m02_w_data[19] m02_w_data[1] m02_w_data[20] m02_w_data[21]
+ m02_w_data[22] m02_w_data[23] m02_w_data[24] m02_w_data[25] m02_w_data[26] m02_w_data[27]
+ m02_w_data[28] m02_w_data[29] m02_w_data[2] m02_w_data[30] m02_w_data[31] m02_w_data[3]
+ m02_w_data[4] m02_w_data[5] m02_w_data[6] m02_w_data[7] m02_w_data[8] m02_w_data[9]
+ m02_w_last m02_w_ready m02_w_strb[0] m02_w_strb[1] m02_w_strb[2] m02_w_strb[3] m02_w_user[-1]
+ m02_w_user[0] m02_w_valid rst_n s00_ar_addr[0] s00_ar_addr[10] s00_ar_addr[11] s00_ar_addr[12]
+ s00_ar_addr[13] s00_ar_addr[14] s00_ar_addr[15] s00_ar_addr[16] s00_ar_addr[17]
+ s00_ar_addr[18] s00_ar_addr[19] s00_ar_addr[1] s00_ar_addr[20] s00_ar_addr[21] s00_ar_addr[22]
+ s00_ar_addr[23] s00_ar_addr[24] s00_ar_addr[25] s00_ar_addr[26] s00_ar_addr[27]
+ s00_ar_addr[28] s00_ar_addr[29] s00_ar_addr[2] s00_ar_addr[30] s00_ar_addr[31] s00_ar_addr[3]
+ s00_ar_addr[4] s00_ar_addr[5] s00_ar_addr[6] s00_ar_addr[7] s00_ar_addr[8] s00_ar_addr[9]
+ s00_ar_burst[0] s00_ar_burst[1] s00_ar_cache[0] s00_ar_cache[1] s00_ar_cache[2]
+ s00_ar_cache[3] s00_ar_id[0] s00_ar_id[1] s00_ar_id[2] s00_ar_id[3] s00_ar_id[4]
+ s00_ar_id[5] s00_ar_id[6] s00_ar_id[7] s00_ar_id[8] s00_ar_id[9] s00_ar_len[0] s00_ar_len[1]
+ s00_ar_len[2] s00_ar_len[3] s00_ar_len[4] s00_ar_len[5] s00_ar_len[6] s00_ar_len[7]
+ s00_ar_lock s00_ar_prot[0] s00_ar_prot[1] s00_ar_prot[2] s00_ar_qos[0] s00_ar_qos[1]
+ s00_ar_qos[2] s00_ar_qos[3] s00_ar_ready s00_ar_region[0] s00_ar_region[1] s00_ar_region[2]
+ s00_ar_region[3] s00_ar_size[0] s00_ar_size[1] s00_ar_size[2] s00_ar_user[-1] s00_ar_user[0]
+ s00_ar_valid s00_aw_addr[0] s00_aw_addr[10] s00_aw_addr[11] s00_aw_addr[12] s00_aw_addr[13]
+ s00_aw_addr[14] s00_aw_addr[15] s00_aw_addr[16] s00_aw_addr[17] s00_aw_addr[18]
+ s00_aw_addr[19] s00_aw_addr[1] s00_aw_addr[20] s00_aw_addr[21] s00_aw_addr[22] s00_aw_addr[23]
+ s00_aw_addr[24] s00_aw_addr[25] s00_aw_addr[26] s00_aw_addr[27] s00_aw_addr[28]
+ s00_aw_addr[29] s00_aw_addr[2] s00_aw_addr[30] s00_aw_addr[31] s00_aw_addr[3] s00_aw_addr[4]
+ s00_aw_addr[5] s00_aw_addr[6] s00_aw_addr[7] s00_aw_addr[8] s00_aw_addr[9] s00_aw_burst[0]
+ s00_aw_burst[1] s00_aw_cache[0] s00_aw_cache[1] s00_aw_cache[2] s00_aw_cache[3]
+ s00_aw_id[0] s00_aw_id[1] s00_aw_id[2] s00_aw_id[3] s00_aw_id[4] s00_aw_id[5] s00_aw_id[6]
+ s00_aw_id[7] s00_aw_id[8] s00_aw_id[9] s00_aw_len[0] s00_aw_len[1] s00_aw_len[2]
+ s00_aw_len[3] s00_aw_len[4] s00_aw_len[5] s00_aw_len[6] s00_aw_len[7] s00_aw_lock
+ s00_aw_prot[0] s00_aw_prot[1] s00_aw_prot[2] s00_aw_qos[0] s00_aw_qos[1] s00_aw_qos[2]
+ s00_aw_qos[3] s00_aw_ready s00_aw_region[0] s00_aw_region[1] s00_aw_region[2] s00_aw_region[3]
+ s00_aw_size[0] s00_aw_size[1] s00_aw_size[2] s00_aw_user[-1] s00_aw_user[0] s00_aw_valid
+ s00_b_id[0] s00_b_id[1] s00_b_id[2] s00_b_id[3] s00_b_id[4] s00_b_id[5] s00_b_id[6]
+ s00_b_id[7] s00_b_id[8] s00_b_id[9] s00_b_ready s00_b_resp[0] s00_b_resp[1] s00_b_user[-1]
+ s00_b_user[0] s00_b_valid s00_r_data[0] s00_r_data[10] s00_r_data[11] s00_r_data[12]
+ s00_r_data[13] s00_r_data[14] s00_r_data[15] s00_r_data[16] s00_r_data[17] s00_r_data[18]
+ s00_r_data[19] s00_r_data[1] s00_r_data[20] s00_r_data[21] s00_r_data[22] s00_r_data[23]
+ s00_r_data[24] s00_r_data[25] s00_r_data[26] s00_r_data[27] s00_r_data[28] s00_r_data[29]
+ s00_r_data[2] s00_r_data[30] s00_r_data[31] s00_r_data[3] s00_r_data[4] s00_r_data[5]
+ s00_r_data[6] s00_r_data[7] s00_r_data[8] s00_r_data[9] s00_r_id[0] s00_r_id[1]
+ s00_r_id[2] s00_r_id[3] s00_r_id[4] s00_r_id[5] s00_r_id[6] s00_r_id[7] s00_r_id[8]
+ s00_r_id[9] s00_r_last s00_r_ready s00_r_resp[0] s00_r_resp[1] s00_r_user[-1] s00_r_user[0]
+ s00_r_valid s00_w_data[0] s00_w_data[10] s00_w_data[11] s00_w_data[12] s00_w_data[13]
+ s00_w_data[14] s00_w_data[15] s00_w_data[16] s00_w_data[17] s00_w_data[18] s00_w_data[19]
+ s00_w_data[1] s00_w_data[20] s00_w_data[21] s00_w_data[22] s00_w_data[23] s00_w_data[24]
+ s00_w_data[25] s00_w_data[26] s00_w_data[27] s00_w_data[28] s00_w_data[29] s00_w_data[2]
+ s00_w_data[30] s00_w_data[31] s00_w_data[3] s00_w_data[4] s00_w_data[5] s00_w_data[6]
+ s00_w_data[7] s00_w_data[8] s00_w_data[9] s00_w_last s00_w_ready s00_w_strb[0] s00_w_strb[1]
+ s00_w_strb[2] s00_w_strb[3] s00_w_user[-1] s00_w_user[0] s00_w_valid s01_ar_addr[0]
+ s01_ar_addr[10] s01_ar_addr[11] s01_ar_addr[12] s01_ar_addr[13] s01_ar_addr[14]
+ s01_ar_addr[15] s01_ar_addr[16] s01_ar_addr[17] s01_ar_addr[18] s01_ar_addr[19]
+ s01_ar_addr[1] s01_ar_addr[20] s01_ar_addr[21] s01_ar_addr[22] s01_ar_addr[23] s01_ar_addr[24]
+ s01_ar_addr[25] s01_ar_addr[26] s01_ar_addr[27] s01_ar_addr[28] s01_ar_addr[29]
+ s01_ar_addr[2] s01_ar_addr[30] s01_ar_addr[31] s01_ar_addr[3] s01_ar_addr[4] s01_ar_addr[5]
+ s01_ar_addr[6] s01_ar_addr[7] s01_ar_addr[8] s01_ar_addr[9] s01_ar_burst[0] s01_ar_burst[1]
+ s01_ar_cache[0] s01_ar_cache[1] s01_ar_cache[2] s01_ar_cache[3] s01_ar_id[0] s01_ar_id[1]
+ s01_ar_id[2] s01_ar_id[3] s01_ar_id[4] s01_ar_id[5] s01_ar_id[6] s01_ar_id[7] s01_ar_id[8]
+ s01_ar_id[9] s01_ar_len[0] s01_ar_len[1] s01_ar_len[2] s01_ar_len[3] s01_ar_len[4]
+ s01_ar_len[5] s01_ar_len[6] s01_ar_len[7] s01_ar_lock s01_ar_prot[0] s01_ar_prot[1]
+ s01_ar_prot[2] s01_ar_qos[0] s01_ar_qos[1] s01_ar_qos[2] s01_ar_qos[3] s01_ar_ready
+ s01_ar_region[0] s01_ar_region[1] s01_ar_region[2] s01_ar_region[3] s01_ar_size[0]
+ s01_ar_size[1] s01_ar_size[2] s01_ar_user[-1] s01_ar_user[0] s01_ar_valid s01_aw_addr[0]
+ s01_aw_addr[10] s01_aw_addr[11] s01_aw_addr[12] s01_aw_addr[13] s01_aw_addr[14]
+ s01_aw_addr[15] s01_aw_addr[16] s01_aw_addr[17] s01_aw_addr[18] s01_aw_addr[19]
+ s01_aw_addr[1] s01_aw_addr[20] s01_aw_addr[21] s01_aw_addr[22] s01_aw_addr[23] s01_aw_addr[24]
+ s01_aw_addr[25] s01_aw_addr[26] s01_aw_addr[27] s01_aw_addr[28] s01_aw_addr[29]
+ s01_aw_addr[2] s01_aw_addr[30] s01_aw_addr[31] s01_aw_addr[3] s01_aw_addr[4] s01_aw_addr[5]
+ s01_aw_addr[6] s01_aw_addr[7] s01_aw_addr[8] s01_aw_addr[9] s01_aw_burst[0] s01_aw_burst[1]
+ s01_aw_cache[0] s01_aw_cache[1] s01_aw_cache[2] s01_aw_cache[3] s01_aw_id[0] s01_aw_id[1]
+ s01_aw_id[2] s01_aw_id[3] s01_aw_id[4] s01_aw_id[5] s01_aw_id[6] s01_aw_id[7] s01_aw_id[8]
+ s01_aw_id[9] s01_aw_len[0] s01_aw_len[1] s01_aw_len[2] s01_aw_len[3] s01_aw_len[4]
+ s01_aw_len[5] s01_aw_len[6] s01_aw_len[7] s01_aw_lock s01_aw_prot[0] s01_aw_prot[1]
+ s01_aw_prot[2] s01_aw_qos[0] s01_aw_qos[1] s01_aw_qos[2] s01_aw_qos[3] s01_aw_ready
+ s01_aw_region[0] s01_aw_region[1] s01_aw_region[2] s01_aw_region[3] s01_aw_size[0]
+ s01_aw_size[1] s01_aw_size[2] s01_aw_user[-1] s01_aw_user[0] s01_aw_valid s01_b_id[0]
+ s01_b_id[1] s01_b_id[2] s01_b_id[3] s01_b_id[4] s01_b_id[5] s01_b_id[6] s01_b_id[7]
+ s01_b_id[8] s01_b_id[9] s01_b_ready s01_b_resp[0] s01_b_resp[1] s01_b_user[-1] s01_b_user[0]
+ s01_b_valid s01_r_data[0] s01_r_data[10] s01_r_data[11] s01_r_data[12] s01_r_data[13]
+ s01_r_data[14] s01_r_data[15] s01_r_data[16] s01_r_data[17] s01_r_data[18] s01_r_data[19]
+ s01_r_data[1] s01_r_data[20] s01_r_data[21] s01_r_data[22] s01_r_data[23] s01_r_data[24]
+ s01_r_data[25] s01_r_data[26] s01_r_data[27] s01_r_data[28] s01_r_data[29] s01_r_data[2]
+ s01_r_data[30] s01_r_data[31] s01_r_data[3] s01_r_data[4] s01_r_data[5] s01_r_data[6]
+ s01_r_data[7] s01_r_data[8] s01_r_data[9] s01_r_id[0] s01_r_id[1] s01_r_id[2] s01_r_id[3]
+ s01_r_id[4] s01_r_id[5] s01_r_id[6] s01_r_id[7] s01_r_id[8] s01_r_id[9] s01_r_last
+ s01_r_ready s01_r_resp[0] s01_r_resp[1] s01_r_user[-1] s01_r_user[0] s01_r_valid
+ s01_w_data[0] s01_w_data[10] s01_w_data[11] s01_w_data[12] s01_w_data[13] s01_w_data[14]
+ s01_w_data[15] s01_w_data[16] s01_w_data[17] s01_w_data[18] s01_w_data[19] s01_w_data[1]
+ s01_w_data[20] s01_w_data[21] s01_w_data[22] s01_w_data[23] s01_w_data[24] s01_w_data[25]
+ s01_w_data[26] s01_w_data[27] s01_w_data[28] s01_w_data[29] s01_w_data[2] s01_w_data[30]
+ s01_w_data[31] s01_w_data[3] s01_w_data[4] s01_w_data[5] s01_w_data[6] s01_w_data[7]
+ s01_w_data[8] s01_w_data[9] s01_w_last s01_w_ready s01_w_strb[0] s01_w_strb[1] s01_w_strb[2]
+ s01_w_strb[3] s01_w_user[-1] s01_w_user[0] s01_w_valid s02_ar_addr[0] s02_ar_addr[10]
+ s02_ar_addr[11] s02_ar_addr[12] s02_ar_addr[13] s02_ar_addr[14] s02_ar_addr[15]
+ s02_ar_addr[16] s02_ar_addr[17] s02_ar_addr[18] s02_ar_addr[19] s02_ar_addr[1] s02_ar_addr[20]
+ s02_ar_addr[21] s02_ar_addr[22] s02_ar_addr[23] s02_ar_addr[24] s02_ar_addr[25]
+ s02_ar_addr[26] s02_ar_addr[27] s02_ar_addr[28] s02_ar_addr[29] s02_ar_addr[2] s02_ar_addr[30]
+ s02_ar_addr[31] s02_ar_addr[3] s02_ar_addr[4] s02_ar_addr[5] s02_ar_addr[6] s02_ar_addr[7]
+ s02_ar_addr[8] s02_ar_addr[9] s02_ar_burst[0] s02_ar_burst[1] s02_ar_cache[0] s02_ar_cache[1]
+ s02_ar_cache[2] s02_ar_cache[3] s02_ar_id[0] s02_ar_id[1] s02_ar_id[2] s02_ar_id[3]
+ s02_ar_id[4] s02_ar_id[5] s02_ar_id[6] s02_ar_id[7] s02_ar_id[8] s02_ar_id[9] s02_ar_len[0]
+ s02_ar_len[1] s02_ar_len[2] s02_ar_len[3] s02_ar_len[4] s02_ar_len[5] s02_ar_len[6]
+ s02_ar_len[7] s02_ar_lock s02_ar_prot[0] s02_ar_prot[1] s02_ar_prot[2] s02_ar_qos[0]
+ s02_ar_qos[1] s02_ar_qos[2] s02_ar_qos[3] s02_ar_ready s02_ar_region[0] s02_ar_region[1]
+ s02_ar_region[2] s02_ar_region[3] s02_ar_size[0] s02_ar_size[1] s02_ar_size[2] s02_ar_user[-1]
+ s02_ar_user[0] s02_ar_valid s02_aw_addr[0] s02_aw_addr[10] s02_aw_addr[11] s02_aw_addr[12]
+ s02_aw_addr[13] s02_aw_addr[14] s02_aw_addr[15] s02_aw_addr[16] s02_aw_addr[17]
+ s02_aw_addr[18] s02_aw_addr[19] s02_aw_addr[1] s02_aw_addr[20] s02_aw_addr[21] s02_aw_addr[22]
+ s02_aw_addr[23] s02_aw_addr[24] s02_aw_addr[25] s02_aw_addr[26] s02_aw_addr[27]
+ s02_aw_addr[28] s02_aw_addr[29] s02_aw_addr[2] s02_aw_addr[30] s02_aw_addr[31] s02_aw_addr[3]
+ s02_aw_addr[4] s02_aw_addr[5] s02_aw_addr[6] s02_aw_addr[7] s02_aw_addr[8] s02_aw_addr[9]
+ s02_aw_burst[0] s02_aw_burst[1] s02_aw_cache[0] s02_aw_cache[1] s02_aw_cache[2]
+ s02_aw_cache[3] s02_aw_id[0] s02_aw_id[1] s02_aw_id[2] s02_aw_id[3] s02_aw_id[4]
+ s02_aw_id[5] s02_aw_id[6] s02_aw_id[7] s02_aw_id[8] s02_aw_id[9] s02_aw_len[0] s02_aw_len[1]
+ s02_aw_len[2] s02_aw_len[3] s02_aw_len[4] s02_aw_len[5] s02_aw_len[6] s02_aw_len[7]
+ s02_aw_lock s02_aw_prot[0] s02_aw_prot[1] s02_aw_prot[2] s02_aw_qos[0] s02_aw_qos[1]
+ s02_aw_qos[2] s02_aw_qos[3] s02_aw_ready s02_aw_region[0] s02_aw_region[1] s02_aw_region[2]
+ s02_aw_region[3] s02_aw_size[0] s02_aw_size[1] s02_aw_size[2] s02_aw_user[-1] s02_aw_user[0]
+ s02_aw_valid s02_b_id[0] s02_b_id[1] s02_b_id[2] s02_b_id[3] s02_b_id[4] s02_b_id[5]
+ s02_b_id[6] s02_b_id[7] s02_b_id[8] s02_b_id[9] s02_b_ready s02_b_resp[0] s02_b_resp[1]
+ s02_b_user[-1] s02_b_user[0] s02_b_valid s02_r_data[0] s02_r_data[10] s02_r_data[11]
+ s02_r_data[12] s02_r_data[13] s02_r_data[14] s02_r_data[15] s02_r_data[16] s02_r_data[17]
+ s02_r_data[18] s02_r_data[19] s02_r_data[1] s02_r_data[20] s02_r_data[21] s02_r_data[22]
+ s02_r_data[23] s02_r_data[24] s02_r_data[25] s02_r_data[26] s02_r_data[27] s02_r_data[28]
+ s02_r_data[29] s02_r_data[2] s02_r_data[30] s02_r_data[31] s02_r_data[3] s02_r_data[4]
+ s02_r_data[5] s02_r_data[6] s02_r_data[7] s02_r_data[8] s02_r_data[9] s02_r_id[0]
+ s02_r_id[1] s02_r_id[2] s02_r_id[3] s02_r_id[4] s02_r_id[5] s02_r_id[6] s02_r_id[7]
+ s02_r_id[8] s02_r_id[9] s02_r_last s02_r_ready s02_r_resp[0] s02_r_resp[1] s02_r_user[-1]
+ s02_r_user[0] s02_r_valid s02_w_data[0] s02_w_data[10] s02_w_data[11] s02_w_data[12]
+ s02_w_data[13] s02_w_data[14] s02_w_data[15] s02_w_data[16] s02_w_data[17] s02_w_data[18]
+ s02_w_data[19] s02_w_data[1] s02_w_data[20] s02_w_data[21] s02_w_data[22] s02_w_data[23]
+ s02_w_data[24] s02_w_data[25] s02_w_data[26] s02_w_data[27] s02_w_data[28] s02_w_data[29]
+ s02_w_data[2] s02_w_data[30] s02_w_data[31] s02_w_data[3] s02_w_data[4] s02_w_data[5]
+ s02_w_data[6] s02_w_data[7] s02_w_data[8] s02_w_data[9] s02_w_last s02_w_ready s02_w_strb[0]
+ s02_w_strb[1] s02_w_strb[2] s02_w_strb[3] s02_w_user[-1] s02_w_user[0] s02_w_valid
+ test_en_i vccd1 vssd1
.ends

* Black-box entry subcircuit for mba_core_region abstract view
.subckt mba_core_region boot_addr_i[0] boot_addr_i[10] boot_addr_i[11] boot_addr_i[12]
+ boot_addr_i[13] boot_addr_i[14] boot_addr_i[15] boot_addr_i[16] boot_addr_i[17]
+ boot_addr_i[18] boot_addr_i[19] boot_addr_i[1] boot_addr_i[20] boot_addr_i[21] boot_addr_i[22]
+ boot_addr_i[23] boot_addr_i[24] boot_addr_i[25] boot_addr_i[26] boot_addr_i[27]
+ boot_addr_i[28] boot_addr_i[29] boot_addr_i[2] boot_addr_i[30] boot_addr_i[31] boot_addr_i[3]
+ boot_addr_i[4] boot_addr_i[5] boot_addr_i[6] boot_addr_i[7] boot_addr_i[8] boot_addr_i[9]
+ clk clock_gating_i core_busy_o core_master_ar_addr[0] core_master_ar_addr[10] core_master_ar_addr[11]
+ core_master_ar_addr[12] core_master_ar_addr[13] core_master_ar_addr[14] core_master_ar_addr[15]
+ core_master_ar_addr[16] core_master_ar_addr[17] core_master_ar_addr[18] core_master_ar_addr[19]
+ core_master_ar_addr[1] core_master_ar_addr[20] core_master_ar_addr[21] core_master_ar_addr[22]
+ core_master_ar_addr[23] core_master_ar_addr[24] core_master_ar_addr[25] core_master_ar_addr[26]
+ core_master_ar_addr[27] core_master_ar_addr[28] core_master_ar_addr[29] core_master_ar_addr[2]
+ core_master_ar_addr[30] core_master_ar_addr[31] core_master_ar_addr[3] core_master_ar_addr[4]
+ core_master_ar_addr[5] core_master_ar_addr[6] core_master_ar_addr[7] core_master_ar_addr[8]
+ core_master_ar_addr[9] core_master_ar_burst[0] core_master_ar_burst[1] core_master_ar_cache[0]
+ core_master_ar_cache[1] core_master_ar_cache[2] core_master_ar_cache[3] core_master_ar_id[0]
+ core_master_ar_id[1] core_master_ar_id[2] core_master_ar_id[3] core_master_ar_id[4]
+ core_master_ar_id[5] core_master_ar_id[6] core_master_ar_id[7] core_master_ar_id[8]
+ core_master_ar_id[9] core_master_ar_len[0] core_master_ar_len[1] core_master_ar_len[2]
+ core_master_ar_len[3] core_master_ar_len[4] core_master_ar_len[5] core_master_ar_len[6]
+ core_master_ar_len[7] core_master_ar_lock core_master_ar_prot[0] core_master_ar_prot[1]
+ core_master_ar_prot[2] core_master_ar_qos[0] core_master_ar_qos[1] core_master_ar_qos[2]
+ core_master_ar_qos[3] core_master_ar_ready core_master_ar_region[0] core_master_ar_region[1]
+ core_master_ar_region[2] core_master_ar_region[3] core_master_ar_size[0] core_master_ar_size[1]
+ core_master_ar_size[2] core_master_ar_user[-1] core_master_ar_user[0] core_master_ar_valid
+ core_master_aw_addr[0] core_master_aw_addr[10] core_master_aw_addr[11] core_master_aw_addr[12]
+ core_master_aw_addr[13] core_master_aw_addr[14] core_master_aw_addr[15] core_master_aw_addr[16]
+ core_master_aw_addr[17] core_master_aw_addr[18] core_master_aw_addr[19] core_master_aw_addr[1]
+ core_master_aw_addr[20] core_master_aw_addr[21] core_master_aw_addr[22] core_master_aw_addr[23]
+ core_master_aw_addr[24] core_master_aw_addr[25] core_master_aw_addr[26] core_master_aw_addr[27]
+ core_master_aw_addr[28] core_master_aw_addr[29] core_master_aw_addr[2] core_master_aw_addr[30]
+ core_master_aw_addr[31] core_master_aw_addr[3] core_master_aw_addr[4] core_master_aw_addr[5]
+ core_master_aw_addr[6] core_master_aw_addr[7] core_master_aw_addr[8] core_master_aw_addr[9]
+ core_master_aw_burst[0] core_master_aw_burst[1] core_master_aw_cache[0] core_master_aw_cache[1]
+ core_master_aw_cache[2] core_master_aw_cache[3] core_master_aw_id[0] core_master_aw_id[1]
+ core_master_aw_id[2] core_master_aw_id[3] core_master_aw_id[4] core_master_aw_id[5]
+ core_master_aw_id[6] core_master_aw_id[7] core_master_aw_id[8] core_master_aw_id[9]
+ core_master_aw_len[0] core_master_aw_len[1] core_master_aw_len[2] core_master_aw_len[3]
+ core_master_aw_len[4] core_master_aw_len[5] core_master_aw_len[6] core_master_aw_len[7]
+ core_master_aw_lock core_master_aw_prot[0] core_master_aw_prot[1] core_master_aw_prot[2]
+ core_master_aw_qos[0] core_master_aw_qos[1] core_master_aw_qos[2] core_master_aw_qos[3]
+ core_master_aw_ready core_master_aw_region[0] core_master_aw_region[1] core_master_aw_region[2]
+ core_master_aw_region[3] core_master_aw_size[0] core_master_aw_size[1] core_master_aw_size[2]
+ core_master_aw_user[-1] core_master_aw_user[0] core_master_aw_valid core_master_b_id[0]
+ core_master_b_id[1] core_master_b_id[2] core_master_b_id[3] core_master_b_id[4]
+ core_master_b_id[5] core_master_b_id[6] core_master_b_id[7] core_master_b_id[8]
+ core_master_b_id[9] core_master_b_ready core_master_b_resp[0] core_master_b_resp[1]
+ core_master_b_user[-1] core_master_b_user[0] core_master_b_valid core_master_r_data[0]
+ core_master_r_data[10] core_master_r_data[11] core_master_r_data[12] core_master_r_data[13]
+ core_master_r_data[14] core_master_r_data[15] core_master_r_data[16] core_master_r_data[17]
+ core_master_r_data[18] core_master_r_data[19] core_master_r_data[1] core_master_r_data[20]
+ core_master_r_data[21] core_master_r_data[22] core_master_r_data[23] core_master_r_data[24]
+ core_master_r_data[25] core_master_r_data[26] core_master_r_data[27] core_master_r_data[28]
+ core_master_r_data[29] core_master_r_data[2] core_master_r_data[30] core_master_r_data[31]
+ core_master_r_data[32] core_master_r_data[33] core_master_r_data[34] core_master_r_data[35]
+ core_master_r_data[36] core_master_r_data[37] core_master_r_data[38] core_master_r_data[39]
+ core_master_r_data[3] core_master_r_data[40] core_master_r_data[41] core_master_r_data[42]
+ core_master_r_data[43] core_master_r_data[44] core_master_r_data[45] core_master_r_data[46]
+ core_master_r_data[47] core_master_r_data[48] core_master_r_data[49] core_master_r_data[4]
+ core_master_r_data[50] core_master_r_data[51] core_master_r_data[52] core_master_r_data[53]
+ core_master_r_data[54] core_master_r_data[55] core_master_r_data[56] core_master_r_data[57]
+ core_master_r_data[58] core_master_r_data[59] core_master_r_data[5] core_master_r_data[60]
+ core_master_r_data[61] core_master_r_data[62] core_master_r_data[63] core_master_r_data[6]
+ core_master_r_data[7] core_master_r_data[8] core_master_r_data[9] core_master_r_id[0]
+ core_master_r_id[1] core_master_r_id[2] core_master_r_id[3] core_master_r_id[4]
+ core_master_r_id[5] core_master_r_id[6] core_master_r_id[7] core_master_r_id[8]
+ core_master_r_id[9] core_master_r_last core_master_r_ready core_master_r_resp[0]
+ core_master_r_resp[1] core_master_r_user[-1] core_master_r_user[0] core_master_r_valid
+ core_master_w_data[0] core_master_w_data[10] core_master_w_data[11] core_master_w_data[12]
+ core_master_w_data[13] core_master_w_data[14] core_master_w_data[15] core_master_w_data[16]
+ core_master_w_data[17] core_master_w_data[18] core_master_w_data[19] core_master_w_data[1]
+ core_master_w_data[20] core_master_w_data[21] core_master_w_data[22] core_master_w_data[23]
+ core_master_w_data[24] core_master_w_data[25] core_master_w_data[26] core_master_w_data[27]
+ core_master_w_data[28] core_master_w_data[29] core_master_w_data[2] core_master_w_data[30]
+ core_master_w_data[31] core_master_w_data[32] core_master_w_data[33] core_master_w_data[34]
+ core_master_w_data[35] core_master_w_data[36] core_master_w_data[37] core_master_w_data[38]
+ core_master_w_data[39] core_master_w_data[3] core_master_w_data[40] core_master_w_data[41]
+ core_master_w_data[42] core_master_w_data[43] core_master_w_data[44] core_master_w_data[45]
+ core_master_w_data[46] core_master_w_data[47] core_master_w_data[48] core_master_w_data[49]
+ core_master_w_data[4] core_master_w_data[50] core_master_w_data[51] core_master_w_data[52]
+ core_master_w_data[53] core_master_w_data[54] core_master_w_data[55] core_master_w_data[56]
+ core_master_w_data[57] core_master_w_data[58] core_master_w_data[59] core_master_w_data[5]
+ core_master_w_data[60] core_master_w_data[61] core_master_w_data[62] core_master_w_data[63]
+ core_master_w_data[6] core_master_w_data[7] core_master_w_data[8] core_master_w_data[9]
+ core_master_w_last core_master_w_ready core_master_w_strb[0] core_master_w_strb[1]
+ core_master_w_strb[2] core_master_w_strb[3] core_master_w_strb[4] core_master_w_strb[5]
+ core_master_w_strb[6] core_master_w_strb[7] core_master_w_user[-1] core_master_w_user[0]
+ core_master_w_valid data_slave_ar_addr[0] data_slave_ar_addr[10] data_slave_ar_addr[11]
+ data_slave_ar_addr[12] data_slave_ar_addr[13] data_slave_ar_addr[14] data_slave_ar_addr[15]
+ data_slave_ar_addr[16] data_slave_ar_addr[17] data_slave_ar_addr[18] data_slave_ar_addr[19]
+ data_slave_ar_addr[1] data_slave_ar_addr[20] data_slave_ar_addr[21] data_slave_ar_addr[22]
+ data_slave_ar_addr[23] data_slave_ar_addr[24] data_slave_ar_addr[25] data_slave_ar_addr[26]
+ data_slave_ar_addr[27] data_slave_ar_addr[28] data_slave_ar_addr[29] data_slave_ar_addr[2]
+ data_slave_ar_addr[30] data_slave_ar_addr[31] data_slave_ar_addr[3] data_slave_ar_addr[4]
+ data_slave_ar_addr[5] data_slave_ar_addr[6] data_slave_ar_addr[7] data_slave_ar_addr[8]
+ data_slave_ar_addr[9] data_slave_ar_burst[0] data_slave_ar_burst[1] data_slave_ar_cache[0]
+ data_slave_ar_cache[1] data_slave_ar_cache[2] data_slave_ar_cache[3] data_slave_ar_id[0]
+ data_slave_ar_id[1] data_slave_ar_id[2] data_slave_ar_id[3] data_slave_ar_id[4]
+ data_slave_ar_id[5] data_slave_ar_id[6] data_slave_ar_id[7] data_slave_ar_id[8]
+ data_slave_ar_id[9] data_slave_ar_len[0] data_slave_ar_len[1] data_slave_ar_len[2]
+ data_slave_ar_len[3] data_slave_ar_len[4] data_slave_ar_len[5] data_slave_ar_len[6]
+ data_slave_ar_len[7] data_slave_ar_lock data_slave_ar_prot[0] data_slave_ar_prot[1]
+ data_slave_ar_prot[2] data_slave_ar_qos[0] data_slave_ar_qos[1] data_slave_ar_qos[2]
+ data_slave_ar_qos[3] data_slave_ar_ready data_slave_ar_region[0] data_slave_ar_region[1]
+ data_slave_ar_region[2] data_slave_ar_region[3] data_slave_ar_size[0] data_slave_ar_size[1]
+ data_slave_ar_size[2] data_slave_ar_user[-1] data_slave_ar_user[0] data_slave_ar_valid
+ data_slave_aw_addr[0] data_slave_aw_addr[10] data_slave_aw_addr[11] data_slave_aw_addr[12]
+ data_slave_aw_addr[13] data_slave_aw_addr[14] data_slave_aw_addr[15] data_slave_aw_addr[16]
+ data_slave_aw_addr[17] data_slave_aw_addr[18] data_slave_aw_addr[19] data_slave_aw_addr[1]
+ data_slave_aw_addr[20] data_slave_aw_addr[21] data_slave_aw_addr[22] data_slave_aw_addr[23]
+ data_slave_aw_addr[24] data_slave_aw_addr[25] data_slave_aw_addr[26] data_slave_aw_addr[27]
+ data_slave_aw_addr[28] data_slave_aw_addr[29] data_slave_aw_addr[2] data_slave_aw_addr[30]
+ data_slave_aw_addr[31] data_slave_aw_addr[3] data_slave_aw_addr[4] data_slave_aw_addr[5]
+ data_slave_aw_addr[6] data_slave_aw_addr[7] data_slave_aw_addr[8] data_slave_aw_addr[9]
+ data_slave_aw_burst[0] data_slave_aw_burst[1] data_slave_aw_cache[0] data_slave_aw_cache[1]
+ data_slave_aw_cache[2] data_slave_aw_cache[3] data_slave_aw_id[0] data_slave_aw_id[1]
+ data_slave_aw_id[2] data_slave_aw_id[3] data_slave_aw_id[4] data_slave_aw_id[5]
+ data_slave_aw_id[6] data_slave_aw_id[7] data_slave_aw_id[8] data_slave_aw_id[9]
+ data_slave_aw_len[0] data_slave_aw_len[1] data_slave_aw_len[2] data_slave_aw_len[3]
+ data_slave_aw_len[4] data_slave_aw_len[5] data_slave_aw_len[6] data_slave_aw_len[7]
+ data_slave_aw_lock data_slave_aw_prot[0] data_slave_aw_prot[1] data_slave_aw_prot[2]
+ data_slave_aw_qos[0] data_slave_aw_qos[1] data_slave_aw_qos[2] data_slave_aw_qos[3]
+ data_slave_aw_ready data_slave_aw_region[0] data_slave_aw_region[1] data_slave_aw_region[2]
+ data_slave_aw_region[3] data_slave_aw_size[0] data_slave_aw_size[1] data_slave_aw_size[2]
+ data_slave_aw_user[-1] data_slave_aw_user[0] data_slave_aw_valid data_slave_b_id[0]
+ data_slave_b_id[1] data_slave_b_id[2] data_slave_b_id[3] data_slave_b_id[4] data_slave_b_id[5]
+ data_slave_b_id[6] data_slave_b_id[7] data_slave_b_id[8] data_slave_b_id[9] data_slave_b_ready
+ data_slave_b_resp[0] data_slave_b_resp[1] data_slave_b_user[-1] data_slave_b_user[0]
+ data_slave_b_valid data_slave_r_data[0] data_slave_r_data[10] data_slave_r_data[11]
+ data_slave_r_data[12] data_slave_r_data[13] data_slave_r_data[14] data_slave_r_data[15]
+ data_slave_r_data[16] data_slave_r_data[17] data_slave_r_data[18] data_slave_r_data[19]
+ data_slave_r_data[1] data_slave_r_data[20] data_slave_r_data[21] data_slave_r_data[22]
+ data_slave_r_data[23] data_slave_r_data[24] data_slave_r_data[25] data_slave_r_data[26]
+ data_slave_r_data[27] data_slave_r_data[28] data_slave_r_data[29] data_slave_r_data[2]
+ data_slave_r_data[30] data_slave_r_data[31] data_slave_r_data[32] data_slave_r_data[33]
+ data_slave_r_data[34] data_slave_r_data[35] data_slave_r_data[36] data_slave_r_data[37]
+ data_slave_r_data[38] data_slave_r_data[39] data_slave_r_data[3] data_slave_r_data[40]
+ data_slave_r_data[41] data_slave_r_data[42] data_slave_r_data[43] data_slave_r_data[44]
+ data_slave_r_data[45] data_slave_r_data[46] data_slave_r_data[47] data_slave_r_data[48]
+ data_slave_r_data[49] data_slave_r_data[4] data_slave_r_data[50] data_slave_r_data[51]
+ data_slave_r_data[52] data_slave_r_data[53] data_slave_r_data[54] data_slave_r_data[55]
+ data_slave_r_data[56] data_slave_r_data[57] data_slave_r_data[58] data_slave_r_data[59]
+ data_slave_r_data[5] data_slave_r_data[60] data_slave_r_data[61] data_slave_r_data[62]
+ data_slave_r_data[63] data_slave_r_data[6] data_slave_r_data[7] data_slave_r_data[8]
+ data_slave_r_data[9] data_slave_r_id[0] data_slave_r_id[1] data_slave_r_id[2] data_slave_r_id[3]
+ data_slave_r_id[4] data_slave_r_id[5] data_slave_r_id[6] data_slave_r_id[7] data_slave_r_id[8]
+ data_slave_r_id[9] data_slave_r_last data_slave_r_ready data_slave_r_resp[0] data_slave_r_resp[1]
+ data_slave_r_user[-1] data_slave_r_user[0] data_slave_r_valid data_slave_w_data[0]
+ data_slave_w_data[10] data_slave_w_data[11] data_slave_w_data[12] data_slave_w_data[13]
+ data_slave_w_data[14] data_slave_w_data[15] data_slave_w_data[16] data_slave_w_data[17]
+ data_slave_w_data[18] data_slave_w_data[19] data_slave_w_data[1] data_slave_w_data[20]
+ data_slave_w_data[21] data_slave_w_data[22] data_slave_w_data[23] data_slave_w_data[24]
+ data_slave_w_data[25] data_slave_w_data[26] data_slave_w_data[27] data_slave_w_data[28]
+ data_slave_w_data[29] data_slave_w_data[2] data_slave_w_data[30] data_slave_w_data[31]
+ data_slave_w_data[32] data_slave_w_data[33] data_slave_w_data[34] data_slave_w_data[35]
+ data_slave_w_data[36] data_slave_w_data[37] data_slave_w_data[38] data_slave_w_data[39]
+ data_slave_w_data[3] data_slave_w_data[40] data_slave_w_data[41] data_slave_w_data[42]
+ data_slave_w_data[43] data_slave_w_data[44] data_slave_w_data[45] data_slave_w_data[46]
+ data_slave_w_data[47] data_slave_w_data[48] data_slave_w_data[49] data_slave_w_data[4]
+ data_slave_w_data[50] data_slave_w_data[51] data_slave_w_data[52] data_slave_w_data[53]
+ data_slave_w_data[54] data_slave_w_data[55] data_slave_w_data[56] data_slave_w_data[57]
+ data_slave_w_data[58] data_slave_w_data[59] data_slave_w_data[5] data_slave_w_data[60]
+ data_slave_w_data[61] data_slave_w_data[62] data_slave_w_data[63] data_slave_w_data[6]
+ data_slave_w_data[7] data_slave_w_data[8] data_slave_w_data[9] data_slave_w_last
+ data_slave_w_ready data_slave_w_strb[0] data_slave_w_strb[1] data_slave_w_strb[2]
+ data_slave_w_strb[3] data_slave_w_strb[4] data_slave_w_strb[5] data_slave_w_strb[6]
+ data_slave_w_strb[7] data_slave_w_user[-1] data_slave_w_user[0] data_slave_w_valid
+ dbg_master_ar_addr[0] dbg_master_ar_addr[10] dbg_master_ar_addr[11] dbg_master_ar_addr[12]
+ dbg_master_ar_addr[13] dbg_master_ar_addr[14] dbg_master_ar_addr[15] dbg_master_ar_addr[16]
+ dbg_master_ar_addr[17] dbg_master_ar_addr[18] dbg_master_ar_addr[19] dbg_master_ar_addr[1]
+ dbg_master_ar_addr[20] dbg_master_ar_addr[21] dbg_master_ar_addr[22] dbg_master_ar_addr[23]
+ dbg_master_ar_addr[24] dbg_master_ar_addr[25] dbg_master_ar_addr[26] dbg_master_ar_addr[27]
+ dbg_master_ar_addr[28] dbg_master_ar_addr[29] dbg_master_ar_addr[2] dbg_master_ar_addr[30]
+ dbg_master_ar_addr[31] dbg_master_ar_addr[3] dbg_master_ar_addr[4] dbg_master_ar_addr[5]
+ dbg_master_ar_addr[6] dbg_master_ar_addr[7] dbg_master_ar_addr[8] dbg_master_ar_addr[9]
+ dbg_master_ar_burst[0] dbg_master_ar_burst[1] dbg_master_ar_cache[0] dbg_master_ar_cache[1]
+ dbg_master_ar_cache[2] dbg_master_ar_cache[3] dbg_master_ar_id[0] dbg_master_ar_id[1]
+ dbg_master_ar_id[2] dbg_master_ar_id[3] dbg_master_ar_id[4] dbg_master_ar_id[5]
+ dbg_master_ar_id[6] dbg_master_ar_id[7] dbg_master_ar_id[8] dbg_master_ar_id[9]
+ dbg_master_ar_len[0] dbg_master_ar_len[1] dbg_master_ar_len[2] dbg_master_ar_len[3]
+ dbg_master_ar_len[4] dbg_master_ar_len[5] dbg_master_ar_len[6] dbg_master_ar_len[7]
+ dbg_master_ar_lock dbg_master_ar_prot[0] dbg_master_ar_prot[1] dbg_master_ar_prot[2]
+ dbg_master_ar_qos[0] dbg_master_ar_qos[1] dbg_master_ar_qos[2] dbg_master_ar_qos[3]
+ dbg_master_ar_ready dbg_master_ar_region[0] dbg_master_ar_region[1] dbg_master_ar_region[2]
+ dbg_master_ar_region[3] dbg_master_ar_size[0] dbg_master_ar_size[1] dbg_master_ar_size[2]
+ dbg_master_ar_user[-1] dbg_master_ar_user[0] dbg_master_ar_valid dbg_master_aw_addr[0]
+ dbg_master_aw_addr[10] dbg_master_aw_addr[11] dbg_master_aw_addr[12] dbg_master_aw_addr[13]
+ dbg_master_aw_addr[14] dbg_master_aw_addr[15] dbg_master_aw_addr[16] dbg_master_aw_addr[17]
+ dbg_master_aw_addr[18] dbg_master_aw_addr[19] dbg_master_aw_addr[1] dbg_master_aw_addr[20]
+ dbg_master_aw_addr[21] dbg_master_aw_addr[22] dbg_master_aw_addr[23] dbg_master_aw_addr[24]
+ dbg_master_aw_addr[25] dbg_master_aw_addr[26] dbg_master_aw_addr[27] dbg_master_aw_addr[28]
+ dbg_master_aw_addr[29] dbg_master_aw_addr[2] dbg_master_aw_addr[30] dbg_master_aw_addr[31]
+ dbg_master_aw_addr[3] dbg_master_aw_addr[4] dbg_master_aw_addr[5] dbg_master_aw_addr[6]
+ dbg_master_aw_addr[7] dbg_master_aw_addr[8] dbg_master_aw_addr[9] dbg_master_aw_burst[0]
+ dbg_master_aw_burst[1] dbg_master_aw_cache[0] dbg_master_aw_cache[1] dbg_master_aw_cache[2]
+ dbg_master_aw_cache[3] dbg_master_aw_id[0] dbg_master_aw_id[1] dbg_master_aw_id[2]
+ dbg_master_aw_id[3] dbg_master_aw_id[4] dbg_master_aw_id[5] dbg_master_aw_id[6]
+ dbg_master_aw_id[7] dbg_master_aw_id[8] dbg_master_aw_id[9] dbg_master_aw_len[0]
+ dbg_master_aw_len[1] dbg_master_aw_len[2] dbg_master_aw_len[3] dbg_master_aw_len[4]
+ dbg_master_aw_len[5] dbg_master_aw_len[6] dbg_master_aw_len[7] dbg_master_aw_lock
+ dbg_master_aw_prot[0] dbg_master_aw_prot[1] dbg_master_aw_prot[2] dbg_master_aw_qos[0]
+ dbg_master_aw_qos[1] dbg_master_aw_qos[2] dbg_master_aw_qos[3] dbg_master_aw_ready
+ dbg_master_aw_region[0] dbg_master_aw_region[1] dbg_master_aw_region[2] dbg_master_aw_region[3]
+ dbg_master_aw_size[0] dbg_master_aw_size[1] dbg_master_aw_size[2] dbg_master_aw_user[-1]
+ dbg_master_aw_user[0] dbg_master_aw_valid dbg_master_b_id[0] dbg_master_b_id[1]
+ dbg_master_b_id[2] dbg_master_b_id[3] dbg_master_b_id[4] dbg_master_b_id[5] dbg_master_b_id[6]
+ dbg_master_b_id[7] dbg_master_b_id[8] dbg_master_b_id[9] dbg_master_b_ready dbg_master_b_resp[0]
+ dbg_master_b_resp[1] dbg_master_b_user[-1] dbg_master_b_user[0] dbg_master_b_valid
+ dbg_master_r_data[0] dbg_master_r_data[10] dbg_master_r_data[11] dbg_master_r_data[12]
+ dbg_master_r_data[13] dbg_master_r_data[14] dbg_master_r_data[15] dbg_master_r_data[16]
+ dbg_master_r_data[17] dbg_master_r_data[18] dbg_master_r_data[19] dbg_master_r_data[1]
+ dbg_master_r_data[20] dbg_master_r_data[21] dbg_master_r_data[22] dbg_master_r_data[23]
+ dbg_master_r_data[24] dbg_master_r_data[25] dbg_master_r_data[26] dbg_master_r_data[27]
+ dbg_master_r_data[28] dbg_master_r_data[29] dbg_master_r_data[2] dbg_master_r_data[30]
+ dbg_master_r_data[31] dbg_master_r_data[32] dbg_master_r_data[33] dbg_master_r_data[34]
+ dbg_master_r_data[35] dbg_master_r_data[36] dbg_master_r_data[37] dbg_master_r_data[38]
+ dbg_master_r_data[39] dbg_master_r_data[3] dbg_master_r_data[40] dbg_master_r_data[41]
+ dbg_master_r_data[42] dbg_master_r_data[43] dbg_master_r_data[44] dbg_master_r_data[45]
+ dbg_master_r_data[46] dbg_master_r_data[47] dbg_master_r_data[48] dbg_master_r_data[49]
+ dbg_master_r_data[4] dbg_master_r_data[50] dbg_master_r_data[51] dbg_master_r_data[52]
+ dbg_master_r_data[53] dbg_master_r_data[54] dbg_master_r_data[55] dbg_master_r_data[56]
+ dbg_master_r_data[57] dbg_master_r_data[58] dbg_master_r_data[59] dbg_master_r_data[5]
+ dbg_master_r_data[60] dbg_master_r_data[61] dbg_master_r_data[62] dbg_master_r_data[63]
+ dbg_master_r_data[6] dbg_master_r_data[7] dbg_master_r_data[8] dbg_master_r_data[9]
+ dbg_master_r_id[0] dbg_master_r_id[1] dbg_master_r_id[2] dbg_master_r_id[3] dbg_master_r_id[4]
+ dbg_master_r_id[5] dbg_master_r_id[6] dbg_master_r_id[7] dbg_master_r_id[8] dbg_master_r_id[9]
+ dbg_master_r_last dbg_master_r_ready dbg_master_r_resp[0] dbg_master_r_resp[1] dbg_master_r_user[-1]
+ dbg_master_r_user[0] dbg_master_r_valid dbg_master_w_data[0] dbg_master_w_data[10]
+ dbg_master_w_data[11] dbg_master_w_data[12] dbg_master_w_data[13] dbg_master_w_data[14]
+ dbg_master_w_data[15] dbg_master_w_data[16] dbg_master_w_data[17] dbg_master_w_data[18]
+ dbg_master_w_data[19] dbg_master_w_data[1] dbg_master_w_data[20] dbg_master_w_data[21]
+ dbg_master_w_data[22] dbg_master_w_data[23] dbg_master_w_data[24] dbg_master_w_data[25]
+ dbg_master_w_data[26] dbg_master_w_data[27] dbg_master_w_data[28] dbg_master_w_data[29]
+ dbg_master_w_data[2] dbg_master_w_data[30] dbg_master_w_data[31] dbg_master_w_data[32]
+ dbg_master_w_data[33] dbg_master_w_data[34] dbg_master_w_data[35] dbg_master_w_data[36]
+ dbg_master_w_data[37] dbg_master_w_data[38] dbg_master_w_data[39] dbg_master_w_data[3]
+ dbg_master_w_data[40] dbg_master_w_data[41] dbg_master_w_data[42] dbg_master_w_data[43]
+ dbg_master_w_data[44] dbg_master_w_data[45] dbg_master_w_data[46] dbg_master_w_data[47]
+ dbg_master_w_data[48] dbg_master_w_data[49] dbg_master_w_data[4] dbg_master_w_data[50]
+ dbg_master_w_data[51] dbg_master_w_data[52] dbg_master_w_data[53] dbg_master_w_data[54]
+ dbg_master_w_data[55] dbg_master_w_data[56] dbg_master_w_data[57] dbg_master_w_data[58]
+ dbg_master_w_data[59] dbg_master_w_data[5] dbg_master_w_data[60] dbg_master_w_data[61]
+ dbg_master_w_data[62] dbg_master_w_data[63] dbg_master_w_data[6] dbg_master_w_data[7]
+ dbg_master_w_data[8] dbg_master_w_data[9] dbg_master_w_last dbg_master_w_ready dbg_master_w_strb[0]
+ dbg_master_w_strb[1] dbg_master_w_strb[2] dbg_master_w_strb[3] dbg_master_w_strb[4]
+ dbg_master_w_strb[5] dbg_master_w_strb[6] dbg_master_w_strb[7] dbg_master_w_user[-1]
+ dbg_master_w_user[0] dbg_master_w_valid debug_addr[0] debug_addr[10] debug_addr[11]
+ debug_addr[12] debug_addr[13] debug_addr[14] debug_addr[1] debug_addr[2] debug_addr[3]
+ debug_addr[4] debug_addr[5] debug_addr[6] debug_addr[7] debug_addr[8] debug_addr[9]
+ debug_gnt debug_rdata[0] debug_rdata[10] debug_rdata[11] debug_rdata[12] debug_rdata[13]
+ debug_rdata[14] debug_rdata[15] debug_rdata[16] debug_rdata[17] debug_rdata[18]
+ debug_rdata[19] debug_rdata[1] debug_rdata[20] debug_rdata[21] debug_rdata[22] debug_rdata[23]
+ debug_rdata[24] debug_rdata[25] debug_rdata[26] debug_rdata[27] debug_rdata[28]
+ debug_rdata[29] debug_rdata[2] debug_rdata[30] debug_rdata[31] debug_rdata[3] debug_rdata[4]
+ debug_rdata[5] debug_rdata[6] debug_rdata[7] debug_rdata[8] debug_rdata[9] debug_req
+ debug_rvalid debug_wdata[0] debug_wdata[10] debug_wdata[11] debug_wdata[12] debug_wdata[13]
+ debug_wdata[14] debug_wdata[15] debug_wdata[16] debug_wdata[17] debug_wdata[18]
+ debug_wdata[19] debug_wdata[1] debug_wdata[20] debug_wdata[21] debug_wdata[22] debug_wdata[23]
+ debug_wdata[24] debug_wdata[25] debug_wdata[26] debug_wdata[27] debug_wdata[28]
+ debug_wdata[29] debug_wdata[2] debug_wdata[30] debug_wdata[31] debug_wdata[3] debug_wdata[4]
+ debug_wdata[5] debug_wdata[6] debug_wdata[7] debug_wdata[8] debug_wdata[9] debug_we
+ fetch_enable_i instr_slave_ar_addr[0] instr_slave_ar_addr[10] instr_slave_ar_addr[11]
+ instr_slave_ar_addr[12] instr_slave_ar_addr[13] instr_slave_ar_addr[14] instr_slave_ar_addr[15]
+ instr_slave_ar_addr[16] instr_slave_ar_addr[17] instr_slave_ar_addr[18] instr_slave_ar_addr[19]
+ instr_slave_ar_addr[1] instr_slave_ar_addr[20] instr_slave_ar_addr[21] instr_slave_ar_addr[22]
+ instr_slave_ar_addr[23] instr_slave_ar_addr[24] instr_slave_ar_addr[25] instr_slave_ar_addr[26]
+ instr_slave_ar_addr[27] instr_slave_ar_addr[28] instr_slave_ar_addr[29] instr_slave_ar_addr[2]
+ instr_slave_ar_addr[30] instr_slave_ar_addr[31] instr_slave_ar_addr[3] instr_slave_ar_addr[4]
+ instr_slave_ar_addr[5] instr_slave_ar_addr[6] instr_slave_ar_addr[7] instr_slave_ar_addr[8]
+ instr_slave_ar_addr[9] instr_slave_ar_burst[0] instr_slave_ar_burst[1] instr_slave_ar_cache[0]
+ instr_slave_ar_cache[1] instr_slave_ar_cache[2] instr_slave_ar_cache[3] instr_slave_ar_id[0]
+ instr_slave_ar_id[1] instr_slave_ar_id[2] instr_slave_ar_id[3] instr_slave_ar_id[4]
+ instr_slave_ar_id[5] instr_slave_ar_id[6] instr_slave_ar_id[7] instr_slave_ar_id[8]
+ instr_slave_ar_id[9] instr_slave_ar_len[0] instr_slave_ar_len[1] instr_slave_ar_len[2]
+ instr_slave_ar_len[3] instr_slave_ar_len[4] instr_slave_ar_len[5] instr_slave_ar_len[6]
+ instr_slave_ar_len[7] instr_slave_ar_lock instr_slave_ar_prot[0] instr_slave_ar_prot[1]
+ instr_slave_ar_prot[2] instr_slave_ar_qos[0] instr_slave_ar_qos[1] instr_slave_ar_qos[2]
+ instr_slave_ar_qos[3] instr_slave_ar_ready instr_slave_ar_region[0] instr_slave_ar_region[1]
+ instr_slave_ar_region[2] instr_slave_ar_region[3] instr_slave_ar_size[0] instr_slave_ar_size[1]
+ instr_slave_ar_size[2] instr_slave_ar_user[-1] instr_slave_ar_user[0] instr_slave_ar_valid
+ instr_slave_aw_addr[0] instr_slave_aw_addr[10] instr_slave_aw_addr[11] instr_slave_aw_addr[12]
+ instr_slave_aw_addr[13] instr_slave_aw_addr[14] instr_slave_aw_addr[15] instr_slave_aw_addr[16]
+ instr_slave_aw_addr[17] instr_slave_aw_addr[18] instr_slave_aw_addr[19] instr_slave_aw_addr[1]
+ instr_slave_aw_addr[20] instr_slave_aw_addr[21] instr_slave_aw_addr[22] instr_slave_aw_addr[23]
+ instr_slave_aw_addr[24] instr_slave_aw_addr[25] instr_slave_aw_addr[26] instr_slave_aw_addr[27]
+ instr_slave_aw_addr[28] instr_slave_aw_addr[29] instr_slave_aw_addr[2] instr_slave_aw_addr[30]
+ instr_slave_aw_addr[31] instr_slave_aw_addr[3] instr_slave_aw_addr[4] instr_slave_aw_addr[5]
+ instr_slave_aw_addr[6] instr_slave_aw_addr[7] instr_slave_aw_addr[8] instr_slave_aw_addr[9]
+ instr_slave_aw_burst[0] instr_slave_aw_burst[1] instr_slave_aw_cache[0] instr_slave_aw_cache[1]
+ instr_slave_aw_cache[2] instr_slave_aw_cache[3] instr_slave_aw_id[0] instr_slave_aw_id[1]
+ instr_slave_aw_id[2] instr_slave_aw_id[3] instr_slave_aw_id[4] instr_slave_aw_id[5]
+ instr_slave_aw_id[6] instr_slave_aw_id[7] instr_slave_aw_id[8] instr_slave_aw_id[9]
+ instr_slave_aw_len[0] instr_slave_aw_len[1] instr_slave_aw_len[2] instr_slave_aw_len[3]
+ instr_slave_aw_len[4] instr_slave_aw_len[5] instr_slave_aw_len[6] instr_slave_aw_len[7]
+ instr_slave_aw_lock instr_slave_aw_prot[0] instr_slave_aw_prot[1] instr_slave_aw_prot[2]
+ instr_slave_aw_qos[0] instr_slave_aw_qos[1] instr_slave_aw_qos[2] instr_slave_aw_qos[3]
+ instr_slave_aw_ready instr_slave_aw_region[0] instr_slave_aw_region[1] instr_slave_aw_region[2]
+ instr_slave_aw_region[3] instr_slave_aw_size[0] instr_slave_aw_size[1] instr_slave_aw_size[2]
+ instr_slave_aw_user[-1] instr_slave_aw_user[0] instr_slave_aw_valid instr_slave_b_id[0]
+ instr_slave_b_id[1] instr_slave_b_id[2] instr_slave_b_id[3] instr_slave_b_id[4]
+ instr_slave_b_id[5] instr_slave_b_id[6] instr_slave_b_id[7] instr_slave_b_id[8]
+ instr_slave_b_id[9] instr_slave_b_ready instr_slave_b_resp[0] instr_slave_b_resp[1]
+ instr_slave_b_user[-1] instr_slave_b_user[0] instr_slave_b_valid instr_slave_r_data[0]
+ instr_slave_r_data[10] instr_slave_r_data[11] instr_slave_r_data[12] instr_slave_r_data[13]
+ instr_slave_r_data[14] instr_slave_r_data[15] instr_slave_r_data[16] instr_slave_r_data[17]
+ instr_slave_r_data[18] instr_slave_r_data[19] instr_slave_r_data[1] instr_slave_r_data[20]
+ instr_slave_r_data[21] instr_slave_r_data[22] instr_slave_r_data[23] instr_slave_r_data[24]
+ instr_slave_r_data[25] instr_slave_r_data[26] instr_slave_r_data[27] instr_slave_r_data[28]
+ instr_slave_r_data[29] instr_slave_r_data[2] instr_slave_r_data[30] instr_slave_r_data[31]
+ instr_slave_r_data[32] instr_slave_r_data[33] instr_slave_r_data[34] instr_slave_r_data[35]
+ instr_slave_r_data[36] instr_slave_r_data[37] instr_slave_r_data[38] instr_slave_r_data[39]
+ instr_slave_r_data[3] instr_slave_r_data[40] instr_slave_r_data[41] instr_slave_r_data[42]
+ instr_slave_r_data[43] instr_slave_r_data[44] instr_slave_r_data[45] instr_slave_r_data[46]
+ instr_slave_r_data[47] instr_slave_r_data[48] instr_slave_r_data[49] instr_slave_r_data[4]
+ instr_slave_r_data[50] instr_slave_r_data[51] instr_slave_r_data[52] instr_slave_r_data[53]
+ instr_slave_r_data[54] instr_slave_r_data[55] instr_slave_r_data[56] instr_slave_r_data[57]
+ instr_slave_r_data[58] instr_slave_r_data[59] instr_slave_r_data[5] instr_slave_r_data[60]
+ instr_slave_r_data[61] instr_slave_r_data[62] instr_slave_r_data[63] instr_slave_r_data[6]
+ instr_slave_r_data[7] instr_slave_r_data[8] instr_slave_r_data[9] instr_slave_r_id[0]
+ instr_slave_r_id[1] instr_slave_r_id[2] instr_slave_r_id[3] instr_slave_r_id[4]
+ instr_slave_r_id[5] instr_slave_r_id[6] instr_slave_r_id[7] instr_slave_r_id[8]
+ instr_slave_r_id[9] instr_slave_r_last instr_slave_r_ready instr_slave_r_resp[0]
+ instr_slave_r_resp[1] instr_slave_r_user[-1] instr_slave_r_user[0] instr_slave_r_valid
+ instr_slave_w_data[0] instr_slave_w_data[10] instr_slave_w_data[11] instr_slave_w_data[12]
+ instr_slave_w_data[13] instr_slave_w_data[14] instr_slave_w_data[15] instr_slave_w_data[16]
+ instr_slave_w_data[17] instr_slave_w_data[18] instr_slave_w_data[19] instr_slave_w_data[1]
+ instr_slave_w_data[20] instr_slave_w_data[21] instr_slave_w_data[22] instr_slave_w_data[23]
+ instr_slave_w_data[24] instr_slave_w_data[25] instr_slave_w_data[26] instr_slave_w_data[27]
+ instr_slave_w_data[28] instr_slave_w_data[29] instr_slave_w_data[2] instr_slave_w_data[30]
+ instr_slave_w_data[31] instr_slave_w_data[32] instr_slave_w_data[33] instr_slave_w_data[34]
+ instr_slave_w_data[35] instr_slave_w_data[36] instr_slave_w_data[37] instr_slave_w_data[38]
+ instr_slave_w_data[39] instr_slave_w_data[3] instr_slave_w_data[40] instr_slave_w_data[41]
+ instr_slave_w_data[42] instr_slave_w_data[43] instr_slave_w_data[44] instr_slave_w_data[45]
+ instr_slave_w_data[46] instr_slave_w_data[47] instr_slave_w_data[48] instr_slave_w_data[49]
+ instr_slave_w_data[4] instr_slave_w_data[50] instr_slave_w_data[51] instr_slave_w_data[52]
+ instr_slave_w_data[53] instr_slave_w_data[54] instr_slave_w_data[55] instr_slave_w_data[56]
+ instr_slave_w_data[57] instr_slave_w_data[58] instr_slave_w_data[59] instr_slave_w_data[5]
+ instr_slave_w_data[60] instr_slave_w_data[61] instr_slave_w_data[62] instr_slave_w_data[63]
+ instr_slave_w_data[6] instr_slave_w_data[7] instr_slave_w_data[8] instr_slave_w_data[9]
+ instr_slave_w_last instr_slave_w_ready instr_slave_w_strb[0] instr_slave_w_strb[1]
+ instr_slave_w_strb[2] instr_slave_w_strb[3] instr_slave_w_strb[4] instr_slave_w_strb[5]
+ instr_slave_w_strb[6] instr_slave_w_strb[7] instr_slave_w_user[-1] instr_slave_w_user[0]
+ instr_slave_w_valid irq_i[0] irq_i[10] irq_i[11] irq_i[12] irq_i[13] irq_i[14] irq_i[15]
+ irq_i[16] irq_i[17] irq_i[18] irq_i[19] irq_i[1] irq_i[20] irq_i[21] irq_i[22] irq_i[23]
+ irq_i[24] irq_i[25] irq_i[26] irq_i[27] irq_i[28] irq_i[29] irq_i[2] irq_i[30] irq_i[31]
+ irq_i[3] irq_i[4] irq_i[5] irq_i[6] irq_i[7] irq_i[8] irq_i[9] mba_data_mem_addr0_o[0]
+ mba_data_mem_addr0_o[10] mba_data_mem_addr0_o[11] mba_data_mem_addr0_o[12] mba_data_mem_addr0_o[13]
+ mba_data_mem_addr0_o[14] mba_data_mem_addr0_o[15] mba_data_mem_addr0_o[16] mba_data_mem_addr0_o[17]
+ mba_data_mem_addr0_o[18] mba_data_mem_addr0_o[19] mba_data_mem_addr0_o[1] mba_data_mem_addr0_o[20]
+ mba_data_mem_addr0_o[21] mba_data_mem_addr0_o[22] mba_data_mem_addr0_o[23] mba_data_mem_addr0_o[24]
+ mba_data_mem_addr0_o[25] mba_data_mem_addr0_o[26] mba_data_mem_addr0_o[27] mba_data_mem_addr0_o[28]
+ mba_data_mem_addr0_o[29] mba_data_mem_addr0_o[2] mba_data_mem_addr0_o[30] mba_data_mem_addr0_o[31]
+ mba_data_mem_addr0_o[3] mba_data_mem_addr0_o[4] mba_data_mem_addr0_o[5] mba_data_mem_addr0_o[6]
+ mba_data_mem_addr0_o[7] mba_data_mem_addr0_o[8] mba_data_mem_addr0_o[9] mba_data_mem_addr1_o[0]
+ mba_data_mem_addr1_o[10] mba_data_mem_addr1_o[11] mba_data_mem_addr1_o[12] mba_data_mem_addr1_o[13]
+ mba_data_mem_addr1_o[14] mba_data_mem_addr1_o[15] mba_data_mem_addr1_o[16] mba_data_mem_addr1_o[17]
+ mba_data_mem_addr1_o[18] mba_data_mem_addr1_o[19] mba_data_mem_addr1_o[1] mba_data_mem_addr1_o[20]
+ mba_data_mem_addr1_o[21] mba_data_mem_addr1_o[22] mba_data_mem_addr1_o[23] mba_data_mem_addr1_o[24]
+ mba_data_mem_addr1_o[25] mba_data_mem_addr1_o[26] mba_data_mem_addr1_o[27] mba_data_mem_addr1_o[28]
+ mba_data_mem_addr1_o[29] mba_data_mem_addr1_o[2] mba_data_mem_addr1_o[30] mba_data_mem_addr1_o[31]
+ mba_data_mem_addr1_o[3] mba_data_mem_addr1_o[4] mba_data_mem_addr1_o[5] mba_data_mem_addr1_o[6]
+ mba_data_mem_addr1_o[7] mba_data_mem_addr1_o[8] mba_data_mem_addr1_o[9] mba_data_mem_csb0_o
+ mba_data_mem_csb1_o mba_data_mem_din0_o[0] mba_data_mem_din0_o[10] mba_data_mem_din0_o[11]
+ mba_data_mem_din0_o[12] mba_data_mem_din0_o[13] mba_data_mem_din0_o[14] mba_data_mem_din0_o[15]
+ mba_data_mem_din0_o[16] mba_data_mem_din0_o[17] mba_data_mem_din0_o[18] mba_data_mem_din0_o[19]
+ mba_data_mem_din0_o[1] mba_data_mem_din0_o[20] mba_data_mem_din0_o[21] mba_data_mem_din0_o[22]
+ mba_data_mem_din0_o[23] mba_data_mem_din0_o[24] mba_data_mem_din0_o[25] mba_data_mem_din0_o[26]
+ mba_data_mem_din0_o[27] mba_data_mem_din0_o[28] mba_data_mem_din0_o[29] mba_data_mem_din0_o[2]
+ mba_data_mem_din0_o[30] mba_data_mem_din0_o[31] mba_data_mem_din0_o[3] mba_data_mem_din0_o[4]
+ mba_data_mem_din0_o[5] mba_data_mem_din0_o[6] mba_data_mem_din0_o[7] mba_data_mem_din0_o[8]
+ mba_data_mem_din0_o[9] mba_data_mem_dout0_i[0] mba_data_mem_dout0_i[10] mba_data_mem_dout0_i[11]
+ mba_data_mem_dout0_i[12] mba_data_mem_dout0_i[13] mba_data_mem_dout0_i[14] mba_data_mem_dout0_i[15]
+ mba_data_mem_dout0_i[16] mba_data_mem_dout0_i[17] mba_data_mem_dout0_i[18] mba_data_mem_dout0_i[19]
+ mba_data_mem_dout0_i[1] mba_data_mem_dout0_i[20] mba_data_mem_dout0_i[21] mba_data_mem_dout0_i[22]
+ mba_data_mem_dout0_i[23] mba_data_mem_dout0_i[24] mba_data_mem_dout0_i[25] mba_data_mem_dout0_i[26]
+ mba_data_mem_dout0_i[27] mba_data_mem_dout0_i[28] mba_data_mem_dout0_i[29] mba_data_mem_dout0_i[2]
+ mba_data_mem_dout0_i[30] mba_data_mem_dout0_i[31] mba_data_mem_dout0_i[3] mba_data_mem_dout0_i[4]
+ mba_data_mem_dout0_i[5] mba_data_mem_dout0_i[6] mba_data_mem_dout0_i[7] mba_data_mem_dout0_i[8]
+ mba_data_mem_dout0_i[9] mba_data_mem_web0_o mba_data_mem_wmask0_o[0] mba_data_mem_wmask0_o[1]
+ mba_data_mem_wmask0_o[2] mba_data_mem_wmask0_o[3] mba_instr_mem_addr0_o[0] mba_instr_mem_addr0_o[10]
+ mba_instr_mem_addr0_o[11] mba_instr_mem_addr0_o[12] mba_instr_mem_addr0_o[13] mba_instr_mem_addr0_o[14]
+ mba_instr_mem_addr0_o[15] mba_instr_mem_addr0_o[16] mba_instr_mem_addr0_o[17] mba_instr_mem_addr0_o[18]
+ mba_instr_mem_addr0_o[19] mba_instr_mem_addr0_o[1] mba_instr_mem_addr0_o[20] mba_instr_mem_addr0_o[21]
+ mba_instr_mem_addr0_o[22] mba_instr_mem_addr0_o[23] mba_instr_mem_addr0_o[24] mba_instr_mem_addr0_o[25]
+ mba_instr_mem_addr0_o[26] mba_instr_mem_addr0_o[27] mba_instr_mem_addr0_o[28] mba_instr_mem_addr0_o[29]
+ mba_instr_mem_addr0_o[2] mba_instr_mem_addr0_o[30] mba_instr_mem_addr0_o[31] mba_instr_mem_addr0_o[3]
+ mba_instr_mem_addr0_o[4] mba_instr_mem_addr0_o[5] mba_instr_mem_addr0_o[6] mba_instr_mem_addr0_o[7]
+ mba_instr_mem_addr0_o[8] mba_instr_mem_addr0_o[9] mba_instr_mem_addr1_o[0] mba_instr_mem_addr1_o[10]
+ mba_instr_mem_addr1_o[11] mba_instr_mem_addr1_o[12] mba_instr_mem_addr1_o[13] mba_instr_mem_addr1_o[14]
+ mba_instr_mem_addr1_o[15] mba_instr_mem_addr1_o[16] mba_instr_mem_addr1_o[17] mba_instr_mem_addr1_o[18]
+ mba_instr_mem_addr1_o[19] mba_instr_mem_addr1_o[1] mba_instr_mem_addr1_o[20] mba_instr_mem_addr1_o[21]
+ mba_instr_mem_addr1_o[22] mba_instr_mem_addr1_o[23] mba_instr_mem_addr1_o[24] mba_instr_mem_addr1_o[25]
+ mba_instr_mem_addr1_o[26] mba_instr_mem_addr1_o[27] mba_instr_mem_addr1_o[28] mba_instr_mem_addr1_o[29]
+ mba_instr_mem_addr1_o[2] mba_instr_mem_addr1_o[30] mba_instr_mem_addr1_o[31] mba_instr_mem_addr1_o[3]
+ mba_instr_mem_addr1_o[4] mba_instr_mem_addr1_o[5] mba_instr_mem_addr1_o[6] mba_instr_mem_addr1_o[7]
+ mba_instr_mem_addr1_o[8] mba_instr_mem_addr1_o[9] mba_instr_mem_csb0_o mba_instr_mem_csb1_o
+ mba_instr_mem_din0_o[0] mba_instr_mem_din0_o[10] mba_instr_mem_din0_o[11] mba_instr_mem_din0_o[12]
+ mba_instr_mem_din0_o[13] mba_instr_mem_din0_o[14] mba_instr_mem_din0_o[15] mba_instr_mem_din0_o[16]
+ mba_instr_mem_din0_o[17] mba_instr_mem_din0_o[18] mba_instr_mem_din0_o[19] mba_instr_mem_din0_o[1]
+ mba_instr_mem_din0_o[20] mba_instr_mem_din0_o[21] mba_instr_mem_din0_o[22] mba_instr_mem_din0_o[23]
+ mba_instr_mem_din0_o[24] mba_instr_mem_din0_o[25] mba_instr_mem_din0_o[26] mba_instr_mem_din0_o[27]
+ mba_instr_mem_din0_o[28] mba_instr_mem_din0_o[29] mba_instr_mem_din0_o[2] mba_instr_mem_din0_o[30]
+ mba_instr_mem_din0_o[31] mba_instr_mem_din0_o[3] mba_instr_mem_din0_o[4] mba_instr_mem_din0_o[5]
+ mba_instr_mem_din0_o[6] mba_instr_mem_din0_o[7] mba_instr_mem_din0_o[8] mba_instr_mem_din0_o[9]
+ mba_instr_mem_dout0_i[0] mba_instr_mem_dout0_i[10] mba_instr_mem_dout0_i[11] mba_instr_mem_dout0_i[12]
+ mba_instr_mem_dout0_i[13] mba_instr_mem_dout0_i[14] mba_instr_mem_dout0_i[15] mba_instr_mem_dout0_i[16]
+ mba_instr_mem_dout0_i[17] mba_instr_mem_dout0_i[18] mba_instr_mem_dout0_i[19] mba_instr_mem_dout0_i[1]
+ mba_instr_mem_dout0_i[20] mba_instr_mem_dout0_i[21] mba_instr_mem_dout0_i[22] mba_instr_mem_dout0_i[23]
+ mba_instr_mem_dout0_i[24] mba_instr_mem_dout0_i[25] mba_instr_mem_dout0_i[26] mba_instr_mem_dout0_i[27]
+ mba_instr_mem_dout0_i[28] mba_instr_mem_dout0_i[29] mba_instr_mem_dout0_i[2] mba_instr_mem_dout0_i[30]
+ mba_instr_mem_dout0_i[31] mba_instr_mem_dout0_i[3] mba_instr_mem_dout0_i[4] mba_instr_mem_dout0_i[5]
+ mba_instr_mem_dout0_i[6] mba_instr_mem_dout0_i[7] mba_instr_mem_dout0_i[8] mba_instr_mem_dout0_i[9]
+ mba_instr_mem_web0_o mba_instr_mem_wmask0_o[0] mba_instr_mem_wmask0_o[1] mba_instr_mem_wmask0_o[2]
+ mba_instr_mem_wmask0_o[3] rst_n tck_i tdi_i tdo_o testmode_i tms_i trstn_i vccd1
+ vssd1
.ends

* Black-box entry subcircuit for sky130_sram_2kbyte_1rw1r_32x512_8 abstract view
.subckt sky130_sram_2kbyte_1rw1r_32x512_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr1[0]
+ addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] addr1[8] csb0 csb1
+ web0 clk0 clk1 wmask0[0] wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4]
+ dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13]
+ dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21]
+ dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29]
+ dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for peripherals abstract view
.subckt peripherals axi_spi_master_ar_addr[0] axi_spi_master_ar_addr[10] axi_spi_master_ar_addr[11]
+ axi_spi_master_ar_addr[12] axi_spi_master_ar_addr[13] axi_spi_master_ar_addr[14]
+ axi_spi_master_ar_addr[15] axi_spi_master_ar_addr[16] axi_spi_master_ar_addr[17]
+ axi_spi_master_ar_addr[18] axi_spi_master_ar_addr[19] axi_spi_master_ar_addr[1]
+ axi_spi_master_ar_addr[20] axi_spi_master_ar_addr[21] axi_spi_master_ar_addr[22]
+ axi_spi_master_ar_addr[23] axi_spi_master_ar_addr[24] axi_spi_master_ar_addr[25]
+ axi_spi_master_ar_addr[26] axi_spi_master_ar_addr[27] axi_spi_master_ar_addr[28]
+ axi_spi_master_ar_addr[29] axi_spi_master_ar_addr[2] axi_spi_master_ar_addr[30]
+ axi_spi_master_ar_addr[31] axi_spi_master_ar_addr[3] axi_spi_master_ar_addr[4] axi_spi_master_ar_addr[5]
+ axi_spi_master_ar_addr[6] axi_spi_master_ar_addr[7] axi_spi_master_ar_addr[8] axi_spi_master_ar_addr[9]
+ axi_spi_master_ar_burst[0] axi_spi_master_ar_burst[1] axi_spi_master_ar_cache[0]
+ axi_spi_master_ar_cache[1] axi_spi_master_ar_cache[2] axi_spi_master_ar_cache[3]
+ axi_spi_master_ar_id[0] axi_spi_master_ar_id[1] axi_spi_master_ar_id[2] axi_spi_master_ar_id[3]
+ axi_spi_master_ar_id[4] axi_spi_master_ar_id[5] axi_spi_master_ar_len[0] axi_spi_master_ar_len[1]
+ axi_spi_master_ar_len[2] axi_spi_master_ar_len[3] axi_spi_master_ar_len[4] axi_spi_master_ar_len[5]
+ axi_spi_master_ar_len[6] axi_spi_master_ar_len[7] axi_spi_master_ar_lock axi_spi_master_ar_prot[0]
+ axi_spi_master_ar_prot[1] axi_spi_master_ar_prot[2] axi_spi_master_ar_qos[0] axi_spi_master_ar_qos[1]
+ axi_spi_master_ar_qos[2] axi_spi_master_ar_qos[3] axi_spi_master_ar_ready axi_spi_master_ar_region[0]
+ axi_spi_master_ar_region[1] axi_spi_master_ar_region[2] axi_spi_master_ar_region[3]
+ axi_spi_master_ar_size[0] axi_spi_master_ar_size[1] axi_spi_master_ar_size[2] axi_spi_master_ar_user[0]
+ axi_spi_master_ar_user[1] axi_spi_master_ar_user[2] axi_spi_master_ar_user[3] axi_spi_master_ar_user[4]
+ axi_spi_master_ar_user[5] axi_spi_master_ar_valid axi_spi_master_aw_addr[0] axi_spi_master_aw_addr[10]
+ axi_spi_master_aw_addr[11] axi_spi_master_aw_addr[12] axi_spi_master_aw_addr[13]
+ axi_spi_master_aw_addr[14] axi_spi_master_aw_addr[15] axi_spi_master_aw_addr[16]
+ axi_spi_master_aw_addr[17] axi_spi_master_aw_addr[18] axi_spi_master_aw_addr[19]
+ axi_spi_master_aw_addr[1] axi_spi_master_aw_addr[20] axi_spi_master_aw_addr[21]
+ axi_spi_master_aw_addr[22] axi_spi_master_aw_addr[23] axi_spi_master_aw_addr[24]
+ axi_spi_master_aw_addr[25] axi_spi_master_aw_addr[26] axi_spi_master_aw_addr[27]
+ axi_spi_master_aw_addr[28] axi_spi_master_aw_addr[29] axi_spi_master_aw_addr[2]
+ axi_spi_master_aw_addr[30] axi_spi_master_aw_addr[31] axi_spi_master_aw_addr[3]
+ axi_spi_master_aw_addr[4] axi_spi_master_aw_addr[5] axi_spi_master_aw_addr[6] axi_spi_master_aw_addr[7]
+ axi_spi_master_aw_addr[8] axi_spi_master_aw_addr[9] axi_spi_master_aw_burst[0] axi_spi_master_aw_burst[1]
+ axi_spi_master_aw_cache[0] axi_spi_master_aw_cache[1] axi_spi_master_aw_cache[2]
+ axi_spi_master_aw_cache[3] axi_spi_master_aw_id[0] axi_spi_master_aw_id[1] axi_spi_master_aw_id[2]
+ axi_spi_master_aw_id[3] axi_spi_master_aw_id[4] axi_spi_master_aw_id[5] axi_spi_master_aw_len[0]
+ axi_spi_master_aw_len[1] axi_spi_master_aw_len[2] axi_spi_master_aw_len[3] axi_spi_master_aw_len[4]
+ axi_spi_master_aw_len[5] axi_spi_master_aw_len[6] axi_spi_master_aw_len[7] axi_spi_master_aw_lock
+ axi_spi_master_aw_prot[0] axi_spi_master_aw_prot[1] axi_spi_master_aw_prot[2] axi_spi_master_aw_qos[0]
+ axi_spi_master_aw_qos[1] axi_spi_master_aw_qos[2] axi_spi_master_aw_qos[3] axi_spi_master_aw_ready
+ axi_spi_master_aw_region[0] axi_spi_master_aw_region[1] axi_spi_master_aw_region[2]
+ axi_spi_master_aw_region[3] axi_spi_master_aw_size[0] axi_spi_master_aw_size[1]
+ axi_spi_master_aw_size[2] axi_spi_master_aw_user[0] axi_spi_master_aw_user[1] axi_spi_master_aw_user[2]
+ axi_spi_master_aw_user[3] axi_spi_master_aw_user[4] axi_spi_master_aw_user[5] axi_spi_master_aw_valid
+ axi_spi_master_b_id[0] axi_spi_master_b_id[1] axi_spi_master_b_id[2] axi_spi_master_b_id[3]
+ axi_spi_master_b_id[4] axi_spi_master_b_id[5] axi_spi_master_b_ready axi_spi_master_b_resp[0]
+ axi_spi_master_b_resp[1] axi_spi_master_b_user[0] axi_spi_master_b_user[1] axi_spi_master_b_user[2]
+ axi_spi_master_b_user[3] axi_spi_master_b_user[4] axi_spi_master_b_user[5] axi_spi_master_b_valid
+ axi_spi_master_r_data[0] axi_spi_master_r_data[10] axi_spi_master_r_data[11] axi_spi_master_r_data[12]
+ axi_spi_master_r_data[13] axi_spi_master_r_data[14] axi_spi_master_r_data[15] axi_spi_master_r_data[16]
+ axi_spi_master_r_data[17] axi_spi_master_r_data[18] axi_spi_master_r_data[19] axi_spi_master_r_data[1]
+ axi_spi_master_r_data[20] axi_spi_master_r_data[21] axi_spi_master_r_data[22] axi_spi_master_r_data[23]
+ axi_spi_master_r_data[24] axi_spi_master_r_data[25] axi_spi_master_r_data[26] axi_spi_master_r_data[27]
+ axi_spi_master_r_data[28] axi_spi_master_r_data[29] axi_spi_master_r_data[2] axi_spi_master_r_data[30]
+ axi_spi_master_r_data[31] axi_spi_master_r_data[32] axi_spi_master_r_data[33] axi_spi_master_r_data[34]
+ axi_spi_master_r_data[35] axi_spi_master_r_data[36] axi_spi_master_r_data[37] axi_spi_master_r_data[38]
+ axi_spi_master_r_data[39] axi_spi_master_r_data[3] axi_spi_master_r_data[40] axi_spi_master_r_data[41]
+ axi_spi_master_r_data[42] axi_spi_master_r_data[43] axi_spi_master_r_data[44] axi_spi_master_r_data[45]
+ axi_spi_master_r_data[46] axi_spi_master_r_data[47] axi_spi_master_r_data[48] axi_spi_master_r_data[49]
+ axi_spi_master_r_data[4] axi_spi_master_r_data[50] axi_spi_master_r_data[51] axi_spi_master_r_data[52]
+ axi_spi_master_r_data[53] axi_spi_master_r_data[54] axi_spi_master_r_data[55] axi_spi_master_r_data[56]
+ axi_spi_master_r_data[57] axi_spi_master_r_data[58] axi_spi_master_r_data[59] axi_spi_master_r_data[5]
+ axi_spi_master_r_data[60] axi_spi_master_r_data[61] axi_spi_master_r_data[62] axi_spi_master_r_data[63]
+ axi_spi_master_r_data[6] axi_spi_master_r_data[7] axi_spi_master_r_data[8] axi_spi_master_r_data[9]
+ axi_spi_master_r_id[0] axi_spi_master_r_id[1] axi_spi_master_r_id[2] axi_spi_master_r_id[3]
+ axi_spi_master_r_id[4] axi_spi_master_r_id[5] axi_spi_master_r_last axi_spi_master_r_ready
+ axi_spi_master_r_resp[0] axi_spi_master_r_resp[1] axi_spi_master_r_user[0] axi_spi_master_r_user[1]
+ axi_spi_master_r_user[2] axi_spi_master_r_user[3] axi_spi_master_r_user[4] axi_spi_master_r_user[5]
+ axi_spi_master_r_valid axi_spi_master_w_data[0] axi_spi_master_w_data[10] axi_spi_master_w_data[11]
+ axi_spi_master_w_data[12] axi_spi_master_w_data[13] axi_spi_master_w_data[14] axi_spi_master_w_data[15]
+ axi_spi_master_w_data[16] axi_spi_master_w_data[17] axi_spi_master_w_data[18] axi_spi_master_w_data[19]
+ axi_spi_master_w_data[1] axi_spi_master_w_data[20] axi_spi_master_w_data[21] axi_spi_master_w_data[22]
+ axi_spi_master_w_data[23] axi_spi_master_w_data[24] axi_spi_master_w_data[25] axi_spi_master_w_data[26]
+ axi_spi_master_w_data[27] axi_spi_master_w_data[28] axi_spi_master_w_data[29] axi_spi_master_w_data[2]
+ axi_spi_master_w_data[30] axi_spi_master_w_data[31] axi_spi_master_w_data[32] axi_spi_master_w_data[33]
+ axi_spi_master_w_data[34] axi_spi_master_w_data[35] axi_spi_master_w_data[36] axi_spi_master_w_data[37]
+ axi_spi_master_w_data[38] axi_spi_master_w_data[39] axi_spi_master_w_data[3] axi_spi_master_w_data[40]
+ axi_spi_master_w_data[41] axi_spi_master_w_data[42] axi_spi_master_w_data[43] axi_spi_master_w_data[44]
+ axi_spi_master_w_data[45] axi_spi_master_w_data[46] axi_spi_master_w_data[47] axi_spi_master_w_data[48]
+ axi_spi_master_w_data[49] axi_spi_master_w_data[4] axi_spi_master_w_data[50] axi_spi_master_w_data[51]
+ axi_spi_master_w_data[52] axi_spi_master_w_data[53] axi_spi_master_w_data[54] axi_spi_master_w_data[55]
+ axi_spi_master_w_data[56] axi_spi_master_w_data[57] axi_spi_master_w_data[58] axi_spi_master_w_data[59]
+ axi_spi_master_w_data[5] axi_spi_master_w_data[60] axi_spi_master_w_data[61] axi_spi_master_w_data[62]
+ axi_spi_master_w_data[63] axi_spi_master_w_data[6] axi_spi_master_w_data[7] axi_spi_master_w_data[8]
+ axi_spi_master_w_data[9] axi_spi_master_w_last axi_spi_master_w_ready axi_spi_master_w_strb[0]
+ axi_spi_master_w_strb[1] axi_spi_master_w_strb[2] axi_spi_master_w_strb[3] axi_spi_master_w_strb[4]
+ axi_spi_master_w_strb[5] axi_spi_master_w_strb[6] axi_spi_master_w_strb[7] axi_spi_master_w_user[0]
+ axi_spi_master_w_user[1] axi_spi_master_w_user[2] axi_spi_master_w_user[3] axi_spi_master_w_user[4]
+ axi_spi_master_w_user[5] axi_spi_master_w_valid boot_addr_o[0] boot_addr_o[10] boot_addr_o[11]
+ boot_addr_o[12] boot_addr_o[13] boot_addr_o[14] boot_addr_o[15] boot_addr_o[16]
+ boot_addr_o[17] boot_addr_o[18] boot_addr_o[19] boot_addr_o[1] boot_addr_o[20] boot_addr_o[21]
+ boot_addr_o[22] boot_addr_o[23] boot_addr_o[24] boot_addr_o[25] boot_addr_o[26]
+ boot_addr_o[27] boot_addr_o[28] boot_addr_o[29] boot_addr_o[2] boot_addr_o[30] boot_addr_o[31]
+ boot_addr_o[3] boot_addr_o[4] boot_addr_o[5] boot_addr_o[6] boot_addr_o[7] boot_addr_o[8]
+ boot_addr_o[9] clk_gate_core_o clk_i clk_i_pll clk_o_pll clk_sel_i_pll clk_standalone_i_pll
+ core_busy_i debug_addr[0] debug_addr[10] debug_addr[11] debug_addr[12] debug_addr[13]
+ debug_addr[14] debug_addr[1] debug_addr[2] debug_addr[3] debug_addr[4] debug_addr[5]
+ debug_addr[6] debug_addr[7] debug_addr[8] debug_addr[9] debug_gnt debug_rdata[0]
+ debug_rdata[10] debug_rdata[11] debug_rdata[12] debug_rdata[13] debug_rdata[14]
+ debug_rdata[15] debug_rdata[16] debug_rdata[17] debug_rdata[18] debug_rdata[19]
+ debug_rdata[1] debug_rdata[20] debug_rdata[21] debug_rdata[22] debug_rdata[23] debug_rdata[24]
+ debug_rdata[25] debug_rdata[26] debug_rdata[27] debug_rdata[28] debug_rdata[29]
+ debug_rdata[2] debug_rdata[30] debug_rdata[31] debug_rdata[3] debug_rdata[4] debug_rdata[5]
+ debug_rdata[6] debug_rdata[7] debug_rdata[8] debug_rdata[9] debug_req debug_rvalid
+ debug_wdata[0] debug_wdata[10] debug_wdata[11] debug_wdata[12] debug_wdata[13] debug_wdata[14]
+ debug_wdata[15] debug_wdata[16] debug_wdata[17] debug_wdata[18] debug_wdata[19]
+ debug_wdata[1] debug_wdata[20] debug_wdata[21] debug_wdata[22] debug_wdata[23] debug_wdata[24]
+ debug_wdata[25] debug_wdata[26] debug_wdata[27] debug_wdata[28] debug_wdata[29]
+ debug_wdata[2] debug_wdata[30] debug_wdata[31] debug_wdata[3] debug_wdata[4] debug_wdata[5]
+ debug_wdata[6] debug_wdata[7] debug_wdata[8] debug_wdata[9] debug_we fetch_enable_i
+ fetch_enable_o fll1_ack_i fll1_add_o[0] fll1_add_o[1] fll1_lock_i fll1_rdata_i[0]
+ fll1_rdata_i[10] fll1_rdata_i[11] fll1_rdata_i[12] fll1_rdata_i[13] fll1_rdata_i[14]
+ fll1_rdata_i[15] fll1_rdata_i[16] fll1_rdata_i[17] fll1_rdata_i[18] fll1_rdata_i[19]
+ fll1_rdata_i[1] fll1_rdata_i[20] fll1_rdata_i[21] fll1_rdata_i[22] fll1_rdata_i[23]
+ fll1_rdata_i[24] fll1_rdata_i[25] fll1_rdata_i[26] fll1_rdata_i[27] fll1_rdata_i[28]
+ fll1_rdata_i[29] fll1_rdata_i[2] fll1_rdata_i[30] fll1_rdata_i[31] fll1_rdata_i[3]
+ fll1_rdata_i[4] fll1_rdata_i[5] fll1_rdata_i[6] fll1_rdata_i[7] fll1_rdata_i[8]
+ fll1_rdata_i[9] fll1_req_o fll1_wdata_o[0] fll1_wdata_o[10] fll1_wdata_o[11] fll1_wdata_o[12]
+ fll1_wdata_o[13] fll1_wdata_o[14] fll1_wdata_o[15] fll1_wdata_o[16] fll1_wdata_o[17]
+ fll1_wdata_o[18] fll1_wdata_o[19] fll1_wdata_o[1] fll1_wdata_o[20] fll1_wdata_o[21]
+ fll1_wdata_o[22] fll1_wdata_o[23] fll1_wdata_o[24] fll1_wdata_o[25] fll1_wdata_o[26]
+ fll1_wdata_o[27] fll1_wdata_o[28] fll1_wdata_o[29] fll1_wdata_o[2] fll1_wdata_o[30]
+ fll1_wdata_o[31] fll1_wdata_o[3] fll1_wdata_o[4] fll1_wdata_o[5] fll1_wdata_o[6]
+ fll1_wdata_o[7] fll1_wdata_o[8] fll1_wdata_o[9] fll1_wrn_o fll_ack_o_pll fll_add_i_pll[0]
+ fll_add_i_pll[1] fll_data_i_pll[0] fll_data_i_pll[10] fll_data_i_pll[11] fll_data_i_pll[12]
+ fll_data_i_pll[13] fll_data_i_pll[14] fll_data_i_pll[15] fll_data_i_pll[16] fll_data_i_pll[17]
+ fll_data_i_pll[18] fll_data_i_pll[19] fll_data_i_pll[1] fll_data_i_pll[20] fll_data_i_pll[21]
+ fll_data_i_pll[22] fll_data_i_pll[23] fll_data_i_pll[24] fll_data_i_pll[25] fll_data_i_pll[26]
+ fll_data_i_pll[27] fll_data_i_pll[28] fll_data_i_pll[29] fll_data_i_pll[2] fll_data_i_pll[30]
+ fll_data_i_pll[31] fll_data_i_pll[3] fll_data_i_pll[4] fll_data_i_pll[5] fll_data_i_pll[6]
+ fll_data_i_pll[7] fll_data_i_pll[8] fll_data_i_pll[9] fll_lock_o_pll fll_r_data_o_pll[0]
+ fll_r_data_o_pll[10] fll_r_data_o_pll[11] fll_r_data_o_pll[12] fll_r_data_o_pll[13]
+ fll_r_data_o_pll[14] fll_r_data_o_pll[15] fll_r_data_o_pll[16] fll_r_data_o_pll[17]
+ fll_r_data_o_pll[18] fll_r_data_o_pll[19] fll_r_data_o_pll[1] fll_r_data_o_pll[20]
+ fll_r_data_o_pll[21] fll_r_data_o_pll[22] fll_r_data_o_pll[23] fll_r_data_o_pll[24]
+ fll_r_data_o_pll[25] fll_r_data_o_pll[26] fll_r_data_o_pll[27] fll_r_data_o_pll[28]
+ fll_r_data_o_pll[29] fll_r_data_o_pll[2] fll_r_data_o_pll[30] fll_r_data_o_pll[31]
+ fll_r_data_o_pll[3] fll_r_data_o_pll[4] fll_r_data_o_pll[5] fll_r_data_o_pll[6]
+ fll_r_data_o_pll[7] fll_r_data_o_pll[8] fll_r_data_o_pll[9] fll_req_i_pll fll_wrn_i_pll
+ gpio_dir[0] gpio_dir[10] gpio_dir[11] gpio_dir[12] gpio_dir[13] gpio_dir[14] gpio_dir[15]
+ gpio_dir[16] gpio_dir[17] gpio_dir[18] gpio_dir[19] gpio_dir[1] gpio_dir[20] gpio_dir[21]
+ gpio_dir[22] gpio_dir[23] gpio_dir[24] gpio_dir[25] gpio_dir[26] gpio_dir[27] gpio_dir[28]
+ gpio_dir[29] gpio_dir[2] gpio_dir[30] gpio_dir[31] gpio_dir[3] gpio_dir[4] gpio_dir[5]
+ gpio_dir[6] gpio_dir[7] gpio_dir[8] gpio_dir[9] gpio_in[0] gpio_in[10] gpio_in[11]
+ gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18]
+ gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24]
+ gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30]
+ gpio_in[31] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15]
+ gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21]
+ gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28]
+ gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[3] gpio_out[4] gpio_out[5]
+ gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] gpio_padcfg[0] gpio_padcfg[100]
+ gpio_padcfg[101] gpio_padcfg[102] gpio_padcfg[103] gpio_padcfg[104] gpio_padcfg[105]
+ gpio_padcfg[106] gpio_padcfg[107] gpio_padcfg[108] gpio_padcfg[109] gpio_padcfg[10]
+ gpio_padcfg[110] gpio_padcfg[111] gpio_padcfg[112] gpio_padcfg[113] gpio_padcfg[114]
+ gpio_padcfg[115] gpio_padcfg[116] gpio_padcfg[117] gpio_padcfg[118] gpio_padcfg[119]
+ gpio_padcfg[11] gpio_padcfg[120] gpio_padcfg[121] gpio_padcfg[122] gpio_padcfg[123]
+ gpio_padcfg[124] gpio_padcfg[125] gpio_padcfg[126] gpio_padcfg[127] gpio_padcfg[128]
+ gpio_padcfg[129] gpio_padcfg[12] gpio_padcfg[130] gpio_padcfg[131] gpio_padcfg[132]
+ gpio_padcfg[133] gpio_padcfg[134] gpio_padcfg[135] gpio_padcfg[136] gpio_padcfg[137]
+ gpio_padcfg[138] gpio_padcfg[139] gpio_padcfg[13] gpio_padcfg[140] gpio_padcfg[141]
+ gpio_padcfg[142] gpio_padcfg[143] gpio_padcfg[144] gpio_padcfg[145] gpio_padcfg[146]
+ gpio_padcfg[147] gpio_padcfg[148] gpio_padcfg[149] gpio_padcfg[14] gpio_padcfg[150]
+ gpio_padcfg[151] gpio_padcfg[152] gpio_padcfg[153] gpio_padcfg[154] gpio_padcfg[155]
+ gpio_padcfg[156] gpio_padcfg[157] gpio_padcfg[158] gpio_padcfg[159] gpio_padcfg[15]
+ gpio_padcfg[160] gpio_padcfg[161] gpio_padcfg[162] gpio_padcfg[163] gpio_padcfg[164]
+ gpio_padcfg[165] gpio_padcfg[166] gpio_padcfg[167] gpio_padcfg[168] gpio_padcfg[169]
+ gpio_padcfg[16] gpio_padcfg[170] gpio_padcfg[171] gpio_padcfg[172] gpio_padcfg[173]
+ gpio_padcfg[174] gpio_padcfg[175] gpio_padcfg[176] gpio_padcfg[177] gpio_padcfg[178]
+ gpio_padcfg[179] gpio_padcfg[17] gpio_padcfg[180] gpio_padcfg[181] gpio_padcfg[182]
+ gpio_padcfg[183] gpio_padcfg[184] gpio_padcfg[185] gpio_padcfg[186] gpio_padcfg[187]
+ gpio_padcfg[188] gpio_padcfg[189] gpio_padcfg[18] gpio_padcfg[190] gpio_padcfg[191]
+ gpio_padcfg[19] gpio_padcfg[1] gpio_padcfg[20] gpio_padcfg[21] gpio_padcfg[22] gpio_padcfg[23]
+ gpio_padcfg[24] gpio_padcfg[25] gpio_padcfg[26] gpio_padcfg[27] gpio_padcfg[28]
+ gpio_padcfg[29] gpio_padcfg[2] gpio_padcfg[30] gpio_padcfg[31] gpio_padcfg[32] gpio_padcfg[33]
+ gpio_padcfg[34] gpio_padcfg[35] gpio_padcfg[36] gpio_padcfg[37] gpio_padcfg[38]
+ gpio_padcfg[39] gpio_padcfg[3] gpio_padcfg[40] gpio_padcfg[41] gpio_padcfg[42] gpio_padcfg[43]
+ gpio_padcfg[44] gpio_padcfg[45] gpio_padcfg[46] gpio_padcfg[47] gpio_padcfg[48]
+ gpio_padcfg[49] gpio_padcfg[4] gpio_padcfg[50] gpio_padcfg[51] gpio_padcfg[52] gpio_padcfg[53]
+ gpio_padcfg[54] gpio_padcfg[55] gpio_padcfg[56] gpio_padcfg[57] gpio_padcfg[58]
+ gpio_padcfg[59] gpio_padcfg[5] gpio_padcfg[60] gpio_padcfg[61] gpio_padcfg[62] gpio_padcfg[63]
+ gpio_padcfg[64] gpio_padcfg[65] gpio_padcfg[66] gpio_padcfg[67] gpio_padcfg[68]
+ gpio_padcfg[69] gpio_padcfg[6] gpio_padcfg[70] gpio_padcfg[71] gpio_padcfg[72] gpio_padcfg[73]
+ gpio_padcfg[74] gpio_padcfg[75] gpio_padcfg[76] gpio_padcfg[77] gpio_padcfg[78]
+ gpio_padcfg[79] gpio_padcfg[7] gpio_padcfg[80] gpio_padcfg[81] gpio_padcfg[82] gpio_padcfg[83]
+ gpio_padcfg[84] gpio_padcfg[85] gpio_padcfg[86] gpio_padcfg[87] gpio_padcfg[88]
+ gpio_padcfg[89] gpio_padcfg[8] gpio_padcfg[90] gpio_padcfg[91] gpio_padcfg[92] gpio_padcfg[93]
+ gpio_padcfg[94] gpio_padcfg[95] gpio_padcfg[96] gpio_padcfg[97] gpio_padcfg[98]
+ gpio_padcfg[99] gpio_padcfg[9] io_oeb_pll[0] io_oeb_pll[10] io_oeb_pll[11] io_oeb_pll[12]
+ io_oeb_pll[13] io_oeb_pll[14] io_oeb_pll[15] io_oeb_pll[16] io_oeb_pll[17] io_oeb_pll[18]
+ io_oeb_pll[19] io_oeb_pll[1] io_oeb_pll[20] io_oeb_pll[21] io_oeb_pll[22] io_oeb_pll[23]
+ io_oeb_pll[24] io_oeb_pll[25] io_oeb_pll[26] io_oeb_pll[27] io_oeb_pll[28] io_oeb_pll[29]
+ io_oeb_pll[2] io_oeb_pll[30] io_oeb_pll[31] io_oeb_pll[32] io_oeb_pll[33] io_oeb_pll[34]
+ io_oeb_pll[35] io_oeb_pll[36] io_oeb_pll[37] io_oeb_pll[3] io_oeb_pll[4] io_oeb_pll[5]
+ io_oeb_pll[6] io_oeb_pll[7] io_oeb_pll[8] io_oeb_pll[9] io_out_pll[0] io_out_pll[10]
+ io_out_pll[11] io_out_pll[12] io_out_pll[13] io_out_pll[14] io_out_pll[15] io_out_pll[16]
+ io_out_pll[17] io_out_pll[18] io_out_pll[19] io_out_pll[1] io_out_pll[20] io_out_pll[21]
+ io_out_pll[22] io_out_pll[23] io_out_pll[24] io_out_pll[25] io_out_pll[2] io_out_pll[3]
+ io_out_pll[4] io_out_pll[5] io_out_pll[6] io_out_pll[7] io_out_pll[8] io_out_pll[9]
+ irq_o[0] irq_o[10] irq_o[11] irq_o[12] irq_o[13] irq_o[14] irq_o[15] irq_o[16] irq_o[17]
+ irq_o[18] irq_o[19] irq_o[1] irq_o[20] irq_o[21] irq_o[22] irq_o[23] irq_o[24] irq_o[25]
+ irq_o[26] irq_o[27] irq_o[28] irq_o[29] irq_o[2] irq_o[30] irq_o[31] irq_o[3] irq_o[4]
+ irq_o[5] irq_o[6] irq_o[7] irq_o[8] irq_o[9] la_data_out_pll[0] la_data_out_pll[10]
+ la_data_out_pll[11] la_data_out_pll[12] la_data_out_pll[13] la_data_out_pll[14]
+ la_data_out_pll[15] la_data_out_pll[16] la_data_out_pll[17] la_data_out_pll[18]
+ la_data_out_pll[19] la_data_out_pll[1] la_data_out_pll[20] la_data_out_pll[21] la_data_out_pll[22]
+ la_data_out_pll[23] la_data_out_pll[24] la_data_out_pll[25] la_data_out_pll[26]
+ la_data_out_pll[27] la_data_out_pll[28] la_data_out_pll[29] la_data_out_pll[2] la_data_out_pll[30]
+ la_data_out_pll[31] la_data_out_pll[32] la_data_out_pll[33] la_data_out_pll[34]
+ la_data_out_pll[35] la_data_out_pll[36] la_data_out_pll[37] la_data_out_pll[38]
+ la_data_out_pll[39] la_data_out_pll[3] la_data_out_pll[40] la_data_out_pll[41] la_data_out_pll[42]
+ la_data_out_pll[43] la_data_out_pll[44] la_data_out_pll[45] la_data_out_pll[46]
+ la_data_out_pll[47] la_data_out_pll[48] la_data_out_pll[49] la_data_out_pll[4] la_data_out_pll[50]
+ la_data_out_pll[51] la_data_out_pll[52] la_data_out_pll[53] la_data_out_pll[54]
+ la_data_out_pll[55] la_data_out_pll[56] la_data_out_pll[57] la_data_out_pll[58]
+ la_data_out_pll[59] la_data_out_pll[5] la_data_out_pll[60] la_data_out_pll[61] la_data_out_pll[62]
+ la_data_out_pll[63] la_data_out_pll[6] la_data_out_pll[7] la_data_out_pll[8] la_data_out_pll[9]
+ rst_n rstn_i_pll rstn_o_pll scan_en_i_pll scan_i_pll scan_o_pll scl_pad_i scl_pad_o
+ scl_padoen_o sda_pad_i sda_pad_o sda_padoen_o slave_ar_addr[0] slave_ar_addr[10]
+ slave_ar_addr[11] slave_ar_addr[12] slave_ar_addr[13] slave_ar_addr[14] slave_ar_addr[15]
+ slave_ar_addr[16] slave_ar_addr[17] slave_ar_addr[18] slave_ar_addr[19] slave_ar_addr[1]
+ slave_ar_addr[20] slave_ar_addr[21] slave_ar_addr[22] slave_ar_addr[23] slave_ar_addr[24]
+ slave_ar_addr[25] slave_ar_addr[26] slave_ar_addr[27] slave_ar_addr[28] slave_ar_addr[29]
+ slave_ar_addr[2] slave_ar_addr[30] slave_ar_addr[31] slave_ar_addr[3] slave_ar_addr[4]
+ slave_ar_addr[5] slave_ar_addr[6] slave_ar_addr[7] slave_ar_addr[8] slave_ar_addr[9]
+ slave_ar_burst[0] slave_ar_burst[1] slave_ar_cache[0] slave_ar_cache[1] slave_ar_cache[2]
+ slave_ar_cache[3] slave_ar_id[0] slave_ar_id[1] slave_ar_id[2] slave_ar_id[3] slave_ar_id[4]
+ slave_ar_id[5] slave_ar_len[0] slave_ar_len[1] slave_ar_len[2] slave_ar_len[3] slave_ar_len[4]
+ slave_ar_len[5] slave_ar_len[6] slave_ar_len[7] slave_ar_lock slave_ar_prot[0] slave_ar_prot[1]
+ slave_ar_prot[2] slave_ar_qos[0] slave_ar_qos[1] slave_ar_qos[2] slave_ar_qos[3]
+ slave_ar_ready slave_ar_region[0] slave_ar_region[1] slave_ar_region[2] slave_ar_region[3]
+ slave_ar_size[0] slave_ar_size[1] slave_ar_size[2] slave_ar_user[0] slave_ar_user[1]
+ slave_ar_user[2] slave_ar_user[3] slave_ar_user[4] slave_ar_user[5] slave_ar_valid
+ slave_aw_addr[0] slave_aw_addr[10] slave_aw_addr[11] slave_aw_addr[12] slave_aw_addr[13]
+ slave_aw_addr[14] slave_aw_addr[15] slave_aw_addr[16] slave_aw_addr[17] slave_aw_addr[18]
+ slave_aw_addr[19] slave_aw_addr[1] slave_aw_addr[20] slave_aw_addr[21] slave_aw_addr[22]
+ slave_aw_addr[23] slave_aw_addr[24] slave_aw_addr[25] slave_aw_addr[26] slave_aw_addr[27]
+ slave_aw_addr[28] slave_aw_addr[29] slave_aw_addr[2] slave_aw_addr[30] slave_aw_addr[31]
+ slave_aw_addr[3] slave_aw_addr[4] slave_aw_addr[5] slave_aw_addr[6] slave_aw_addr[7]
+ slave_aw_addr[8] slave_aw_addr[9] slave_aw_burst[0] slave_aw_burst[1] slave_aw_cache[0]
+ slave_aw_cache[1] slave_aw_cache[2] slave_aw_cache[3] slave_aw_id[0] slave_aw_id[1]
+ slave_aw_id[2] slave_aw_id[3] slave_aw_id[4] slave_aw_id[5] slave_aw_len[0] slave_aw_len[1]
+ slave_aw_len[2] slave_aw_len[3] slave_aw_len[4] slave_aw_len[5] slave_aw_len[6]
+ slave_aw_len[7] slave_aw_lock slave_aw_prot[0] slave_aw_prot[1] slave_aw_prot[2]
+ slave_aw_qos[0] slave_aw_qos[1] slave_aw_qos[2] slave_aw_qos[3] slave_aw_ready slave_aw_region[0]
+ slave_aw_region[1] slave_aw_region[2] slave_aw_region[3] slave_aw_size[0] slave_aw_size[1]
+ slave_aw_size[2] slave_aw_user[0] slave_aw_user[1] slave_aw_user[2] slave_aw_user[3]
+ slave_aw_user[4] slave_aw_user[5] slave_aw_valid slave_b_id[0] slave_b_id[1] slave_b_id[2]
+ slave_b_id[3] slave_b_id[4] slave_b_id[5] slave_b_ready slave_b_resp[0] slave_b_resp[1]
+ slave_b_user[0] slave_b_user[1] slave_b_user[2] slave_b_user[3] slave_b_user[4]
+ slave_b_user[5] slave_b_valid slave_r_data[0] slave_r_data[10] slave_r_data[11]
+ slave_r_data[12] slave_r_data[13] slave_r_data[14] slave_r_data[15] slave_r_data[16]
+ slave_r_data[17] slave_r_data[18] slave_r_data[19] slave_r_data[1] slave_r_data[20]
+ slave_r_data[21] slave_r_data[22] slave_r_data[23] slave_r_data[24] slave_r_data[25]
+ slave_r_data[26] slave_r_data[27] slave_r_data[28] slave_r_data[29] slave_r_data[2]
+ slave_r_data[30] slave_r_data[31] slave_r_data[32] slave_r_data[33] slave_r_data[34]
+ slave_r_data[35] slave_r_data[36] slave_r_data[37] slave_r_data[38] slave_r_data[39]
+ slave_r_data[3] slave_r_data[40] slave_r_data[41] slave_r_data[42] slave_r_data[43]
+ slave_r_data[44] slave_r_data[45] slave_r_data[46] slave_r_data[47] slave_r_data[48]
+ slave_r_data[49] slave_r_data[4] slave_r_data[50] slave_r_data[51] slave_r_data[52]
+ slave_r_data[53] slave_r_data[54] slave_r_data[55] slave_r_data[56] slave_r_data[57]
+ slave_r_data[58] slave_r_data[59] slave_r_data[5] slave_r_data[60] slave_r_data[61]
+ slave_r_data[62] slave_r_data[63] slave_r_data[6] slave_r_data[7] slave_r_data[8]
+ slave_r_data[9] slave_r_id[0] slave_r_id[1] slave_r_id[2] slave_r_id[3] slave_r_id[4]
+ slave_r_id[5] slave_r_last slave_r_ready slave_r_resp[0] slave_r_resp[1] slave_r_user[0]
+ slave_r_user[1] slave_r_user[2] slave_r_user[3] slave_r_user[4] slave_r_user[5]
+ slave_r_valid slave_w_data[0] slave_w_data[10] slave_w_data[11] slave_w_data[12]
+ slave_w_data[13] slave_w_data[14] slave_w_data[15] slave_w_data[16] slave_w_data[17]
+ slave_w_data[18] slave_w_data[19] slave_w_data[1] slave_w_data[20] slave_w_data[21]
+ slave_w_data[22] slave_w_data[23] slave_w_data[24] slave_w_data[25] slave_w_data[26]
+ slave_w_data[27] slave_w_data[28] slave_w_data[29] slave_w_data[2] slave_w_data[30]
+ slave_w_data[31] slave_w_data[32] slave_w_data[33] slave_w_data[34] slave_w_data[35]
+ slave_w_data[36] slave_w_data[37] slave_w_data[38] slave_w_data[39] slave_w_data[3]
+ slave_w_data[40] slave_w_data[41] slave_w_data[42] slave_w_data[43] slave_w_data[44]
+ slave_w_data[45] slave_w_data[46] slave_w_data[47] slave_w_data[48] slave_w_data[49]
+ slave_w_data[4] slave_w_data[50] slave_w_data[51] slave_w_data[52] slave_w_data[53]
+ slave_w_data[54] slave_w_data[55] slave_w_data[56] slave_w_data[57] slave_w_data[58]
+ slave_w_data[59] slave_w_data[5] slave_w_data[60] slave_w_data[61] slave_w_data[62]
+ slave_w_data[63] slave_w_data[6] slave_w_data[7] slave_w_data[8] slave_w_data[9]
+ slave_w_last slave_w_ready slave_w_strb[0] slave_w_strb[1] slave_w_strb[2] slave_w_strb[3]
+ slave_w_strb[4] slave_w_strb[5] slave_w_strb[6] slave_w_strb[7] slave_w_user[0]
+ slave_w_user[1] slave_w_user[2] slave_w_user[3] slave_w_user[4] slave_w_user[5]
+ slave_w_valid spi_clk_i spi_cs_i spi_master_clk spi_master_csn0 spi_master_csn1
+ spi_master_csn2 spi_master_csn3 spi_master_mode[0] spi_master_mode[1] spi_master_sdi0
+ spi_master_sdi1 spi_master_sdi2 spi_master_sdi3 spi_master_sdo0 spi_master_sdo1
+ spi_master_sdo2 spi_master_sdo3 spi_mode_o[0] spi_mode_o[1] spi_sdi0_i spi_sdi1_i
+ spi_sdi2_i spi_sdi3_i spi_sdo0_o spi_sdo1_o spi_sdo2_o spi_sdo3_o testmode_i testmode_i_pll
+ uart_cts uart_dsr uart_dtr uart_rts uart_rx uart_tx user_irq_pll[0] user_irq_pll[1]
+ user_irq_pll[2] vccd1 vssd1 wbs_ack_o_pll wbs_dat_o_pll[0] wbs_dat_o_pll[10] wbs_dat_o_pll[11]
+ wbs_dat_o_pll[12] wbs_dat_o_pll[13] wbs_dat_o_pll[14] wbs_dat_o_pll[15] wbs_dat_o_pll[16]
+ wbs_dat_o_pll[17] wbs_dat_o_pll[18] wbs_dat_o_pll[19] wbs_dat_o_pll[1] wbs_dat_o_pll[20]
+ wbs_dat_o_pll[21] wbs_dat_o_pll[22] wbs_dat_o_pll[23] wbs_dat_o_pll[24] wbs_dat_o_pll[25]
+ wbs_dat_o_pll[26] wbs_dat_o_pll[27] wbs_dat_o_pll[28] wbs_dat_o_pll[29] wbs_dat_o_pll[2]
+ wbs_dat_o_pll[30] wbs_dat_o_pll[31] wbs_dat_o_pll[3] wbs_dat_o_pll[4] wbs_dat_o_pll[5]
+ wbs_dat_o_pll[6] wbs_dat_o_pll[7] wbs_dat_o_pll[8] wbs_dat_o_pll[9]
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xaxi_interconnect_i data_ram/clk0 axi_interconnect_i/m00_ar_addr[0] axi_interconnect_i/m00_ar_addr[10]
+ axi_interconnect_i/m00_ar_addr[11] axi_interconnect_i/m00_ar_addr[12] axi_interconnect_i/m00_ar_addr[13]
+ axi_interconnect_i/m00_ar_addr[14] axi_interconnect_i/m00_ar_addr[15] axi_interconnect_i/m00_ar_addr[16]
+ axi_interconnect_i/m00_ar_addr[17] axi_interconnect_i/m00_ar_addr[18] axi_interconnect_i/m00_ar_addr[19]
+ axi_interconnect_i/m00_ar_addr[1] axi_interconnect_i/m00_ar_addr[20] axi_interconnect_i/m00_ar_addr[21]
+ axi_interconnect_i/m00_ar_addr[22] axi_interconnect_i/m00_ar_addr[23] axi_interconnect_i/m00_ar_addr[24]
+ axi_interconnect_i/m00_ar_addr[25] axi_interconnect_i/m00_ar_addr[26] axi_interconnect_i/m00_ar_addr[27]
+ axi_interconnect_i/m00_ar_addr[28] axi_interconnect_i/m00_ar_addr[29] axi_interconnect_i/m00_ar_addr[2]
+ axi_interconnect_i/m00_ar_addr[30] axi_interconnect_i/m00_ar_addr[31] axi_interconnect_i/m00_ar_addr[3]
+ axi_interconnect_i/m00_ar_addr[4] axi_interconnect_i/m00_ar_addr[5] axi_interconnect_i/m00_ar_addr[6]
+ axi_interconnect_i/m00_ar_addr[7] axi_interconnect_i/m00_ar_addr[8] axi_interconnect_i/m00_ar_addr[9]
+ axi_interconnect_i/m00_ar_burst[0] axi_interconnect_i/m00_ar_burst[1] axi_interconnect_i/m00_ar_cache[0]
+ axi_interconnect_i/m00_ar_cache[1] axi_interconnect_i/m00_ar_cache[2] axi_interconnect_i/m00_ar_cache[3]
+ axi_interconnect_i/m00_ar_id[0] axi_interconnect_i/m00_ar_id[10] axi_interconnect_i/m00_ar_id[11]
+ axi_interconnect_i/m00_ar_id[1] axi_interconnect_i/m00_ar_id[2] axi_interconnect_i/m00_ar_id[3]
+ axi_interconnect_i/m00_ar_id[4] axi_interconnect_i/m00_ar_id[5] axi_interconnect_i/m00_ar_id[6]
+ axi_interconnect_i/m00_ar_id[7] axi_interconnect_i/m00_ar_id[8] axi_interconnect_i/m00_ar_id[9]
+ axi_interconnect_i/m00_ar_len[0] axi_interconnect_i/m00_ar_len[1] axi_interconnect_i/m00_ar_len[2]
+ axi_interconnect_i/m00_ar_len[3] axi_interconnect_i/m00_ar_len[4] axi_interconnect_i/m00_ar_len[5]
+ axi_interconnect_i/m00_ar_len[6] axi_interconnect_i/m00_ar_len[7] axi_interconnect_i/m00_ar_lock
+ axi_interconnect_i/m00_ar_prot[0] axi_interconnect_i/m00_ar_prot[1] axi_interconnect_i/m00_ar_prot[2]
+ axi_interconnect_i/m00_ar_qos[0] axi_interconnect_i/m00_ar_qos[1] axi_interconnect_i/m00_ar_qos[2]
+ axi_interconnect_i/m00_ar_qos[3] axi_interconnect_i/m00_ar_ready axi_interconnect_i/m00_ar_region[0]
+ axi_interconnect_i/m00_ar_region[1] axi_interconnect_i/m00_ar_region[2] axi_interconnect_i/m00_ar_region[3]
+ axi_interconnect_i/m00_ar_size[0] axi_interconnect_i/m00_ar_size[1] axi_interconnect_i/m00_ar_size[2]
+ axi_interconnect_i/m00_ar_user[-1] axi_interconnect_i/m00_ar_user[0] axi_interconnect_i/m00_ar_valid
+ axi_interconnect_i/m00_aw_addr[0] axi_interconnect_i/m00_aw_addr[10] axi_interconnect_i/m00_aw_addr[11]
+ axi_interconnect_i/m00_aw_addr[12] axi_interconnect_i/m00_aw_addr[13] axi_interconnect_i/m00_aw_addr[14]
+ axi_interconnect_i/m00_aw_addr[15] axi_interconnect_i/m00_aw_addr[16] axi_interconnect_i/m00_aw_addr[17]
+ axi_interconnect_i/m00_aw_addr[18] axi_interconnect_i/m00_aw_addr[19] axi_interconnect_i/m00_aw_addr[1]
+ axi_interconnect_i/m00_aw_addr[20] axi_interconnect_i/m00_aw_addr[21] axi_interconnect_i/m00_aw_addr[22]
+ axi_interconnect_i/m00_aw_addr[23] axi_interconnect_i/m00_aw_addr[24] axi_interconnect_i/m00_aw_addr[25]
+ axi_interconnect_i/m00_aw_addr[26] axi_interconnect_i/m00_aw_addr[27] axi_interconnect_i/m00_aw_addr[28]
+ axi_interconnect_i/m00_aw_addr[29] axi_interconnect_i/m00_aw_addr[2] axi_interconnect_i/m00_aw_addr[30]
+ axi_interconnect_i/m00_aw_addr[31] axi_interconnect_i/m00_aw_addr[3] axi_interconnect_i/m00_aw_addr[4]
+ axi_interconnect_i/m00_aw_addr[5] axi_interconnect_i/m00_aw_addr[6] axi_interconnect_i/m00_aw_addr[7]
+ axi_interconnect_i/m00_aw_addr[8] axi_interconnect_i/m00_aw_addr[9] axi_interconnect_i/m00_aw_burst[0]
+ axi_interconnect_i/m00_aw_burst[1] axi_interconnect_i/m00_aw_cache[0] axi_interconnect_i/m00_aw_cache[1]
+ axi_interconnect_i/m00_aw_cache[2] axi_interconnect_i/m00_aw_cache[3] axi_interconnect_i/m00_aw_id[0]
+ axi_interconnect_i/m00_aw_id[10] axi_interconnect_i/m00_aw_id[11] axi_interconnect_i/m00_aw_id[1]
+ axi_interconnect_i/m00_aw_id[2] axi_interconnect_i/m00_aw_id[3] axi_interconnect_i/m00_aw_id[4]
+ axi_interconnect_i/m00_aw_id[5] axi_interconnect_i/m00_aw_id[6] axi_interconnect_i/m00_aw_id[7]
+ axi_interconnect_i/m00_aw_id[8] axi_interconnect_i/m00_aw_id[9] axi_interconnect_i/m00_aw_len[0]
+ axi_interconnect_i/m00_aw_len[1] axi_interconnect_i/m00_aw_len[2] axi_interconnect_i/m00_aw_len[3]
+ axi_interconnect_i/m00_aw_len[4] axi_interconnect_i/m00_aw_len[5] axi_interconnect_i/m00_aw_len[6]
+ axi_interconnect_i/m00_aw_len[7] axi_interconnect_i/m00_aw_lock axi_interconnect_i/m00_aw_prot[0]
+ axi_interconnect_i/m00_aw_prot[1] axi_interconnect_i/m00_aw_prot[2] axi_interconnect_i/m00_aw_qos[0]
+ axi_interconnect_i/m00_aw_qos[1] axi_interconnect_i/m00_aw_qos[2] axi_interconnect_i/m00_aw_qos[3]
+ axi_interconnect_i/m00_aw_ready axi_interconnect_i/m00_aw_region[0] axi_interconnect_i/m00_aw_region[1]
+ axi_interconnect_i/m00_aw_region[2] axi_interconnect_i/m00_aw_region[3] axi_interconnect_i/m00_aw_size[0]
+ axi_interconnect_i/m00_aw_size[1] axi_interconnect_i/m00_aw_size[2] axi_interconnect_i/m00_aw_user[-1]
+ axi_interconnect_i/m00_aw_user[0] axi_interconnect_i/m00_aw_valid axi_interconnect_i/m00_b_id[0]
+ axi_interconnect_i/m00_b_id[10] axi_interconnect_i/m00_b_id[11] axi_interconnect_i/m00_b_id[1]
+ axi_interconnect_i/m00_b_id[2] axi_interconnect_i/m00_b_id[3] axi_interconnect_i/m00_b_id[4]
+ axi_interconnect_i/m00_b_id[5] axi_interconnect_i/m00_b_id[6] axi_interconnect_i/m00_b_id[7]
+ axi_interconnect_i/m00_b_id[8] axi_interconnect_i/m00_b_id[9] axi_interconnect_i/m00_b_ready
+ axi_interconnect_i/m00_b_resp[0] axi_interconnect_i/m00_b_resp[1] axi_interconnect_i/m00_b_user[-1]
+ axi_interconnect_i/m00_b_user[0] axi_interconnect_i/m00_b_valid axi_interconnect_i/m00_r_data[0]
+ axi_interconnect_i/m00_r_data[10] axi_interconnect_i/m00_r_data[11] axi_interconnect_i/m00_r_data[12]
+ axi_interconnect_i/m00_r_data[13] axi_interconnect_i/m00_r_data[14] axi_interconnect_i/m00_r_data[15]
+ axi_interconnect_i/m00_r_data[16] axi_interconnect_i/m00_r_data[17] axi_interconnect_i/m00_r_data[18]
+ axi_interconnect_i/m00_r_data[19] axi_interconnect_i/m00_r_data[1] axi_interconnect_i/m00_r_data[20]
+ axi_interconnect_i/m00_r_data[21] axi_interconnect_i/m00_r_data[22] axi_interconnect_i/m00_r_data[23]
+ axi_interconnect_i/m00_r_data[24] axi_interconnect_i/m00_r_data[25] axi_interconnect_i/m00_r_data[26]
+ axi_interconnect_i/m00_r_data[27] axi_interconnect_i/m00_r_data[28] axi_interconnect_i/m00_r_data[29]
+ axi_interconnect_i/m00_r_data[2] axi_interconnect_i/m00_r_data[30] axi_interconnect_i/m00_r_data[31]
+ axi_interconnect_i/m00_r_data[3] axi_interconnect_i/m00_r_data[4] axi_interconnect_i/m00_r_data[5]
+ axi_interconnect_i/m00_r_data[6] axi_interconnect_i/m00_r_data[7] axi_interconnect_i/m00_r_data[8]
+ axi_interconnect_i/m00_r_data[9] axi_interconnect_i/m00_r_id[0] axi_interconnect_i/m00_r_id[10]
+ axi_interconnect_i/m00_r_id[11] axi_interconnect_i/m00_r_id[1] axi_interconnect_i/m00_r_id[2]
+ axi_interconnect_i/m00_r_id[3] axi_interconnect_i/m00_r_id[4] axi_interconnect_i/m00_r_id[5]
+ axi_interconnect_i/m00_r_id[6] axi_interconnect_i/m00_r_id[7] axi_interconnect_i/m00_r_id[8]
+ axi_interconnect_i/m00_r_id[9] axi_interconnect_i/m00_r_last axi_interconnect_i/m00_r_ready
+ axi_interconnect_i/m00_r_resp[0] axi_interconnect_i/m00_r_resp[1] axi_interconnect_i/m00_r_user[-1]
+ axi_interconnect_i/m00_r_user[0] axi_interconnect_i/m00_r_valid axi_interconnect_i/m00_w_data[0]
+ axi_interconnect_i/m00_w_data[10] axi_interconnect_i/m00_w_data[11] axi_interconnect_i/m00_w_data[12]
+ axi_interconnect_i/m00_w_data[13] axi_interconnect_i/m00_w_data[14] axi_interconnect_i/m00_w_data[15]
+ axi_interconnect_i/m00_w_data[16] axi_interconnect_i/m00_w_data[17] axi_interconnect_i/m00_w_data[18]
+ axi_interconnect_i/m00_w_data[19] axi_interconnect_i/m00_w_data[1] axi_interconnect_i/m00_w_data[20]
+ axi_interconnect_i/m00_w_data[21] axi_interconnect_i/m00_w_data[22] axi_interconnect_i/m00_w_data[23]
+ axi_interconnect_i/m00_w_data[24] axi_interconnect_i/m00_w_data[25] axi_interconnect_i/m00_w_data[26]
+ axi_interconnect_i/m00_w_data[27] axi_interconnect_i/m00_w_data[28] axi_interconnect_i/m00_w_data[29]
+ axi_interconnect_i/m00_w_data[2] axi_interconnect_i/m00_w_data[30] axi_interconnect_i/m00_w_data[31]
+ axi_interconnect_i/m00_w_data[3] axi_interconnect_i/m00_w_data[4] axi_interconnect_i/m00_w_data[5]
+ axi_interconnect_i/m00_w_data[6] axi_interconnect_i/m00_w_data[7] axi_interconnect_i/m00_w_data[8]
+ axi_interconnect_i/m00_w_data[9] axi_interconnect_i/m00_w_last axi_interconnect_i/m00_w_ready
+ axi_interconnect_i/m00_w_strb[0] axi_interconnect_i/m00_w_strb[1] axi_interconnect_i/m00_w_strb[2]
+ axi_interconnect_i/m00_w_strb[3] axi_interconnect_i/m00_w_user[-1] axi_interconnect_i/m00_w_user[0]
+ axi_interconnect_i/m00_w_valid axi_interconnect_i/m01_ar_addr[0] axi_interconnect_i/m01_ar_addr[10]
+ axi_interconnect_i/m01_ar_addr[11] axi_interconnect_i/m01_ar_addr[12] axi_interconnect_i/m01_ar_addr[13]
+ axi_interconnect_i/m01_ar_addr[14] axi_interconnect_i/m01_ar_addr[15] axi_interconnect_i/m01_ar_addr[16]
+ axi_interconnect_i/m01_ar_addr[17] axi_interconnect_i/m01_ar_addr[18] axi_interconnect_i/m01_ar_addr[19]
+ axi_interconnect_i/m01_ar_addr[1] axi_interconnect_i/m01_ar_addr[20] axi_interconnect_i/m01_ar_addr[21]
+ axi_interconnect_i/m01_ar_addr[22] axi_interconnect_i/m01_ar_addr[23] axi_interconnect_i/m01_ar_addr[24]
+ axi_interconnect_i/m01_ar_addr[25] axi_interconnect_i/m01_ar_addr[26] axi_interconnect_i/m01_ar_addr[27]
+ axi_interconnect_i/m01_ar_addr[28] axi_interconnect_i/m01_ar_addr[29] axi_interconnect_i/m01_ar_addr[2]
+ axi_interconnect_i/m01_ar_addr[30] axi_interconnect_i/m01_ar_addr[31] axi_interconnect_i/m01_ar_addr[3]
+ axi_interconnect_i/m01_ar_addr[4] axi_interconnect_i/m01_ar_addr[5] axi_interconnect_i/m01_ar_addr[6]
+ axi_interconnect_i/m01_ar_addr[7] axi_interconnect_i/m01_ar_addr[8] axi_interconnect_i/m01_ar_addr[9]
+ axi_interconnect_i/m01_ar_burst[0] axi_interconnect_i/m01_ar_burst[1] axi_interconnect_i/m01_ar_cache[0]
+ axi_interconnect_i/m01_ar_cache[1] axi_interconnect_i/m01_ar_cache[2] axi_interconnect_i/m01_ar_cache[3]
+ axi_interconnect_i/m01_ar_id[0] axi_interconnect_i/m01_ar_id[10] axi_interconnect_i/m01_ar_id[11]
+ axi_interconnect_i/m01_ar_id[1] axi_interconnect_i/m01_ar_id[2] axi_interconnect_i/m01_ar_id[3]
+ axi_interconnect_i/m01_ar_id[4] axi_interconnect_i/m01_ar_id[5] axi_interconnect_i/m01_ar_id[6]
+ axi_interconnect_i/m01_ar_id[7] axi_interconnect_i/m01_ar_id[8] axi_interconnect_i/m01_ar_id[9]
+ axi_interconnect_i/m01_ar_len[0] axi_interconnect_i/m01_ar_len[1] axi_interconnect_i/m01_ar_len[2]
+ axi_interconnect_i/m01_ar_len[3] axi_interconnect_i/m01_ar_len[4] axi_interconnect_i/m01_ar_len[5]
+ axi_interconnect_i/m01_ar_len[6] axi_interconnect_i/m01_ar_len[7] axi_interconnect_i/m01_ar_lock
+ axi_interconnect_i/m01_ar_prot[0] axi_interconnect_i/m01_ar_prot[1] axi_interconnect_i/m01_ar_prot[2]
+ axi_interconnect_i/m01_ar_qos[0] axi_interconnect_i/m01_ar_qos[1] axi_interconnect_i/m01_ar_qos[2]
+ axi_interconnect_i/m01_ar_qos[3] axi_interconnect_i/m01_ar_ready axi_interconnect_i/m01_ar_region[0]
+ axi_interconnect_i/m01_ar_region[1] axi_interconnect_i/m01_ar_region[2] axi_interconnect_i/m01_ar_region[3]
+ axi_interconnect_i/m01_ar_size[0] axi_interconnect_i/m01_ar_size[1] axi_interconnect_i/m01_ar_size[2]
+ axi_interconnect_i/m01_ar_user[-1] axi_interconnect_i/m01_ar_user[0] axi_interconnect_i/m01_ar_valid
+ axi_interconnect_i/m01_aw_addr[0] axi_interconnect_i/m01_aw_addr[10] axi_interconnect_i/m01_aw_addr[11]
+ axi_interconnect_i/m01_aw_addr[12] axi_interconnect_i/m01_aw_addr[13] axi_interconnect_i/m01_aw_addr[14]
+ axi_interconnect_i/m01_aw_addr[15] axi_interconnect_i/m01_aw_addr[16] axi_interconnect_i/m01_aw_addr[17]
+ axi_interconnect_i/m01_aw_addr[18] axi_interconnect_i/m01_aw_addr[19] axi_interconnect_i/m01_aw_addr[1]
+ axi_interconnect_i/m01_aw_addr[20] axi_interconnect_i/m01_aw_addr[21] axi_interconnect_i/m01_aw_addr[22]
+ axi_interconnect_i/m01_aw_addr[23] axi_interconnect_i/m01_aw_addr[24] axi_interconnect_i/m01_aw_addr[25]
+ axi_interconnect_i/m01_aw_addr[26] axi_interconnect_i/m01_aw_addr[27] axi_interconnect_i/m01_aw_addr[28]
+ axi_interconnect_i/m01_aw_addr[29] axi_interconnect_i/m01_aw_addr[2] axi_interconnect_i/m01_aw_addr[30]
+ axi_interconnect_i/m01_aw_addr[31] axi_interconnect_i/m01_aw_addr[3] axi_interconnect_i/m01_aw_addr[4]
+ axi_interconnect_i/m01_aw_addr[5] axi_interconnect_i/m01_aw_addr[6] axi_interconnect_i/m01_aw_addr[7]
+ axi_interconnect_i/m01_aw_addr[8] axi_interconnect_i/m01_aw_addr[9] axi_interconnect_i/m01_aw_burst[0]
+ axi_interconnect_i/m01_aw_burst[1] axi_interconnect_i/m01_aw_cache[0] axi_interconnect_i/m01_aw_cache[1]
+ axi_interconnect_i/m01_aw_cache[2] axi_interconnect_i/m01_aw_cache[3] axi_interconnect_i/m01_aw_id[0]
+ axi_interconnect_i/m01_aw_id[10] axi_interconnect_i/m01_aw_id[11] axi_interconnect_i/m01_aw_id[1]
+ axi_interconnect_i/m01_aw_id[2] axi_interconnect_i/m01_aw_id[3] axi_interconnect_i/m01_aw_id[4]
+ axi_interconnect_i/m01_aw_id[5] axi_interconnect_i/m01_aw_id[6] axi_interconnect_i/m01_aw_id[7]
+ axi_interconnect_i/m01_aw_id[8] axi_interconnect_i/m01_aw_id[9] axi_interconnect_i/m01_aw_len[0]
+ axi_interconnect_i/m01_aw_len[1] axi_interconnect_i/m01_aw_len[2] axi_interconnect_i/m01_aw_len[3]
+ axi_interconnect_i/m01_aw_len[4] axi_interconnect_i/m01_aw_len[5] axi_interconnect_i/m01_aw_len[6]
+ axi_interconnect_i/m01_aw_len[7] axi_interconnect_i/m01_aw_lock axi_interconnect_i/m01_aw_prot[0]
+ axi_interconnect_i/m01_aw_prot[1] axi_interconnect_i/m01_aw_prot[2] axi_interconnect_i/m01_aw_qos[0]
+ axi_interconnect_i/m01_aw_qos[1] axi_interconnect_i/m01_aw_qos[2] axi_interconnect_i/m01_aw_qos[3]
+ axi_interconnect_i/m01_aw_ready axi_interconnect_i/m01_aw_region[0] axi_interconnect_i/m01_aw_region[1]
+ axi_interconnect_i/m01_aw_region[2] axi_interconnect_i/m01_aw_region[3] axi_interconnect_i/m01_aw_size[0]
+ axi_interconnect_i/m01_aw_size[1] axi_interconnect_i/m01_aw_size[2] axi_interconnect_i/m01_aw_user[-1]
+ axi_interconnect_i/m01_aw_user[0] axi_interconnect_i/m01_aw_valid axi_interconnect_i/m01_b_id[0]
+ axi_interconnect_i/m01_b_id[10] axi_interconnect_i/m01_b_id[11] axi_interconnect_i/m01_b_id[1]
+ axi_interconnect_i/m01_b_id[2] axi_interconnect_i/m01_b_id[3] axi_interconnect_i/m01_b_id[4]
+ axi_interconnect_i/m01_b_id[5] axi_interconnect_i/m01_b_id[6] axi_interconnect_i/m01_b_id[7]
+ axi_interconnect_i/m01_b_id[8] axi_interconnect_i/m01_b_id[9] axi_interconnect_i/m01_b_ready
+ axi_interconnect_i/m01_b_resp[0] axi_interconnect_i/m01_b_resp[1] axi_interconnect_i/m01_b_user[-1]
+ axi_interconnect_i/m01_b_user[0] axi_interconnect_i/m01_b_valid axi_interconnect_i/m01_r_data[0]
+ axi_interconnect_i/m01_r_data[10] axi_interconnect_i/m01_r_data[11] axi_interconnect_i/m01_r_data[12]
+ axi_interconnect_i/m01_r_data[13] axi_interconnect_i/m01_r_data[14] axi_interconnect_i/m01_r_data[15]
+ axi_interconnect_i/m01_r_data[16] axi_interconnect_i/m01_r_data[17] axi_interconnect_i/m01_r_data[18]
+ axi_interconnect_i/m01_r_data[19] axi_interconnect_i/m01_r_data[1] axi_interconnect_i/m01_r_data[20]
+ axi_interconnect_i/m01_r_data[21] axi_interconnect_i/m01_r_data[22] axi_interconnect_i/m01_r_data[23]
+ axi_interconnect_i/m01_r_data[24] axi_interconnect_i/m01_r_data[25] axi_interconnect_i/m01_r_data[26]
+ axi_interconnect_i/m01_r_data[27] axi_interconnect_i/m01_r_data[28] axi_interconnect_i/m01_r_data[29]
+ axi_interconnect_i/m01_r_data[2] axi_interconnect_i/m01_r_data[30] axi_interconnect_i/m01_r_data[31]
+ axi_interconnect_i/m01_r_data[3] axi_interconnect_i/m01_r_data[4] axi_interconnect_i/m01_r_data[5]
+ axi_interconnect_i/m01_r_data[6] axi_interconnect_i/m01_r_data[7] axi_interconnect_i/m01_r_data[8]
+ axi_interconnect_i/m01_r_data[9] axi_interconnect_i/m01_r_id[0] axi_interconnect_i/m01_r_id[10]
+ axi_interconnect_i/m01_r_id[11] axi_interconnect_i/m01_r_id[1] axi_interconnect_i/m01_r_id[2]
+ axi_interconnect_i/m01_r_id[3] axi_interconnect_i/m01_r_id[4] axi_interconnect_i/m01_r_id[5]
+ axi_interconnect_i/m01_r_id[6] axi_interconnect_i/m01_r_id[7] axi_interconnect_i/m01_r_id[8]
+ axi_interconnect_i/m01_r_id[9] axi_interconnect_i/m01_r_last axi_interconnect_i/m01_r_ready
+ axi_interconnect_i/m01_r_resp[0] axi_interconnect_i/m01_r_resp[1] axi_interconnect_i/m01_r_user[-1]
+ axi_interconnect_i/m01_r_user[0] axi_interconnect_i/m01_r_valid axi_interconnect_i/m01_w_data[0]
+ axi_interconnect_i/m01_w_data[10] axi_interconnect_i/m01_w_data[11] axi_interconnect_i/m01_w_data[12]
+ axi_interconnect_i/m01_w_data[13] axi_interconnect_i/m01_w_data[14] axi_interconnect_i/m01_w_data[15]
+ axi_interconnect_i/m01_w_data[16] axi_interconnect_i/m01_w_data[17] axi_interconnect_i/m01_w_data[18]
+ axi_interconnect_i/m01_w_data[19] axi_interconnect_i/m01_w_data[1] axi_interconnect_i/m01_w_data[20]
+ axi_interconnect_i/m01_w_data[21] axi_interconnect_i/m01_w_data[22] axi_interconnect_i/m01_w_data[23]
+ axi_interconnect_i/m01_w_data[24] axi_interconnect_i/m01_w_data[25] axi_interconnect_i/m01_w_data[26]
+ axi_interconnect_i/m01_w_data[27] axi_interconnect_i/m01_w_data[28] axi_interconnect_i/m01_w_data[29]
+ axi_interconnect_i/m01_w_data[2] axi_interconnect_i/m01_w_data[30] axi_interconnect_i/m01_w_data[31]
+ axi_interconnect_i/m01_w_data[3] axi_interconnect_i/m01_w_data[4] axi_interconnect_i/m01_w_data[5]
+ axi_interconnect_i/m01_w_data[6] axi_interconnect_i/m01_w_data[7] axi_interconnect_i/m01_w_data[8]
+ axi_interconnect_i/m01_w_data[9] axi_interconnect_i/m01_w_last axi_interconnect_i/m01_w_ready
+ axi_interconnect_i/m01_w_strb[0] axi_interconnect_i/m01_w_strb[1] axi_interconnect_i/m01_w_strb[2]
+ axi_interconnect_i/m01_w_strb[3] axi_interconnect_i/m01_w_user[-1] axi_interconnect_i/m01_w_user[0]
+ axi_interconnect_i/m01_w_valid peripherals_i/slave_ar_addr[0] peripherals_i/slave_ar_addr[10]
+ peripherals_i/slave_ar_addr[11] peripherals_i/slave_ar_addr[12] peripherals_i/slave_ar_addr[13]
+ peripherals_i/slave_ar_addr[14] peripherals_i/slave_ar_addr[15] peripherals_i/slave_ar_addr[16]
+ peripherals_i/slave_ar_addr[17] peripherals_i/slave_ar_addr[18] peripherals_i/slave_ar_addr[19]
+ peripherals_i/slave_ar_addr[1] peripherals_i/slave_ar_addr[20] peripherals_i/slave_ar_addr[21]
+ peripherals_i/slave_ar_addr[22] peripherals_i/slave_ar_addr[23] peripherals_i/slave_ar_addr[24]
+ peripherals_i/slave_ar_addr[25] peripherals_i/slave_ar_addr[26] peripherals_i/slave_ar_addr[27]
+ peripherals_i/slave_ar_addr[28] peripherals_i/slave_ar_addr[29] peripherals_i/slave_ar_addr[2]
+ peripherals_i/slave_ar_addr[30] peripherals_i/slave_ar_addr[31] peripherals_i/slave_ar_addr[3]
+ peripherals_i/slave_ar_addr[4] peripherals_i/slave_ar_addr[5] peripherals_i/slave_ar_addr[6]
+ peripherals_i/slave_ar_addr[7] peripherals_i/slave_ar_addr[8] peripherals_i/slave_ar_addr[9]
+ peripherals_i/slave_ar_burst[0] peripherals_i/slave_ar_burst[1] peripherals_i/slave_ar_cache[0]
+ peripherals_i/slave_ar_cache[1] peripherals_i/slave_ar_cache[2] peripherals_i/slave_ar_cache[3]
+ axi_interconnect_i/m02_ar_id[0] axi_interconnect_i/m02_ar_id[10] axi_interconnect_i/m02_ar_id[11]
+ axi_interconnect_i/m02_ar_id[1] axi_interconnect_i/m02_ar_id[2] axi_interconnect_i/m02_ar_id[3]
+ axi_interconnect_i/m02_ar_id[4] axi_interconnect_i/m02_ar_id[5] axi_interconnect_i/m02_ar_id[6]
+ axi_interconnect_i/m02_ar_id[7] axi_interconnect_i/m02_ar_id[8] axi_interconnect_i/m02_ar_id[9]
+ peripherals_i/slave_ar_len[0] peripherals_i/slave_ar_len[1] peripherals_i/slave_ar_len[2]
+ peripherals_i/slave_ar_len[3] peripherals_i/slave_ar_len[4] peripherals_i/slave_ar_len[5]
+ peripherals_i/slave_ar_len[6] peripherals_i/slave_ar_len[7] peripherals_i/slave_ar_lock
+ peripherals_i/slave_ar_prot[0] peripherals_i/slave_ar_prot[1] peripherals_i/slave_ar_prot[2]
+ peripherals_i/slave_ar_qos[0] peripherals_i/slave_ar_qos[1] peripherals_i/slave_ar_qos[2]
+ peripherals_i/slave_ar_qos[3] peripherals_i/slave_ar_ready peripherals_i/slave_ar_region[0]
+ peripherals_i/slave_ar_region[1] peripherals_i/slave_ar_region[2] peripherals_i/slave_ar_region[3]
+ peripherals_i/slave_ar_size[0] peripherals_i/slave_ar_size[1] peripherals_i/slave_ar_size[2]
+ axi_interconnect_i/m02_ar_user[-1] axi_interconnect_i/m02_ar_user[0] peripherals_i/slave_ar_valid
+ peripherals_i/slave_aw_addr[0] peripherals_i/slave_aw_addr[10] peripherals_i/slave_aw_addr[11]
+ peripherals_i/slave_aw_addr[12] peripherals_i/slave_aw_addr[13] peripherals_i/slave_aw_addr[14]
+ peripherals_i/slave_aw_addr[15] peripherals_i/slave_aw_addr[16] peripherals_i/slave_aw_addr[17]
+ peripherals_i/slave_aw_addr[18] peripherals_i/slave_aw_addr[19] peripherals_i/slave_aw_addr[1]
+ peripherals_i/slave_aw_addr[20] peripherals_i/slave_aw_addr[21] peripherals_i/slave_aw_addr[22]
+ peripherals_i/slave_aw_addr[23] peripherals_i/slave_aw_addr[24] peripherals_i/slave_aw_addr[25]
+ peripherals_i/slave_aw_addr[26] peripherals_i/slave_aw_addr[27] peripherals_i/slave_aw_addr[28]
+ peripherals_i/slave_aw_addr[29] peripherals_i/slave_aw_addr[2] peripherals_i/slave_aw_addr[30]
+ peripherals_i/slave_aw_addr[31] peripherals_i/slave_aw_addr[3] peripherals_i/slave_aw_addr[4]
+ peripherals_i/slave_aw_addr[5] peripherals_i/slave_aw_addr[6] peripherals_i/slave_aw_addr[7]
+ peripherals_i/slave_aw_addr[8] peripherals_i/slave_aw_addr[9] peripherals_i/slave_aw_burst[0]
+ peripherals_i/slave_aw_burst[1] peripherals_i/slave_aw_cache[0] peripherals_i/slave_aw_cache[1]
+ peripherals_i/slave_aw_cache[2] peripherals_i/slave_aw_cache[3] axi_interconnect_i/m02_aw_id[0]
+ axi_interconnect_i/m02_aw_id[10] axi_interconnect_i/m02_aw_id[11] axi_interconnect_i/m02_aw_id[1]
+ axi_interconnect_i/m02_aw_id[2] axi_interconnect_i/m02_aw_id[3] axi_interconnect_i/m02_aw_id[4]
+ axi_interconnect_i/m02_aw_id[5] axi_interconnect_i/m02_aw_id[6] axi_interconnect_i/m02_aw_id[7]
+ axi_interconnect_i/m02_aw_id[8] axi_interconnect_i/m02_aw_id[9] peripherals_i/slave_aw_len[0]
+ peripherals_i/slave_aw_len[1] peripherals_i/slave_aw_len[2] peripherals_i/slave_aw_len[3]
+ peripherals_i/slave_aw_len[4] peripherals_i/slave_aw_len[5] peripherals_i/slave_aw_len[6]
+ peripherals_i/slave_aw_len[7] peripherals_i/slave_aw_lock peripherals_i/slave_aw_prot[0]
+ peripherals_i/slave_aw_prot[1] peripherals_i/slave_aw_prot[2] peripherals_i/slave_aw_qos[0]
+ peripherals_i/slave_aw_qos[1] peripherals_i/slave_aw_qos[2] peripherals_i/slave_aw_qos[3]
+ peripherals_i/slave_aw_ready peripherals_i/slave_aw_region[0] peripherals_i/slave_aw_region[1]
+ peripherals_i/slave_aw_region[2] peripherals_i/slave_aw_region[3] peripherals_i/slave_aw_size[0]
+ peripherals_i/slave_aw_size[1] peripherals_i/slave_aw_size[2] axi_interconnect_i/m02_aw_user[-1]
+ axi_interconnect_i/m02_aw_user[0] peripherals_i/slave_aw_valid axi_interconnect_i/m02_b_id[0]
+ axi_interconnect_i/m02_b_id[10] axi_interconnect_i/m02_b_id[11] axi_interconnect_i/m02_b_id[1]
+ axi_interconnect_i/m02_b_id[2] axi_interconnect_i/m02_b_id[3] axi_interconnect_i/m02_b_id[4]
+ axi_interconnect_i/m02_b_id[5] axi_interconnect_i/m02_b_id[6] axi_interconnect_i/m02_b_id[7]
+ axi_interconnect_i/m02_b_id[8] axi_interconnect_i/m02_b_id[9] peripherals_i/slave_b_ready
+ peripherals_i/slave_b_resp[0] peripherals_i/slave_b_resp[1] axi_interconnect_i/m02_b_user[-1]
+ axi_interconnect_i/m02_b_user[0] peripherals_i/slave_b_valid axi_interconnect_i/m02_r_data[0]
+ axi_interconnect_i/m02_r_data[10] axi_interconnect_i/m02_r_data[11] axi_interconnect_i/m02_r_data[12]
+ axi_interconnect_i/m02_r_data[13] axi_interconnect_i/m02_r_data[14] axi_interconnect_i/m02_r_data[15]
+ axi_interconnect_i/m02_r_data[16] axi_interconnect_i/m02_r_data[17] axi_interconnect_i/m02_r_data[18]
+ axi_interconnect_i/m02_r_data[19] axi_interconnect_i/m02_r_data[1] axi_interconnect_i/m02_r_data[20]
+ axi_interconnect_i/m02_r_data[21] axi_interconnect_i/m02_r_data[22] axi_interconnect_i/m02_r_data[23]
+ axi_interconnect_i/m02_r_data[24] axi_interconnect_i/m02_r_data[25] axi_interconnect_i/m02_r_data[26]
+ axi_interconnect_i/m02_r_data[27] axi_interconnect_i/m02_r_data[28] axi_interconnect_i/m02_r_data[29]
+ axi_interconnect_i/m02_r_data[2] axi_interconnect_i/m02_r_data[30] axi_interconnect_i/m02_r_data[31]
+ axi_interconnect_i/m02_r_data[3] axi_interconnect_i/m02_r_data[4] axi_interconnect_i/m02_r_data[5]
+ axi_interconnect_i/m02_r_data[6] axi_interconnect_i/m02_r_data[7] axi_interconnect_i/m02_r_data[8]
+ axi_interconnect_i/m02_r_data[9] axi_interconnect_i/m02_r_id[0] axi_interconnect_i/m02_r_id[10]
+ axi_interconnect_i/m02_r_id[11] axi_interconnect_i/m02_r_id[1] axi_interconnect_i/m02_r_id[2]
+ axi_interconnect_i/m02_r_id[3] axi_interconnect_i/m02_r_id[4] axi_interconnect_i/m02_r_id[5]
+ axi_interconnect_i/m02_r_id[6] axi_interconnect_i/m02_r_id[7] axi_interconnect_i/m02_r_id[8]
+ axi_interconnect_i/m02_r_id[9] peripherals_i/slave_r_last peripherals_i/slave_r_ready
+ peripherals_i/slave_r_resp[0] peripherals_i/slave_r_resp[1] axi_interconnect_i/m02_r_user[-1]
+ axi_interconnect_i/m02_r_user[0] peripherals_i/slave_r_valid axi_interconnect_i/m02_w_data[0]
+ axi_interconnect_i/m02_w_data[10] axi_interconnect_i/m02_w_data[11] axi_interconnect_i/m02_w_data[12]
+ axi_interconnect_i/m02_w_data[13] axi_interconnect_i/m02_w_data[14] axi_interconnect_i/m02_w_data[15]
+ axi_interconnect_i/m02_w_data[16] axi_interconnect_i/m02_w_data[17] axi_interconnect_i/m02_w_data[18]
+ axi_interconnect_i/m02_w_data[19] axi_interconnect_i/m02_w_data[1] axi_interconnect_i/m02_w_data[20]
+ axi_interconnect_i/m02_w_data[21] axi_interconnect_i/m02_w_data[22] axi_interconnect_i/m02_w_data[23]
+ axi_interconnect_i/m02_w_data[24] axi_interconnect_i/m02_w_data[25] axi_interconnect_i/m02_w_data[26]
+ axi_interconnect_i/m02_w_data[27] axi_interconnect_i/m02_w_data[28] axi_interconnect_i/m02_w_data[29]
+ axi_interconnect_i/m02_w_data[2] axi_interconnect_i/m02_w_data[30] axi_interconnect_i/m02_w_data[31]
+ axi_interconnect_i/m02_w_data[3] axi_interconnect_i/m02_w_data[4] axi_interconnect_i/m02_w_data[5]
+ axi_interconnect_i/m02_w_data[6] axi_interconnect_i/m02_w_data[7] axi_interconnect_i/m02_w_data[8]
+ axi_interconnect_i/m02_w_data[9] peripherals_i/slave_w_last peripherals_i/slave_w_ready
+ axi_interconnect_i/m02_w_strb[0] axi_interconnect_i/m02_w_strb[1] axi_interconnect_i/m02_w_strb[2]
+ axi_interconnect_i/m02_w_strb[3] axi_interconnect_i/m02_w_user[-1] axi_interconnect_i/m02_w_user[0]
+ peripherals_i/slave_w_valid peripherals_i/rst_n axi_interconnect_i/s00_ar_addr[0]
+ axi_interconnect_i/s00_ar_addr[10] axi_interconnect_i/s00_ar_addr[11] axi_interconnect_i/s00_ar_addr[12]
+ axi_interconnect_i/s00_ar_addr[13] axi_interconnect_i/s00_ar_addr[14] axi_interconnect_i/s00_ar_addr[15]
+ axi_interconnect_i/s00_ar_addr[16] axi_interconnect_i/s00_ar_addr[17] axi_interconnect_i/s00_ar_addr[18]
+ axi_interconnect_i/s00_ar_addr[19] axi_interconnect_i/s00_ar_addr[1] axi_interconnect_i/s00_ar_addr[20]
+ axi_interconnect_i/s00_ar_addr[21] axi_interconnect_i/s00_ar_addr[22] axi_interconnect_i/s00_ar_addr[23]
+ axi_interconnect_i/s00_ar_addr[24] axi_interconnect_i/s00_ar_addr[25] axi_interconnect_i/s00_ar_addr[26]
+ axi_interconnect_i/s00_ar_addr[27] axi_interconnect_i/s00_ar_addr[28] axi_interconnect_i/s00_ar_addr[29]
+ axi_interconnect_i/s00_ar_addr[2] axi_interconnect_i/s00_ar_addr[30] axi_interconnect_i/s00_ar_addr[31]
+ axi_interconnect_i/s00_ar_addr[3] axi_interconnect_i/s00_ar_addr[4] axi_interconnect_i/s00_ar_addr[5]
+ axi_interconnect_i/s00_ar_addr[6] axi_interconnect_i/s00_ar_addr[7] axi_interconnect_i/s00_ar_addr[8]
+ axi_interconnect_i/s00_ar_addr[9] axi_interconnect_i/s00_ar_burst[0] axi_interconnect_i/s00_ar_burst[1]
+ axi_interconnect_i/s00_ar_cache[0] axi_interconnect_i/s00_ar_cache[1] axi_interconnect_i/s00_ar_cache[2]
+ axi_interconnect_i/s00_ar_cache[3] axi_interconnect_i/s00_ar_id[0] axi_interconnect_i/s00_ar_id[1]
+ axi_interconnect_i/s00_ar_id[2] axi_interconnect_i/s00_ar_id[3] axi_interconnect_i/s00_ar_id[4]
+ axi_interconnect_i/s00_ar_id[5] axi_interconnect_i/s00_ar_id[6] axi_interconnect_i/s00_ar_id[7]
+ axi_interconnect_i/s00_ar_id[8] axi_interconnect_i/s00_ar_id[9] axi_interconnect_i/s00_ar_len[0]
+ axi_interconnect_i/s00_ar_len[1] axi_interconnect_i/s00_ar_len[2] axi_interconnect_i/s00_ar_len[3]
+ axi_interconnect_i/s00_ar_len[4] axi_interconnect_i/s00_ar_len[5] axi_interconnect_i/s00_ar_len[6]
+ axi_interconnect_i/s00_ar_len[7] axi_interconnect_i/s00_ar_lock axi_interconnect_i/s00_ar_prot[0]
+ axi_interconnect_i/s00_ar_prot[1] axi_interconnect_i/s00_ar_prot[2] axi_interconnect_i/s00_ar_qos[0]
+ axi_interconnect_i/s00_ar_qos[1] axi_interconnect_i/s00_ar_qos[2] axi_interconnect_i/s00_ar_qos[3]
+ axi_interconnect_i/s00_ar_ready axi_interconnect_i/s00_ar_region[0] axi_interconnect_i/s00_ar_region[1]
+ axi_interconnect_i/s00_ar_region[2] axi_interconnect_i/s00_ar_region[3] axi_interconnect_i/s00_ar_size[0]
+ axi_interconnect_i/s00_ar_size[1] axi_interconnect_i/s00_ar_size[2] axi_interconnect_i/s00_ar_user[-1]
+ axi_interconnect_i/s00_ar_user[0] axi_interconnect_i/s00_ar_valid axi_interconnect_i/s00_aw_addr[0]
+ axi_interconnect_i/s00_aw_addr[10] axi_interconnect_i/s00_aw_addr[11] axi_interconnect_i/s00_aw_addr[12]
+ axi_interconnect_i/s00_aw_addr[13] axi_interconnect_i/s00_aw_addr[14] axi_interconnect_i/s00_aw_addr[15]
+ axi_interconnect_i/s00_aw_addr[16] axi_interconnect_i/s00_aw_addr[17] axi_interconnect_i/s00_aw_addr[18]
+ axi_interconnect_i/s00_aw_addr[19] axi_interconnect_i/s00_aw_addr[1] axi_interconnect_i/s00_aw_addr[20]
+ axi_interconnect_i/s00_aw_addr[21] axi_interconnect_i/s00_aw_addr[22] axi_interconnect_i/s00_aw_addr[23]
+ axi_interconnect_i/s00_aw_addr[24] axi_interconnect_i/s00_aw_addr[25] axi_interconnect_i/s00_aw_addr[26]
+ axi_interconnect_i/s00_aw_addr[27] axi_interconnect_i/s00_aw_addr[28] axi_interconnect_i/s00_aw_addr[29]
+ axi_interconnect_i/s00_aw_addr[2] axi_interconnect_i/s00_aw_addr[30] axi_interconnect_i/s00_aw_addr[31]
+ axi_interconnect_i/s00_aw_addr[3] axi_interconnect_i/s00_aw_addr[4] axi_interconnect_i/s00_aw_addr[5]
+ axi_interconnect_i/s00_aw_addr[6] axi_interconnect_i/s00_aw_addr[7] axi_interconnect_i/s00_aw_addr[8]
+ axi_interconnect_i/s00_aw_addr[9] axi_interconnect_i/s00_aw_burst[0] axi_interconnect_i/s00_aw_burst[1]
+ axi_interconnect_i/s00_aw_cache[0] axi_interconnect_i/s00_aw_cache[1] axi_interconnect_i/s00_aw_cache[2]
+ axi_interconnect_i/s00_aw_cache[3] axi_interconnect_i/s00_aw_id[0] axi_interconnect_i/s00_aw_id[1]
+ axi_interconnect_i/s00_aw_id[2] axi_interconnect_i/s00_aw_id[3] axi_interconnect_i/s00_aw_id[4]
+ axi_interconnect_i/s00_aw_id[5] axi_interconnect_i/s00_aw_id[6] axi_interconnect_i/s00_aw_id[7]
+ axi_interconnect_i/s00_aw_id[8] axi_interconnect_i/s00_aw_id[9] axi_interconnect_i/s00_aw_len[0]
+ axi_interconnect_i/s00_aw_len[1] axi_interconnect_i/s00_aw_len[2] axi_interconnect_i/s00_aw_len[3]
+ axi_interconnect_i/s00_aw_len[4] axi_interconnect_i/s00_aw_len[5] axi_interconnect_i/s00_aw_len[6]
+ axi_interconnect_i/s00_aw_len[7] axi_interconnect_i/s00_aw_lock axi_interconnect_i/s00_aw_prot[0]
+ axi_interconnect_i/s00_aw_prot[1] axi_interconnect_i/s00_aw_prot[2] axi_interconnect_i/s00_aw_qos[0]
+ axi_interconnect_i/s00_aw_qos[1] axi_interconnect_i/s00_aw_qos[2] axi_interconnect_i/s00_aw_qos[3]
+ axi_interconnect_i/s00_aw_ready axi_interconnect_i/s00_aw_region[0] axi_interconnect_i/s00_aw_region[1]
+ axi_interconnect_i/s00_aw_region[2] axi_interconnect_i/s00_aw_region[3] axi_interconnect_i/s00_aw_size[0]
+ axi_interconnect_i/s00_aw_size[1] axi_interconnect_i/s00_aw_size[2] axi_interconnect_i/s00_aw_user[-1]
+ axi_interconnect_i/s00_aw_user[0] axi_interconnect_i/s00_aw_valid axi_interconnect_i/s00_b_id[0]
+ axi_interconnect_i/s00_b_id[1] axi_interconnect_i/s00_b_id[2] axi_interconnect_i/s00_b_id[3]
+ axi_interconnect_i/s00_b_id[4] axi_interconnect_i/s00_b_id[5] axi_interconnect_i/s00_b_id[6]
+ axi_interconnect_i/s00_b_id[7] axi_interconnect_i/s00_b_id[8] axi_interconnect_i/s00_b_id[9]
+ axi_interconnect_i/s00_b_ready axi_interconnect_i/s00_b_resp[0] axi_interconnect_i/s00_b_resp[1]
+ axi_interconnect_i/s00_b_user[-1] axi_interconnect_i/s00_b_user[0] axi_interconnect_i/s00_b_valid
+ axi_interconnect_i/s00_r_data[0] axi_interconnect_i/s00_r_data[10] axi_interconnect_i/s00_r_data[11]
+ axi_interconnect_i/s00_r_data[12] axi_interconnect_i/s00_r_data[13] axi_interconnect_i/s00_r_data[14]
+ axi_interconnect_i/s00_r_data[15] axi_interconnect_i/s00_r_data[16] axi_interconnect_i/s00_r_data[17]
+ axi_interconnect_i/s00_r_data[18] axi_interconnect_i/s00_r_data[19] axi_interconnect_i/s00_r_data[1]
+ axi_interconnect_i/s00_r_data[20] axi_interconnect_i/s00_r_data[21] axi_interconnect_i/s00_r_data[22]
+ axi_interconnect_i/s00_r_data[23] axi_interconnect_i/s00_r_data[24] axi_interconnect_i/s00_r_data[25]
+ axi_interconnect_i/s00_r_data[26] axi_interconnect_i/s00_r_data[27] axi_interconnect_i/s00_r_data[28]
+ axi_interconnect_i/s00_r_data[29] axi_interconnect_i/s00_r_data[2] axi_interconnect_i/s00_r_data[30]
+ axi_interconnect_i/s00_r_data[31] axi_interconnect_i/s00_r_data[3] axi_interconnect_i/s00_r_data[4]
+ axi_interconnect_i/s00_r_data[5] axi_interconnect_i/s00_r_data[6] axi_interconnect_i/s00_r_data[7]
+ axi_interconnect_i/s00_r_data[8] axi_interconnect_i/s00_r_data[9] axi_interconnect_i/s00_r_id[0]
+ axi_interconnect_i/s00_r_id[1] axi_interconnect_i/s00_r_id[2] axi_interconnect_i/s00_r_id[3]
+ axi_interconnect_i/s00_r_id[4] axi_interconnect_i/s00_r_id[5] axi_interconnect_i/s00_r_id[6]
+ axi_interconnect_i/s00_r_id[7] axi_interconnect_i/s00_r_id[8] axi_interconnect_i/s00_r_id[9]
+ axi_interconnect_i/s00_r_last axi_interconnect_i/s00_r_ready axi_interconnect_i/s00_r_resp[0]
+ axi_interconnect_i/s00_r_resp[1] axi_interconnect_i/s00_r_user[-1] axi_interconnect_i/s00_r_user[0]
+ axi_interconnect_i/s00_r_valid axi_interconnect_i/s00_w_data[0] axi_interconnect_i/s00_w_data[10]
+ axi_interconnect_i/s00_w_data[11] axi_interconnect_i/s00_w_data[12] axi_interconnect_i/s00_w_data[13]
+ axi_interconnect_i/s00_w_data[14] axi_interconnect_i/s00_w_data[15] axi_interconnect_i/s00_w_data[16]
+ axi_interconnect_i/s00_w_data[17] axi_interconnect_i/s00_w_data[18] axi_interconnect_i/s00_w_data[19]
+ axi_interconnect_i/s00_w_data[1] axi_interconnect_i/s00_w_data[20] axi_interconnect_i/s00_w_data[21]
+ axi_interconnect_i/s00_w_data[22] axi_interconnect_i/s00_w_data[23] axi_interconnect_i/s00_w_data[24]
+ axi_interconnect_i/s00_w_data[25] axi_interconnect_i/s00_w_data[26] axi_interconnect_i/s00_w_data[27]
+ axi_interconnect_i/s00_w_data[28] axi_interconnect_i/s00_w_data[29] axi_interconnect_i/s00_w_data[2]
+ axi_interconnect_i/s00_w_data[30] axi_interconnect_i/s00_w_data[31] axi_interconnect_i/s00_w_data[3]
+ axi_interconnect_i/s00_w_data[4] axi_interconnect_i/s00_w_data[5] axi_interconnect_i/s00_w_data[6]
+ axi_interconnect_i/s00_w_data[7] axi_interconnect_i/s00_w_data[8] axi_interconnect_i/s00_w_data[9]
+ axi_interconnect_i/s00_w_last axi_interconnect_i/s00_w_ready axi_interconnect_i/s00_w_strb[0]
+ axi_interconnect_i/s00_w_strb[1] axi_interconnect_i/s00_w_strb[2] axi_interconnect_i/s00_w_strb[3]
+ axi_interconnect_i/s00_w_user[-1] axi_interconnect_i/s00_w_user[0] axi_interconnect_i/s00_w_valid
+ axi_interconnect_i/s01_ar_addr[0] axi_interconnect_i/s01_ar_addr[10] axi_interconnect_i/s01_ar_addr[11]
+ axi_interconnect_i/s01_ar_addr[12] axi_interconnect_i/s01_ar_addr[13] axi_interconnect_i/s01_ar_addr[14]
+ axi_interconnect_i/s01_ar_addr[15] axi_interconnect_i/s01_ar_addr[16] axi_interconnect_i/s01_ar_addr[17]
+ axi_interconnect_i/s01_ar_addr[18] axi_interconnect_i/s01_ar_addr[19] axi_interconnect_i/s01_ar_addr[1]
+ axi_interconnect_i/s01_ar_addr[20] axi_interconnect_i/s01_ar_addr[21] axi_interconnect_i/s01_ar_addr[22]
+ axi_interconnect_i/s01_ar_addr[23] axi_interconnect_i/s01_ar_addr[24] axi_interconnect_i/s01_ar_addr[25]
+ axi_interconnect_i/s01_ar_addr[26] axi_interconnect_i/s01_ar_addr[27] axi_interconnect_i/s01_ar_addr[28]
+ axi_interconnect_i/s01_ar_addr[29] axi_interconnect_i/s01_ar_addr[2] axi_interconnect_i/s01_ar_addr[30]
+ axi_interconnect_i/s01_ar_addr[31] axi_interconnect_i/s01_ar_addr[3] axi_interconnect_i/s01_ar_addr[4]
+ axi_interconnect_i/s01_ar_addr[5] axi_interconnect_i/s01_ar_addr[6] axi_interconnect_i/s01_ar_addr[7]
+ axi_interconnect_i/s01_ar_addr[8] axi_interconnect_i/s01_ar_addr[9] axi_interconnect_i/s01_ar_burst[0]
+ axi_interconnect_i/s01_ar_burst[1] axi_interconnect_i/s01_ar_cache[0] axi_interconnect_i/s01_ar_cache[1]
+ axi_interconnect_i/s01_ar_cache[2] axi_interconnect_i/s01_ar_cache[3] axi_interconnect_i/s01_ar_id[0]
+ axi_interconnect_i/s01_ar_id[1] axi_interconnect_i/s01_ar_id[2] axi_interconnect_i/s01_ar_id[3]
+ axi_interconnect_i/s01_ar_id[4] axi_interconnect_i/s01_ar_id[5] axi_interconnect_i/s01_ar_id[6]
+ axi_interconnect_i/s01_ar_id[7] axi_interconnect_i/s01_ar_id[8] axi_interconnect_i/s01_ar_id[9]
+ axi_interconnect_i/s01_ar_len[0] axi_interconnect_i/s01_ar_len[1] axi_interconnect_i/s01_ar_len[2]
+ axi_interconnect_i/s01_ar_len[3] axi_interconnect_i/s01_ar_len[4] axi_interconnect_i/s01_ar_len[5]
+ axi_interconnect_i/s01_ar_len[6] axi_interconnect_i/s01_ar_len[7] axi_interconnect_i/s01_ar_lock
+ axi_interconnect_i/s01_ar_prot[0] axi_interconnect_i/s01_ar_prot[1] axi_interconnect_i/s01_ar_prot[2]
+ axi_interconnect_i/s01_ar_qos[0] axi_interconnect_i/s01_ar_qos[1] axi_interconnect_i/s01_ar_qos[2]
+ axi_interconnect_i/s01_ar_qos[3] axi_interconnect_i/s01_ar_ready axi_interconnect_i/s01_ar_region[0]
+ axi_interconnect_i/s01_ar_region[1] axi_interconnect_i/s01_ar_region[2] axi_interconnect_i/s01_ar_region[3]
+ axi_interconnect_i/s01_ar_size[0] axi_interconnect_i/s01_ar_size[1] axi_interconnect_i/s01_ar_size[2]
+ axi_interconnect_i/s01_ar_user[-1] axi_interconnect_i/s01_ar_user[0] axi_interconnect_i/s01_ar_valid
+ axi_interconnect_i/s01_aw_addr[0] axi_interconnect_i/s01_aw_addr[10] axi_interconnect_i/s01_aw_addr[11]
+ axi_interconnect_i/s01_aw_addr[12] axi_interconnect_i/s01_aw_addr[13] axi_interconnect_i/s01_aw_addr[14]
+ axi_interconnect_i/s01_aw_addr[15] axi_interconnect_i/s01_aw_addr[16] axi_interconnect_i/s01_aw_addr[17]
+ axi_interconnect_i/s01_aw_addr[18] axi_interconnect_i/s01_aw_addr[19] axi_interconnect_i/s01_aw_addr[1]
+ axi_interconnect_i/s01_aw_addr[20] axi_interconnect_i/s01_aw_addr[21] axi_interconnect_i/s01_aw_addr[22]
+ axi_interconnect_i/s01_aw_addr[23] axi_interconnect_i/s01_aw_addr[24] axi_interconnect_i/s01_aw_addr[25]
+ axi_interconnect_i/s01_aw_addr[26] axi_interconnect_i/s01_aw_addr[27] axi_interconnect_i/s01_aw_addr[28]
+ axi_interconnect_i/s01_aw_addr[29] axi_interconnect_i/s01_aw_addr[2] axi_interconnect_i/s01_aw_addr[30]
+ axi_interconnect_i/s01_aw_addr[31] axi_interconnect_i/s01_aw_addr[3] axi_interconnect_i/s01_aw_addr[4]
+ axi_interconnect_i/s01_aw_addr[5] axi_interconnect_i/s01_aw_addr[6] axi_interconnect_i/s01_aw_addr[7]
+ axi_interconnect_i/s01_aw_addr[8] axi_interconnect_i/s01_aw_addr[9] axi_interconnect_i/s01_aw_burst[0]
+ axi_interconnect_i/s01_aw_burst[1] axi_interconnect_i/s01_aw_cache[0] axi_interconnect_i/s01_aw_cache[1]
+ axi_interconnect_i/s01_aw_cache[2] axi_interconnect_i/s01_aw_cache[3] axi_interconnect_i/s01_aw_id[0]
+ axi_interconnect_i/s01_aw_id[1] axi_interconnect_i/s01_aw_id[2] axi_interconnect_i/s01_aw_id[3]
+ axi_interconnect_i/s01_aw_id[4] axi_interconnect_i/s01_aw_id[5] axi_interconnect_i/s01_aw_id[6]
+ axi_interconnect_i/s01_aw_id[7] axi_interconnect_i/s01_aw_id[8] axi_interconnect_i/s01_aw_id[9]
+ axi_interconnect_i/s01_aw_len[0] axi_interconnect_i/s01_aw_len[1] axi_interconnect_i/s01_aw_len[2]
+ axi_interconnect_i/s01_aw_len[3] axi_interconnect_i/s01_aw_len[4] axi_interconnect_i/s01_aw_len[5]
+ axi_interconnect_i/s01_aw_len[6] axi_interconnect_i/s01_aw_len[7] axi_interconnect_i/s01_aw_lock
+ axi_interconnect_i/s01_aw_prot[0] axi_interconnect_i/s01_aw_prot[1] axi_interconnect_i/s01_aw_prot[2]
+ axi_interconnect_i/s01_aw_qos[0] axi_interconnect_i/s01_aw_qos[1] axi_interconnect_i/s01_aw_qos[2]
+ axi_interconnect_i/s01_aw_qos[3] axi_interconnect_i/s01_aw_ready axi_interconnect_i/s01_aw_region[0]
+ axi_interconnect_i/s01_aw_region[1] axi_interconnect_i/s01_aw_region[2] axi_interconnect_i/s01_aw_region[3]
+ axi_interconnect_i/s01_aw_size[0] axi_interconnect_i/s01_aw_size[1] axi_interconnect_i/s01_aw_size[2]
+ axi_interconnect_i/s01_aw_user[-1] axi_interconnect_i/s01_aw_user[0] axi_interconnect_i/s01_aw_valid
+ axi_interconnect_i/s01_b_id[0] axi_interconnect_i/s01_b_id[1] axi_interconnect_i/s01_b_id[2]
+ axi_interconnect_i/s01_b_id[3] axi_interconnect_i/s01_b_id[4] axi_interconnect_i/s01_b_id[5]
+ axi_interconnect_i/s01_b_id[6] axi_interconnect_i/s01_b_id[7] axi_interconnect_i/s01_b_id[8]
+ axi_interconnect_i/s01_b_id[9] axi_interconnect_i/s01_b_ready axi_interconnect_i/s01_b_resp[0]
+ axi_interconnect_i/s01_b_resp[1] axi_interconnect_i/s01_b_user[-1] axi_interconnect_i/s01_b_user[0]
+ axi_interconnect_i/s01_b_valid axi_interconnect_i/s01_r_data[0] axi_interconnect_i/s01_r_data[10]
+ axi_interconnect_i/s01_r_data[11] axi_interconnect_i/s01_r_data[12] axi_interconnect_i/s01_r_data[13]
+ axi_interconnect_i/s01_r_data[14] axi_interconnect_i/s01_r_data[15] axi_interconnect_i/s01_r_data[16]
+ axi_interconnect_i/s01_r_data[17] axi_interconnect_i/s01_r_data[18] axi_interconnect_i/s01_r_data[19]
+ axi_interconnect_i/s01_r_data[1] axi_interconnect_i/s01_r_data[20] axi_interconnect_i/s01_r_data[21]
+ axi_interconnect_i/s01_r_data[22] axi_interconnect_i/s01_r_data[23] axi_interconnect_i/s01_r_data[24]
+ axi_interconnect_i/s01_r_data[25] axi_interconnect_i/s01_r_data[26] axi_interconnect_i/s01_r_data[27]
+ axi_interconnect_i/s01_r_data[28] axi_interconnect_i/s01_r_data[29] axi_interconnect_i/s01_r_data[2]
+ axi_interconnect_i/s01_r_data[30] axi_interconnect_i/s01_r_data[31] axi_interconnect_i/s01_r_data[3]
+ axi_interconnect_i/s01_r_data[4] axi_interconnect_i/s01_r_data[5] axi_interconnect_i/s01_r_data[6]
+ axi_interconnect_i/s01_r_data[7] axi_interconnect_i/s01_r_data[8] axi_interconnect_i/s01_r_data[9]
+ axi_interconnect_i/s01_r_id[0] axi_interconnect_i/s01_r_id[1] axi_interconnect_i/s01_r_id[2]
+ axi_interconnect_i/s01_r_id[3] axi_interconnect_i/s01_r_id[4] axi_interconnect_i/s01_r_id[5]
+ axi_interconnect_i/s01_r_id[6] axi_interconnect_i/s01_r_id[7] axi_interconnect_i/s01_r_id[8]
+ axi_interconnect_i/s01_r_id[9] axi_interconnect_i/s01_r_last axi_interconnect_i/s01_r_ready
+ axi_interconnect_i/s01_r_resp[0] axi_interconnect_i/s01_r_resp[1] axi_interconnect_i/s01_r_user[-1]
+ axi_interconnect_i/s01_r_user[0] axi_interconnect_i/s01_r_valid axi_interconnect_i/s01_w_data[0]
+ axi_interconnect_i/s01_w_data[10] axi_interconnect_i/s01_w_data[11] axi_interconnect_i/s01_w_data[12]
+ axi_interconnect_i/s01_w_data[13] axi_interconnect_i/s01_w_data[14] axi_interconnect_i/s01_w_data[15]
+ axi_interconnect_i/s01_w_data[16] axi_interconnect_i/s01_w_data[17] axi_interconnect_i/s01_w_data[18]
+ axi_interconnect_i/s01_w_data[19] axi_interconnect_i/s01_w_data[1] axi_interconnect_i/s01_w_data[20]
+ axi_interconnect_i/s01_w_data[21] axi_interconnect_i/s01_w_data[22] axi_interconnect_i/s01_w_data[23]
+ axi_interconnect_i/s01_w_data[24] axi_interconnect_i/s01_w_data[25] axi_interconnect_i/s01_w_data[26]
+ axi_interconnect_i/s01_w_data[27] axi_interconnect_i/s01_w_data[28] axi_interconnect_i/s01_w_data[29]
+ axi_interconnect_i/s01_w_data[2] axi_interconnect_i/s01_w_data[30] axi_interconnect_i/s01_w_data[31]
+ axi_interconnect_i/s01_w_data[3] axi_interconnect_i/s01_w_data[4] axi_interconnect_i/s01_w_data[5]
+ axi_interconnect_i/s01_w_data[6] axi_interconnect_i/s01_w_data[7] axi_interconnect_i/s01_w_data[8]
+ axi_interconnect_i/s01_w_data[9] axi_interconnect_i/s01_w_last axi_interconnect_i/s01_w_ready
+ axi_interconnect_i/s01_w_strb[0] axi_interconnect_i/s01_w_strb[1] axi_interconnect_i/s01_w_strb[2]
+ axi_interconnect_i/s01_w_strb[3] axi_interconnect_i/s01_w_user[-1] axi_interconnect_i/s01_w_user[0]
+ axi_interconnect_i/s01_w_valid axi_interconnect_i/s02_ar_addr[0] axi_interconnect_i/s02_ar_addr[10]
+ axi_interconnect_i/s02_ar_addr[11] axi_interconnect_i/s02_ar_addr[12] axi_interconnect_i/s02_ar_addr[13]
+ axi_interconnect_i/s02_ar_addr[14] axi_interconnect_i/s02_ar_addr[15] axi_interconnect_i/s02_ar_addr[16]
+ axi_interconnect_i/s02_ar_addr[17] axi_interconnect_i/s02_ar_addr[18] axi_interconnect_i/s02_ar_addr[19]
+ axi_interconnect_i/s02_ar_addr[1] axi_interconnect_i/s02_ar_addr[20] axi_interconnect_i/s02_ar_addr[21]
+ axi_interconnect_i/s02_ar_addr[22] axi_interconnect_i/s02_ar_addr[23] axi_interconnect_i/s02_ar_addr[24]
+ axi_interconnect_i/s02_ar_addr[25] axi_interconnect_i/s02_ar_addr[26] axi_interconnect_i/s02_ar_addr[27]
+ axi_interconnect_i/s02_ar_addr[28] axi_interconnect_i/s02_ar_addr[29] axi_interconnect_i/s02_ar_addr[2]
+ axi_interconnect_i/s02_ar_addr[30] axi_interconnect_i/s02_ar_addr[31] axi_interconnect_i/s02_ar_addr[3]
+ axi_interconnect_i/s02_ar_addr[4] axi_interconnect_i/s02_ar_addr[5] axi_interconnect_i/s02_ar_addr[6]
+ axi_interconnect_i/s02_ar_addr[7] axi_interconnect_i/s02_ar_addr[8] axi_interconnect_i/s02_ar_addr[9]
+ axi_interconnect_i/s02_ar_burst[0] axi_interconnect_i/s02_ar_burst[1] axi_interconnect_i/s02_ar_cache[0]
+ axi_interconnect_i/s02_ar_cache[1] axi_interconnect_i/s02_ar_cache[2] axi_interconnect_i/s02_ar_cache[3]
+ axi_interconnect_i/s02_ar_id[0] axi_interconnect_i/s02_ar_id[1] axi_interconnect_i/s02_ar_id[2]
+ axi_interconnect_i/s02_ar_id[3] axi_interconnect_i/s02_ar_id[4] axi_interconnect_i/s02_ar_id[5]
+ axi_interconnect_i/s02_ar_id[6] axi_interconnect_i/s02_ar_id[7] axi_interconnect_i/s02_ar_id[8]
+ axi_interconnect_i/s02_ar_id[9] axi_interconnect_i/s02_ar_len[0] axi_interconnect_i/s02_ar_len[1]
+ axi_interconnect_i/s02_ar_len[2] axi_interconnect_i/s02_ar_len[3] axi_interconnect_i/s02_ar_len[4]
+ axi_interconnect_i/s02_ar_len[5] axi_interconnect_i/s02_ar_len[6] axi_interconnect_i/s02_ar_len[7]
+ axi_interconnect_i/s02_ar_lock axi_interconnect_i/s02_ar_prot[0] axi_interconnect_i/s02_ar_prot[1]
+ axi_interconnect_i/s02_ar_prot[2] axi_interconnect_i/s02_ar_qos[0] axi_interconnect_i/s02_ar_qos[1]
+ axi_interconnect_i/s02_ar_qos[2] axi_interconnect_i/s02_ar_qos[3] axi_interconnect_i/s02_ar_ready
+ axi_interconnect_i/s02_ar_region[0] axi_interconnect_i/s02_ar_region[1] axi_interconnect_i/s02_ar_region[2]
+ axi_interconnect_i/s02_ar_region[3] axi_interconnect_i/s02_ar_size[0] axi_interconnect_i/s02_ar_size[1]
+ axi_interconnect_i/s02_ar_size[2] axi_interconnect_i/s02_ar_user[-1] axi_interconnect_i/s02_ar_user[0]
+ axi_interconnect_i/s02_ar_valid axi_interconnect_i/s02_aw_addr[0] axi_interconnect_i/s02_aw_addr[10]
+ axi_interconnect_i/s02_aw_addr[11] axi_interconnect_i/s02_aw_addr[12] axi_interconnect_i/s02_aw_addr[13]
+ axi_interconnect_i/s02_aw_addr[14] axi_interconnect_i/s02_aw_addr[15] axi_interconnect_i/s02_aw_addr[16]
+ axi_interconnect_i/s02_aw_addr[17] axi_interconnect_i/s02_aw_addr[18] axi_interconnect_i/s02_aw_addr[19]
+ axi_interconnect_i/s02_aw_addr[1] axi_interconnect_i/s02_aw_addr[20] axi_interconnect_i/s02_aw_addr[21]
+ axi_interconnect_i/s02_aw_addr[22] axi_interconnect_i/s02_aw_addr[23] axi_interconnect_i/s02_aw_addr[24]
+ axi_interconnect_i/s02_aw_addr[25] axi_interconnect_i/s02_aw_addr[26] axi_interconnect_i/s02_aw_addr[27]
+ axi_interconnect_i/s02_aw_addr[28] axi_interconnect_i/s02_aw_addr[29] axi_interconnect_i/s02_aw_addr[2]
+ axi_interconnect_i/s02_aw_addr[30] axi_interconnect_i/s02_aw_addr[31] axi_interconnect_i/s02_aw_addr[3]
+ axi_interconnect_i/s02_aw_addr[4] axi_interconnect_i/s02_aw_addr[5] axi_interconnect_i/s02_aw_addr[6]
+ axi_interconnect_i/s02_aw_addr[7] axi_interconnect_i/s02_aw_addr[8] axi_interconnect_i/s02_aw_addr[9]
+ axi_interconnect_i/s02_aw_burst[0] axi_interconnect_i/s02_aw_burst[1] axi_interconnect_i/s02_aw_cache[0]
+ axi_interconnect_i/s02_aw_cache[1] axi_interconnect_i/s02_aw_cache[2] axi_interconnect_i/s02_aw_cache[3]
+ axi_interconnect_i/s02_aw_id[0] axi_interconnect_i/s02_aw_id[1] axi_interconnect_i/s02_aw_id[2]
+ axi_interconnect_i/s02_aw_id[3] axi_interconnect_i/s02_aw_id[4] axi_interconnect_i/s02_aw_id[5]
+ axi_interconnect_i/s02_aw_id[6] axi_interconnect_i/s02_aw_id[7] axi_interconnect_i/s02_aw_id[8]
+ axi_interconnect_i/s02_aw_id[9] axi_interconnect_i/s02_aw_len[0] axi_interconnect_i/s02_aw_len[1]
+ axi_interconnect_i/s02_aw_len[2] axi_interconnect_i/s02_aw_len[3] axi_interconnect_i/s02_aw_len[4]
+ axi_interconnect_i/s02_aw_len[5] axi_interconnect_i/s02_aw_len[6] axi_interconnect_i/s02_aw_len[7]
+ axi_interconnect_i/s02_aw_lock axi_interconnect_i/s02_aw_prot[0] axi_interconnect_i/s02_aw_prot[1]
+ axi_interconnect_i/s02_aw_prot[2] axi_interconnect_i/s02_aw_qos[0] axi_interconnect_i/s02_aw_qos[1]
+ axi_interconnect_i/s02_aw_qos[2] axi_interconnect_i/s02_aw_qos[3] axi_interconnect_i/s02_aw_ready
+ axi_interconnect_i/s02_aw_region[0] axi_interconnect_i/s02_aw_region[1] axi_interconnect_i/s02_aw_region[2]
+ axi_interconnect_i/s02_aw_region[3] axi_interconnect_i/s02_aw_size[0] axi_interconnect_i/s02_aw_size[1]
+ axi_interconnect_i/s02_aw_size[2] axi_interconnect_i/s02_aw_user[-1] axi_interconnect_i/s02_aw_user[0]
+ axi_interconnect_i/s02_aw_valid axi_interconnect_i/s02_b_id[0] axi_interconnect_i/s02_b_id[1]
+ axi_interconnect_i/s02_b_id[2] axi_interconnect_i/s02_b_id[3] axi_interconnect_i/s02_b_id[4]
+ axi_interconnect_i/s02_b_id[5] axi_interconnect_i/s02_b_id[6] axi_interconnect_i/s02_b_id[7]
+ axi_interconnect_i/s02_b_id[8] axi_interconnect_i/s02_b_id[9] axi_interconnect_i/s02_b_ready
+ axi_interconnect_i/s02_b_resp[0] axi_interconnect_i/s02_b_resp[1] axi_interconnect_i/s02_b_user[-1]
+ axi_interconnect_i/s02_b_user[0] axi_interconnect_i/s02_b_valid axi_interconnect_i/s02_r_data[0]
+ axi_interconnect_i/s02_r_data[10] axi_interconnect_i/s02_r_data[11] axi_interconnect_i/s02_r_data[12]
+ axi_interconnect_i/s02_r_data[13] axi_interconnect_i/s02_r_data[14] axi_interconnect_i/s02_r_data[15]
+ axi_interconnect_i/s02_r_data[16] axi_interconnect_i/s02_r_data[17] axi_interconnect_i/s02_r_data[18]
+ axi_interconnect_i/s02_r_data[19] axi_interconnect_i/s02_r_data[1] axi_interconnect_i/s02_r_data[20]
+ axi_interconnect_i/s02_r_data[21] axi_interconnect_i/s02_r_data[22] axi_interconnect_i/s02_r_data[23]
+ axi_interconnect_i/s02_r_data[24] axi_interconnect_i/s02_r_data[25] axi_interconnect_i/s02_r_data[26]
+ axi_interconnect_i/s02_r_data[27] axi_interconnect_i/s02_r_data[28] axi_interconnect_i/s02_r_data[29]
+ axi_interconnect_i/s02_r_data[2] axi_interconnect_i/s02_r_data[30] axi_interconnect_i/s02_r_data[31]
+ axi_interconnect_i/s02_r_data[3] axi_interconnect_i/s02_r_data[4] axi_interconnect_i/s02_r_data[5]
+ axi_interconnect_i/s02_r_data[6] axi_interconnect_i/s02_r_data[7] axi_interconnect_i/s02_r_data[8]
+ axi_interconnect_i/s02_r_data[9] axi_interconnect_i/s02_r_id[0] axi_interconnect_i/s02_r_id[1]
+ axi_interconnect_i/s02_r_id[2] axi_interconnect_i/s02_r_id[3] axi_interconnect_i/s02_r_id[4]
+ axi_interconnect_i/s02_r_id[5] axi_interconnect_i/s02_r_id[6] axi_interconnect_i/s02_r_id[7]
+ axi_interconnect_i/s02_r_id[8] axi_interconnect_i/s02_r_id[9] axi_interconnect_i/s02_r_last
+ axi_interconnect_i/s02_r_ready axi_interconnect_i/s02_r_resp[0] axi_interconnect_i/s02_r_resp[1]
+ axi_interconnect_i/s02_r_user[-1] axi_interconnect_i/s02_r_user[0] axi_interconnect_i/s02_r_valid
+ axi_interconnect_i/s02_w_data[0] axi_interconnect_i/s02_w_data[10] axi_interconnect_i/s02_w_data[11]
+ axi_interconnect_i/s02_w_data[12] axi_interconnect_i/s02_w_data[13] axi_interconnect_i/s02_w_data[14]
+ axi_interconnect_i/s02_w_data[15] axi_interconnect_i/s02_w_data[16] axi_interconnect_i/s02_w_data[17]
+ axi_interconnect_i/s02_w_data[18] axi_interconnect_i/s02_w_data[19] axi_interconnect_i/s02_w_data[1]
+ axi_interconnect_i/s02_w_data[20] axi_interconnect_i/s02_w_data[21] axi_interconnect_i/s02_w_data[22]
+ axi_interconnect_i/s02_w_data[23] axi_interconnect_i/s02_w_data[24] axi_interconnect_i/s02_w_data[25]
+ axi_interconnect_i/s02_w_data[26] axi_interconnect_i/s02_w_data[27] axi_interconnect_i/s02_w_data[28]
+ axi_interconnect_i/s02_w_data[29] axi_interconnect_i/s02_w_data[2] axi_interconnect_i/s02_w_data[30]
+ axi_interconnect_i/s02_w_data[31] axi_interconnect_i/s02_w_data[3] axi_interconnect_i/s02_w_data[4]
+ axi_interconnect_i/s02_w_data[5] axi_interconnect_i/s02_w_data[6] axi_interconnect_i/s02_w_data[7]
+ axi_interconnect_i/s02_w_data[8] axi_interconnect_i/s02_w_data[9] axi_interconnect_i/s02_w_last
+ axi_interconnect_i/s02_w_ready axi_interconnect_i/s02_w_strb[0] axi_interconnect_i/s02_w_strb[1]
+ axi_interconnect_i/s02_w_strb[2] axi_interconnect_i/s02_w_strb[3] axi_interconnect_i/s02_w_user[-1]
+ axi_interconnect_i/s02_w_user[0] axi_interconnect_i/s02_w_valid la_data_in[2] vccd1
+ vssd1 axi_node_intf_wrap
Xcore_region_i peripherals_i/boot_addr_o[0] peripherals_i/boot_addr_o[10] peripherals_i/boot_addr_o[11]
+ peripherals_i/boot_addr_o[12] peripherals_i/boot_addr_o[13] peripherals_i/boot_addr_o[14]
+ peripherals_i/boot_addr_o[15] peripherals_i/boot_addr_o[16] peripherals_i/boot_addr_o[17]
+ peripherals_i/boot_addr_o[18] peripherals_i/boot_addr_o[19] peripherals_i/boot_addr_o[1]
+ peripherals_i/boot_addr_o[20] peripherals_i/boot_addr_o[21] peripherals_i/boot_addr_o[22]
+ peripherals_i/boot_addr_o[23] peripherals_i/boot_addr_o[24] peripherals_i/boot_addr_o[25]
+ peripherals_i/boot_addr_o[26] peripherals_i/boot_addr_o[27] peripherals_i/boot_addr_o[28]
+ peripherals_i/boot_addr_o[29] peripherals_i/boot_addr_o[2] peripherals_i/boot_addr_o[30]
+ peripherals_i/boot_addr_o[31] peripherals_i/boot_addr_o[3] peripherals_i/boot_addr_o[4]
+ peripherals_i/boot_addr_o[5] peripherals_i/boot_addr_o[6] peripherals_i/boot_addr_o[7]
+ peripherals_i/boot_addr_o[8] peripherals_i/boot_addr_o[9] data_ram/clk0 core_region_i/clock_gating_i
+ peripherals_i/core_busy_i axi_interconnect_i/s00_ar_addr[0] axi_interconnect_i/s00_ar_addr[10]
+ axi_interconnect_i/s00_ar_addr[11] axi_interconnect_i/s00_ar_addr[12] axi_interconnect_i/s00_ar_addr[13]
+ axi_interconnect_i/s00_ar_addr[14] axi_interconnect_i/s00_ar_addr[15] axi_interconnect_i/s00_ar_addr[16]
+ axi_interconnect_i/s00_ar_addr[17] axi_interconnect_i/s00_ar_addr[18] axi_interconnect_i/s00_ar_addr[19]
+ axi_interconnect_i/s00_ar_addr[1] axi_interconnect_i/s00_ar_addr[20] axi_interconnect_i/s00_ar_addr[21]
+ axi_interconnect_i/s00_ar_addr[22] axi_interconnect_i/s00_ar_addr[23] axi_interconnect_i/s00_ar_addr[24]
+ axi_interconnect_i/s00_ar_addr[25] axi_interconnect_i/s00_ar_addr[26] axi_interconnect_i/s00_ar_addr[27]
+ axi_interconnect_i/s00_ar_addr[28] axi_interconnect_i/s00_ar_addr[29] axi_interconnect_i/s00_ar_addr[2]
+ axi_interconnect_i/s00_ar_addr[30] axi_interconnect_i/s00_ar_addr[31] axi_interconnect_i/s00_ar_addr[3]
+ axi_interconnect_i/s00_ar_addr[4] axi_interconnect_i/s00_ar_addr[5] axi_interconnect_i/s00_ar_addr[6]
+ axi_interconnect_i/s00_ar_addr[7] axi_interconnect_i/s00_ar_addr[8] axi_interconnect_i/s00_ar_addr[9]
+ axi_interconnect_i/s00_ar_burst[0] axi_interconnect_i/s00_ar_burst[1] axi_interconnect_i/s00_ar_cache[0]
+ axi_interconnect_i/s00_ar_cache[1] axi_interconnect_i/s00_ar_cache[2] axi_interconnect_i/s00_ar_cache[3]
+ core_region_i/core_master_ar_id[0] core_region_i/core_master_ar_id[1] core_region_i/core_master_ar_id[2]
+ core_region_i/core_master_ar_id[3] core_region_i/core_master_ar_id[4] core_region_i/core_master_ar_id[5]
+ core_region_i/core_master_ar_id[6] core_region_i/core_master_ar_id[7] core_region_i/core_master_ar_id[8]
+ core_region_i/core_master_ar_id[9] axi_interconnect_i/s00_ar_len[0] axi_interconnect_i/s00_ar_len[1]
+ axi_interconnect_i/s00_ar_len[2] axi_interconnect_i/s00_ar_len[3] axi_interconnect_i/s00_ar_len[4]
+ axi_interconnect_i/s00_ar_len[5] axi_interconnect_i/s00_ar_len[6] axi_interconnect_i/s00_ar_len[7]
+ axi_interconnect_i/s00_ar_lock axi_interconnect_i/s00_ar_prot[0] axi_interconnect_i/s00_ar_prot[1]
+ axi_interconnect_i/s00_ar_prot[2] axi_interconnect_i/s00_ar_qos[0] axi_interconnect_i/s00_ar_qos[1]
+ axi_interconnect_i/s00_ar_qos[2] axi_interconnect_i/s00_ar_qos[3] axi_interconnect_i/s00_ar_ready
+ axi_interconnect_i/s00_ar_region[0] axi_interconnect_i/s00_ar_region[1] axi_interconnect_i/s00_ar_region[2]
+ axi_interconnect_i/s00_ar_region[3] axi_interconnect_i/s00_ar_size[0] axi_interconnect_i/s00_ar_size[1]
+ axi_interconnect_i/s00_ar_size[2] core_region_i/core_master_ar_user[-1] core_region_i/core_master_ar_user[0]
+ axi_interconnect_i/s00_ar_valid axi_interconnect_i/s00_aw_addr[0] axi_interconnect_i/s00_aw_addr[10]
+ axi_interconnect_i/s00_aw_addr[11] axi_interconnect_i/s00_aw_addr[12] axi_interconnect_i/s00_aw_addr[13]
+ axi_interconnect_i/s00_aw_addr[14] axi_interconnect_i/s00_aw_addr[15] axi_interconnect_i/s00_aw_addr[16]
+ axi_interconnect_i/s00_aw_addr[17] axi_interconnect_i/s00_aw_addr[18] axi_interconnect_i/s00_aw_addr[19]
+ axi_interconnect_i/s00_aw_addr[1] axi_interconnect_i/s00_aw_addr[20] axi_interconnect_i/s00_aw_addr[21]
+ axi_interconnect_i/s00_aw_addr[22] axi_interconnect_i/s00_aw_addr[23] axi_interconnect_i/s00_aw_addr[24]
+ axi_interconnect_i/s00_aw_addr[25] axi_interconnect_i/s00_aw_addr[26] axi_interconnect_i/s00_aw_addr[27]
+ axi_interconnect_i/s00_aw_addr[28] axi_interconnect_i/s00_aw_addr[29] axi_interconnect_i/s00_aw_addr[2]
+ axi_interconnect_i/s00_aw_addr[30] axi_interconnect_i/s00_aw_addr[31] axi_interconnect_i/s00_aw_addr[3]
+ axi_interconnect_i/s00_aw_addr[4] axi_interconnect_i/s00_aw_addr[5] axi_interconnect_i/s00_aw_addr[6]
+ axi_interconnect_i/s00_aw_addr[7] axi_interconnect_i/s00_aw_addr[8] axi_interconnect_i/s00_aw_addr[9]
+ axi_interconnect_i/s00_aw_burst[0] axi_interconnect_i/s00_aw_burst[1] axi_interconnect_i/s00_aw_cache[0]
+ axi_interconnect_i/s00_aw_cache[1] axi_interconnect_i/s00_aw_cache[2] axi_interconnect_i/s00_aw_cache[3]
+ core_region_i/core_master_aw_id[0] core_region_i/core_master_aw_id[1] core_region_i/core_master_aw_id[2]
+ core_region_i/core_master_aw_id[3] core_region_i/core_master_aw_id[4] core_region_i/core_master_aw_id[5]
+ core_region_i/core_master_aw_id[6] core_region_i/core_master_aw_id[7] core_region_i/core_master_aw_id[8]
+ core_region_i/core_master_aw_id[9] axi_interconnect_i/s00_aw_len[0] axi_interconnect_i/s00_aw_len[1]
+ axi_interconnect_i/s00_aw_len[2] axi_interconnect_i/s00_aw_len[3] axi_interconnect_i/s00_aw_len[4]
+ axi_interconnect_i/s00_aw_len[5] axi_interconnect_i/s00_aw_len[6] axi_interconnect_i/s00_aw_len[7]
+ axi_interconnect_i/s00_aw_lock axi_interconnect_i/s00_aw_prot[0] axi_interconnect_i/s00_aw_prot[1]
+ axi_interconnect_i/s00_aw_prot[2] axi_interconnect_i/s00_aw_qos[0] axi_interconnect_i/s00_aw_qos[1]
+ axi_interconnect_i/s00_aw_qos[2] axi_interconnect_i/s00_aw_qos[3] axi_interconnect_i/s00_aw_ready
+ axi_interconnect_i/s00_aw_region[0] axi_interconnect_i/s00_aw_region[1] axi_interconnect_i/s00_aw_region[2]
+ axi_interconnect_i/s00_aw_region[3] axi_interconnect_i/s00_aw_size[0] axi_interconnect_i/s00_aw_size[1]
+ axi_interconnect_i/s00_aw_size[2] core_region_i/core_master_aw_user[-1] core_region_i/core_master_aw_user[0]
+ axi_interconnect_i/s00_aw_valid core_region_i/core_master_b_id[0] core_region_i/core_master_b_id[1]
+ core_region_i/core_master_b_id[2] core_region_i/core_master_b_id[3] core_region_i/core_master_b_id[4]
+ core_region_i/core_master_b_id[5] core_region_i/core_master_b_id[6] core_region_i/core_master_b_id[7]
+ core_region_i/core_master_b_id[8] core_region_i/core_master_b_id[9] axi_interconnect_i/s00_b_ready
+ axi_interconnect_i/s00_b_resp[0] axi_interconnect_i/s00_b_resp[1] core_region_i/core_master_b_user[-1]
+ core_region_i/core_master_b_user[0] axi_interconnect_i/s00_b_valid core_region_i/core_master_r_data[0]
+ core_region_i/core_master_r_data[10] core_region_i/core_master_r_data[11] core_region_i/core_master_r_data[12]
+ core_region_i/core_master_r_data[13] core_region_i/core_master_r_data[14] core_region_i/core_master_r_data[15]
+ core_region_i/core_master_r_data[16] core_region_i/core_master_r_data[17] core_region_i/core_master_r_data[18]
+ core_region_i/core_master_r_data[19] core_region_i/core_master_r_data[1] core_region_i/core_master_r_data[20]
+ core_region_i/core_master_r_data[21] core_region_i/core_master_r_data[22] core_region_i/core_master_r_data[23]
+ core_region_i/core_master_r_data[24] core_region_i/core_master_r_data[25] core_region_i/core_master_r_data[26]
+ core_region_i/core_master_r_data[27] core_region_i/core_master_r_data[28] core_region_i/core_master_r_data[29]
+ core_region_i/core_master_r_data[2] core_region_i/core_master_r_data[30] core_region_i/core_master_r_data[31]
+ core_region_i/core_master_r_data[32] core_region_i/core_master_r_data[33] core_region_i/core_master_r_data[34]
+ core_region_i/core_master_r_data[35] core_region_i/core_master_r_data[36] core_region_i/core_master_r_data[37]
+ core_region_i/core_master_r_data[38] core_region_i/core_master_r_data[39] core_region_i/core_master_r_data[3]
+ core_region_i/core_master_r_data[40] core_region_i/core_master_r_data[41] core_region_i/core_master_r_data[42]
+ core_region_i/core_master_r_data[43] core_region_i/core_master_r_data[44] core_region_i/core_master_r_data[45]
+ core_region_i/core_master_r_data[46] core_region_i/core_master_r_data[47] core_region_i/core_master_r_data[48]
+ core_region_i/core_master_r_data[49] core_region_i/core_master_r_data[4] core_region_i/core_master_r_data[50]
+ core_region_i/core_master_r_data[51] core_region_i/core_master_r_data[52] core_region_i/core_master_r_data[53]
+ core_region_i/core_master_r_data[54] core_region_i/core_master_r_data[55] core_region_i/core_master_r_data[56]
+ core_region_i/core_master_r_data[57] core_region_i/core_master_r_data[58] core_region_i/core_master_r_data[59]
+ core_region_i/core_master_r_data[5] core_region_i/core_master_r_data[60] core_region_i/core_master_r_data[61]
+ core_region_i/core_master_r_data[62] core_region_i/core_master_r_data[63] core_region_i/core_master_r_data[6]
+ core_region_i/core_master_r_data[7] core_region_i/core_master_r_data[8] core_region_i/core_master_r_data[9]
+ core_region_i/core_master_r_id[0] core_region_i/core_master_r_id[1] core_region_i/core_master_r_id[2]
+ core_region_i/core_master_r_id[3] core_region_i/core_master_r_id[4] core_region_i/core_master_r_id[5]
+ core_region_i/core_master_r_id[6] core_region_i/core_master_r_id[7] core_region_i/core_master_r_id[8]
+ core_region_i/core_master_r_id[9] axi_interconnect_i/s00_r_last axi_interconnect_i/s00_r_ready
+ axi_interconnect_i/s00_r_resp[0] axi_interconnect_i/s00_r_resp[1] core_region_i/core_master_r_user[-1]
+ core_region_i/core_master_r_user[0] axi_interconnect_i/s00_r_valid core_region_i/core_master_w_data[0]
+ core_region_i/core_master_w_data[10] core_region_i/core_master_w_data[11] core_region_i/core_master_w_data[12]
+ core_region_i/core_master_w_data[13] core_region_i/core_master_w_data[14] core_region_i/core_master_w_data[15]
+ core_region_i/core_master_w_data[16] core_region_i/core_master_w_data[17] core_region_i/core_master_w_data[18]
+ core_region_i/core_master_w_data[19] core_region_i/core_master_w_data[1] core_region_i/core_master_w_data[20]
+ core_region_i/core_master_w_data[21] core_region_i/core_master_w_data[22] core_region_i/core_master_w_data[23]
+ core_region_i/core_master_w_data[24] core_region_i/core_master_w_data[25] core_region_i/core_master_w_data[26]
+ core_region_i/core_master_w_data[27] core_region_i/core_master_w_data[28] core_region_i/core_master_w_data[29]
+ core_region_i/core_master_w_data[2] core_region_i/core_master_w_data[30] core_region_i/core_master_w_data[31]
+ core_region_i/core_master_w_data[32] core_region_i/core_master_w_data[33] core_region_i/core_master_w_data[34]
+ core_region_i/core_master_w_data[35] core_region_i/core_master_w_data[36] core_region_i/core_master_w_data[37]
+ core_region_i/core_master_w_data[38] core_region_i/core_master_w_data[39] core_region_i/core_master_w_data[3]
+ core_region_i/core_master_w_data[40] core_region_i/core_master_w_data[41] core_region_i/core_master_w_data[42]
+ core_region_i/core_master_w_data[43] core_region_i/core_master_w_data[44] core_region_i/core_master_w_data[45]
+ core_region_i/core_master_w_data[46] core_region_i/core_master_w_data[47] core_region_i/core_master_w_data[48]
+ core_region_i/core_master_w_data[49] core_region_i/core_master_w_data[4] core_region_i/core_master_w_data[50]
+ core_region_i/core_master_w_data[51] core_region_i/core_master_w_data[52] core_region_i/core_master_w_data[53]
+ core_region_i/core_master_w_data[54] core_region_i/core_master_w_data[55] core_region_i/core_master_w_data[56]
+ core_region_i/core_master_w_data[57] core_region_i/core_master_w_data[58] core_region_i/core_master_w_data[59]
+ core_region_i/core_master_w_data[5] core_region_i/core_master_w_data[60] core_region_i/core_master_w_data[61]
+ core_region_i/core_master_w_data[62] core_region_i/core_master_w_data[63] core_region_i/core_master_w_data[6]
+ core_region_i/core_master_w_data[7] core_region_i/core_master_w_data[8] core_region_i/core_master_w_data[9]
+ axi_interconnect_i/s00_w_last axi_interconnect_i/s00_w_ready core_region_i/core_master_w_strb[0]
+ core_region_i/core_master_w_strb[1] core_region_i/core_master_w_strb[2] core_region_i/core_master_w_strb[3]
+ core_region_i/core_master_w_strb[4] core_region_i/core_master_w_strb[5] core_region_i/core_master_w_strb[6]
+ core_region_i/core_master_w_strb[7] core_region_i/core_master_w_user[-1] core_region_i/core_master_w_user[0]
+ axi_interconnect_i/s00_w_valid axi_interconnect_i/m01_ar_addr[0] axi_interconnect_i/m01_ar_addr[10]
+ axi_interconnect_i/m01_ar_addr[11] axi_interconnect_i/m01_ar_addr[12] axi_interconnect_i/m01_ar_addr[13]
+ axi_interconnect_i/m01_ar_addr[14] axi_interconnect_i/m01_ar_addr[15] axi_interconnect_i/m01_ar_addr[16]
+ axi_interconnect_i/m01_ar_addr[17] axi_interconnect_i/m01_ar_addr[18] axi_interconnect_i/m01_ar_addr[19]
+ axi_interconnect_i/m01_ar_addr[1] axi_interconnect_i/m01_ar_addr[20] axi_interconnect_i/m01_ar_addr[21]
+ axi_interconnect_i/m01_ar_addr[22] axi_interconnect_i/m01_ar_addr[23] axi_interconnect_i/m01_ar_addr[24]
+ axi_interconnect_i/m01_ar_addr[25] axi_interconnect_i/m01_ar_addr[26] axi_interconnect_i/m01_ar_addr[27]
+ axi_interconnect_i/m01_ar_addr[28] axi_interconnect_i/m01_ar_addr[29] axi_interconnect_i/m01_ar_addr[2]
+ axi_interconnect_i/m01_ar_addr[30] axi_interconnect_i/m01_ar_addr[31] axi_interconnect_i/m01_ar_addr[3]
+ axi_interconnect_i/m01_ar_addr[4] axi_interconnect_i/m01_ar_addr[5] axi_interconnect_i/m01_ar_addr[6]
+ axi_interconnect_i/m01_ar_addr[7] axi_interconnect_i/m01_ar_addr[8] axi_interconnect_i/m01_ar_addr[9]
+ axi_interconnect_i/m01_ar_burst[0] axi_interconnect_i/m01_ar_burst[1] axi_interconnect_i/m01_ar_cache[0]
+ axi_interconnect_i/m01_ar_cache[1] axi_interconnect_i/m01_ar_cache[2] axi_interconnect_i/m01_ar_cache[3]
+ core_region_i/data_slave_ar_id[0] core_region_i/data_slave_ar_id[1] core_region_i/data_slave_ar_id[2]
+ core_region_i/data_slave_ar_id[3] core_region_i/data_slave_ar_id[4] core_region_i/data_slave_ar_id[5]
+ core_region_i/data_slave_ar_id[6] core_region_i/data_slave_ar_id[7] core_region_i/data_slave_ar_id[8]
+ core_region_i/data_slave_ar_id[9] axi_interconnect_i/m01_ar_len[0] axi_interconnect_i/m01_ar_len[1]
+ axi_interconnect_i/m01_ar_len[2] axi_interconnect_i/m01_ar_len[3] axi_interconnect_i/m01_ar_len[4]
+ axi_interconnect_i/m01_ar_len[5] axi_interconnect_i/m01_ar_len[6] axi_interconnect_i/m01_ar_len[7]
+ axi_interconnect_i/m01_ar_lock axi_interconnect_i/m01_ar_prot[0] axi_interconnect_i/m01_ar_prot[1]
+ axi_interconnect_i/m01_ar_prot[2] axi_interconnect_i/m01_ar_qos[0] axi_interconnect_i/m01_ar_qos[1]
+ axi_interconnect_i/m01_ar_qos[2] axi_interconnect_i/m01_ar_qos[3] axi_interconnect_i/m01_ar_ready
+ axi_interconnect_i/m01_ar_region[0] axi_interconnect_i/m01_ar_region[1] axi_interconnect_i/m01_ar_region[2]
+ axi_interconnect_i/m01_ar_region[3] axi_interconnect_i/m01_ar_size[0] axi_interconnect_i/m01_ar_size[1]
+ axi_interconnect_i/m01_ar_size[2] core_region_i/data_slave_ar_user[-1] core_region_i/data_slave_ar_user[0]
+ axi_interconnect_i/m01_ar_valid axi_interconnect_i/m01_aw_addr[0] axi_interconnect_i/m01_aw_addr[10]
+ axi_interconnect_i/m01_aw_addr[11] axi_interconnect_i/m01_aw_addr[12] axi_interconnect_i/m01_aw_addr[13]
+ axi_interconnect_i/m01_aw_addr[14] axi_interconnect_i/m01_aw_addr[15] axi_interconnect_i/m01_aw_addr[16]
+ axi_interconnect_i/m01_aw_addr[17] axi_interconnect_i/m01_aw_addr[18] axi_interconnect_i/m01_aw_addr[19]
+ axi_interconnect_i/m01_aw_addr[1] axi_interconnect_i/m01_aw_addr[20] axi_interconnect_i/m01_aw_addr[21]
+ axi_interconnect_i/m01_aw_addr[22] axi_interconnect_i/m01_aw_addr[23] axi_interconnect_i/m01_aw_addr[24]
+ axi_interconnect_i/m01_aw_addr[25] axi_interconnect_i/m01_aw_addr[26] axi_interconnect_i/m01_aw_addr[27]
+ axi_interconnect_i/m01_aw_addr[28] axi_interconnect_i/m01_aw_addr[29] axi_interconnect_i/m01_aw_addr[2]
+ axi_interconnect_i/m01_aw_addr[30] axi_interconnect_i/m01_aw_addr[31] axi_interconnect_i/m01_aw_addr[3]
+ axi_interconnect_i/m01_aw_addr[4] axi_interconnect_i/m01_aw_addr[5] axi_interconnect_i/m01_aw_addr[6]
+ axi_interconnect_i/m01_aw_addr[7] axi_interconnect_i/m01_aw_addr[8] axi_interconnect_i/m01_aw_addr[9]
+ axi_interconnect_i/m01_aw_burst[0] axi_interconnect_i/m01_aw_burst[1] axi_interconnect_i/m01_aw_cache[0]
+ axi_interconnect_i/m01_aw_cache[1] axi_interconnect_i/m01_aw_cache[2] axi_interconnect_i/m01_aw_cache[3]
+ core_region_i/data_slave_aw_id[0] core_region_i/data_slave_aw_id[1] core_region_i/data_slave_aw_id[2]
+ core_region_i/data_slave_aw_id[3] core_region_i/data_slave_aw_id[4] core_region_i/data_slave_aw_id[5]
+ core_region_i/data_slave_aw_id[6] core_region_i/data_slave_aw_id[7] core_region_i/data_slave_aw_id[8]
+ core_region_i/data_slave_aw_id[9] axi_interconnect_i/m01_aw_len[0] axi_interconnect_i/m01_aw_len[1]
+ axi_interconnect_i/m01_aw_len[2] axi_interconnect_i/m01_aw_len[3] axi_interconnect_i/m01_aw_len[4]
+ axi_interconnect_i/m01_aw_len[5] axi_interconnect_i/m01_aw_len[6] axi_interconnect_i/m01_aw_len[7]
+ axi_interconnect_i/m01_aw_lock axi_interconnect_i/m01_aw_prot[0] axi_interconnect_i/m01_aw_prot[1]
+ axi_interconnect_i/m01_aw_prot[2] axi_interconnect_i/m01_aw_qos[0] axi_interconnect_i/m01_aw_qos[1]
+ axi_interconnect_i/m01_aw_qos[2] axi_interconnect_i/m01_aw_qos[3] axi_interconnect_i/m01_aw_ready
+ axi_interconnect_i/m01_aw_region[0] axi_interconnect_i/m01_aw_region[1] axi_interconnect_i/m01_aw_region[2]
+ axi_interconnect_i/m01_aw_region[3] axi_interconnect_i/m01_aw_size[0] axi_interconnect_i/m01_aw_size[1]
+ axi_interconnect_i/m01_aw_size[2] core_region_i/data_slave_aw_user[-1] core_region_i/data_slave_aw_user[0]
+ axi_interconnect_i/m01_aw_valid core_region_i/data_slave_b_id[0] core_region_i/data_slave_b_id[1]
+ core_region_i/data_slave_b_id[2] core_region_i/data_slave_b_id[3] core_region_i/data_slave_b_id[4]
+ core_region_i/data_slave_b_id[5] core_region_i/data_slave_b_id[6] core_region_i/data_slave_b_id[7]
+ core_region_i/data_slave_b_id[8] core_region_i/data_slave_b_id[9] axi_interconnect_i/m01_b_ready
+ axi_interconnect_i/m01_b_resp[0] axi_interconnect_i/m01_b_resp[1] core_region_i/data_slave_b_user[-1]
+ core_region_i/data_slave_b_user[0] axi_interconnect_i/m01_b_valid core_region_i/data_slave_r_data[0]
+ core_region_i/data_slave_r_data[10] core_region_i/data_slave_r_data[11] core_region_i/data_slave_r_data[12]
+ core_region_i/data_slave_r_data[13] core_region_i/data_slave_r_data[14] core_region_i/data_slave_r_data[15]
+ core_region_i/data_slave_r_data[16] core_region_i/data_slave_r_data[17] core_region_i/data_slave_r_data[18]
+ core_region_i/data_slave_r_data[19] core_region_i/data_slave_r_data[1] core_region_i/data_slave_r_data[20]
+ core_region_i/data_slave_r_data[21] core_region_i/data_slave_r_data[22] core_region_i/data_slave_r_data[23]
+ core_region_i/data_slave_r_data[24] core_region_i/data_slave_r_data[25] core_region_i/data_slave_r_data[26]
+ core_region_i/data_slave_r_data[27] core_region_i/data_slave_r_data[28] core_region_i/data_slave_r_data[29]
+ core_region_i/data_slave_r_data[2] core_region_i/data_slave_r_data[30] core_region_i/data_slave_r_data[31]
+ core_region_i/data_slave_r_data[32] core_region_i/data_slave_r_data[33] core_region_i/data_slave_r_data[34]
+ core_region_i/data_slave_r_data[35] core_region_i/data_slave_r_data[36] core_region_i/data_slave_r_data[37]
+ core_region_i/data_slave_r_data[38] core_region_i/data_slave_r_data[39] core_region_i/data_slave_r_data[3]
+ core_region_i/data_slave_r_data[40] core_region_i/data_slave_r_data[41] core_region_i/data_slave_r_data[42]
+ core_region_i/data_slave_r_data[43] core_region_i/data_slave_r_data[44] core_region_i/data_slave_r_data[45]
+ core_region_i/data_slave_r_data[46] core_region_i/data_slave_r_data[47] core_region_i/data_slave_r_data[48]
+ core_region_i/data_slave_r_data[49] core_region_i/data_slave_r_data[4] core_region_i/data_slave_r_data[50]
+ core_region_i/data_slave_r_data[51] core_region_i/data_slave_r_data[52] core_region_i/data_slave_r_data[53]
+ core_region_i/data_slave_r_data[54] core_region_i/data_slave_r_data[55] core_region_i/data_slave_r_data[56]
+ core_region_i/data_slave_r_data[57] core_region_i/data_slave_r_data[58] core_region_i/data_slave_r_data[59]
+ core_region_i/data_slave_r_data[5] core_region_i/data_slave_r_data[60] core_region_i/data_slave_r_data[61]
+ core_region_i/data_slave_r_data[62] core_region_i/data_slave_r_data[63] core_region_i/data_slave_r_data[6]
+ core_region_i/data_slave_r_data[7] core_region_i/data_slave_r_data[8] core_region_i/data_slave_r_data[9]
+ core_region_i/data_slave_r_id[0] core_region_i/data_slave_r_id[1] core_region_i/data_slave_r_id[2]
+ core_region_i/data_slave_r_id[3] core_region_i/data_slave_r_id[4] core_region_i/data_slave_r_id[5]
+ core_region_i/data_slave_r_id[6] core_region_i/data_slave_r_id[7] core_region_i/data_slave_r_id[8]
+ core_region_i/data_slave_r_id[9] axi_interconnect_i/m01_r_last axi_interconnect_i/m01_r_ready
+ axi_interconnect_i/m01_r_resp[0] axi_interconnect_i/m01_r_resp[1] core_region_i/data_slave_r_user[-1]
+ core_region_i/data_slave_r_user[0] axi_interconnect_i/m01_r_valid core_region_i/data_slave_w_data[0]
+ core_region_i/data_slave_w_data[10] core_region_i/data_slave_w_data[11] core_region_i/data_slave_w_data[12]
+ core_region_i/data_slave_w_data[13] core_region_i/data_slave_w_data[14] core_region_i/data_slave_w_data[15]
+ core_region_i/data_slave_w_data[16] core_region_i/data_slave_w_data[17] core_region_i/data_slave_w_data[18]
+ core_region_i/data_slave_w_data[19] core_region_i/data_slave_w_data[1] core_region_i/data_slave_w_data[20]
+ core_region_i/data_slave_w_data[21] core_region_i/data_slave_w_data[22] core_region_i/data_slave_w_data[23]
+ core_region_i/data_slave_w_data[24] core_region_i/data_slave_w_data[25] core_region_i/data_slave_w_data[26]
+ core_region_i/data_slave_w_data[27] core_region_i/data_slave_w_data[28] core_region_i/data_slave_w_data[29]
+ core_region_i/data_slave_w_data[2] core_region_i/data_slave_w_data[30] core_region_i/data_slave_w_data[31]
+ core_region_i/data_slave_w_data[32] core_region_i/data_slave_w_data[33] core_region_i/data_slave_w_data[34]
+ core_region_i/data_slave_w_data[35] core_region_i/data_slave_w_data[36] core_region_i/data_slave_w_data[37]
+ core_region_i/data_slave_w_data[38] core_region_i/data_slave_w_data[39] core_region_i/data_slave_w_data[3]
+ core_region_i/data_slave_w_data[40] core_region_i/data_slave_w_data[41] core_region_i/data_slave_w_data[42]
+ core_region_i/data_slave_w_data[43] core_region_i/data_slave_w_data[44] core_region_i/data_slave_w_data[45]
+ core_region_i/data_slave_w_data[46] core_region_i/data_slave_w_data[47] core_region_i/data_slave_w_data[48]
+ core_region_i/data_slave_w_data[49] core_region_i/data_slave_w_data[4] core_region_i/data_slave_w_data[50]
+ core_region_i/data_slave_w_data[51] core_region_i/data_slave_w_data[52] core_region_i/data_slave_w_data[53]
+ core_region_i/data_slave_w_data[54] core_region_i/data_slave_w_data[55] core_region_i/data_slave_w_data[56]
+ core_region_i/data_slave_w_data[57] core_region_i/data_slave_w_data[58] core_region_i/data_slave_w_data[59]
+ core_region_i/data_slave_w_data[5] core_region_i/data_slave_w_data[60] core_region_i/data_slave_w_data[61]
+ core_region_i/data_slave_w_data[62] core_region_i/data_slave_w_data[63] core_region_i/data_slave_w_data[6]
+ core_region_i/data_slave_w_data[7] core_region_i/data_slave_w_data[8] core_region_i/data_slave_w_data[9]
+ axi_interconnect_i/m01_w_last axi_interconnect_i/m01_w_ready core_region_i/data_slave_w_strb[0]
+ core_region_i/data_slave_w_strb[1] core_region_i/data_slave_w_strb[2] core_region_i/data_slave_w_strb[3]
+ core_region_i/data_slave_w_strb[4] core_region_i/data_slave_w_strb[5] core_region_i/data_slave_w_strb[6]
+ core_region_i/data_slave_w_strb[7] core_region_i/data_slave_w_user[-1] core_region_i/data_slave_w_user[0]
+ axi_interconnect_i/m01_w_valid axi_interconnect_i/s01_ar_addr[0] axi_interconnect_i/s01_ar_addr[10]
+ axi_interconnect_i/s01_ar_addr[11] axi_interconnect_i/s01_ar_addr[12] axi_interconnect_i/s01_ar_addr[13]
+ axi_interconnect_i/s01_ar_addr[14] axi_interconnect_i/s01_ar_addr[15] axi_interconnect_i/s01_ar_addr[16]
+ axi_interconnect_i/s01_ar_addr[17] axi_interconnect_i/s01_ar_addr[18] axi_interconnect_i/s01_ar_addr[19]
+ axi_interconnect_i/s01_ar_addr[1] axi_interconnect_i/s01_ar_addr[20] axi_interconnect_i/s01_ar_addr[21]
+ axi_interconnect_i/s01_ar_addr[22] axi_interconnect_i/s01_ar_addr[23] axi_interconnect_i/s01_ar_addr[24]
+ axi_interconnect_i/s01_ar_addr[25] axi_interconnect_i/s01_ar_addr[26] axi_interconnect_i/s01_ar_addr[27]
+ axi_interconnect_i/s01_ar_addr[28] axi_interconnect_i/s01_ar_addr[29] axi_interconnect_i/s01_ar_addr[2]
+ axi_interconnect_i/s01_ar_addr[30] axi_interconnect_i/s01_ar_addr[31] axi_interconnect_i/s01_ar_addr[3]
+ axi_interconnect_i/s01_ar_addr[4] axi_interconnect_i/s01_ar_addr[5] axi_interconnect_i/s01_ar_addr[6]
+ axi_interconnect_i/s01_ar_addr[7] axi_interconnect_i/s01_ar_addr[8] axi_interconnect_i/s01_ar_addr[9]
+ axi_interconnect_i/s01_ar_burst[0] axi_interconnect_i/s01_ar_burst[1] axi_interconnect_i/s01_ar_cache[0]
+ axi_interconnect_i/s01_ar_cache[1] axi_interconnect_i/s01_ar_cache[2] axi_interconnect_i/s01_ar_cache[3]
+ core_region_i/dbg_master_ar_id[0] core_region_i/dbg_master_ar_id[1] core_region_i/dbg_master_ar_id[2]
+ core_region_i/dbg_master_ar_id[3] core_region_i/dbg_master_ar_id[4] core_region_i/dbg_master_ar_id[5]
+ core_region_i/dbg_master_ar_id[6] core_region_i/dbg_master_ar_id[7] core_region_i/dbg_master_ar_id[8]
+ core_region_i/dbg_master_ar_id[9] axi_interconnect_i/s01_ar_len[0] axi_interconnect_i/s01_ar_len[1]
+ axi_interconnect_i/s01_ar_len[2] axi_interconnect_i/s01_ar_len[3] axi_interconnect_i/s01_ar_len[4]
+ axi_interconnect_i/s01_ar_len[5] axi_interconnect_i/s01_ar_len[6] axi_interconnect_i/s01_ar_len[7]
+ axi_interconnect_i/s01_ar_lock axi_interconnect_i/s01_ar_prot[0] axi_interconnect_i/s01_ar_prot[1]
+ axi_interconnect_i/s01_ar_prot[2] axi_interconnect_i/s01_ar_qos[0] axi_interconnect_i/s01_ar_qos[1]
+ axi_interconnect_i/s01_ar_qos[2] axi_interconnect_i/s01_ar_qos[3] axi_interconnect_i/s01_ar_ready
+ axi_interconnect_i/s01_ar_region[0] axi_interconnect_i/s01_ar_region[1] axi_interconnect_i/s01_ar_region[2]
+ axi_interconnect_i/s01_ar_region[3] axi_interconnect_i/s01_ar_size[0] axi_interconnect_i/s01_ar_size[1]
+ axi_interconnect_i/s01_ar_size[2] core_region_i/dbg_master_ar_user[-1] core_region_i/dbg_master_ar_user[0]
+ axi_interconnect_i/s01_ar_valid axi_interconnect_i/s01_aw_addr[0] axi_interconnect_i/s01_aw_addr[10]
+ axi_interconnect_i/s01_aw_addr[11] axi_interconnect_i/s01_aw_addr[12] axi_interconnect_i/s01_aw_addr[13]
+ axi_interconnect_i/s01_aw_addr[14] axi_interconnect_i/s01_aw_addr[15] axi_interconnect_i/s01_aw_addr[16]
+ axi_interconnect_i/s01_aw_addr[17] axi_interconnect_i/s01_aw_addr[18] axi_interconnect_i/s01_aw_addr[19]
+ axi_interconnect_i/s01_aw_addr[1] axi_interconnect_i/s01_aw_addr[20] axi_interconnect_i/s01_aw_addr[21]
+ axi_interconnect_i/s01_aw_addr[22] axi_interconnect_i/s01_aw_addr[23] axi_interconnect_i/s01_aw_addr[24]
+ axi_interconnect_i/s01_aw_addr[25] axi_interconnect_i/s01_aw_addr[26] axi_interconnect_i/s01_aw_addr[27]
+ axi_interconnect_i/s01_aw_addr[28] axi_interconnect_i/s01_aw_addr[29] axi_interconnect_i/s01_aw_addr[2]
+ axi_interconnect_i/s01_aw_addr[30] axi_interconnect_i/s01_aw_addr[31] axi_interconnect_i/s01_aw_addr[3]
+ axi_interconnect_i/s01_aw_addr[4] axi_interconnect_i/s01_aw_addr[5] axi_interconnect_i/s01_aw_addr[6]
+ axi_interconnect_i/s01_aw_addr[7] axi_interconnect_i/s01_aw_addr[8] axi_interconnect_i/s01_aw_addr[9]
+ axi_interconnect_i/s01_aw_burst[0] axi_interconnect_i/s01_aw_burst[1] axi_interconnect_i/s01_aw_cache[0]
+ axi_interconnect_i/s01_aw_cache[1] axi_interconnect_i/s01_aw_cache[2] axi_interconnect_i/s01_aw_cache[3]
+ core_region_i/dbg_master_aw_id[0] core_region_i/dbg_master_aw_id[1] core_region_i/dbg_master_aw_id[2]
+ core_region_i/dbg_master_aw_id[3] core_region_i/dbg_master_aw_id[4] core_region_i/dbg_master_aw_id[5]
+ core_region_i/dbg_master_aw_id[6] core_region_i/dbg_master_aw_id[7] core_region_i/dbg_master_aw_id[8]
+ core_region_i/dbg_master_aw_id[9] axi_interconnect_i/s01_aw_len[0] axi_interconnect_i/s01_aw_len[1]
+ axi_interconnect_i/s01_aw_len[2] axi_interconnect_i/s01_aw_len[3] axi_interconnect_i/s01_aw_len[4]
+ axi_interconnect_i/s01_aw_len[5] axi_interconnect_i/s01_aw_len[6] axi_interconnect_i/s01_aw_len[7]
+ axi_interconnect_i/s01_aw_lock axi_interconnect_i/s01_aw_prot[0] axi_interconnect_i/s01_aw_prot[1]
+ axi_interconnect_i/s01_aw_prot[2] axi_interconnect_i/s01_aw_qos[0] axi_interconnect_i/s01_aw_qos[1]
+ axi_interconnect_i/s01_aw_qos[2] axi_interconnect_i/s01_aw_qos[3] axi_interconnect_i/s01_aw_ready
+ axi_interconnect_i/s01_aw_region[0] axi_interconnect_i/s01_aw_region[1] axi_interconnect_i/s01_aw_region[2]
+ axi_interconnect_i/s01_aw_region[3] axi_interconnect_i/s01_aw_size[0] axi_interconnect_i/s01_aw_size[1]
+ axi_interconnect_i/s01_aw_size[2] core_region_i/dbg_master_aw_user[-1] core_region_i/dbg_master_aw_user[0]
+ axi_interconnect_i/s01_aw_valid core_region_i/dbg_master_b_id[0] core_region_i/dbg_master_b_id[1]
+ core_region_i/dbg_master_b_id[2] core_region_i/dbg_master_b_id[3] core_region_i/dbg_master_b_id[4]
+ core_region_i/dbg_master_b_id[5] core_region_i/dbg_master_b_id[6] core_region_i/dbg_master_b_id[7]
+ core_region_i/dbg_master_b_id[8] core_region_i/dbg_master_b_id[9] axi_interconnect_i/s01_b_ready
+ axi_interconnect_i/s01_b_resp[0] axi_interconnect_i/s01_b_resp[1] core_region_i/dbg_master_b_user[-1]
+ core_region_i/dbg_master_b_user[0] axi_interconnect_i/s01_b_valid core_region_i/dbg_master_r_data[0]
+ core_region_i/dbg_master_r_data[10] core_region_i/dbg_master_r_data[11] core_region_i/dbg_master_r_data[12]
+ core_region_i/dbg_master_r_data[13] core_region_i/dbg_master_r_data[14] core_region_i/dbg_master_r_data[15]
+ core_region_i/dbg_master_r_data[16] core_region_i/dbg_master_r_data[17] core_region_i/dbg_master_r_data[18]
+ core_region_i/dbg_master_r_data[19] core_region_i/dbg_master_r_data[1] core_region_i/dbg_master_r_data[20]
+ core_region_i/dbg_master_r_data[21] core_region_i/dbg_master_r_data[22] core_region_i/dbg_master_r_data[23]
+ core_region_i/dbg_master_r_data[24] core_region_i/dbg_master_r_data[25] core_region_i/dbg_master_r_data[26]
+ core_region_i/dbg_master_r_data[27] core_region_i/dbg_master_r_data[28] core_region_i/dbg_master_r_data[29]
+ core_region_i/dbg_master_r_data[2] core_region_i/dbg_master_r_data[30] core_region_i/dbg_master_r_data[31]
+ core_region_i/dbg_master_r_data[32] core_region_i/dbg_master_r_data[33] core_region_i/dbg_master_r_data[34]
+ core_region_i/dbg_master_r_data[35] core_region_i/dbg_master_r_data[36] core_region_i/dbg_master_r_data[37]
+ core_region_i/dbg_master_r_data[38] core_region_i/dbg_master_r_data[39] core_region_i/dbg_master_r_data[3]
+ core_region_i/dbg_master_r_data[40] core_region_i/dbg_master_r_data[41] core_region_i/dbg_master_r_data[42]
+ core_region_i/dbg_master_r_data[43] core_region_i/dbg_master_r_data[44] core_region_i/dbg_master_r_data[45]
+ core_region_i/dbg_master_r_data[46] core_region_i/dbg_master_r_data[47] core_region_i/dbg_master_r_data[48]
+ core_region_i/dbg_master_r_data[49] core_region_i/dbg_master_r_data[4] core_region_i/dbg_master_r_data[50]
+ core_region_i/dbg_master_r_data[51] core_region_i/dbg_master_r_data[52] core_region_i/dbg_master_r_data[53]
+ core_region_i/dbg_master_r_data[54] core_region_i/dbg_master_r_data[55] core_region_i/dbg_master_r_data[56]
+ core_region_i/dbg_master_r_data[57] core_region_i/dbg_master_r_data[58] core_region_i/dbg_master_r_data[59]
+ core_region_i/dbg_master_r_data[5] core_region_i/dbg_master_r_data[60] core_region_i/dbg_master_r_data[61]
+ core_region_i/dbg_master_r_data[62] core_region_i/dbg_master_r_data[63] core_region_i/dbg_master_r_data[6]
+ core_region_i/dbg_master_r_data[7] core_region_i/dbg_master_r_data[8] core_region_i/dbg_master_r_data[9]
+ core_region_i/dbg_master_r_id[0] core_region_i/dbg_master_r_id[1] core_region_i/dbg_master_r_id[2]
+ core_region_i/dbg_master_r_id[3] core_region_i/dbg_master_r_id[4] core_region_i/dbg_master_r_id[5]
+ core_region_i/dbg_master_r_id[6] core_region_i/dbg_master_r_id[7] core_region_i/dbg_master_r_id[8]
+ core_region_i/dbg_master_r_id[9] axi_interconnect_i/s01_r_last axi_interconnect_i/s01_r_ready
+ axi_interconnect_i/s01_r_resp[0] axi_interconnect_i/s01_r_resp[1] core_region_i/dbg_master_r_user[-1]
+ core_region_i/dbg_master_r_user[0] axi_interconnect_i/s01_r_valid core_region_i/dbg_master_w_data[0]
+ core_region_i/dbg_master_w_data[10] core_region_i/dbg_master_w_data[11] core_region_i/dbg_master_w_data[12]
+ core_region_i/dbg_master_w_data[13] core_region_i/dbg_master_w_data[14] core_region_i/dbg_master_w_data[15]
+ core_region_i/dbg_master_w_data[16] core_region_i/dbg_master_w_data[17] core_region_i/dbg_master_w_data[18]
+ core_region_i/dbg_master_w_data[19] core_region_i/dbg_master_w_data[1] core_region_i/dbg_master_w_data[20]
+ core_region_i/dbg_master_w_data[21] core_region_i/dbg_master_w_data[22] core_region_i/dbg_master_w_data[23]
+ core_region_i/dbg_master_w_data[24] core_region_i/dbg_master_w_data[25] core_region_i/dbg_master_w_data[26]
+ core_region_i/dbg_master_w_data[27] core_region_i/dbg_master_w_data[28] core_region_i/dbg_master_w_data[29]
+ core_region_i/dbg_master_w_data[2] core_region_i/dbg_master_w_data[30] core_region_i/dbg_master_w_data[31]
+ core_region_i/dbg_master_w_data[32] core_region_i/dbg_master_w_data[33] core_region_i/dbg_master_w_data[34]
+ core_region_i/dbg_master_w_data[35] core_region_i/dbg_master_w_data[36] core_region_i/dbg_master_w_data[37]
+ core_region_i/dbg_master_w_data[38] core_region_i/dbg_master_w_data[39] core_region_i/dbg_master_w_data[3]
+ core_region_i/dbg_master_w_data[40] core_region_i/dbg_master_w_data[41] core_region_i/dbg_master_w_data[42]
+ core_region_i/dbg_master_w_data[43] core_region_i/dbg_master_w_data[44] core_region_i/dbg_master_w_data[45]
+ core_region_i/dbg_master_w_data[46] core_region_i/dbg_master_w_data[47] core_region_i/dbg_master_w_data[48]
+ core_region_i/dbg_master_w_data[49] core_region_i/dbg_master_w_data[4] core_region_i/dbg_master_w_data[50]
+ core_region_i/dbg_master_w_data[51] core_region_i/dbg_master_w_data[52] core_region_i/dbg_master_w_data[53]
+ core_region_i/dbg_master_w_data[54] core_region_i/dbg_master_w_data[55] core_region_i/dbg_master_w_data[56]
+ core_region_i/dbg_master_w_data[57] core_region_i/dbg_master_w_data[58] core_region_i/dbg_master_w_data[59]
+ core_region_i/dbg_master_w_data[5] core_region_i/dbg_master_w_data[60] core_region_i/dbg_master_w_data[61]
+ core_region_i/dbg_master_w_data[62] core_region_i/dbg_master_w_data[63] core_region_i/dbg_master_w_data[6]
+ core_region_i/dbg_master_w_data[7] core_region_i/dbg_master_w_data[8] core_region_i/dbg_master_w_data[9]
+ axi_interconnect_i/s01_w_last axi_interconnect_i/s01_w_ready core_region_i/dbg_master_w_strb[0]
+ core_region_i/dbg_master_w_strb[1] core_region_i/dbg_master_w_strb[2] core_region_i/dbg_master_w_strb[3]
+ core_region_i/dbg_master_w_strb[4] core_region_i/dbg_master_w_strb[5] core_region_i/dbg_master_w_strb[6]
+ core_region_i/dbg_master_w_strb[7] core_region_i/dbg_master_w_user[-1] core_region_i/dbg_master_w_user[0]
+ axi_interconnect_i/s01_w_valid peripherals_i/debug_addr[0] peripherals_i/debug_addr[10]
+ peripherals_i/debug_addr[11] peripherals_i/debug_addr[12] peripherals_i/debug_addr[13]
+ peripherals_i/debug_addr[14] peripherals_i/debug_addr[1] peripherals_i/debug_addr[2]
+ peripherals_i/debug_addr[3] peripherals_i/debug_addr[4] peripherals_i/debug_addr[5]
+ peripherals_i/debug_addr[6] peripherals_i/debug_addr[7] peripherals_i/debug_addr[8]
+ peripherals_i/debug_addr[9] peripherals_i/debug_gnt peripherals_i/debug_rdata[0]
+ peripherals_i/debug_rdata[10] peripherals_i/debug_rdata[11] peripherals_i/debug_rdata[12]
+ peripherals_i/debug_rdata[13] peripherals_i/debug_rdata[14] peripherals_i/debug_rdata[15]
+ peripherals_i/debug_rdata[16] peripherals_i/debug_rdata[17] peripherals_i/debug_rdata[18]
+ peripherals_i/debug_rdata[19] peripherals_i/debug_rdata[1] peripherals_i/debug_rdata[20]
+ peripherals_i/debug_rdata[21] peripherals_i/debug_rdata[22] peripherals_i/debug_rdata[23]
+ peripherals_i/debug_rdata[24] peripherals_i/debug_rdata[25] peripherals_i/debug_rdata[26]
+ peripherals_i/debug_rdata[27] peripherals_i/debug_rdata[28] peripherals_i/debug_rdata[29]
+ peripherals_i/debug_rdata[2] peripherals_i/debug_rdata[30] peripherals_i/debug_rdata[31]
+ peripherals_i/debug_rdata[3] peripherals_i/debug_rdata[4] peripherals_i/debug_rdata[5]
+ peripherals_i/debug_rdata[6] peripherals_i/debug_rdata[7] peripherals_i/debug_rdata[8]
+ peripherals_i/debug_rdata[9] peripherals_i/debug_req peripherals_i/debug_rvalid
+ peripherals_i/debug_wdata[0] peripherals_i/debug_wdata[10] peripherals_i/debug_wdata[11]
+ peripherals_i/debug_wdata[12] peripherals_i/debug_wdata[13] peripherals_i/debug_wdata[14]
+ peripherals_i/debug_wdata[15] peripherals_i/debug_wdata[16] peripherals_i/debug_wdata[17]
+ peripherals_i/debug_wdata[18] peripherals_i/debug_wdata[19] peripherals_i/debug_wdata[1]
+ peripherals_i/debug_wdata[20] peripherals_i/debug_wdata[21] peripherals_i/debug_wdata[22]
+ peripherals_i/debug_wdata[23] peripherals_i/debug_wdata[24] peripherals_i/debug_wdata[25]
+ peripherals_i/debug_wdata[26] peripherals_i/debug_wdata[27] peripherals_i/debug_wdata[28]
+ peripherals_i/debug_wdata[29] peripherals_i/debug_wdata[2] peripherals_i/debug_wdata[30]
+ peripherals_i/debug_wdata[31] peripherals_i/debug_wdata[3] peripherals_i/debug_wdata[4]
+ peripherals_i/debug_wdata[5] peripherals_i/debug_wdata[6] peripherals_i/debug_wdata[7]
+ peripherals_i/debug_wdata[8] peripherals_i/debug_wdata[9] peripherals_i/debug_we
+ peripherals_i/fetch_enable_o axi_interconnect_i/m00_ar_addr[0] axi_interconnect_i/m00_ar_addr[10]
+ axi_interconnect_i/m00_ar_addr[11] axi_interconnect_i/m00_ar_addr[12] axi_interconnect_i/m00_ar_addr[13]
+ axi_interconnect_i/m00_ar_addr[14] axi_interconnect_i/m00_ar_addr[15] axi_interconnect_i/m00_ar_addr[16]
+ axi_interconnect_i/m00_ar_addr[17] axi_interconnect_i/m00_ar_addr[18] axi_interconnect_i/m00_ar_addr[19]
+ axi_interconnect_i/m00_ar_addr[1] axi_interconnect_i/m00_ar_addr[20] axi_interconnect_i/m00_ar_addr[21]
+ axi_interconnect_i/m00_ar_addr[22] axi_interconnect_i/m00_ar_addr[23] axi_interconnect_i/m00_ar_addr[24]
+ axi_interconnect_i/m00_ar_addr[25] axi_interconnect_i/m00_ar_addr[26] axi_interconnect_i/m00_ar_addr[27]
+ axi_interconnect_i/m00_ar_addr[28] axi_interconnect_i/m00_ar_addr[29] axi_interconnect_i/m00_ar_addr[2]
+ axi_interconnect_i/m00_ar_addr[30] axi_interconnect_i/m00_ar_addr[31] axi_interconnect_i/m00_ar_addr[3]
+ axi_interconnect_i/m00_ar_addr[4] axi_interconnect_i/m00_ar_addr[5] axi_interconnect_i/m00_ar_addr[6]
+ axi_interconnect_i/m00_ar_addr[7] axi_interconnect_i/m00_ar_addr[8] axi_interconnect_i/m00_ar_addr[9]
+ axi_interconnect_i/m00_ar_burst[0] axi_interconnect_i/m00_ar_burst[1] axi_interconnect_i/m00_ar_cache[0]
+ axi_interconnect_i/m00_ar_cache[1] axi_interconnect_i/m00_ar_cache[2] axi_interconnect_i/m00_ar_cache[3]
+ core_region_i/instr_slave_ar_id[0] core_region_i/instr_slave_ar_id[1] core_region_i/instr_slave_ar_id[2]
+ core_region_i/instr_slave_ar_id[3] core_region_i/instr_slave_ar_id[4] core_region_i/instr_slave_ar_id[5]
+ core_region_i/instr_slave_ar_id[6] core_region_i/instr_slave_ar_id[7] core_region_i/instr_slave_ar_id[8]
+ core_region_i/instr_slave_ar_id[9] axi_interconnect_i/m00_ar_len[0] axi_interconnect_i/m00_ar_len[1]
+ axi_interconnect_i/m00_ar_len[2] axi_interconnect_i/m00_ar_len[3] axi_interconnect_i/m00_ar_len[4]
+ axi_interconnect_i/m00_ar_len[5] axi_interconnect_i/m00_ar_len[6] axi_interconnect_i/m00_ar_len[7]
+ axi_interconnect_i/m00_ar_lock axi_interconnect_i/m00_ar_prot[0] axi_interconnect_i/m00_ar_prot[1]
+ axi_interconnect_i/m00_ar_prot[2] axi_interconnect_i/m00_ar_qos[0] axi_interconnect_i/m00_ar_qos[1]
+ axi_interconnect_i/m00_ar_qos[2] axi_interconnect_i/m00_ar_qos[3] axi_interconnect_i/m00_ar_ready
+ axi_interconnect_i/m00_ar_region[0] axi_interconnect_i/m00_ar_region[1] axi_interconnect_i/m00_ar_region[2]
+ axi_interconnect_i/m00_ar_region[3] axi_interconnect_i/m00_ar_size[0] axi_interconnect_i/m00_ar_size[1]
+ axi_interconnect_i/m00_ar_size[2] core_region_i/instr_slave_ar_user[-1] core_region_i/instr_slave_ar_user[0]
+ axi_interconnect_i/m00_ar_valid axi_interconnect_i/m00_aw_addr[0] axi_interconnect_i/m00_aw_addr[10]
+ axi_interconnect_i/m00_aw_addr[11] axi_interconnect_i/m00_aw_addr[12] axi_interconnect_i/m00_aw_addr[13]
+ axi_interconnect_i/m00_aw_addr[14] axi_interconnect_i/m00_aw_addr[15] axi_interconnect_i/m00_aw_addr[16]
+ axi_interconnect_i/m00_aw_addr[17] axi_interconnect_i/m00_aw_addr[18] axi_interconnect_i/m00_aw_addr[19]
+ axi_interconnect_i/m00_aw_addr[1] axi_interconnect_i/m00_aw_addr[20] axi_interconnect_i/m00_aw_addr[21]
+ axi_interconnect_i/m00_aw_addr[22] axi_interconnect_i/m00_aw_addr[23] axi_interconnect_i/m00_aw_addr[24]
+ axi_interconnect_i/m00_aw_addr[25] axi_interconnect_i/m00_aw_addr[26] axi_interconnect_i/m00_aw_addr[27]
+ axi_interconnect_i/m00_aw_addr[28] axi_interconnect_i/m00_aw_addr[29] axi_interconnect_i/m00_aw_addr[2]
+ axi_interconnect_i/m00_aw_addr[30] axi_interconnect_i/m00_aw_addr[31] axi_interconnect_i/m00_aw_addr[3]
+ axi_interconnect_i/m00_aw_addr[4] axi_interconnect_i/m00_aw_addr[5] axi_interconnect_i/m00_aw_addr[6]
+ axi_interconnect_i/m00_aw_addr[7] axi_interconnect_i/m00_aw_addr[8] axi_interconnect_i/m00_aw_addr[9]
+ axi_interconnect_i/m00_aw_burst[0] axi_interconnect_i/m00_aw_burst[1] axi_interconnect_i/m00_aw_cache[0]
+ axi_interconnect_i/m00_aw_cache[1] axi_interconnect_i/m00_aw_cache[2] axi_interconnect_i/m00_aw_cache[3]
+ core_region_i/instr_slave_aw_id[0] core_region_i/instr_slave_aw_id[1] core_region_i/instr_slave_aw_id[2]
+ core_region_i/instr_slave_aw_id[3] core_region_i/instr_slave_aw_id[4] core_region_i/instr_slave_aw_id[5]
+ core_region_i/instr_slave_aw_id[6] core_region_i/instr_slave_aw_id[7] core_region_i/instr_slave_aw_id[8]
+ core_region_i/instr_slave_aw_id[9] axi_interconnect_i/m00_aw_len[0] axi_interconnect_i/m00_aw_len[1]
+ axi_interconnect_i/m00_aw_len[2] axi_interconnect_i/m00_aw_len[3] axi_interconnect_i/m00_aw_len[4]
+ axi_interconnect_i/m00_aw_len[5] axi_interconnect_i/m00_aw_len[6] axi_interconnect_i/m00_aw_len[7]
+ axi_interconnect_i/m00_aw_lock axi_interconnect_i/m00_aw_prot[0] axi_interconnect_i/m00_aw_prot[1]
+ axi_interconnect_i/m00_aw_prot[2] axi_interconnect_i/m00_aw_qos[0] axi_interconnect_i/m00_aw_qos[1]
+ axi_interconnect_i/m00_aw_qos[2] axi_interconnect_i/m00_aw_qos[3] axi_interconnect_i/m00_aw_ready
+ axi_interconnect_i/m00_aw_region[0] axi_interconnect_i/m00_aw_region[1] axi_interconnect_i/m00_aw_region[2]
+ axi_interconnect_i/m00_aw_region[3] axi_interconnect_i/m00_aw_size[0] axi_interconnect_i/m00_aw_size[1]
+ axi_interconnect_i/m00_aw_size[2] core_region_i/instr_slave_aw_user[-1] core_region_i/instr_slave_aw_user[0]
+ axi_interconnect_i/m00_aw_valid core_region_i/instr_slave_b_id[0] core_region_i/instr_slave_b_id[1]
+ core_region_i/instr_slave_b_id[2] core_region_i/instr_slave_b_id[3] core_region_i/instr_slave_b_id[4]
+ core_region_i/instr_slave_b_id[5] core_region_i/instr_slave_b_id[6] core_region_i/instr_slave_b_id[7]
+ core_region_i/instr_slave_b_id[8] core_region_i/instr_slave_b_id[9] axi_interconnect_i/m00_b_ready
+ axi_interconnect_i/m00_b_resp[0] axi_interconnect_i/m00_b_resp[1] core_region_i/instr_slave_b_user[-1]
+ core_region_i/instr_slave_b_user[0] axi_interconnect_i/m00_b_valid core_region_i/instr_slave_r_data[0]
+ core_region_i/instr_slave_r_data[10] core_region_i/instr_slave_r_data[11] core_region_i/instr_slave_r_data[12]
+ core_region_i/instr_slave_r_data[13] core_region_i/instr_slave_r_data[14] core_region_i/instr_slave_r_data[15]
+ core_region_i/instr_slave_r_data[16] core_region_i/instr_slave_r_data[17] core_region_i/instr_slave_r_data[18]
+ core_region_i/instr_slave_r_data[19] core_region_i/instr_slave_r_data[1] core_region_i/instr_slave_r_data[20]
+ core_region_i/instr_slave_r_data[21] core_region_i/instr_slave_r_data[22] core_region_i/instr_slave_r_data[23]
+ core_region_i/instr_slave_r_data[24] core_region_i/instr_slave_r_data[25] core_region_i/instr_slave_r_data[26]
+ core_region_i/instr_slave_r_data[27] core_region_i/instr_slave_r_data[28] core_region_i/instr_slave_r_data[29]
+ core_region_i/instr_slave_r_data[2] core_region_i/instr_slave_r_data[30] core_region_i/instr_slave_r_data[31]
+ core_region_i/instr_slave_r_data[32] core_region_i/instr_slave_r_data[33] core_region_i/instr_slave_r_data[34]
+ core_region_i/instr_slave_r_data[35] core_region_i/instr_slave_r_data[36] core_region_i/instr_slave_r_data[37]
+ core_region_i/instr_slave_r_data[38] core_region_i/instr_slave_r_data[39] core_region_i/instr_slave_r_data[3]
+ core_region_i/instr_slave_r_data[40] core_region_i/instr_slave_r_data[41] core_region_i/instr_slave_r_data[42]
+ core_region_i/instr_slave_r_data[43] core_region_i/instr_slave_r_data[44] core_region_i/instr_slave_r_data[45]
+ core_region_i/instr_slave_r_data[46] core_region_i/instr_slave_r_data[47] core_region_i/instr_slave_r_data[48]
+ core_region_i/instr_slave_r_data[49] core_region_i/instr_slave_r_data[4] core_region_i/instr_slave_r_data[50]
+ core_region_i/instr_slave_r_data[51] core_region_i/instr_slave_r_data[52] core_region_i/instr_slave_r_data[53]
+ core_region_i/instr_slave_r_data[54] core_region_i/instr_slave_r_data[55] core_region_i/instr_slave_r_data[56]
+ core_region_i/instr_slave_r_data[57] core_region_i/instr_slave_r_data[58] core_region_i/instr_slave_r_data[59]
+ core_region_i/instr_slave_r_data[5] core_region_i/instr_slave_r_data[60] core_region_i/instr_slave_r_data[61]
+ core_region_i/instr_slave_r_data[62] core_region_i/instr_slave_r_data[63] core_region_i/instr_slave_r_data[6]
+ core_region_i/instr_slave_r_data[7] core_region_i/instr_slave_r_data[8] core_region_i/instr_slave_r_data[9]
+ core_region_i/instr_slave_r_id[0] core_region_i/instr_slave_r_id[1] core_region_i/instr_slave_r_id[2]
+ core_region_i/instr_slave_r_id[3] core_region_i/instr_slave_r_id[4] core_region_i/instr_slave_r_id[5]
+ core_region_i/instr_slave_r_id[6] core_region_i/instr_slave_r_id[7] core_region_i/instr_slave_r_id[8]
+ core_region_i/instr_slave_r_id[9] axi_interconnect_i/m00_r_last axi_interconnect_i/m00_r_ready
+ axi_interconnect_i/m00_r_resp[0] axi_interconnect_i/m00_r_resp[1] core_region_i/instr_slave_r_user[-1]
+ core_region_i/instr_slave_r_user[0] axi_interconnect_i/m00_r_valid core_region_i/instr_slave_w_data[0]
+ core_region_i/instr_slave_w_data[10] core_region_i/instr_slave_w_data[11] core_region_i/instr_slave_w_data[12]
+ core_region_i/instr_slave_w_data[13] core_region_i/instr_slave_w_data[14] core_region_i/instr_slave_w_data[15]
+ core_region_i/instr_slave_w_data[16] core_region_i/instr_slave_w_data[17] core_region_i/instr_slave_w_data[18]
+ core_region_i/instr_slave_w_data[19] core_region_i/instr_slave_w_data[1] core_region_i/instr_slave_w_data[20]
+ core_region_i/instr_slave_w_data[21] core_region_i/instr_slave_w_data[22] core_region_i/instr_slave_w_data[23]
+ core_region_i/instr_slave_w_data[24] core_region_i/instr_slave_w_data[25] core_region_i/instr_slave_w_data[26]
+ core_region_i/instr_slave_w_data[27] core_region_i/instr_slave_w_data[28] core_region_i/instr_slave_w_data[29]
+ core_region_i/instr_slave_w_data[2] core_region_i/instr_slave_w_data[30] core_region_i/instr_slave_w_data[31]
+ core_region_i/instr_slave_w_data[32] core_region_i/instr_slave_w_data[33] core_region_i/instr_slave_w_data[34]
+ core_region_i/instr_slave_w_data[35] core_region_i/instr_slave_w_data[36] core_region_i/instr_slave_w_data[37]
+ core_region_i/instr_slave_w_data[38] core_region_i/instr_slave_w_data[39] core_region_i/instr_slave_w_data[3]
+ core_region_i/instr_slave_w_data[40] core_region_i/instr_slave_w_data[41] core_region_i/instr_slave_w_data[42]
+ core_region_i/instr_slave_w_data[43] core_region_i/instr_slave_w_data[44] core_region_i/instr_slave_w_data[45]
+ core_region_i/instr_slave_w_data[46] core_region_i/instr_slave_w_data[47] core_region_i/instr_slave_w_data[48]
+ core_region_i/instr_slave_w_data[49] core_region_i/instr_slave_w_data[4] core_region_i/instr_slave_w_data[50]
+ core_region_i/instr_slave_w_data[51] core_region_i/instr_slave_w_data[52] core_region_i/instr_slave_w_data[53]
+ core_region_i/instr_slave_w_data[54] core_region_i/instr_slave_w_data[55] core_region_i/instr_slave_w_data[56]
+ core_region_i/instr_slave_w_data[57] core_region_i/instr_slave_w_data[58] core_region_i/instr_slave_w_data[59]
+ core_region_i/instr_slave_w_data[5] core_region_i/instr_slave_w_data[60] core_region_i/instr_slave_w_data[61]
+ core_region_i/instr_slave_w_data[62] core_region_i/instr_slave_w_data[63] core_region_i/instr_slave_w_data[6]
+ core_region_i/instr_slave_w_data[7] core_region_i/instr_slave_w_data[8] core_region_i/instr_slave_w_data[9]
+ axi_interconnect_i/m00_w_last axi_interconnect_i/m00_w_ready core_region_i/instr_slave_w_strb[0]
+ core_region_i/instr_slave_w_strb[1] core_region_i/instr_slave_w_strb[2] core_region_i/instr_slave_w_strb[3]
+ core_region_i/instr_slave_w_strb[4] core_region_i/instr_slave_w_strb[5] core_region_i/instr_slave_w_strb[6]
+ core_region_i/instr_slave_w_strb[7] core_region_i/instr_slave_w_user[-1] core_region_i/instr_slave_w_user[0]
+ axi_interconnect_i/m00_w_valid peripherals_i/irq_o[0] peripherals_i/irq_o[10] peripherals_i/irq_o[11]
+ peripherals_i/irq_o[12] peripherals_i/irq_o[13] peripherals_i/irq_o[14] peripherals_i/irq_o[15]
+ peripherals_i/irq_o[16] peripherals_i/irq_o[17] peripherals_i/irq_o[18] peripherals_i/irq_o[19]
+ peripherals_i/irq_o[1] peripherals_i/irq_o[20] peripherals_i/irq_o[21] peripherals_i/irq_o[22]
+ peripherals_i/irq_o[23] peripherals_i/irq_o[24] peripherals_i/irq_o[25] peripherals_i/irq_o[26]
+ peripherals_i/irq_o[27] peripherals_i/irq_o[28] peripherals_i/irq_o[29] peripherals_i/irq_o[2]
+ peripherals_i/irq_o[30] peripherals_i/irq_o[31] peripherals_i/irq_o[3] peripherals_i/irq_o[4]
+ peripherals_i/irq_o[5] peripherals_i/irq_o[6] peripherals_i/irq_o[7] peripherals_i/irq_o[8]
+ peripherals_i/irq_o[9] core_region_i/mba_data_mem_addr0_o[0] data_ram/addr0[8] core_region_i/mba_data_mem_addr0_o[11]
+ core_region_i/mba_data_mem_addr0_o[12] core_region_i/mba_data_mem_addr0_o[13] core_region_i/mba_data_mem_addr0_o[14]
+ core_region_i/mba_data_mem_addr0_o[15] core_region_i/mba_data_mem_addr0_o[16] core_region_i/mba_data_mem_addr0_o[17]
+ core_region_i/mba_data_mem_addr0_o[18] core_region_i/mba_data_mem_addr0_o[19] core_region_i/mba_data_mem_addr0_o[1]
+ core_region_i/mba_data_mem_addr0_o[20] core_region_i/mba_data_mem_addr0_o[21] core_region_i/mba_data_mem_addr0_o[22]
+ core_region_i/mba_data_mem_addr0_o[23] core_region_i/mba_data_mem_addr0_o[24] core_region_i/mba_data_mem_addr0_o[25]
+ core_region_i/mba_data_mem_addr0_o[26] core_region_i/mba_data_mem_addr0_o[27] core_region_i/mba_data_mem_addr0_o[28]
+ core_region_i/mba_data_mem_addr0_o[29] data_ram/addr0[0] core_region_i/mba_data_mem_addr0_o[30]
+ core_region_i/mba_data_mem_addr0_o[31] data_ram/addr0[1] data_ram/addr0[2] data_ram/addr0[3]
+ data_ram/addr0[4] data_ram/addr0[5] data_ram/addr0[6] data_ram/addr0[7] core_region_i/mba_data_mem_addr1_o[0]
+ data_ram/addr1[8] core_region_i/mba_data_mem_addr1_o[11] core_region_i/mba_data_mem_addr1_o[12]
+ core_region_i/mba_data_mem_addr1_o[13] core_region_i/mba_data_mem_addr1_o[14] core_region_i/mba_data_mem_addr1_o[15]
+ core_region_i/mba_data_mem_addr1_o[16] core_region_i/mba_data_mem_addr1_o[17] core_region_i/mba_data_mem_addr1_o[18]
+ core_region_i/mba_data_mem_addr1_o[19] core_region_i/mba_data_mem_addr1_o[1] core_region_i/mba_data_mem_addr1_o[20]
+ core_region_i/mba_data_mem_addr1_o[21] core_region_i/mba_data_mem_addr1_o[22] core_region_i/mba_data_mem_addr1_o[23]
+ core_region_i/mba_data_mem_addr1_o[24] core_region_i/mba_data_mem_addr1_o[25] core_region_i/mba_data_mem_addr1_o[26]
+ core_region_i/mba_data_mem_addr1_o[27] core_region_i/mba_data_mem_addr1_o[28] core_region_i/mba_data_mem_addr1_o[29]
+ data_ram/addr1[0] core_region_i/mba_data_mem_addr1_o[30] core_region_i/mba_data_mem_addr1_o[31]
+ data_ram/addr1[1] data_ram/addr1[2] data_ram/addr1[3] data_ram/addr1[4] data_ram/addr1[5]
+ data_ram/addr1[6] data_ram/addr1[7] data_ram/csb0 data_ram/csb1 data_ram/din0[0]
+ data_ram/din0[10] data_ram/din0[11] data_ram/din0[12] data_ram/din0[13] data_ram/din0[14]
+ data_ram/din0[15] data_ram/din0[16] data_ram/din0[17] data_ram/din0[18] data_ram/din0[19]
+ data_ram/din0[1] data_ram/din0[20] data_ram/din0[21] data_ram/din0[22] data_ram/din0[23]
+ data_ram/din0[24] data_ram/din0[25] data_ram/din0[26] data_ram/din0[27] data_ram/din0[28]
+ data_ram/din0[29] data_ram/din0[2] data_ram/din0[30] data_ram/din0[31] data_ram/din0[3]
+ data_ram/din0[4] data_ram/din0[5] data_ram/din0[6] data_ram/din0[7] data_ram/din0[8]
+ data_ram/din0[9] data_ram/dout0[0] data_ram/dout0[10] data_ram/dout0[11] data_ram/dout0[12]
+ data_ram/dout0[13] data_ram/dout0[14] data_ram/dout0[15] data_ram/dout0[16] data_ram/dout0[17]
+ data_ram/dout0[18] data_ram/dout0[19] data_ram/dout0[1] data_ram/dout0[20] data_ram/dout0[21]
+ data_ram/dout0[22] data_ram/dout0[23] data_ram/dout0[24] data_ram/dout0[25] data_ram/dout0[26]
+ data_ram/dout0[27] data_ram/dout0[28] data_ram/dout0[29] data_ram/dout0[2] data_ram/dout0[30]
+ data_ram/dout0[31] data_ram/dout0[3] data_ram/dout0[4] data_ram/dout0[5] data_ram/dout0[6]
+ data_ram/dout0[7] data_ram/dout0[8] data_ram/dout0[9] data_ram/web0 data_ram/wmask0[0]
+ data_ram/wmask0[1] data_ram/wmask0[2] data_ram/wmask0[3] core_region_i/mba_instr_mem_addr0_o[0]
+ instr_ram/addr0[8] core_region_i/mba_instr_mem_addr0_o[11] core_region_i/mba_instr_mem_addr0_o[12]
+ core_region_i/mba_instr_mem_addr0_o[13] core_region_i/mba_instr_mem_addr0_o[14]
+ core_region_i/mba_instr_mem_addr0_o[15] core_region_i/mba_instr_mem_addr0_o[16]
+ core_region_i/mba_instr_mem_addr0_o[17] core_region_i/mba_instr_mem_addr0_o[18]
+ core_region_i/mba_instr_mem_addr0_o[19] core_region_i/mba_instr_mem_addr0_o[1] core_region_i/mba_instr_mem_addr0_o[20]
+ core_region_i/mba_instr_mem_addr0_o[21] core_region_i/mba_instr_mem_addr0_o[22]
+ core_region_i/mba_instr_mem_addr0_o[23] core_region_i/mba_instr_mem_addr0_o[24]
+ core_region_i/mba_instr_mem_addr0_o[25] core_region_i/mba_instr_mem_addr0_o[26]
+ core_region_i/mba_instr_mem_addr0_o[27] core_region_i/mba_instr_mem_addr0_o[28]
+ core_region_i/mba_instr_mem_addr0_o[29] instr_ram/addr0[0] core_region_i/mba_instr_mem_addr0_o[30]
+ core_region_i/mba_instr_mem_addr0_o[31] instr_ram/addr0[1] instr_ram/addr0[2] instr_ram/addr0[3]
+ instr_ram/addr0[4] instr_ram/addr0[5] instr_ram/addr0[6] instr_ram/addr0[7] core_region_i/mba_instr_mem_addr1_o[0]
+ instr_ram/addr1[8] core_region_i/mba_instr_mem_addr1_o[11] core_region_i/mba_instr_mem_addr1_o[12]
+ core_region_i/mba_instr_mem_addr1_o[13] core_region_i/mba_instr_mem_addr1_o[14]
+ core_region_i/mba_instr_mem_addr1_o[15] core_region_i/mba_instr_mem_addr1_o[16]
+ core_region_i/mba_instr_mem_addr1_o[17] core_region_i/mba_instr_mem_addr1_o[18]
+ core_region_i/mba_instr_mem_addr1_o[19] core_region_i/mba_instr_mem_addr1_o[1] core_region_i/mba_instr_mem_addr1_o[20]
+ core_region_i/mba_instr_mem_addr1_o[21] core_region_i/mba_instr_mem_addr1_o[22]
+ core_region_i/mba_instr_mem_addr1_o[23] core_region_i/mba_instr_mem_addr1_o[24]
+ core_region_i/mba_instr_mem_addr1_o[25] core_region_i/mba_instr_mem_addr1_o[26]
+ core_region_i/mba_instr_mem_addr1_o[27] core_region_i/mba_instr_mem_addr1_o[28]
+ core_region_i/mba_instr_mem_addr1_o[29] instr_ram/addr1[0] core_region_i/mba_instr_mem_addr1_o[30]
+ core_region_i/mba_instr_mem_addr1_o[31] instr_ram/addr1[1] instr_ram/addr1[2] instr_ram/addr1[3]
+ instr_ram/addr1[4] instr_ram/addr1[5] instr_ram/addr1[6] instr_ram/addr1[7] instr_ram/csb0
+ instr_ram/csb1 instr_ram/din0[0] instr_ram/din0[10] instr_ram/din0[11] instr_ram/din0[12]
+ instr_ram/din0[13] instr_ram/din0[14] instr_ram/din0[15] instr_ram/din0[16] instr_ram/din0[17]
+ instr_ram/din0[18] instr_ram/din0[19] instr_ram/din0[1] instr_ram/din0[20] instr_ram/din0[21]
+ instr_ram/din0[22] instr_ram/din0[23] instr_ram/din0[24] instr_ram/din0[25] instr_ram/din0[26]
+ instr_ram/din0[27] instr_ram/din0[28] instr_ram/din0[29] instr_ram/din0[2] instr_ram/din0[30]
+ instr_ram/din0[31] instr_ram/din0[3] instr_ram/din0[4] instr_ram/din0[5] instr_ram/din0[6]
+ instr_ram/din0[7] instr_ram/din0[8] instr_ram/din0[9] instr_ram/dout0[0] instr_ram/dout0[10]
+ instr_ram/dout0[11] instr_ram/dout0[12] instr_ram/dout0[13] instr_ram/dout0[14]
+ instr_ram/dout0[15] instr_ram/dout0[16] instr_ram/dout0[17] instr_ram/dout0[18]
+ instr_ram/dout0[19] instr_ram/dout0[1] instr_ram/dout0[20] instr_ram/dout0[21] instr_ram/dout0[22]
+ instr_ram/dout0[23] instr_ram/dout0[24] instr_ram/dout0[25] instr_ram/dout0[26]
+ instr_ram/dout0[27] instr_ram/dout0[28] instr_ram/dout0[29] instr_ram/dout0[2] instr_ram/dout0[30]
+ instr_ram/dout0[31] instr_ram/dout0[3] instr_ram/dout0[4] instr_ram/dout0[5] instr_ram/dout0[6]
+ instr_ram/dout0[7] instr_ram/dout0[8] instr_ram/dout0[9] instr_ram/web0 instr_ram/wmask0[0]
+ instr_ram/wmask0[1] instr_ram/wmask0[2] instr_ram/wmask0[3] peripherals_i/rst_n
+ io_in[12] io_in[15] io_out[26] la_data_in[2] io_in[14] io_in[13] vccd1 vssd1 mba_core_region
Xdata_ram data_ram/din0[0] data_ram/din0[1] data_ram/din0[2] data_ram/din0[3] data_ram/din0[4]
+ data_ram/din0[5] data_ram/din0[6] data_ram/din0[7] data_ram/din0[8] data_ram/din0[9]
+ data_ram/din0[10] data_ram/din0[11] data_ram/din0[12] data_ram/din0[13] data_ram/din0[14]
+ data_ram/din0[15] data_ram/din0[16] data_ram/din0[17] data_ram/din0[18] data_ram/din0[19]
+ data_ram/din0[20] data_ram/din0[21] data_ram/din0[22] data_ram/din0[23] data_ram/din0[24]
+ data_ram/din0[25] data_ram/din0[26] data_ram/din0[27] data_ram/din0[28] data_ram/din0[29]
+ data_ram/din0[30] data_ram/din0[31] data_ram/addr0[0] data_ram/addr0[1] data_ram/addr0[2]
+ data_ram/addr0[3] data_ram/addr0[4] data_ram/addr0[5] data_ram/addr0[6] data_ram/addr0[7]
+ data_ram/addr0[8] data_ram/addr1[0] data_ram/addr1[1] data_ram/addr1[2] data_ram/addr1[3]
+ data_ram/addr1[4] data_ram/addr1[5] data_ram/addr1[6] data_ram/addr1[7] data_ram/addr1[8]
+ data_ram/csb0 data_ram/csb1 data_ram/web0 data_ram/clk0 io_in[21] data_ram/wmask0[0]
+ data_ram/wmask0[1] data_ram/wmask0[2] data_ram/wmask0[3] data_ram/dout0[0] data_ram/dout0[1]
+ data_ram/dout0[2] data_ram/dout0[3] data_ram/dout0[4] data_ram/dout0[5] data_ram/dout0[6]
+ data_ram/dout0[7] data_ram/dout0[8] data_ram/dout0[9] data_ram/dout0[10] data_ram/dout0[11]
+ data_ram/dout0[12] data_ram/dout0[13] data_ram/dout0[14] data_ram/dout0[15] data_ram/dout0[16]
+ data_ram/dout0[17] data_ram/dout0[18] data_ram/dout0[19] data_ram/dout0[20] data_ram/dout0[21]
+ data_ram/dout0[22] data_ram/dout0[23] data_ram/dout0[24] data_ram/dout0[25] data_ram/dout0[26]
+ data_ram/dout0[27] data_ram/dout0[28] data_ram/dout0[29] data_ram/dout0[30] data_ram/dout0[31]
+ data_ram/dout1[0] data_ram/dout1[1] data_ram/dout1[2] data_ram/dout1[3] data_ram/dout1[4]
+ data_ram/dout1[5] data_ram/dout1[6] data_ram/dout1[7] data_ram/dout1[8] data_ram/dout1[9]
+ data_ram/dout1[10] data_ram/dout1[11] data_ram/dout1[12] data_ram/dout1[13] data_ram/dout1[14]
+ data_ram/dout1[15] data_ram/dout1[16] data_ram/dout1[17] data_ram/dout1[18] data_ram/dout1[19]
+ data_ram/dout1[20] data_ram/dout1[21] data_ram/dout1[22] data_ram/dout1[23] data_ram/dout1[24]
+ data_ram/dout1[25] data_ram/dout1[26] data_ram/dout1[27] data_ram/dout1[28] data_ram/dout1[29]
+ data_ram/dout1[30] data_ram/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xinstr_ram instr_ram/din0[0] instr_ram/din0[1] instr_ram/din0[2] instr_ram/din0[3]
+ instr_ram/din0[4] instr_ram/din0[5] instr_ram/din0[6] instr_ram/din0[7] instr_ram/din0[8]
+ instr_ram/din0[9] instr_ram/din0[10] instr_ram/din0[11] instr_ram/din0[12] instr_ram/din0[13]
+ instr_ram/din0[14] instr_ram/din0[15] instr_ram/din0[16] instr_ram/din0[17] instr_ram/din0[18]
+ instr_ram/din0[19] instr_ram/din0[20] instr_ram/din0[21] instr_ram/din0[22] instr_ram/din0[23]
+ instr_ram/din0[24] instr_ram/din0[25] instr_ram/din0[26] instr_ram/din0[27] instr_ram/din0[28]
+ instr_ram/din0[29] instr_ram/din0[30] instr_ram/din0[31] instr_ram/addr0[0] instr_ram/addr0[1]
+ instr_ram/addr0[2] instr_ram/addr0[3] instr_ram/addr0[4] instr_ram/addr0[5] instr_ram/addr0[6]
+ instr_ram/addr0[7] instr_ram/addr0[8] instr_ram/addr1[0] instr_ram/addr1[1] instr_ram/addr1[2]
+ instr_ram/addr1[3] instr_ram/addr1[4] instr_ram/addr1[5] instr_ram/addr1[6] instr_ram/addr1[7]
+ instr_ram/addr1[8] instr_ram/csb0 instr_ram/csb1 instr_ram/web0 data_ram/clk0 io_in[21]
+ instr_ram/wmask0[0] instr_ram/wmask0[1] instr_ram/wmask0[2] instr_ram/wmask0[3]
+ instr_ram/dout0[0] instr_ram/dout0[1] instr_ram/dout0[2] instr_ram/dout0[3] instr_ram/dout0[4]
+ instr_ram/dout0[5] instr_ram/dout0[6] instr_ram/dout0[7] instr_ram/dout0[8] instr_ram/dout0[9]
+ instr_ram/dout0[10] instr_ram/dout0[11] instr_ram/dout0[12] instr_ram/dout0[13]
+ instr_ram/dout0[14] instr_ram/dout0[15] instr_ram/dout0[16] instr_ram/dout0[17]
+ instr_ram/dout0[18] instr_ram/dout0[19] instr_ram/dout0[20] instr_ram/dout0[21]
+ instr_ram/dout0[22] instr_ram/dout0[23] instr_ram/dout0[24] instr_ram/dout0[25]
+ instr_ram/dout0[26] instr_ram/dout0[27] instr_ram/dout0[28] instr_ram/dout0[29]
+ instr_ram/dout0[30] instr_ram/dout0[31] instr_ram/dout1[0] instr_ram/dout1[1] instr_ram/dout1[2]
+ instr_ram/dout1[3] instr_ram/dout1[4] instr_ram/dout1[5] instr_ram/dout1[6] instr_ram/dout1[7]
+ instr_ram/dout1[8] instr_ram/dout1[9] instr_ram/dout1[10] instr_ram/dout1[11] instr_ram/dout1[12]
+ instr_ram/dout1[13] instr_ram/dout1[14] instr_ram/dout1[15] instr_ram/dout1[16]
+ instr_ram/dout1[17] instr_ram/dout1[18] instr_ram/dout1[19] instr_ram/dout1[20]
+ instr_ram/dout1[21] instr_ram/dout1[22] instr_ram/dout1[23] instr_ram/dout1[24]
+ instr_ram/dout1[25] instr_ram/dout1[26] instr_ram/dout1[27] instr_ram/dout1[28]
+ instr_ram/dout1[29] instr_ram/dout1[30] instr_ram/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xperipherals_i axi_interconnect_i/s02_ar_addr[0] axi_interconnect_i/s02_ar_addr[10]
+ axi_interconnect_i/s02_ar_addr[11] axi_interconnect_i/s02_ar_addr[12] axi_interconnect_i/s02_ar_addr[13]
+ axi_interconnect_i/s02_ar_addr[14] axi_interconnect_i/s02_ar_addr[15] axi_interconnect_i/s02_ar_addr[16]
+ axi_interconnect_i/s02_ar_addr[17] axi_interconnect_i/s02_ar_addr[18] axi_interconnect_i/s02_ar_addr[19]
+ axi_interconnect_i/s02_ar_addr[1] axi_interconnect_i/s02_ar_addr[20] axi_interconnect_i/s02_ar_addr[21]
+ axi_interconnect_i/s02_ar_addr[22] axi_interconnect_i/s02_ar_addr[23] axi_interconnect_i/s02_ar_addr[24]
+ axi_interconnect_i/s02_ar_addr[25] axi_interconnect_i/s02_ar_addr[26] axi_interconnect_i/s02_ar_addr[27]
+ axi_interconnect_i/s02_ar_addr[28] axi_interconnect_i/s02_ar_addr[29] axi_interconnect_i/s02_ar_addr[2]
+ axi_interconnect_i/s02_ar_addr[30] axi_interconnect_i/s02_ar_addr[31] axi_interconnect_i/s02_ar_addr[3]
+ axi_interconnect_i/s02_ar_addr[4] axi_interconnect_i/s02_ar_addr[5] axi_interconnect_i/s02_ar_addr[6]
+ axi_interconnect_i/s02_ar_addr[7] axi_interconnect_i/s02_ar_addr[8] axi_interconnect_i/s02_ar_addr[9]
+ axi_interconnect_i/s02_ar_burst[0] axi_interconnect_i/s02_ar_burst[1] axi_interconnect_i/s02_ar_cache[0]
+ axi_interconnect_i/s02_ar_cache[1] axi_interconnect_i/s02_ar_cache[2] axi_interconnect_i/s02_ar_cache[3]
+ peripherals_i/axi_spi_master_ar_id[0] peripherals_i/axi_spi_master_ar_id[1] peripherals_i/axi_spi_master_ar_id[2]
+ peripherals_i/axi_spi_master_ar_id[3] peripherals_i/axi_spi_master_ar_id[4] peripherals_i/axi_spi_master_ar_id[5]
+ axi_interconnect_i/s02_ar_len[0] axi_interconnect_i/s02_ar_len[1] axi_interconnect_i/s02_ar_len[2]
+ axi_interconnect_i/s02_ar_len[3] axi_interconnect_i/s02_ar_len[4] axi_interconnect_i/s02_ar_len[5]
+ axi_interconnect_i/s02_ar_len[6] axi_interconnect_i/s02_ar_len[7] axi_interconnect_i/s02_ar_lock
+ axi_interconnect_i/s02_ar_prot[0] axi_interconnect_i/s02_ar_prot[1] axi_interconnect_i/s02_ar_prot[2]
+ axi_interconnect_i/s02_ar_qos[0] axi_interconnect_i/s02_ar_qos[1] axi_interconnect_i/s02_ar_qos[2]
+ axi_interconnect_i/s02_ar_qos[3] axi_interconnect_i/s02_ar_ready axi_interconnect_i/s02_ar_region[0]
+ axi_interconnect_i/s02_ar_region[1] axi_interconnect_i/s02_ar_region[2] axi_interconnect_i/s02_ar_region[3]
+ axi_interconnect_i/s02_ar_size[0] axi_interconnect_i/s02_ar_size[1] axi_interconnect_i/s02_ar_size[2]
+ peripherals_i/axi_spi_master_ar_user[0] peripherals_i/axi_spi_master_ar_user[1]
+ peripherals_i/axi_spi_master_ar_user[2] peripherals_i/axi_spi_master_ar_user[3]
+ peripherals_i/axi_spi_master_ar_user[4] peripherals_i/axi_spi_master_ar_user[5]
+ axi_interconnect_i/s02_ar_valid axi_interconnect_i/s02_aw_addr[0] axi_interconnect_i/s02_aw_addr[10]
+ axi_interconnect_i/s02_aw_addr[11] axi_interconnect_i/s02_aw_addr[12] axi_interconnect_i/s02_aw_addr[13]
+ axi_interconnect_i/s02_aw_addr[14] axi_interconnect_i/s02_aw_addr[15] axi_interconnect_i/s02_aw_addr[16]
+ axi_interconnect_i/s02_aw_addr[17] axi_interconnect_i/s02_aw_addr[18] axi_interconnect_i/s02_aw_addr[19]
+ axi_interconnect_i/s02_aw_addr[1] axi_interconnect_i/s02_aw_addr[20] axi_interconnect_i/s02_aw_addr[21]
+ axi_interconnect_i/s02_aw_addr[22] axi_interconnect_i/s02_aw_addr[23] axi_interconnect_i/s02_aw_addr[24]
+ axi_interconnect_i/s02_aw_addr[25] axi_interconnect_i/s02_aw_addr[26] axi_interconnect_i/s02_aw_addr[27]
+ axi_interconnect_i/s02_aw_addr[28] axi_interconnect_i/s02_aw_addr[29] axi_interconnect_i/s02_aw_addr[2]
+ axi_interconnect_i/s02_aw_addr[30] axi_interconnect_i/s02_aw_addr[31] axi_interconnect_i/s02_aw_addr[3]
+ axi_interconnect_i/s02_aw_addr[4] axi_interconnect_i/s02_aw_addr[5] axi_interconnect_i/s02_aw_addr[6]
+ axi_interconnect_i/s02_aw_addr[7] axi_interconnect_i/s02_aw_addr[8] axi_interconnect_i/s02_aw_addr[9]
+ axi_interconnect_i/s02_aw_burst[0] axi_interconnect_i/s02_aw_burst[1] axi_interconnect_i/s02_aw_cache[0]
+ axi_interconnect_i/s02_aw_cache[1] axi_interconnect_i/s02_aw_cache[2] axi_interconnect_i/s02_aw_cache[3]
+ peripherals_i/axi_spi_master_aw_id[0] peripherals_i/axi_spi_master_aw_id[1] peripherals_i/axi_spi_master_aw_id[2]
+ peripherals_i/axi_spi_master_aw_id[3] peripherals_i/axi_spi_master_aw_id[4] peripherals_i/axi_spi_master_aw_id[5]
+ axi_interconnect_i/s02_aw_len[0] axi_interconnect_i/s02_aw_len[1] axi_interconnect_i/s02_aw_len[2]
+ axi_interconnect_i/s02_aw_len[3] axi_interconnect_i/s02_aw_len[4] axi_interconnect_i/s02_aw_len[5]
+ axi_interconnect_i/s02_aw_len[6] axi_interconnect_i/s02_aw_len[7] axi_interconnect_i/s02_aw_lock
+ axi_interconnect_i/s02_aw_prot[0] axi_interconnect_i/s02_aw_prot[1] axi_interconnect_i/s02_aw_prot[2]
+ axi_interconnect_i/s02_aw_qos[0] axi_interconnect_i/s02_aw_qos[1] axi_interconnect_i/s02_aw_qos[2]
+ axi_interconnect_i/s02_aw_qos[3] axi_interconnect_i/s02_aw_ready axi_interconnect_i/s02_aw_region[0]
+ axi_interconnect_i/s02_aw_region[1] axi_interconnect_i/s02_aw_region[2] axi_interconnect_i/s02_aw_region[3]
+ axi_interconnect_i/s02_aw_size[0] axi_interconnect_i/s02_aw_size[1] axi_interconnect_i/s02_aw_size[2]
+ peripherals_i/axi_spi_master_aw_user[0] peripherals_i/axi_spi_master_aw_user[1]
+ peripherals_i/axi_spi_master_aw_user[2] peripherals_i/axi_spi_master_aw_user[3]
+ peripherals_i/axi_spi_master_aw_user[4] peripherals_i/axi_spi_master_aw_user[5]
+ axi_interconnect_i/s02_aw_valid peripherals_i/axi_spi_master_b_id[0] peripherals_i/axi_spi_master_b_id[1]
+ peripherals_i/axi_spi_master_b_id[2] peripherals_i/axi_spi_master_b_id[3] peripherals_i/axi_spi_master_b_id[4]
+ peripherals_i/axi_spi_master_b_id[5] axi_interconnect_i/s02_b_ready axi_interconnect_i/s02_b_resp[0]
+ axi_interconnect_i/s02_b_resp[1] peripherals_i/axi_spi_master_b_user[0] peripherals_i/axi_spi_master_b_user[1]
+ peripherals_i/axi_spi_master_b_user[2] peripherals_i/axi_spi_master_b_user[3] peripherals_i/axi_spi_master_b_user[4]
+ peripherals_i/axi_spi_master_b_user[5] axi_interconnect_i/s02_b_valid peripherals_i/axi_spi_master_r_data[0]
+ peripherals_i/axi_spi_master_r_data[10] peripherals_i/axi_spi_master_r_data[11]
+ peripherals_i/axi_spi_master_r_data[12] peripherals_i/axi_spi_master_r_data[13]
+ peripherals_i/axi_spi_master_r_data[14] peripherals_i/axi_spi_master_r_data[15]
+ peripherals_i/axi_spi_master_r_data[16] peripherals_i/axi_spi_master_r_data[17]
+ peripherals_i/axi_spi_master_r_data[18] peripherals_i/axi_spi_master_r_data[19]
+ peripherals_i/axi_spi_master_r_data[1] peripherals_i/axi_spi_master_r_data[20] peripherals_i/axi_spi_master_r_data[21]
+ peripherals_i/axi_spi_master_r_data[22] peripherals_i/axi_spi_master_r_data[23]
+ peripherals_i/axi_spi_master_r_data[24] peripherals_i/axi_spi_master_r_data[25]
+ peripherals_i/axi_spi_master_r_data[26] peripherals_i/axi_spi_master_r_data[27]
+ peripherals_i/axi_spi_master_r_data[28] peripherals_i/axi_spi_master_r_data[29]
+ peripherals_i/axi_spi_master_r_data[2] peripherals_i/axi_spi_master_r_data[30] peripherals_i/axi_spi_master_r_data[31]
+ peripherals_i/axi_spi_master_r_data[32] peripherals_i/axi_spi_master_r_data[33]
+ peripherals_i/axi_spi_master_r_data[34] peripherals_i/axi_spi_master_r_data[35]
+ peripherals_i/axi_spi_master_r_data[36] peripherals_i/axi_spi_master_r_data[37]
+ peripherals_i/axi_spi_master_r_data[38] peripherals_i/axi_spi_master_r_data[39]
+ peripherals_i/axi_spi_master_r_data[3] peripherals_i/axi_spi_master_r_data[40] peripherals_i/axi_spi_master_r_data[41]
+ peripherals_i/axi_spi_master_r_data[42] peripherals_i/axi_spi_master_r_data[43]
+ peripherals_i/axi_spi_master_r_data[44] peripherals_i/axi_spi_master_r_data[45]
+ peripherals_i/axi_spi_master_r_data[46] peripherals_i/axi_spi_master_r_data[47]
+ peripherals_i/axi_spi_master_r_data[48] peripherals_i/axi_spi_master_r_data[49]
+ peripherals_i/axi_spi_master_r_data[4] peripherals_i/axi_spi_master_r_data[50] peripherals_i/axi_spi_master_r_data[51]
+ peripherals_i/axi_spi_master_r_data[52] peripherals_i/axi_spi_master_r_data[53]
+ peripherals_i/axi_spi_master_r_data[54] peripherals_i/axi_spi_master_r_data[55]
+ peripherals_i/axi_spi_master_r_data[56] peripherals_i/axi_spi_master_r_data[57]
+ peripherals_i/axi_spi_master_r_data[58] peripherals_i/axi_spi_master_r_data[59]
+ peripherals_i/axi_spi_master_r_data[5] peripherals_i/axi_spi_master_r_data[60] peripherals_i/axi_spi_master_r_data[61]
+ peripherals_i/axi_spi_master_r_data[62] peripherals_i/axi_spi_master_r_data[63]
+ peripherals_i/axi_spi_master_r_data[6] peripherals_i/axi_spi_master_r_data[7] peripherals_i/axi_spi_master_r_data[8]
+ peripherals_i/axi_spi_master_r_data[9] peripherals_i/axi_spi_master_r_id[0] peripherals_i/axi_spi_master_r_id[1]
+ peripherals_i/axi_spi_master_r_id[2] peripherals_i/axi_spi_master_r_id[3] peripherals_i/axi_spi_master_r_id[4]
+ peripherals_i/axi_spi_master_r_id[5] axi_interconnect_i/s02_r_last axi_interconnect_i/s02_r_ready
+ axi_interconnect_i/s02_r_resp[0] axi_interconnect_i/s02_r_resp[1] peripherals_i/axi_spi_master_r_user[0]
+ peripherals_i/axi_spi_master_r_user[1] peripherals_i/axi_spi_master_r_user[2] peripherals_i/axi_spi_master_r_user[3]
+ peripherals_i/axi_spi_master_r_user[4] peripherals_i/axi_spi_master_r_user[5] axi_interconnect_i/s02_r_valid
+ peripherals_i/axi_spi_master_w_data[0] peripherals_i/axi_spi_master_w_data[10] peripherals_i/axi_spi_master_w_data[11]
+ peripherals_i/axi_spi_master_w_data[12] peripherals_i/axi_spi_master_w_data[13]
+ peripherals_i/axi_spi_master_w_data[14] peripherals_i/axi_spi_master_w_data[15]
+ peripherals_i/axi_spi_master_w_data[16] peripherals_i/axi_spi_master_w_data[17]
+ peripherals_i/axi_spi_master_w_data[18] peripherals_i/axi_spi_master_w_data[19]
+ peripherals_i/axi_spi_master_w_data[1] peripherals_i/axi_spi_master_w_data[20] peripherals_i/axi_spi_master_w_data[21]
+ peripherals_i/axi_spi_master_w_data[22] peripherals_i/axi_spi_master_w_data[23]
+ peripherals_i/axi_spi_master_w_data[24] peripherals_i/axi_spi_master_w_data[25]
+ peripherals_i/axi_spi_master_w_data[26] peripherals_i/axi_spi_master_w_data[27]
+ peripherals_i/axi_spi_master_w_data[28] peripherals_i/axi_spi_master_w_data[29]
+ peripherals_i/axi_spi_master_w_data[2] peripherals_i/axi_spi_master_w_data[30] peripherals_i/axi_spi_master_w_data[31]
+ peripherals_i/axi_spi_master_w_data[32] peripherals_i/axi_spi_master_w_data[33]
+ peripherals_i/axi_spi_master_w_data[34] peripherals_i/axi_spi_master_w_data[35]
+ peripherals_i/axi_spi_master_w_data[36] peripherals_i/axi_spi_master_w_data[37]
+ peripherals_i/axi_spi_master_w_data[38] peripherals_i/axi_spi_master_w_data[39]
+ peripherals_i/axi_spi_master_w_data[3] peripherals_i/axi_spi_master_w_data[40] peripherals_i/axi_spi_master_w_data[41]
+ peripherals_i/axi_spi_master_w_data[42] peripherals_i/axi_spi_master_w_data[43]
+ peripherals_i/axi_spi_master_w_data[44] peripherals_i/axi_spi_master_w_data[45]
+ peripherals_i/axi_spi_master_w_data[46] peripherals_i/axi_spi_master_w_data[47]
+ peripherals_i/axi_spi_master_w_data[48] peripherals_i/axi_spi_master_w_data[49]
+ peripherals_i/axi_spi_master_w_data[4] peripherals_i/axi_spi_master_w_data[50] peripherals_i/axi_spi_master_w_data[51]
+ peripherals_i/axi_spi_master_w_data[52] peripherals_i/axi_spi_master_w_data[53]
+ peripherals_i/axi_spi_master_w_data[54] peripherals_i/axi_spi_master_w_data[55]
+ peripherals_i/axi_spi_master_w_data[56] peripherals_i/axi_spi_master_w_data[57]
+ peripherals_i/axi_spi_master_w_data[58] peripherals_i/axi_spi_master_w_data[59]
+ peripherals_i/axi_spi_master_w_data[5] peripherals_i/axi_spi_master_w_data[60] peripherals_i/axi_spi_master_w_data[61]
+ peripherals_i/axi_spi_master_w_data[62] peripherals_i/axi_spi_master_w_data[63]
+ peripherals_i/axi_spi_master_w_data[6] peripherals_i/axi_spi_master_w_data[7] peripherals_i/axi_spi_master_w_data[8]
+ peripherals_i/axi_spi_master_w_data[9] axi_interconnect_i/s02_w_last axi_interconnect_i/s02_w_ready
+ peripherals_i/axi_spi_master_w_strb[0] peripherals_i/axi_spi_master_w_strb[1] peripherals_i/axi_spi_master_w_strb[2]
+ peripherals_i/axi_spi_master_w_strb[3] peripherals_i/axi_spi_master_w_strb[4] peripherals_i/axi_spi_master_w_strb[5]
+ peripherals_i/axi_spi_master_w_strb[6] peripherals_i/axi_spi_master_w_strb[7] peripherals_i/axi_spi_master_w_user[0]
+ peripherals_i/axi_spi_master_w_user[1] peripherals_i/axi_spi_master_w_user[2] peripherals_i/axi_spi_master_w_user[3]
+ peripherals_i/axi_spi_master_w_user[4] peripherals_i/axi_spi_master_w_user[5] axi_interconnect_i/s02_w_valid
+ peripherals_i/boot_addr_o[0] peripherals_i/boot_addr_o[10] peripherals_i/boot_addr_o[11]
+ peripherals_i/boot_addr_o[12] peripherals_i/boot_addr_o[13] peripherals_i/boot_addr_o[14]
+ peripherals_i/boot_addr_o[15] peripherals_i/boot_addr_o[16] peripherals_i/boot_addr_o[17]
+ peripherals_i/boot_addr_o[18] peripherals_i/boot_addr_o[19] peripherals_i/boot_addr_o[1]
+ peripherals_i/boot_addr_o[20] peripherals_i/boot_addr_o[21] peripherals_i/boot_addr_o[22]
+ peripherals_i/boot_addr_o[23] peripherals_i/boot_addr_o[24] peripherals_i/boot_addr_o[25]
+ peripherals_i/boot_addr_o[26] peripherals_i/boot_addr_o[27] peripherals_i/boot_addr_o[28]
+ peripherals_i/boot_addr_o[29] peripherals_i/boot_addr_o[2] peripherals_i/boot_addr_o[30]
+ peripherals_i/boot_addr_o[31] peripherals_i/boot_addr_o[3] peripherals_i/boot_addr_o[4]
+ peripherals_i/boot_addr_o[5] peripherals_i/boot_addr_o[6] peripherals_i/boot_addr_o[7]
+ peripherals_i/boot_addr_o[8] peripherals_i/boot_addr_o[9] core_region_i/clock_gating_i
+ data_ram/clk0 user_clock2 data_ram/clk0 la_data_in[0] la_data_in[1] peripherals_i/core_busy_i
+ peripherals_i/debug_addr[0] peripherals_i/debug_addr[10] peripherals_i/debug_addr[11]
+ peripherals_i/debug_addr[12] peripherals_i/debug_addr[13] peripherals_i/debug_addr[14]
+ peripherals_i/debug_addr[1] peripherals_i/debug_addr[2] peripherals_i/debug_addr[3]
+ peripherals_i/debug_addr[4] peripherals_i/debug_addr[5] peripherals_i/debug_addr[6]
+ peripherals_i/debug_addr[7] peripherals_i/debug_addr[8] peripherals_i/debug_addr[9]
+ peripherals_i/debug_gnt peripherals_i/debug_rdata[0] peripherals_i/debug_rdata[10]
+ peripherals_i/debug_rdata[11] peripherals_i/debug_rdata[12] peripherals_i/debug_rdata[13]
+ peripherals_i/debug_rdata[14] peripherals_i/debug_rdata[15] peripherals_i/debug_rdata[16]
+ peripherals_i/debug_rdata[17] peripherals_i/debug_rdata[18] peripherals_i/debug_rdata[19]
+ peripherals_i/debug_rdata[1] peripherals_i/debug_rdata[20] peripherals_i/debug_rdata[21]
+ peripherals_i/debug_rdata[22] peripherals_i/debug_rdata[23] peripherals_i/debug_rdata[24]
+ peripherals_i/debug_rdata[25] peripherals_i/debug_rdata[26] peripherals_i/debug_rdata[27]
+ peripherals_i/debug_rdata[28] peripherals_i/debug_rdata[29] peripherals_i/debug_rdata[2]
+ peripherals_i/debug_rdata[30] peripherals_i/debug_rdata[31] peripherals_i/debug_rdata[3]
+ peripherals_i/debug_rdata[4] peripherals_i/debug_rdata[5] peripherals_i/debug_rdata[6]
+ peripherals_i/debug_rdata[7] peripherals_i/debug_rdata[8] peripherals_i/debug_rdata[9]
+ peripherals_i/debug_req peripherals_i/debug_rvalid peripherals_i/debug_wdata[0]
+ peripherals_i/debug_wdata[10] peripherals_i/debug_wdata[11] peripherals_i/debug_wdata[12]
+ peripherals_i/debug_wdata[13] peripherals_i/debug_wdata[14] peripherals_i/debug_wdata[15]
+ peripherals_i/debug_wdata[16] peripherals_i/debug_wdata[17] peripherals_i/debug_wdata[18]
+ peripherals_i/debug_wdata[19] peripherals_i/debug_wdata[1] peripherals_i/debug_wdata[20]
+ peripherals_i/debug_wdata[21] peripherals_i/debug_wdata[22] peripherals_i/debug_wdata[23]
+ peripherals_i/debug_wdata[24] peripherals_i/debug_wdata[25] peripherals_i/debug_wdata[26]
+ peripherals_i/debug_wdata[27] peripherals_i/debug_wdata[28] peripherals_i/debug_wdata[29]
+ peripherals_i/debug_wdata[2] peripherals_i/debug_wdata[30] peripherals_i/debug_wdata[31]
+ peripherals_i/debug_wdata[3] peripherals_i/debug_wdata[4] peripherals_i/debug_wdata[5]
+ peripherals_i/debug_wdata[6] peripherals_i/debug_wdata[7] peripherals_i/debug_wdata[8]
+ peripherals_i/debug_wdata[9] peripherals_i/debug_we la_data_in[6] peripherals_i/fetch_enable_o
+ peripherals_i/fll1_ack_i peripherals_i/fll1_add_o[0] peripherals_i/fll1_add_o[1]
+ peripherals_i/fll1_lock_i peripherals_i/fll1_rdata_i[0] peripherals_i/fll1_rdata_i[10]
+ peripherals_i/fll1_rdata_i[11] peripherals_i/fll1_rdata_i[12] peripherals_i/fll1_rdata_i[13]
+ peripherals_i/fll1_rdata_i[14] peripherals_i/fll1_rdata_i[15] peripherals_i/fll1_rdata_i[16]
+ peripherals_i/fll1_rdata_i[17] peripherals_i/fll1_rdata_i[18] peripherals_i/fll1_rdata_i[19]
+ peripherals_i/fll1_rdata_i[1] peripherals_i/fll1_rdata_i[20] peripherals_i/fll1_rdata_i[21]
+ peripherals_i/fll1_rdata_i[22] peripherals_i/fll1_rdata_i[23] peripherals_i/fll1_rdata_i[24]
+ peripherals_i/fll1_rdata_i[25] peripherals_i/fll1_rdata_i[26] peripherals_i/fll1_rdata_i[27]
+ peripherals_i/fll1_rdata_i[28] peripherals_i/fll1_rdata_i[29] peripherals_i/fll1_rdata_i[2]
+ peripherals_i/fll1_rdata_i[30] peripherals_i/fll1_rdata_i[31] peripherals_i/fll1_rdata_i[3]
+ peripherals_i/fll1_rdata_i[4] peripherals_i/fll1_rdata_i[5] peripherals_i/fll1_rdata_i[6]
+ peripherals_i/fll1_rdata_i[7] peripherals_i/fll1_rdata_i[8] peripherals_i/fll1_rdata_i[9]
+ peripherals_i/fll1_req_o peripherals_i/fll1_wdata_o[0] peripherals_i/fll1_wdata_o[10]
+ peripherals_i/fll1_wdata_o[11] peripherals_i/fll1_wdata_o[12] peripherals_i/fll1_wdata_o[13]
+ peripherals_i/fll1_wdata_o[14] peripherals_i/fll1_wdata_o[15] peripherals_i/fll1_wdata_o[16]
+ peripherals_i/fll1_wdata_o[17] peripherals_i/fll1_wdata_o[18] peripherals_i/fll1_wdata_o[19]
+ peripherals_i/fll1_wdata_o[1] peripherals_i/fll1_wdata_o[20] peripherals_i/fll1_wdata_o[21]
+ peripherals_i/fll1_wdata_o[22] peripherals_i/fll1_wdata_o[23] peripherals_i/fll1_wdata_o[24]
+ peripherals_i/fll1_wdata_o[25] peripherals_i/fll1_wdata_o[26] peripherals_i/fll1_wdata_o[27]
+ peripherals_i/fll1_wdata_o[28] peripherals_i/fll1_wdata_o[29] peripherals_i/fll1_wdata_o[2]
+ peripherals_i/fll1_wdata_o[30] peripherals_i/fll1_wdata_o[31] peripherals_i/fll1_wdata_o[3]
+ peripherals_i/fll1_wdata_o[4] peripherals_i/fll1_wdata_o[5] peripherals_i/fll1_wdata_o[6]
+ peripherals_i/fll1_wdata_o[7] peripherals_i/fll1_wdata_o[8] peripherals_i/fll1_wdata_o[9]
+ peripherals_i/fll1_wrn_o peripherals_i/fll1_ack_i peripherals_i/fll1_add_o[0] peripherals_i/fll1_add_o[1]
+ peripherals_i/fll1_wdata_o[0] peripherals_i/fll1_wdata_o[10] peripherals_i/fll1_wdata_o[11]
+ peripherals_i/fll1_wdata_o[12] peripherals_i/fll1_wdata_o[13] peripherals_i/fll1_wdata_o[14]
+ peripherals_i/fll1_wdata_o[15] peripherals_i/fll1_wdata_o[16] peripherals_i/fll1_wdata_o[17]
+ peripherals_i/fll1_wdata_o[18] peripherals_i/fll1_wdata_o[19] peripherals_i/fll1_wdata_o[1]
+ peripherals_i/fll1_wdata_o[20] peripherals_i/fll1_wdata_o[21] peripherals_i/fll1_wdata_o[22]
+ peripherals_i/fll1_wdata_o[23] peripherals_i/fll1_wdata_o[24] peripherals_i/fll1_wdata_o[25]
+ peripherals_i/fll1_wdata_o[26] peripherals_i/fll1_wdata_o[27] peripherals_i/fll1_wdata_o[28]
+ peripherals_i/fll1_wdata_o[29] peripherals_i/fll1_wdata_o[2] peripherals_i/fll1_wdata_o[30]
+ peripherals_i/fll1_wdata_o[31] peripherals_i/fll1_wdata_o[3] peripherals_i/fll1_wdata_o[4]
+ peripherals_i/fll1_wdata_o[5] peripherals_i/fll1_wdata_o[6] peripherals_i/fll1_wdata_o[7]
+ peripherals_i/fll1_wdata_o[8] peripherals_i/fll1_wdata_o[9] peripherals_i/fll1_lock_i
+ peripherals_i/fll1_rdata_i[0] peripherals_i/fll1_rdata_i[10] peripherals_i/fll1_rdata_i[11]
+ peripherals_i/fll1_rdata_i[12] peripherals_i/fll1_rdata_i[13] peripherals_i/fll1_rdata_i[14]
+ peripherals_i/fll1_rdata_i[15] peripherals_i/fll1_rdata_i[16] peripherals_i/fll1_rdata_i[17]
+ peripherals_i/fll1_rdata_i[18] peripherals_i/fll1_rdata_i[19] peripherals_i/fll1_rdata_i[1]
+ peripherals_i/fll1_rdata_i[20] peripherals_i/fll1_rdata_i[21] peripherals_i/fll1_rdata_i[22]
+ peripherals_i/fll1_rdata_i[23] peripherals_i/fll1_rdata_i[24] peripherals_i/fll1_rdata_i[25]
+ peripherals_i/fll1_rdata_i[26] peripherals_i/fll1_rdata_i[27] peripherals_i/fll1_rdata_i[28]
+ peripherals_i/fll1_rdata_i[29] peripherals_i/fll1_rdata_i[2] peripherals_i/fll1_rdata_i[30]
+ peripherals_i/fll1_rdata_i[31] peripherals_i/fll1_rdata_i[3] peripherals_i/fll1_rdata_i[4]
+ peripherals_i/fll1_rdata_i[5] peripherals_i/fll1_rdata_i[6] peripherals_i/fll1_rdata_i[7]
+ peripherals_i/fll1_rdata_i[8] peripherals_i/fll1_rdata_i[9] peripherals_i/fll1_req_o
+ peripherals_i/fll1_wrn_o la_data_out[96] la_data_out[106] la_data_out[107] la_data_out[108]
+ la_data_out[109] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[97] la_data_out[116] la_data_out[117]
+ la_data_out[118] la_data_out[119] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[98] la_data_out[126]
+ la_data_out[127] la_data_out[99] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_in[7] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[8] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[9] la_data_in[37] la_data_in[38] la_data_in[10]
+ la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_out[64] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[65] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[66] la_data_out[94] la_data_out[95]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] peripherals_i/gpio_padcfg[0] peripherals_i/gpio_padcfg[100]
+ peripherals_i/gpio_padcfg[101] peripherals_i/gpio_padcfg[102] peripherals_i/gpio_padcfg[103]
+ peripherals_i/gpio_padcfg[104] peripherals_i/gpio_padcfg[105] peripherals_i/gpio_padcfg[106]
+ peripherals_i/gpio_padcfg[107] peripherals_i/gpio_padcfg[108] peripherals_i/gpio_padcfg[109]
+ peripherals_i/gpio_padcfg[10] peripherals_i/gpio_padcfg[110] peripherals_i/gpio_padcfg[111]
+ peripherals_i/gpio_padcfg[112] peripherals_i/gpio_padcfg[113] peripherals_i/gpio_padcfg[114]
+ peripherals_i/gpio_padcfg[115] peripherals_i/gpio_padcfg[116] peripherals_i/gpio_padcfg[117]
+ peripherals_i/gpio_padcfg[118] peripherals_i/gpio_padcfg[119] peripherals_i/gpio_padcfg[11]
+ peripherals_i/gpio_padcfg[120] peripherals_i/gpio_padcfg[121] peripherals_i/gpio_padcfg[122]
+ peripherals_i/gpio_padcfg[123] peripherals_i/gpio_padcfg[124] peripherals_i/gpio_padcfg[125]
+ peripherals_i/gpio_padcfg[126] peripherals_i/gpio_padcfg[127] peripherals_i/gpio_padcfg[128]
+ peripherals_i/gpio_padcfg[129] peripherals_i/gpio_padcfg[12] peripherals_i/gpio_padcfg[130]
+ peripherals_i/gpio_padcfg[131] peripherals_i/gpio_padcfg[132] peripherals_i/gpio_padcfg[133]
+ peripherals_i/gpio_padcfg[134] peripherals_i/gpio_padcfg[135] peripherals_i/gpio_padcfg[136]
+ peripherals_i/gpio_padcfg[137] peripherals_i/gpio_padcfg[138] peripherals_i/gpio_padcfg[139]
+ peripherals_i/gpio_padcfg[13] peripherals_i/gpio_padcfg[140] peripherals_i/gpio_padcfg[141]
+ peripherals_i/gpio_padcfg[142] peripherals_i/gpio_padcfg[143] peripherals_i/gpio_padcfg[144]
+ peripherals_i/gpio_padcfg[145] peripherals_i/gpio_padcfg[146] peripherals_i/gpio_padcfg[147]
+ peripherals_i/gpio_padcfg[148] peripherals_i/gpio_padcfg[149] peripherals_i/gpio_padcfg[14]
+ peripherals_i/gpio_padcfg[150] peripherals_i/gpio_padcfg[151] peripherals_i/gpio_padcfg[152]
+ peripherals_i/gpio_padcfg[153] peripherals_i/gpio_padcfg[154] peripherals_i/gpio_padcfg[155]
+ peripherals_i/gpio_padcfg[156] peripherals_i/gpio_padcfg[157] peripherals_i/gpio_padcfg[158]
+ peripherals_i/gpio_padcfg[159] peripherals_i/gpio_padcfg[15] peripherals_i/gpio_padcfg[160]
+ peripherals_i/gpio_padcfg[161] peripherals_i/gpio_padcfg[162] peripherals_i/gpio_padcfg[163]
+ peripherals_i/gpio_padcfg[164] peripherals_i/gpio_padcfg[165] peripherals_i/gpio_padcfg[166]
+ peripherals_i/gpio_padcfg[167] peripherals_i/gpio_padcfg[168] peripherals_i/gpio_padcfg[169]
+ peripherals_i/gpio_padcfg[16] peripherals_i/gpio_padcfg[170] peripherals_i/gpio_padcfg[171]
+ peripherals_i/gpio_padcfg[172] peripherals_i/gpio_padcfg[173] peripherals_i/gpio_padcfg[174]
+ peripherals_i/gpio_padcfg[175] peripherals_i/gpio_padcfg[176] peripherals_i/gpio_padcfg[177]
+ peripherals_i/gpio_padcfg[178] peripherals_i/gpio_padcfg[179] peripherals_i/gpio_padcfg[17]
+ peripherals_i/gpio_padcfg[180] peripherals_i/gpio_padcfg[181] peripherals_i/gpio_padcfg[182]
+ peripherals_i/gpio_padcfg[183] peripherals_i/gpio_padcfg[184] peripherals_i/gpio_padcfg[185]
+ peripherals_i/gpio_padcfg[186] peripherals_i/gpio_padcfg[187] peripherals_i/gpio_padcfg[188]
+ peripherals_i/gpio_padcfg[189] peripherals_i/gpio_padcfg[18] peripherals_i/gpio_padcfg[190]
+ peripherals_i/gpio_padcfg[191] peripherals_i/gpio_padcfg[19] peripherals_i/gpio_padcfg[1]
+ peripherals_i/gpio_padcfg[20] peripherals_i/gpio_padcfg[21] peripherals_i/gpio_padcfg[22]
+ peripherals_i/gpio_padcfg[23] peripherals_i/gpio_padcfg[24] peripherals_i/gpio_padcfg[25]
+ peripherals_i/gpio_padcfg[26] peripherals_i/gpio_padcfg[27] peripherals_i/gpio_padcfg[28]
+ peripherals_i/gpio_padcfg[29] peripherals_i/gpio_padcfg[2] peripherals_i/gpio_padcfg[30]
+ peripherals_i/gpio_padcfg[31] peripherals_i/gpio_padcfg[32] peripherals_i/gpio_padcfg[33]
+ peripherals_i/gpio_padcfg[34] peripherals_i/gpio_padcfg[35] peripherals_i/gpio_padcfg[36]
+ peripherals_i/gpio_padcfg[37] peripherals_i/gpio_padcfg[38] peripherals_i/gpio_padcfg[39]
+ peripherals_i/gpio_padcfg[3] peripherals_i/gpio_padcfg[40] peripherals_i/gpio_padcfg[41]
+ peripherals_i/gpio_padcfg[42] peripherals_i/gpio_padcfg[43] peripherals_i/gpio_padcfg[44]
+ peripherals_i/gpio_padcfg[45] peripherals_i/gpio_padcfg[46] peripherals_i/gpio_padcfg[47]
+ peripherals_i/gpio_padcfg[48] peripherals_i/gpio_padcfg[49] peripherals_i/gpio_padcfg[4]
+ peripherals_i/gpio_padcfg[50] peripherals_i/gpio_padcfg[51] peripherals_i/gpio_padcfg[52]
+ peripherals_i/gpio_padcfg[53] peripherals_i/gpio_padcfg[54] peripherals_i/gpio_padcfg[55]
+ peripherals_i/gpio_padcfg[56] peripherals_i/gpio_padcfg[57] peripherals_i/gpio_padcfg[58]
+ peripherals_i/gpio_padcfg[59] peripherals_i/gpio_padcfg[5] peripherals_i/gpio_padcfg[60]
+ peripherals_i/gpio_padcfg[61] peripherals_i/gpio_padcfg[62] peripherals_i/gpio_padcfg[63]
+ peripherals_i/gpio_padcfg[64] peripherals_i/gpio_padcfg[65] peripherals_i/gpio_padcfg[66]
+ peripherals_i/gpio_padcfg[67] peripherals_i/gpio_padcfg[68] peripherals_i/gpio_padcfg[69]
+ peripherals_i/gpio_padcfg[6] peripherals_i/gpio_padcfg[70] peripherals_i/gpio_padcfg[71]
+ peripherals_i/gpio_padcfg[72] peripherals_i/gpio_padcfg[73] peripherals_i/gpio_padcfg[74]
+ peripherals_i/gpio_padcfg[75] peripherals_i/gpio_padcfg[76] peripherals_i/gpio_padcfg[77]
+ peripherals_i/gpio_padcfg[78] peripherals_i/gpio_padcfg[79] peripherals_i/gpio_padcfg[7]
+ peripherals_i/gpio_padcfg[80] peripherals_i/gpio_padcfg[81] peripherals_i/gpio_padcfg[82]
+ peripherals_i/gpio_padcfg[83] peripherals_i/gpio_padcfg[84] peripherals_i/gpio_padcfg[85]
+ peripherals_i/gpio_padcfg[86] peripherals_i/gpio_padcfg[87] peripherals_i/gpio_padcfg[88]
+ peripherals_i/gpio_padcfg[89] peripherals_i/gpio_padcfg[8] peripherals_i/gpio_padcfg[90]
+ peripherals_i/gpio_padcfg[91] peripherals_i/gpio_padcfg[92] peripherals_i/gpio_padcfg[93]
+ peripherals_i/gpio_padcfg[94] peripherals_i/gpio_padcfg[95] peripherals_i/gpio_padcfg[96]
+ peripherals_i/gpio_padcfg[97] peripherals_i/gpio_padcfg[98] peripherals_i/gpio_padcfg[99]
+ peripherals_i/gpio_padcfg[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] peripherals_i/irq_o[0] peripherals_i/irq_o[10] peripherals_i/irq_o[11]
+ peripherals_i/irq_o[12] peripherals_i/irq_o[13] peripherals_i/irq_o[14] peripherals_i/irq_o[15]
+ peripherals_i/irq_o[16] peripherals_i/irq_o[17] peripherals_i/irq_o[18] peripherals_i/irq_o[19]
+ peripherals_i/irq_o[1] peripherals_i/irq_o[20] peripherals_i/irq_o[21] peripherals_i/irq_o[22]
+ peripherals_i/irq_o[23] peripherals_i/irq_o[24] peripherals_i/irq_o[25] peripherals_i/irq_o[26]
+ peripherals_i/irq_o[27] peripherals_i/irq_o[28] peripherals_i/irq_o[29] peripherals_i/irq_o[2]
+ peripherals_i/irq_o[30] peripherals_i/irq_o[31] peripherals_i/irq_o[3] peripherals_i/irq_o[4]
+ peripherals_i/irq_o[5] peripherals_i/irq_o[6] peripherals_i/irq_o[7] peripherals_i/irq_o[8]
+ peripherals_i/irq_o[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] peripherals_i/rst_n
+ wb_rst_i peripherals_i/rst_n la_data_in[3] io_in[21] peripherals_i/scan_o_pll io_in[22]
+ io_out[28] peripherals_i/scl_padoen_o io_in[23] io_out[27] peripherals_i/sda_padoen_o
+ peripherals_i/slave_ar_addr[0] peripherals_i/slave_ar_addr[10] peripherals_i/slave_ar_addr[11]
+ peripherals_i/slave_ar_addr[12] peripherals_i/slave_ar_addr[13] peripherals_i/slave_ar_addr[14]
+ peripherals_i/slave_ar_addr[15] peripherals_i/slave_ar_addr[16] peripherals_i/slave_ar_addr[17]
+ peripherals_i/slave_ar_addr[18] peripherals_i/slave_ar_addr[19] peripherals_i/slave_ar_addr[1]
+ peripherals_i/slave_ar_addr[20] peripherals_i/slave_ar_addr[21] peripherals_i/slave_ar_addr[22]
+ peripherals_i/slave_ar_addr[23] peripherals_i/slave_ar_addr[24] peripherals_i/slave_ar_addr[25]
+ peripherals_i/slave_ar_addr[26] peripherals_i/slave_ar_addr[27] peripherals_i/slave_ar_addr[28]
+ peripherals_i/slave_ar_addr[29] peripherals_i/slave_ar_addr[2] peripherals_i/slave_ar_addr[30]
+ peripherals_i/slave_ar_addr[31] peripherals_i/slave_ar_addr[3] peripherals_i/slave_ar_addr[4]
+ peripherals_i/slave_ar_addr[5] peripherals_i/slave_ar_addr[6] peripherals_i/slave_ar_addr[7]
+ peripherals_i/slave_ar_addr[8] peripherals_i/slave_ar_addr[9] peripherals_i/slave_ar_burst[0]
+ peripherals_i/slave_ar_burst[1] peripherals_i/slave_ar_cache[0] peripherals_i/slave_ar_cache[1]
+ peripherals_i/slave_ar_cache[2] peripherals_i/slave_ar_cache[3] peripherals_i/slave_ar_id[0]
+ peripherals_i/slave_ar_id[1] peripherals_i/slave_ar_id[2] peripherals_i/slave_ar_id[3]
+ peripherals_i/slave_ar_id[4] peripherals_i/slave_ar_id[5] peripherals_i/slave_ar_len[0]
+ peripherals_i/slave_ar_len[1] peripherals_i/slave_ar_len[2] peripherals_i/slave_ar_len[3]
+ peripherals_i/slave_ar_len[4] peripherals_i/slave_ar_len[5] peripherals_i/slave_ar_len[6]
+ peripherals_i/slave_ar_len[7] peripherals_i/slave_ar_lock peripherals_i/slave_ar_prot[0]
+ peripherals_i/slave_ar_prot[1] peripherals_i/slave_ar_prot[2] peripherals_i/slave_ar_qos[0]
+ peripherals_i/slave_ar_qos[1] peripherals_i/slave_ar_qos[2] peripherals_i/slave_ar_qos[3]
+ peripherals_i/slave_ar_ready peripherals_i/slave_ar_region[0] peripherals_i/slave_ar_region[1]
+ peripherals_i/slave_ar_region[2] peripherals_i/slave_ar_region[3] peripherals_i/slave_ar_size[0]
+ peripherals_i/slave_ar_size[1] peripherals_i/slave_ar_size[2] peripherals_i/slave_ar_user[0]
+ peripherals_i/slave_ar_user[1] peripherals_i/slave_ar_user[2] peripherals_i/slave_ar_user[3]
+ peripherals_i/slave_ar_user[4] peripherals_i/slave_ar_user[5] peripherals_i/slave_ar_valid
+ peripherals_i/slave_aw_addr[0] peripherals_i/slave_aw_addr[10] peripherals_i/slave_aw_addr[11]
+ peripherals_i/slave_aw_addr[12] peripherals_i/slave_aw_addr[13] peripherals_i/slave_aw_addr[14]
+ peripherals_i/slave_aw_addr[15] peripherals_i/slave_aw_addr[16] peripherals_i/slave_aw_addr[17]
+ peripherals_i/slave_aw_addr[18] peripherals_i/slave_aw_addr[19] peripherals_i/slave_aw_addr[1]
+ peripherals_i/slave_aw_addr[20] peripherals_i/slave_aw_addr[21] peripherals_i/slave_aw_addr[22]
+ peripherals_i/slave_aw_addr[23] peripherals_i/slave_aw_addr[24] peripherals_i/slave_aw_addr[25]
+ peripherals_i/slave_aw_addr[26] peripherals_i/slave_aw_addr[27] peripherals_i/slave_aw_addr[28]
+ peripherals_i/slave_aw_addr[29] peripherals_i/slave_aw_addr[2] peripherals_i/slave_aw_addr[30]
+ peripherals_i/slave_aw_addr[31] peripherals_i/slave_aw_addr[3] peripherals_i/slave_aw_addr[4]
+ peripherals_i/slave_aw_addr[5] peripherals_i/slave_aw_addr[6] peripherals_i/slave_aw_addr[7]
+ peripherals_i/slave_aw_addr[8] peripherals_i/slave_aw_addr[9] peripherals_i/slave_aw_burst[0]
+ peripherals_i/slave_aw_burst[1] peripherals_i/slave_aw_cache[0] peripherals_i/slave_aw_cache[1]
+ peripherals_i/slave_aw_cache[2] peripherals_i/slave_aw_cache[3] peripherals_i/slave_aw_id[0]
+ peripherals_i/slave_aw_id[1] peripherals_i/slave_aw_id[2] peripherals_i/slave_aw_id[3]
+ peripherals_i/slave_aw_id[4] peripherals_i/slave_aw_id[5] peripherals_i/slave_aw_len[0]
+ peripherals_i/slave_aw_len[1] peripherals_i/slave_aw_len[2] peripherals_i/slave_aw_len[3]
+ peripherals_i/slave_aw_len[4] peripherals_i/slave_aw_len[5] peripherals_i/slave_aw_len[6]
+ peripherals_i/slave_aw_len[7] peripherals_i/slave_aw_lock peripherals_i/slave_aw_prot[0]
+ peripherals_i/slave_aw_prot[1] peripherals_i/slave_aw_prot[2] peripherals_i/slave_aw_qos[0]
+ peripherals_i/slave_aw_qos[1] peripherals_i/slave_aw_qos[2] peripherals_i/slave_aw_qos[3]
+ peripherals_i/slave_aw_ready peripherals_i/slave_aw_region[0] peripherals_i/slave_aw_region[1]
+ peripherals_i/slave_aw_region[2] peripherals_i/slave_aw_region[3] peripherals_i/slave_aw_size[0]
+ peripherals_i/slave_aw_size[1] peripherals_i/slave_aw_size[2] peripherals_i/slave_aw_user[0]
+ peripherals_i/slave_aw_user[1] peripherals_i/slave_aw_user[2] peripherals_i/slave_aw_user[3]
+ peripherals_i/slave_aw_user[4] peripherals_i/slave_aw_user[5] peripherals_i/slave_aw_valid
+ peripherals_i/slave_b_id[0] peripherals_i/slave_b_id[1] peripherals_i/slave_b_id[2]
+ peripherals_i/slave_b_id[3] peripherals_i/slave_b_id[4] peripherals_i/slave_b_id[5]
+ peripherals_i/slave_b_ready peripherals_i/slave_b_resp[0] peripherals_i/slave_b_resp[1]
+ peripherals_i/slave_b_user[0] peripherals_i/slave_b_user[1] peripherals_i/slave_b_user[2]
+ peripherals_i/slave_b_user[3] peripherals_i/slave_b_user[4] peripherals_i/slave_b_user[5]
+ peripherals_i/slave_b_valid peripherals_i/slave_r_data[0] peripherals_i/slave_r_data[10]
+ peripherals_i/slave_r_data[11] peripherals_i/slave_r_data[12] peripherals_i/slave_r_data[13]
+ peripherals_i/slave_r_data[14] peripherals_i/slave_r_data[15] peripherals_i/slave_r_data[16]
+ peripherals_i/slave_r_data[17] peripherals_i/slave_r_data[18] peripherals_i/slave_r_data[19]
+ peripherals_i/slave_r_data[1] peripherals_i/slave_r_data[20] peripherals_i/slave_r_data[21]
+ peripherals_i/slave_r_data[22] peripherals_i/slave_r_data[23] peripherals_i/slave_r_data[24]
+ peripherals_i/slave_r_data[25] peripherals_i/slave_r_data[26] peripherals_i/slave_r_data[27]
+ peripherals_i/slave_r_data[28] peripherals_i/slave_r_data[29] peripherals_i/slave_r_data[2]
+ peripherals_i/slave_r_data[30] peripherals_i/slave_r_data[31] peripherals_i/slave_r_data[32]
+ peripherals_i/slave_r_data[33] peripherals_i/slave_r_data[34] peripherals_i/slave_r_data[35]
+ peripherals_i/slave_r_data[36] peripherals_i/slave_r_data[37] peripherals_i/slave_r_data[38]
+ peripherals_i/slave_r_data[39] peripherals_i/slave_r_data[3] peripherals_i/slave_r_data[40]
+ peripherals_i/slave_r_data[41] peripherals_i/slave_r_data[42] peripherals_i/slave_r_data[43]
+ peripherals_i/slave_r_data[44] peripherals_i/slave_r_data[45] peripherals_i/slave_r_data[46]
+ peripherals_i/slave_r_data[47] peripherals_i/slave_r_data[48] peripherals_i/slave_r_data[49]
+ peripherals_i/slave_r_data[4] peripherals_i/slave_r_data[50] peripherals_i/slave_r_data[51]
+ peripherals_i/slave_r_data[52] peripherals_i/slave_r_data[53] peripherals_i/slave_r_data[54]
+ peripherals_i/slave_r_data[55] peripherals_i/slave_r_data[56] peripherals_i/slave_r_data[57]
+ peripherals_i/slave_r_data[58] peripherals_i/slave_r_data[59] peripherals_i/slave_r_data[5]
+ peripherals_i/slave_r_data[60] peripherals_i/slave_r_data[61] peripherals_i/slave_r_data[62]
+ peripherals_i/slave_r_data[63] peripherals_i/slave_r_data[6] peripherals_i/slave_r_data[7]
+ peripherals_i/slave_r_data[8] peripherals_i/slave_r_data[9] peripherals_i/slave_r_id[0]
+ peripherals_i/slave_r_id[1] peripherals_i/slave_r_id[2] peripherals_i/slave_r_id[3]
+ peripherals_i/slave_r_id[4] peripherals_i/slave_r_id[5] peripherals_i/slave_r_last
+ peripherals_i/slave_r_ready peripherals_i/slave_r_resp[0] peripherals_i/slave_r_resp[1]
+ peripherals_i/slave_r_user[0] peripherals_i/slave_r_user[1] peripherals_i/slave_r_user[2]
+ peripherals_i/slave_r_user[3] peripherals_i/slave_r_user[4] peripherals_i/slave_r_user[5]
+ peripherals_i/slave_r_valid peripherals_i/slave_w_data[0] peripherals_i/slave_w_data[10]
+ peripherals_i/slave_w_data[11] peripherals_i/slave_w_data[12] peripherals_i/slave_w_data[13]
+ peripherals_i/slave_w_data[14] peripherals_i/slave_w_data[15] peripherals_i/slave_w_data[16]
+ peripherals_i/slave_w_data[17] peripherals_i/slave_w_data[18] peripherals_i/slave_w_data[19]
+ peripherals_i/slave_w_data[1] peripherals_i/slave_w_data[20] peripherals_i/slave_w_data[21]
+ peripherals_i/slave_w_data[22] peripherals_i/slave_w_data[23] peripherals_i/slave_w_data[24]
+ peripherals_i/slave_w_data[25] peripherals_i/slave_w_data[26] peripherals_i/slave_w_data[27]
+ peripherals_i/slave_w_data[28] peripherals_i/slave_w_data[29] peripherals_i/slave_w_data[2]
+ peripherals_i/slave_w_data[30] peripherals_i/slave_w_data[31] peripherals_i/slave_w_data[32]
+ peripherals_i/slave_w_data[33] peripherals_i/slave_w_data[34] peripherals_i/slave_w_data[35]
+ peripherals_i/slave_w_data[36] peripherals_i/slave_w_data[37] peripherals_i/slave_w_data[38]
+ peripherals_i/slave_w_data[39] peripherals_i/slave_w_data[3] peripherals_i/slave_w_data[40]
+ peripherals_i/slave_w_data[41] peripherals_i/slave_w_data[42] peripherals_i/slave_w_data[43]
+ peripherals_i/slave_w_data[44] peripherals_i/slave_w_data[45] peripherals_i/slave_w_data[46]
+ peripherals_i/slave_w_data[47] peripherals_i/slave_w_data[48] peripherals_i/slave_w_data[49]
+ peripherals_i/slave_w_data[4] peripherals_i/slave_w_data[50] peripherals_i/slave_w_data[51]
+ peripherals_i/slave_w_data[52] peripherals_i/slave_w_data[53] peripherals_i/slave_w_data[54]
+ peripherals_i/slave_w_data[55] peripherals_i/slave_w_data[56] peripherals_i/slave_w_data[57]
+ peripherals_i/slave_w_data[58] peripherals_i/slave_w_data[59] peripherals_i/slave_w_data[5]
+ peripherals_i/slave_w_data[60] peripherals_i/slave_w_data[61] peripherals_i/slave_w_data[62]
+ peripherals_i/slave_w_data[63] peripherals_i/slave_w_data[6] peripherals_i/slave_w_data[7]
+ peripherals_i/slave_w_data[8] peripherals_i/slave_w_data[9] peripherals_i/slave_w_last
+ peripherals_i/slave_w_ready peripherals_i/slave_w_strb[0] peripherals_i/slave_w_strb[1]
+ peripherals_i/slave_w_strb[2] peripherals_i/slave_w_strb[3] peripherals_i/slave_w_strb[4]
+ peripherals_i/slave_w_strb[5] peripherals_i/slave_w_strb[6] peripherals_i/slave_w_strb[7]
+ peripherals_i/slave_w_user[0] peripherals_i/slave_w_user[1] peripherals_i/slave_w_user[2]
+ peripherals_i/slave_w_user[3] peripherals_i/slave_w_user[4] peripherals_i/slave_w_user[5]
+ peripherals_i/slave_w_valid io_in[17] io_in[18] io_out[33] io_out[32] peripherals_i/spi_master_csn1
+ peripherals_i/spi_master_csn2 peripherals_i/spi_master_csn3 io_out[30] io_out[31]
+ io_in[21] io_in[21] io_in[21] io_in[21] io_out[29] peripherals_i/spi_master_sdo1
+ peripherals_i/spi_master_sdo2 peripherals_i/spi_master_sdo3 io_out[36] io_out[37]
+ io_in[19] io_in[21] io_in[21] io_in[21] io_out[35] peripherals_i/spi_sdo1_o peripherals_i/spi_sdo2_o
+ peripherals_i/spi_sdo3_o la_data_in[2] la_data_in[2] la_data_in[4] la_data_in[5]
+ peripherals_i/uart_dtr peripherals_i/uart_rts io_in[20] io_out[34] user_irq[0] user_irq[1]
+ user_irq[2] vccd1 vssd1 wbs_ack_o wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12]
+ wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18]
+ wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23]
+ wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29]
+ wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5]
+ wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] peripherals
.ends

