magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 891 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 531 47 561 177
rect 615 47 645 177
rect 699 47 729 177
rect 783 47 813 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 531 297 561 497
rect 615 297 645 497
rect 699 297 729 497
rect 783 297 813 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 421 177
rect 365 61 375 95
rect 409 61 421 95
rect 365 47 421 61
rect 475 95 531 177
rect 475 61 487 95
rect 521 61 531 95
rect 475 47 531 61
rect 561 163 615 177
rect 561 129 571 163
rect 605 129 615 163
rect 561 95 615 129
rect 561 61 571 95
rect 605 61 615 95
rect 561 47 615 61
rect 645 95 699 177
rect 645 61 655 95
rect 689 61 699 95
rect 645 47 699 61
rect 729 163 783 177
rect 729 129 739 163
rect 773 129 783 163
rect 729 95 783 129
rect 729 61 739 95
rect 773 61 783 95
rect 729 47 783 61
rect 813 95 865 177
rect 813 61 823 95
rect 857 61 865 95
rect 813 47 865 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 409 335 443
rect 281 375 291 409
rect 325 375 335 409
rect 281 297 335 375
rect 365 409 421 497
rect 365 375 375 409
rect 409 375 421 409
rect 365 341 421 375
rect 365 307 375 341
rect 409 307 421 341
rect 365 297 421 307
rect 475 409 531 497
rect 475 375 487 409
rect 521 375 531 409
rect 475 341 531 375
rect 475 307 487 341
rect 521 307 531 341
rect 475 297 531 307
rect 561 477 615 497
rect 561 443 571 477
rect 605 443 615 477
rect 561 409 615 443
rect 561 375 571 409
rect 605 375 615 409
rect 561 297 615 375
rect 645 477 699 497
rect 645 443 655 477
rect 689 443 699 477
rect 645 409 699 443
rect 645 375 655 409
rect 689 375 699 409
rect 645 341 699 375
rect 645 307 655 341
rect 689 307 699 341
rect 645 297 699 307
rect 729 409 783 497
rect 729 375 739 409
rect 773 375 783 409
rect 729 341 783 375
rect 729 307 739 341
rect 773 307 783 341
rect 729 297 783 307
rect 813 477 865 497
rect 813 443 823 477
rect 857 443 865 477
rect 813 409 865 443
rect 813 375 823 409
rect 857 375 865 409
rect 813 297 865 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 487 61 521 95
rect 571 129 605 163
rect 571 61 605 95
rect 655 61 689 95
rect 739 129 773 163
rect 739 61 773 95
rect 823 61 857 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 443 325 477
rect 291 375 325 409
rect 375 375 409 409
rect 375 307 409 341
rect 487 375 521 409
rect 487 307 521 341
rect 571 443 605 477
rect 571 375 605 409
rect 655 443 689 477
rect 655 375 689 409
rect 655 307 689 341
rect 739 375 773 409
rect 739 307 773 341
rect 823 443 857 477
rect 823 375 857 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 531 497 561 523
rect 615 497 645 523
rect 699 497 729 523
rect 783 497 813 523
rect 83 265 113 297
rect 167 265 197 297
rect 83 249 197 265
rect 83 215 112 249
rect 146 215 197 249
rect 83 199 197 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 265 281 297
rect 335 265 365 297
rect 251 249 365 265
rect 251 215 288 249
rect 322 215 365 249
rect 251 199 365 215
rect 251 177 281 199
rect 335 177 365 199
rect 531 265 561 297
rect 615 265 645 297
rect 531 249 645 265
rect 531 215 571 249
rect 605 215 645 249
rect 531 199 645 215
rect 531 177 561 199
rect 615 177 645 199
rect 699 265 729 297
rect 783 265 813 297
rect 699 249 813 265
rect 699 215 735 249
rect 769 215 813 249
rect 699 199 813 215
rect 699 177 729 199
rect 783 177 813 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 531 21 561 47
rect 615 21 645 47
rect 699 21 729 47
rect 783 21 813 47
<< polycont >>
rect 112 215 146 249
rect 288 215 322 249
rect 571 215 605 249
rect 735 215 769 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 30 307 39 341
rect 73 325 81 341
rect 199 341 249 375
rect 283 477 613 493
rect 283 443 291 477
rect 325 459 571 477
rect 325 443 333 459
rect 283 409 333 443
rect 563 443 571 459
rect 605 443 613 477
rect 283 375 291 409
rect 325 375 333 409
rect 283 359 333 375
rect 367 409 417 425
rect 367 375 375 409
rect 409 375 417 409
rect 199 325 207 341
rect 73 307 207 325
rect 241 325 249 341
rect 367 341 417 375
rect 367 325 375 341
rect 241 307 375 325
rect 409 307 417 341
rect 30 291 417 307
rect 479 409 529 425
rect 479 375 487 409
rect 521 375 529 409
rect 479 341 529 375
rect 563 409 613 443
rect 563 375 571 409
rect 605 375 613 409
rect 563 359 613 375
rect 647 477 865 493
rect 647 443 655 477
rect 689 459 823 477
rect 689 443 697 459
rect 647 409 697 443
rect 815 443 823 459
rect 857 443 865 477
rect 647 375 655 409
rect 689 375 697 409
rect 479 307 487 341
rect 521 325 529 341
rect 647 341 697 375
rect 647 325 655 341
rect 521 307 655 325
rect 689 307 697 341
rect 479 291 697 307
rect 731 409 781 425
rect 731 375 739 409
rect 773 375 781 409
rect 731 341 781 375
rect 815 409 865 443
rect 815 375 823 409
rect 857 375 865 409
rect 815 359 865 375
rect 731 307 739 341
rect 773 325 781 341
rect 773 307 903 325
rect 731 291 903 307
rect 40 249 193 257
rect 40 215 112 249
rect 146 215 193 249
rect 227 249 388 257
rect 227 215 288 249
rect 322 215 388 249
rect 442 249 621 257
rect 442 215 571 249
rect 605 215 621 249
rect 668 249 785 257
rect 668 215 735 249
rect 769 215 785 249
rect 836 181 903 291
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 903 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 571 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 555 129 571 145
rect 605 145 739 163
rect 605 129 621 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 521 111
rect 409 61 487 95
rect 375 17 521 61
rect 555 95 621 129
rect 723 129 739 145
rect 773 145 903 163
rect 773 129 789 145
rect 555 61 571 95
rect 605 61 621 95
rect 555 51 621 61
rect 655 95 689 111
rect 655 17 689 61
rect 723 95 789 129
rect 723 61 739 95
rect 773 61 789 95
rect 723 51 789 61
rect 823 95 881 111
rect 857 61 881 95
rect 823 17 881 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 494 221 528 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 862 153 896 187 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1159106
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1151456
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
