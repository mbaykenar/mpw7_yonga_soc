VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clk_rst_gen
  CLASS BLOCK ;
  FOREIGN clk_rst_gen ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 150.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 74.840 250.000 75.440 ;
    END
  END clk_i
  PIN clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END clk_o
  PIN clk_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 146.000 22.910 150.000 ;
    END
  END clk_sel_i
  PIN clk_standalone_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END clk_standalone_i
  PIN fll_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END fll_ack_o
  PIN fll_add_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 146.240 250.000 146.840 ;
    END
  END fll_add_i[0]
  PIN fll_add_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END fll_add_i[1]
  PIN fll_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 146.000 84.090 150.000 ;
    END
  END fll_data_i[0]
  PIN fll_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END fll_data_i[10]
  PIN fll_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 150.000 ;
    END
  END fll_data_i[11]
  PIN fll_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 105.440 250.000 106.040 ;
    END
  END fll_data_i[12]
  PIN fll_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END fll_data_i[13]
  PIN fll_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 146.000 164.590 150.000 ;
    END
  END fll_data_i[14]
  PIN fll_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 146.000 71.210 150.000 ;
    END
  END fll_data_i[15]
  PIN fll_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 40.840 250.000 41.440 ;
    END
  END fll_data_i[16]
  PIN fll_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END fll_data_i[17]
  PIN fll_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END fll_data_i[18]
  PIN fll_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 146.000 158.150 150.000 ;
    END
  END fll_data_i[19]
  PIN fll_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 146.000 135.610 150.000 ;
    END
  END fll_data_i[1]
  PIN fll_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END fll_data_i[20]
  PIN fll_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 51.040 250.000 51.640 ;
    END
  END fll_data_i[21]
  PIN fll_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END fll_data_i[22]
  PIN fll_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END fll_data_i[23]
  PIN fll_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 54.440 250.000 55.040 ;
    END
  END fll_data_i[24]
  PIN fll_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 146.000 196.790 150.000 ;
    END
  END fll_data_i[25]
  PIN fll_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END fll_data_i[26]
  PIN fll_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 146.000 222.550 150.000 ;
    END
  END fll_data_i[27]
  PIN fll_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 146.000 13.250 150.000 ;
    END
  END fll_data_i[28]
  PIN fll_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END fll_data_i[29]
  PIN fll_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END fll_data_i[2]
  PIN fll_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END fll_data_i[30]
  PIN fll_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 27.240 250.000 27.840 ;
    END
  END fll_data_i[31]
  PIN fll_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 146.000 87.310 150.000 ;
    END
  END fll_data_i[3]
  PIN fll_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END fll_data_i[4]
  PIN fll_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END fll_data_i[5]
  PIN fll_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END fll_data_i[6]
  PIN fll_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END fll_data_i[7]
  PIN fll_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 146.000 148.490 150.000 ;
    END
  END fll_data_i[8]
  PIN fll_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END fll_data_i[9]
  PIN fll_lock_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END fll_lock_o
  PIN fll_r_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 61.240 250.000 61.840 ;
    END
  END fll_r_data_o[0]
  PIN fll_r_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END fll_r_data_o[10]
  PIN fll_r_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 146.000 26.130 150.000 ;
    END
  END fll_r_data_o[11]
  PIN fll_r_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 146.000 154.930 150.000 ;
    END
  END fll_r_data_o[12]
  PIN fll_r_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 23.840 250.000 24.440 ;
    END
  END fll_r_data_o[13]
  PIN fll_r_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 20.440 250.000 21.040 ;
    END
  END fll_r_data_o[14]
  PIN fll_r_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 78.240 250.000 78.840 ;
    END
  END fll_r_data_o[15]
  PIN fll_r_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END fll_r_data_o[16]
  PIN fll_r_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 146.000 232.210 150.000 ;
    END
  END fll_r_data_o[17]
  PIN fll_r_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END fll_r_data_o[18]
  PIN fll_r_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 85.040 250.000 85.640 ;
    END
  END fll_r_data_o[19]
  PIN fll_r_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 146.000 132.390 150.000 ;
    END
  END fll_r_data_o[1]
  PIN fll_r_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 150.000 ;
    END
  END fll_r_data_o[20]
  PIN fll_r_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 146.000 32.570 150.000 ;
    END
  END fll_r_data_o[21]
  PIN fll_r_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END fll_r_data_o[22]
  PIN fll_r_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 146.000 216.110 150.000 ;
    END
  END fll_r_data_o[23]
  PIN fll_r_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END fll_r_data_o[24]
  PIN fll_r_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END fll_r_data_o[25]
  PIN fll_r_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 132.640 250.000 133.240 ;
    END
  END fll_r_data_o[26]
  PIN fll_r_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 146.000 10.030 150.000 ;
    END
  END fll_r_data_o[27]
  PIN fll_r_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 146.000 206.450 150.000 ;
    END
  END fll_r_data_o[28]
  PIN fll_r_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.000 103.410 150.000 ;
    END
  END fll_r_data_o[29]
  PIN fll_r_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 119.040 250.000 119.640 ;
    END
  END fll_r_data_o[2]
  PIN fll_r_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 146.000 161.370 150.000 ;
    END
  END fll_r_data_o[30]
  PIN fll_r_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 47.640 250.000 48.240 ;
    END
  END fll_r_data_o[31]
  PIN fll_r_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END fll_r_data_o[3]
  PIN fll_r_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END fll_r_data_o[4]
  PIN fll_r_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END fll_r_data_o[5]
  PIN fll_r_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 102.040 250.000 102.640 ;
    END
  END fll_r_data_o[6]
  PIN fll_r_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.000 55.110 150.000 ;
    END
  END fll_r_data_o[7]
  PIN fll_r_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END fll_r_data_o[8]
  PIN fll_r_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 146.000 90.530 150.000 ;
    END
  END fll_r_data_o[9]
  PIN fll_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 146.000 212.890 150.000 ;
    END
  END fll_req_i
  PIN fll_wrn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END fll_wrn_i
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 146.000 145.270 150.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 146.000 177.470 150.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 146.000 174.250 150.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 146.000 203.230 150.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 146.000 6.810 150.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 129.240 250.000 129.840 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 13.640 250.000 14.240 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 146.000 109.850 150.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 57.840 250.000 58.440 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 146.000 228.990 150.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 3.440 250.000 4.040 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 146.000 116.290 150.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 146.000 238.650 150.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 146.000 167.810 150.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 150.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 34.040 250.000 34.640 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 150.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.000 58.330 150.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 146.000 138.830 150.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 136.040 250.000 136.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.000 113.070 150.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 146.000 119.510 150.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.040 4.000 0.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 91.840 250.000 92.440 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 146.000 142.050 150.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 146.000 248.310 150.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.000 48.670 150.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_out[25]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 146.000 64.770 150.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.000 61.550 150.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 146.000 235.430 150.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 146.000 245.090 150.000 ;
    END
  END io_out[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 142.840 250.000 143.440 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 146.000 193.570 150.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 17.040 250.000 17.640 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 146.000 122.730 150.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 0.040 250.000 0.640 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 125.840 250.000 126.440 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 81.640 250.000 82.240 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 146.000 74.430 150.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 146.000 180.690 150.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 146.000 209.670 150.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 6.840 250.000 7.440 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 71.440 250.000 72.040 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 115.640 250.000 116.240 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 146.000 29.350 150.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 122.440 250.000 123.040 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 150.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 146.000 190.350 150.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 68.040 250.000 68.640 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 150.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 146.000 106.630 150.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 146.000 100.190 150.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 146.000 39.010 150.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 30.640 250.000 31.240 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 112.240 250.000 112.840 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 146.000 45.450 150.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 64.640 250.000 65.240 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 139.440 250.000 140.040 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 146.000 151.710 150.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END la_data_out[9]
  PIN rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 10.240 250.000 10.840 ;
    END
  END rstn_i
  PIN rstn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 146.000 241.870 150.000 ;
    END
  END rstn_o
  PIN scan_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 98.640 250.000 99.240 ;
    END
  END scan_en_i
  PIN scan_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END scan_i
  PIN scan_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END scan_o
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 37.440 250.000 38.040 ;
    END
  END testmode_i
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 108.840 250.000 109.440 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 146.000 225.770 150.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 34.590 10.640 36.190 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.330 10.640 95.930 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.070 10.640 155.670 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.810 10.640 215.410 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 64.460 10.640 66.060 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.200 10.640 125.800 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.940 10.640 185.540 138.960 ;
    END
  END vssd1
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 146.000 219.330 150.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 146.000 51.890 150.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 146.000 129.170 150.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 146.000 171.030 150.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 146.000 125.950 150.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 146.000 200.010 150.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 146.000 0.370 150.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 95.240 250.000 95.840 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 88.440 250.000 89.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 146.000 187.130 150.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 146.000 183.910 150.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 146.000 42.230 150.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 146.000 77.650 150.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 146.000 19.690 150.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 44.240 250.000 44.840 ;
    END
  END wbs_dat_o[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 138.805 ;
      LAYER met1 ;
        RECT 0.070 10.640 248.330 138.960 ;
      LAYER met2 ;
        RECT 0.650 145.720 3.030 146.725 ;
        RECT 3.870 145.720 6.250 146.725 ;
        RECT 7.090 145.720 9.470 146.725 ;
        RECT 10.310 145.720 12.690 146.725 ;
        RECT 13.530 145.720 15.910 146.725 ;
        RECT 16.750 145.720 19.130 146.725 ;
        RECT 19.970 145.720 22.350 146.725 ;
        RECT 23.190 145.720 25.570 146.725 ;
        RECT 26.410 145.720 28.790 146.725 ;
        RECT 29.630 145.720 32.010 146.725 ;
        RECT 32.850 145.720 35.230 146.725 ;
        RECT 36.070 145.720 38.450 146.725 ;
        RECT 39.290 145.720 41.670 146.725 ;
        RECT 42.510 145.720 44.890 146.725 ;
        RECT 45.730 145.720 48.110 146.725 ;
        RECT 48.950 145.720 51.330 146.725 ;
        RECT 52.170 145.720 54.550 146.725 ;
        RECT 55.390 145.720 57.770 146.725 ;
        RECT 58.610 145.720 60.990 146.725 ;
        RECT 61.830 145.720 64.210 146.725 ;
        RECT 65.050 145.720 67.430 146.725 ;
        RECT 68.270 145.720 70.650 146.725 ;
        RECT 71.490 145.720 73.870 146.725 ;
        RECT 74.710 145.720 77.090 146.725 ;
        RECT 77.930 145.720 80.310 146.725 ;
        RECT 81.150 145.720 83.530 146.725 ;
        RECT 84.370 145.720 86.750 146.725 ;
        RECT 87.590 145.720 89.970 146.725 ;
        RECT 90.810 145.720 93.190 146.725 ;
        RECT 94.030 145.720 96.410 146.725 ;
        RECT 97.250 145.720 99.630 146.725 ;
        RECT 100.470 145.720 102.850 146.725 ;
        RECT 103.690 145.720 106.070 146.725 ;
        RECT 106.910 145.720 109.290 146.725 ;
        RECT 110.130 145.720 112.510 146.725 ;
        RECT 113.350 145.720 115.730 146.725 ;
        RECT 116.570 145.720 118.950 146.725 ;
        RECT 119.790 145.720 122.170 146.725 ;
        RECT 123.010 145.720 125.390 146.725 ;
        RECT 126.230 145.720 128.610 146.725 ;
        RECT 129.450 145.720 131.830 146.725 ;
        RECT 132.670 145.720 135.050 146.725 ;
        RECT 135.890 145.720 138.270 146.725 ;
        RECT 139.110 145.720 141.490 146.725 ;
        RECT 142.330 145.720 144.710 146.725 ;
        RECT 145.550 145.720 147.930 146.725 ;
        RECT 148.770 145.720 151.150 146.725 ;
        RECT 151.990 145.720 154.370 146.725 ;
        RECT 155.210 145.720 157.590 146.725 ;
        RECT 158.430 145.720 160.810 146.725 ;
        RECT 161.650 145.720 164.030 146.725 ;
        RECT 164.870 145.720 167.250 146.725 ;
        RECT 168.090 145.720 170.470 146.725 ;
        RECT 171.310 145.720 173.690 146.725 ;
        RECT 174.530 145.720 176.910 146.725 ;
        RECT 177.750 145.720 180.130 146.725 ;
        RECT 180.970 145.720 183.350 146.725 ;
        RECT 184.190 145.720 186.570 146.725 ;
        RECT 187.410 145.720 189.790 146.725 ;
        RECT 190.630 145.720 193.010 146.725 ;
        RECT 193.850 145.720 196.230 146.725 ;
        RECT 197.070 145.720 199.450 146.725 ;
        RECT 200.290 145.720 202.670 146.725 ;
        RECT 203.510 145.720 205.890 146.725 ;
        RECT 206.730 145.720 209.110 146.725 ;
        RECT 209.950 145.720 212.330 146.725 ;
        RECT 213.170 145.720 215.550 146.725 ;
        RECT 216.390 145.720 218.770 146.725 ;
        RECT 219.610 145.720 221.990 146.725 ;
        RECT 222.830 145.720 225.210 146.725 ;
        RECT 226.050 145.720 228.430 146.725 ;
        RECT 229.270 145.720 231.650 146.725 ;
        RECT 232.490 145.720 234.870 146.725 ;
        RECT 235.710 145.720 238.090 146.725 ;
        RECT 238.930 145.720 241.310 146.725 ;
        RECT 242.150 145.720 244.530 146.725 ;
        RECT 245.370 145.720 247.750 146.725 ;
        RECT 0.100 4.280 248.300 145.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
      LAYER met3 ;
        RECT 4.400 145.840 245.600 146.705 ;
        RECT 4.000 143.840 246.000 145.840 ;
        RECT 4.400 142.440 245.600 143.840 ;
        RECT 4.000 140.440 246.000 142.440 ;
        RECT 4.400 139.040 245.600 140.440 ;
        RECT 4.000 137.040 246.000 139.040 ;
        RECT 4.400 135.640 245.600 137.040 ;
        RECT 4.000 133.640 246.000 135.640 ;
        RECT 4.400 132.240 245.600 133.640 ;
        RECT 4.000 130.240 246.000 132.240 ;
        RECT 4.400 128.840 245.600 130.240 ;
        RECT 4.000 126.840 246.000 128.840 ;
        RECT 4.400 125.440 245.600 126.840 ;
        RECT 4.000 123.440 246.000 125.440 ;
        RECT 4.400 122.040 245.600 123.440 ;
        RECT 4.000 120.040 246.000 122.040 ;
        RECT 4.400 118.640 245.600 120.040 ;
        RECT 4.000 116.640 246.000 118.640 ;
        RECT 4.400 115.240 245.600 116.640 ;
        RECT 4.000 113.240 246.000 115.240 ;
        RECT 4.400 111.840 245.600 113.240 ;
        RECT 4.000 109.840 246.000 111.840 ;
        RECT 4.400 108.440 245.600 109.840 ;
        RECT 4.000 106.440 246.000 108.440 ;
        RECT 4.400 105.040 245.600 106.440 ;
        RECT 4.000 103.040 246.000 105.040 ;
        RECT 4.400 101.640 245.600 103.040 ;
        RECT 4.000 99.640 246.000 101.640 ;
        RECT 4.400 98.240 245.600 99.640 ;
        RECT 4.000 96.240 246.000 98.240 ;
        RECT 4.400 94.840 245.600 96.240 ;
        RECT 4.000 92.840 246.000 94.840 ;
        RECT 4.400 91.440 245.600 92.840 ;
        RECT 4.000 89.440 246.000 91.440 ;
        RECT 4.400 88.040 245.600 89.440 ;
        RECT 4.000 86.040 246.000 88.040 ;
        RECT 4.400 84.640 245.600 86.040 ;
        RECT 4.000 82.640 246.000 84.640 ;
        RECT 4.400 81.240 245.600 82.640 ;
        RECT 4.000 79.240 246.000 81.240 ;
        RECT 4.400 77.840 245.600 79.240 ;
        RECT 4.000 75.840 246.000 77.840 ;
        RECT 4.400 74.440 245.600 75.840 ;
        RECT 4.000 72.440 246.000 74.440 ;
        RECT 4.400 71.040 245.600 72.440 ;
        RECT 4.000 69.040 246.000 71.040 ;
        RECT 4.400 67.640 245.600 69.040 ;
        RECT 4.000 65.640 246.000 67.640 ;
        RECT 4.400 64.240 245.600 65.640 ;
        RECT 4.000 62.240 246.000 64.240 ;
        RECT 4.400 60.840 245.600 62.240 ;
        RECT 4.000 58.840 246.000 60.840 ;
        RECT 4.400 57.440 245.600 58.840 ;
        RECT 4.000 55.440 246.000 57.440 ;
        RECT 4.400 54.040 245.600 55.440 ;
        RECT 4.000 52.040 246.000 54.040 ;
        RECT 4.400 50.640 245.600 52.040 ;
        RECT 4.000 48.640 246.000 50.640 ;
        RECT 4.400 47.240 245.600 48.640 ;
        RECT 4.000 45.240 246.000 47.240 ;
        RECT 4.400 43.840 245.600 45.240 ;
        RECT 4.000 41.840 246.000 43.840 ;
        RECT 4.400 40.440 245.600 41.840 ;
        RECT 4.000 38.440 246.000 40.440 ;
        RECT 4.400 37.040 245.600 38.440 ;
        RECT 4.000 35.040 246.000 37.040 ;
        RECT 4.400 33.640 245.600 35.040 ;
        RECT 4.000 31.640 246.000 33.640 ;
        RECT 4.400 30.240 245.600 31.640 ;
        RECT 4.000 28.240 246.000 30.240 ;
        RECT 4.400 26.840 245.600 28.240 ;
        RECT 4.000 24.840 246.000 26.840 ;
        RECT 4.400 23.440 245.600 24.840 ;
        RECT 4.000 21.440 246.000 23.440 ;
        RECT 4.400 20.040 245.600 21.440 ;
        RECT 4.000 18.040 246.000 20.040 ;
        RECT 4.400 16.640 245.600 18.040 ;
        RECT 4.000 14.640 246.000 16.640 ;
        RECT 4.400 13.240 245.600 14.640 ;
        RECT 4.000 11.240 246.000 13.240 ;
        RECT 4.400 9.840 245.600 11.240 ;
        RECT 4.000 7.840 246.000 9.840 ;
        RECT 4.400 6.440 245.600 7.840 ;
        RECT 4.000 4.440 246.000 6.440 ;
        RECT 4.400 3.040 245.600 4.440 ;
        RECT 4.000 1.040 246.000 3.040 ;
        RECT 4.400 0.175 245.600 1.040 ;
  END
END clk_rst_gen
END LIBRARY

