magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< metal2 >>
rect -4079 12127 -689 12502
rect -4079 11871 -3966 12127
rect -3710 11871 -3442 12127
rect -3186 11871 -2888 12127
rect -2632 11871 -2334 12127
rect -2078 11871 -1810 12127
rect -1554 11871 -689 12127
rect -4079 11633 -689 11871
rect -4079 11377 -3966 11633
rect -3710 11377 -3442 11633
rect -3186 11377 -2888 11633
rect -2632 11377 -2334 11633
rect -2078 11377 -1810 11633
rect -1554 11377 -689 11633
rect -4079 11002 -689 11377
tri -689 11002 811 12502 sw
tri -1311 9000 691 11002 ne
rect 691 10500 811 11002
tri 811 10500 1313 11002 sw
rect 691 10124 4024 10500
rect 691 9868 1511 10124
rect 1767 9868 2035 10124
rect 2291 9868 2589 10124
rect 2845 9868 3143 10124
rect 3399 9868 3667 10124
rect 3923 9868 4024 10124
rect 691 9630 4024 9868
rect 691 9374 1511 9630
rect 1767 9374 2035 9630
rect 2291 9374 2589 9630
rect 2845 9374 3143 9630
rect 3399 9374 3667 9630
rect 3923 9374 4024 9630
rect 691 9000 4024 9374
rect 6408 375 15500 750
rect 6408 119 6552 375
rect 6808 119 7076 375
rect 7332 119 7630 375
rect 7886 119 15500 375
rect 6408 -119 15500 119
rect 6408 -375 6552 -119
rect 6808 -375 7076 -119
rect 7332 -375 7630 -119
rect 7886 -375 15500 -119
rect 6408 -750 15500 -375
tri -1311 -13004 691 -11002 se
rect 691 -11377 3925 -11002
rect 691 -11633 1410 -11377
rect 1666 -11633 1934 -11377
rect 2190 -11633 2488 -11377
rect 2744 -11633 3042 -11377
rect 3298 -11633 3566 -11377
rect 3822 -11633 3925 -11377
rect 691 -11871 3925 -11633
rect 691 -12127 1410 -11871
rect 1666 -12127 1934 -11871
rect 2190 -12127 2488 -11871
rect 2744 -12127 3042 -11871
rect 3298 -12127 3566 -11871
rect 3822 -12127 3925 -11871
rect 691 -12502 3925 -12127
rect 691 -13004 811 -12502
tri 811 -13004 1313 -12502 nw
rect -4123 -13377 -689 -13004
rect -4123 -13633 -4024 -13377
rect -3768 -13633 -3500 -13377
rect -3244 -13633 -2946 -13377
rect -2690 -13633 -2392 -13377
rect -2136 -13633 -1868 -13377
rect -1612 -13633 -689 -13377
rect -4123 -13871 -689 -13633
rect -4123 -14127 -4024 -13871
rect -3768 -14127 -3500 -13871
rect -3244 -14127 -2946 -13871
rect -2690 -14127 -2392 -13871
rect -2136 -14127 -1868 -13871
rect -1612 -14127 -689 -13871
rect -4123 -14504 -689 -14127
tri -689 -14504 811 -13004 nw
<< via2 >>
rect -3966 11871 -3710 12127
rect -3442 11871 -3186 12127
rect -2888 11871 -2632 12127
rect -2334 11871 -2078 12127
rect -1810 11871 -1554 12127
rect -3966 11377 -3710 11633
rect -3442 11377 -3186 11633
rect -2888 11377 -2632 11633
rect -2334 11377 -2078 11633
rect -1810 11377 -1554 11633
rect 1511 9868 1767 10124
rect 2035 9868 2291 10124
rect 2589 9868 2845 10124
rect 3143 9868 3399 10124
rect 3667 9868 3923 10124
rect 1511 9374 1767 9630
rect 2035 9374 2291 9630
rect 2589 9374 2845 9630
rect 3143 9374 3399 9630
rect 3667 9374 3923 9630
rect 6552 119 6808 375
rect 7076 119 7332 375
rect 7630 119 7886 375
rect 6552 -375 6808 -119
rect 7076 -375 7332 -119
rect 7630 -375 7886 -119
rect 1410 -11633 1666 -11377
rect 1934 -11633 2190 -11377
rect 2488 -11633 2744 -11377
rect 3042 -11633 3298 -11377
rect 3566 -11633 3822 -11377
rect 1410 -12127 1666 -11871
rect 1934 -12127 2190 -11871
rect 2488 -12127 2744 -11871
rect 3042 -12127 3298 -11871
rect 3566 -12127 3822 -11871
rect -4024 -13633 -3768 -13377
rect -3500 -13633 -3244 -13377
rect -2946 -13633 -2690 -13377
rect -2392 -13633 -2136 -13377
rect -1868 -13633 -1612 -13377
rect -4024 -14127 -3768 -13871
rect -3500 -14127 -3244 -13871
rect -2946 -14127 -2690 -13871
rect -2392 -14127 -2136 -13871
rect -1868 -14127 -1612 -13871
<< metal3 >>
tri -7509 13004 -6009 14504 se
rect -6009 14497 6009 14504
tri 6009 14497 6016 14504 sw
rect -6009 13004 6016 14497
tri 6016 13004 7509 14497 sw
tri -8131 12382 -7509 13004 se
rect -7509 12502 -5889 13004
tri -5889 12502 -5387 13004 nw
tri 5387 12502 5889 13004 ne
rect 5889 12502 7509 13004
rect -7509 12382 -6009 12502
tri -6009 12382 -5889 12502 nw
tri -5300 12382 -5180 12502 se
rect -5180 12382 -1739 12502
tri -1739 12382 -1619 12502 sw
tri 569 12382 689 12502 se
rect 689 12382 5180 12502
tri -8138 12375 -8131 12382 se
rect -8131 12375 -6016 12382
tri -6016 12375 -6009 12382 nw
tri -5307 12375 -5300 12382 se
rect -5300 12375 -1619 12382
tri -1619 12375 -1612 12382 sw
tri 562 12375 569 12382 se
rect 569 12375 5180 12382
tri 5180 12375 5307 12502 sw
tri 5889 12375 6016 12502 ne
rect 6016 12375 7509 12502
tri 7509 12375 8138 13004 sw
tri -8386 12127 -8138 12375 se
rect -8138 12127 -6264 12375
tri -6264 12127 -6016 12375 nw
tri -5555 12127 -5307 12375 se
rect -5307 12228 -1612 12375
tri -1612 12228 -1465 12375 sw
tri 415 12228 562 12375 se
rect 562 12255 5307 12375
tri 5307 12255 5427 12375 sw
tri 6016 12255 6136 12375 ne
rect 6136 12255 8138 12375
rect 562 12228 5427 12255
rect -5307 12127 -1453 12228
tri -8642 11871 -8386 12127 se
rect -8386 11871 -6520 12127
tri -6520 11871 -6264 12127 nw
tri -5811 11871 -5555 12127 se
rect -5555 11871 -3966 12127
rect -3710 11871 -3442 12127
rect -3186 11871 -2888 12127
rect -2632 11871 -2334 12127
rect -2078 11871 -1810 12127
rect -1554 11871 -1453 12127
tri -8880 11633 -8642 11871 se
rect -8642 11666 -6725 11871
tri -6725 11666 -6520 11871 nw
tri -6016 11666 -5811 11871 se
rect -5811 11666 -1453 11871
rect -8642 11633 -6758 11666
tri -6758 11633 -6725 11666 nw
tri -6049 11633 -6016 11666 se
rect -6016 11633 -1453 11666
tri -9136 11377 -8880 11633 se
rect -8880 11377 -7014 11633
tri -7014 11377 -6758 11633 nw
tri -6305 11377 -6049 11633 se
rect -6049 11377 -3966 11633
rect -3710 11377 -3442 11633
rect -3186 11377 -2888 11633
rect -2632 11377 -2334 11633
rect -2078 11377 -1810 11633
rect -1554 11377 -1453 11633
tri -10133 10380 -9136 11377 se
rect -9136 11089 -7302 11377
tri -7302 11089 -7014 11377 nw
tri -6593 11089 -6305 11377 se
rect -6305 11276 -1453 11377
tri -537 11276 415 12228 se
rect 415 11546 5427 12228
tri 5427 11546 6136 12255 sw
tri 6136 11546 6845 12255 ne
rect 6845 11546 8138 12255
tri 8138 11546 8967 12375 sw
rect 415 11276 6136 11546
rect -6305 11089 -1739 11276
rect -9136 10380 -8011 11089
tri -8011 10380 -7302 11089 nw
tri -7182 10500 -6593 11089 se
rect -6593 11002 -1739 11089
tri -1739 11002 -1465 11276 nw
tri -811 11002 -537 11276 se
rect -537 11002 6136 11276
tri 6136 11002 6680 11546 sw
tri 6845 11002 7389 11546 ne
rect 7389 11002 8967 11546
rect -6593 10500 -5060 11002
tri -5060 10500 -4558 11002 nw
tri -1313 10500 -811 11002 se
rect -811 10500 809 11002
tri 809 10500 1311 11002 nw
tri 4558 10500 5060 11002 ne
rect 5060 10837 6680 11002
tri 6680 10837 6845 11002 sw
tri 7389 10837 7554 11002 ne
rect 7554 10837 8967 11002
rect 5060 10500 6845 10837
tri 6845 10500 7182 10837 sw
tri 7554 10500 7891 10837 ne
rect 7891 10500 8967 10837
tri -7302 10380 -7182 10500 se
rect -7182 10380 -5180 10500
tri -5180 10380 -5060 10500 nw
tri -4471 10380 -4351 10500 se
rect -4351 10380 569 10500
tri -10253 10260 -10133 10380 se
rect -10133 10260 -8131 10380
tri -8131 10260 -8011 10380 nw
tri -7422 10260 -7302 10380 se
rect -7302 10260 -5436 10380
tri -10260 10253 -10253 10260 se
rect -10253 10253 -8138 10260
tri -8138 10253 -8131 10260 nw
tri -7429 10253 -7422 10260 se
rect -7422 10253 -5436 10260
tri -10389 10124 -10260 10253 se
rect -10260 10124 -8267 10253
tri -8267 10124 -8138 10253 nw
tri -7558 10124 -7429 10253 se
rect -7429 10124 -5436 10253
tri -5436 10124 -5180 10380 nw
tri -4727 10124 -4471 10380 se
rect -4471 10260 569 10380
tri 569 10260 809 10500 nw
tri 1444 10260 1684 10500 se
rect 1684 10260 4351 10500
tri 4351 10260 4591 10500 sw
tri 5060 10260 5300 10500 ne
rect 5300 10260 7182 10500
tri 7182 10260 7422 10500 sw
tri 7891 10260 8131 10500 ne
rect 8131 10260 8967 10500
rect -4471 10253 562 10260
tri 562 10253 569 10260 nw
tri 1437 10253 1444 10260 se
rect 1444 10253 4591 10260
tri 4591 10253 4598 10260 sw
tri 5300 10253 5307 10260 ne
rect 5307 10253 7422 10260
tri 7422 10253 7429 10260 sw
tri 8131 10253 8138 10260 ne
rect 8138 10253 8967 10260
tri 8967 10253 10260 11546 sw
rect -4471 10124 433 10253
tri 433 10124 562 10253 nw
tri 1410 10226 1437 10253 se
rect 1437 10226 4598 10253
rect 1410 10124 4598 10226
tri -10645 9868 -10389 10124 se
rect -10389 9868 -8523 10124
tri -8523 9868 -8267 10124 nw
tri -7814 9868 -7558 10124 se
rect -7558 9868 -5692 10124
tri -5692 9868 -5436 10124 nw
tri -4983 9868 -4727 10124 se
rect -4727 9868 177 10124
tri 177 9868 433 10124 nw
rect 1410 9868 1511 10124
rect 1767 9868 2035 10124
rect 2291 9868 2589 10124
rect 2845 9868 3143 10124
rect 3399 9868 3667 10124
rect 3923 9868 4598 10124
tri -10883 9630 -10645 9868 se
rect -10645 9630 -8761 9868
tri -8761 9630 -8523 9868 nw
tri -8052 9630 -7814 9868 se
rect -7814 9671 -5889 9868
tri -5889 9671 -5692 9868 nw
tri -5180 9671 -4983 9868 se
rect -4983 9671 -61 9868
rect -7814 9630 -5930 9671
tri -5930 9630 -5889 9671 nw
tri -5221 9630 -5180 9671 se
rect -5180 9630 -61 9671
tri -61 9630 177 9868 nw
rect 1410 9630 4598 9868
tri -11139 9374 -10883 9630 se
rect -10883 9544 -8847 9630
tri -8847 9544 -8761 9630 nw
tri -8138 9544 -8052 9630 se
rect -8052 9544 -6186 9630
rect -10883 9374 -9017 9544
tri -9017 9374 -8847 9544 nw
tri -8308 9374 -8138 9544 se
rect -8138 9374 -6186 9544
tri -6186 9374 -5930 9630 nw
tri -5477 9374 -5221 9630 se
rect -5221 9374 -317 9630
tri -317 9374 -61 9630 nw
rect 1410 9374 1511 9630
rect 1767 9374 2035 9630
rect 2291 9374 2589 9630
rect 2845 9374 3143 9630
rect 3399 9374 3667 9630
rect 3923 9544 4598 9630
tri 4598 9544 5307 10253 sw
tri 5307 9544 6016 10253 ne
rect 6016 10133 7429 10253
tri 7429 10133 7549 10253 sw
tri 8138 10133 8258 10253 ne
rect 8258 10133 10260 10253
rect 6016 9544 7549 10133
rect 3923 9424 5307 9544
tri 5307 9424 5427 9544 sw
tri 6016 9424 6136 9544 ne
rect 6136 9424 7549 9544
tri 7549 9424 8258 10133 sw
tri 8258 9424 8967 10133 ne
rect 8967 9424 10260 10133
tri 10260 9424 11089 10253 sw
rect 3923 9374 5427 9424
tri -12255 8258 -11139 9374 se
rect -11139 8967 -9424 9374
tri -9424 8967 -9017 9374 nw
tri -8715 8967 -8308 9374 se
rect -8308 9087 -6473 9374
tri -6473 9087 -6186 9374 nw
tri -5764 9087 -5477 9374 se
rect -5477 9087 -691 9374
rect -8308 9000 -6560 9087
tri -6560 9000 -6473 9087 nw
tri -5851 9000 -5764 9087 se
rect -5764 9000 -691 9087
tri -691 9000 -317 9374 nw
rect 1410 9304 5427 9374
tri 5427 9304 5547 9424 sw
tri 6136 9304 6256 9424 ne
rect 6256 9304 8258 9424
rect 1410 9274 5547 9304
tri 1410 9000 1684 9274 ne
rect 1684 9000 5547 9274
tri 5547 9000 5851 9304 sw
tri 6256 9000 6560 9304 ne
rect 6560 9000 8258 9304
tri 8258 9000 8682 9424 sw
tri 8967 9000 9391 9424 ne
rect 9391 9000 11089 9424
rect -8308 8967 -7182 9000
rect -11139 8258 -10133 8967
tri -10133 8258 -9424 8967 nw
tri -9424 8258 -8715 8967 se
rect -8715 8378 -7182 8967
tri -7182 8378 -6560 9000 nw
tri -6256 8595 -5851 9000 se
rect -5851 8595 -4134 9000
tri -4134 8595 -3729 9000 nw
tri 3729 8595 4134 9000 ne
rect 4134 8595 5851 9000
tri 5851 8595 6256 9000 sw
tri 6560 8595 6965 9000 ne
rect 6965 8715 8682 9000
tri 8682 8715 8967 9000 sw
tri 9391 8715 9676 9000 ne
rect 9676 8715 11089 9000
rect 6965 8595 8967 8715
tri -6473 8378 -6256 8595 se
rect -6256 8378 -4351 8595
tri -4351 8378 -4134 8595 nw
tri 4134 8378 4351 8595 ne
rect 4351 8378 6256 8595
rect -8715 8258 -7302 8378
tri -7302 8258 -7182 8378 nw
tri -6593 8258 -6473 8378 se
rect -6473 8258 -4471 8378
tri -4471 8258 -4351 8378 nw
tri 4351 8258 4471 8378 ne
rect 4471 8258 6256 8378
tri 6256 8258 6593 8595 sw
tri 6965 8258 7302 8595 ne
rect 7302 8258 8967 8595
tri -12375 8138 -12255 8258 se
rect -12255 8138 -10253 8258
tri -10253 8138 -10133 8258 nw
tri -9544 8138 -9424 8258 se
rect -9424 8138 -7422 8258
tri -7422 8138 -7302 8258 nw
tri -6713 8138 -6593 8258 se
rect -6593 8138 -4591 8258
tri -4591 8138 -4471 8258 nw
tri 4471 8138 4591 8258 ne
rect 4591 8138 6593 8258
tri 6593 8138 6713 8258 sw
tri 7302 8138 7422 8258 ne
rect 7422 8138 8967 8258
tri 8967 8138 9544 8715 sw
tri 9676 8138 10253 8715 ne
rect 10253 8138 11089 8715
tri -12382 8131 -12375 8138 se
rect -12375 8131 -10260 8138
tri -10260 8131 -10253 8138 nw
tri -9551 8131 -9544 8138 se
rect -9544 8131 -7429 8138
tri -7429 8131 -7422 8138 nw
tri -6720 8131 -6713 8138 se
rect -6713 8131 -4598 8138
tri -4598 8131 -4591 8138 nw
tri 4591 8131 4598 8138 ne
rect 4598 8131 6713 8138
tri 6713 8131 6720 8138 sw
tri 7422 8131 7429 8138 ne
rect 7429 8131 9544 8138
tri 9544 8131 9551 8138 sw
tri 10253 8131 10260 8138 ne
rect 10260 8131 11089 8138
tri 11089 8131 12382 9424 sw
tri -14377 6136 -12382 8131 se
rect -12382 7422 -10969 8131
tri -10969 7422 -10260 8131 nw
tri -10260 7422 -9551 8131 se
rect -9551 7422 -8138 8131
tri -8138 7422 -7429 8131 nw
tri -7429 7422 -6720 8131 se
rect -6720 7422 -5427 8131
rect -12382 6845 -11546 7422
tri -11546 6845 -10969 7422 nw
tri -10837 6845 -10260 7422 se
rect -10260 7302 -8258 7422
tri -8258 7302 -8138 7422 nw
tri -7549 7302 -7429 7422 se
rect -7429 7302 -5427 7422
tri -5427 7302 -4598 8131 nw
tri 4598 7302 5427 8131 ne
rect 5427 7422 6720 8131
tri 6720 7422 7429 8131 sw
tri 7429 7422 8138 8131 ne
rect 8138 8011 9551 8131
tri 9551 8011 9671 8131 sw
tri 10260 8011 10380 8131 ne
rect 10380 8011 12382 8131
rect 8138 7422 9671 8011
rect 5427 7302 7429 7422
tri 7429 7302 7549 7422 sw
tri 8138 7302 8258 7422 ne
rect 8258 7302 9671 7422
tri 9671 7302 10380 8011 sw
tri 10380 7302 11089 8011 ne
rect 11089 7302 12382 8011
tri 12382 7302 13211 8131 sw
rect -10260 6965 -8595 7302
tri -8595 6965 -8258 7302 nw
tri -7886 6965 -7549 7302 se
rect -7549 6965 -6256 7302
rect -10260 6845 -9304 6965
rect -12382 6136 -12255 6845
tri -12255 6136 -11546 6845 nw
tri -11546 6136 -10837 6845 se
rect -10837 6256 -9304 6845
tri -9304 6256 -8595 6965 nw
tri -8378 6473 -7886 6965 se
rect -7886 6473 -6256 6965
tri -6256 6473 -5427 7302 nw
tri 5427 6473 6256 7302 ne
rect 6256 7182 7549 7302
tri 7549 7182 7669 7302 sw
tri 8258 7182 8378 7302 ne
rect 8378 7182 10380 7302
rect 6256 6473 7669 7182
tri 7669 6473 8378 7182 sw
tri 8378 6473 9087 7182 ne
rect 9087 6593 10380 7182
tri 10380 6593 11089 7302 sw
tri 11089 6593 11798 7302 ne
rect 11798 6593 13211 7302
rect 9087 6473 11089 6593
tri -8595 6256 -8378 6473 se
rect -8378 6256 -6473 6473
tri -6473 6256 -6256 6473 nw
tri 6256 6256 6473 6473 ne
rect 6473 6256 8378 6473
rect -10837 6136 -9424 6256
tri -9424 6136 -9304 6256 nw
tri -8715 6136 -8595 6256 se
rect -8595 6136 -6593 6256
tri -6593 6136 -6473 6256 nw
tri 6473 6136 6593 6256 ne
rect 6593 6136 8378 6256
tri 8378 6136 8715 6473 sw
tri 9087 6136 9424 6473 ne
rect 9424 6136 11089 6473
tri -14497 6016 -14377 6136 se
rect -14377 6016 -12375 6136
tri -12375 6016 -12255 6136 nw
tri -11666 6016 -11546 6136 se
rect -11546 6016 -9544 6136
tri -9544 6016 -9424 6136 nw
tri -8835 6016 -8715 6136 se
rect -8715 6016 -6713 6136
tri -6713 6016 -6593 6136 nw
tri 6593 6016 6713 6136 ne
rect 6713 6016 8715 6136
tri 8715 6016 8835 6136 sw
tri 9424 6016 9544 6136 ne
rect 9544 6016 11089 6136
tri 11089 6016 11666 6593 sw
tri 11798 6016 12375 6593 ne
rect 12375 6016 13211 6593
tri -14504 6009 -14497 6016 se
rect -14497 6009 -12382 6016
tri -12382 6009 -12375 6016 nw
tri -11673 6009 -11666 6016 se
rect -11666 6009 -9551 6016
tri -9551 6009 -9544 6016 nw
tri -8842 6009 -8835 6016 se
rect -8835 6009 -6720 6016
tri -6720 6009 -6713 6016 nw
tri 6713 6009 6720 6016 ne
rect 6720 6009 8835 6016
tri 8835 6009 8842 6016 sw
tri 9544 6009 9551 6016 ne
rect 9551 6009 11666 6016
tri 11666 6009 11673 6016 sw
tri 12375 6009 12382 6016 ne
rect 12382 6009 13211 6016
tri 13211 6009 14504 7302 sw
rect -14504 5889 -12502 6009
tri -12502 5889 -12382 6009 nw
tri -11793 5889 -11673 6009 se
rect -11673 5889 -10173 6009
rect -14504 -5889 -13004 5889
tri -13004 5387 -12502 5889 nw
tri -12295 5387 -11793 5889 se
rect -11793 5387 -10173 5889
tri -10173 5387 -9551 6009 nw
tri -9464 5387 -8842 6009 se
rect -8842 5387 -7342 6009
tri -7342 5387 -6720 6009 nw
tri 6720 5387 7342 6009 ne
rect 7342 5387 8842 6009
tri 8842 5387 9464 6009 sw
tri 9551 5387 10173 6009 ne
rect 10173 5889 11673 6009
tri 11673 5889 11793 6009 sw
tri 12382 5889 12502 6009 ne
rect 12502 5889 14504 6009
rect 10173 5387 11793 5889
tri 11793 5387 12295 5889 sw
tri 12502 5387 13004 5889 ne
tri -12502 5180 -12295 5387 se
rect -12295 5180 -10380 5387
tri -10380 5180 -10173 5387 nw
tri -9671 5180 -9464 5387 se
rect -9464 5180 -7549 5387
tri -7549 5180 -7342 5387 nw
tri 7342 5180 7549 5387 ne
rect 7549 5180 9464 5387
tri 9464 5180 9671 5387 sw
tri 10173 5180 10380 5387 ne
rect 10380 5180 12295 5387
tri 12295 5180 12502 5387 sw
rect -12502 5060 -10500 5180
tri -10500 5060 -10380 5180 nw
tri -9791 5060 -9671 5180 se
rect -9671 5060 -8171 5180
rect -12502 -5060 -11002 5060
tri -11002 4558 -10500 5060 nw
tri -10293 4558 -9791 5060 se
rect -9791 4558 -8171 5060
tri -8171 4558 -7549 5180 nw
tri 7549 4558 8171 5180 ne
rect 8171 5060 9671 5180
tri 9671 5060 9791 5180 sw
tri 10380 5060 10500 5180 ne
rect 10500 5060 12502 5180
rect 8171 4558 9791 5060
tri 9791 4558 10293 5060 sw
tri 10500 4558 11002 5060 ne
tri -10500 4351 -10293 4558 se
rect -10293 4351 -8378 4558
tri -8378 4351 -8171 4558 nw
tri 8171 4351 8378 4558 ne
rect 8378 4351 10293 4558
tri 10293 4351 10500 4558 sw
rect -10500 750 -9000 4351
tri -9000 3729 -8378 4351 nw
tri 8378 3729 9000 4351 ne
rect -10500 375 8000 750
rect -10500 119 6552 375
rect 6808 119 7076 375
rect 7332 119 7630 375
rect 7886 119 8000 375
rect -10500 -119 8000 119
rect -10500 -375 6552 -119
rect 6808 -375 7076 -119
rect 7332 -375 7630 -119
rect 7886 -375 8000 -119
rect -10500 -750 8000 -375
rect -10500 -4351 -9000 -750
tri -9000 -4351 -8378 -3729 sw
tri 8378 -4351 9000 -3729 se
rect 9000 -4351 10500 4351
tri -10500 -4558 -10293 -4351 ne
rect -10293 -4558 -8378 -4351
tri -8378 -4558 -8171 -4351 sw
tri 8171 -4558 8378 -4351 se
rect 8378 -4558 10293 -4351
tri 10293 -4558 10500 -4351 nw
tri -11002 -5060 -10500 -4558 sw
tri -10293 -5060 -9791 -4558 ne
rect -9791 -5060 -8171 -4558
rect -12502 -5180 -10500 -5060
tri -10500 -5180 -10380 -5060 sw
tri -9791 -5180 -9671 -5060 ne
rect -9671 -5180 -8171 -5060
tri -8171 -5180 -7549 -4558 sw
tri 7549 -5180 8171 -4558 se
rect 8171 -5060 9791 -4558
tri 9791 -5060 10293 -4558 nw
tri 10500 -5060 11002 -4558 se
rect 11002 -5060 12502 5060
rect 13004 3250 14504 5889
rect 13004 1750 15500 3250
rect 8171 -5180 9671 -5060
tri 9671 -5180 9791 -5060 nw
tri 10380 -5180 10500 -5060 se
rect 10500 -5180 12502 -5060
tri -12502 -5387 -12295 -5180 ne
rect -12295 -5387 -10380 -5180
tri -10380 -5387 -10173 -5180 sw
tri -9671 -5387 -9464 -5180 ne
rect -9464 -5387 -7549 -5180
tri -7549 -5387 -7342 -5180 sw
tri 7342 -5387 7549 -5180 se
rect 7549 -5387 9464 -5180
tri 9464 -5387 9671 -5180 nw
tri 10173 -5387 10380 -5180 se
rect 10380 -5387 12295 -5180
tri 12295 -5387 12502 -5180 nw
rect 13004 -3250 15500 -1750
tri -13004 -5889 -12502 -5387 sw
tri -12295 -5889 -11793 -5387 ne
rect -11793 -5889 -10173 -5387
rect -14504 -6009 -12502 -5889
tri -12502 -6009 -12382 -5889 sw
tri -11793 -6009 -11673 -5889 ne
rect -11673 -6009 -10173 -5889
tri -10173 -6009 -9551 -5387 sw
tri -9464 -6009 -8842 -5387 ne
rect -8842 -6009 -7342 -5387
tri -7342 -6009 -6720 -5387 sw
tri 6720 -6009 7342 -5387 se
rect 7342 -6009 8842 -5387
tri 8842 -6009 9464 -5387 nw
tri 9551 -6009 10173 -5387 se
rect 10173 -5889 11793 -5387
tri 11793 -5889 12295 -5387 nw
tri 12502 -5889 13004 -5387 se
rect 13004 -5889 14504 -3250
rect 10173 -6009 11673 -5889
tri 11673 -6009 11793 -5889 nw
tri 12382 -6009 12502 -5889 se
rect 12502 -6009 14504 -5889
tri -14504 -6016 -14497 -6009 ne
rect -14497 -6016 -12382 -6009
tri -12382 -6016 -12375 -6009 sw
tri -11673 -6016 -11666 -6009 ne
rect -11666 -6016 -9551 -6009
tri -9551 -6016 -9544 -6009 sw
tri -8842 -6016 -8835 -6009 ne
rect -8835 -6016 -6720 -6009
tri -6720 -6016 -6713 -6009 sw
tri 6713 -6016 6720 -6009 se
rect 6720 -6016 8835 -6009
tri 8835 -6016 8842 -6009 nw
tri 9544 -6016 9551 -6009 se
rect 9551 -6016 11666 -6009
tri 11666 -6016 11673 -6009 nw
tri 12375 -6016 12382 -6009 se
rect 12382 -6016 14497 -6009
tri 14497 -6016 14504 -6009 nw
tri -14497 -7302 -13211 -6016 ne
rect -13211 -6593 -12375 -6016
tri -12375 -6593 -11798 -6016 sw
tri -11666 -6593 -11089 -6016 ne
rect -11089 -6136 -9544 -6016
tri -9544 -6136 -9424 -6016 sw
tri -8835 -6136 -8715 -6016 ne
rect -8715 -6136 -6713 -6016
tri -6713 -6136 -6593 -6016 sw
tri 6593 -6136 6713 -6016 se
rect 6713 -6136 8715 -6016
tri 8715 -6136 8835 -6016 nw
tri 9424 -6136 9544 -6016 se
rect 9544 -6136 11546 -6016
tri 11546 -6136 11666 -6016 nw
tri 12255 -6136 12375 -6016 se
rect 12375 -6136 14377 -6016
tri 14377 -6136 14497 -6016 nw
rect -11089 -6473 -9424 -6136
tri -9424 -6473 -9087 -6136 sw
tri -8715 -6256 -8595 -6136 ne
rect -8595 -6256 -6593 -6136
tri -6593 -6256 -6473 -6136 sw
tri 6473 -6256 6593 -6136 se
rect 6593 -6256 8595 -6136
tri 8595 -6256 8715 -6136 nw
tri 9304 -6256 9424 -6136 se
rect 9424 -6256 10837 -6136
tri -8595 -6473 -8378 -6256 ne
rect -8378 -6473 -6473 -6256
tri -6473 -6473 -6256 -6256 sw
tri 6256 -6473 6473 -6256 se
rect 6473 -6473 7886 -6256
rect -11089 -6593 -9087 -6473
rect -13211 -7302 -11798 -6593
tri -11798 -7302 -11089 -6593 sw
tri -11089 -7302 -10380 -6593 ne
rect -10380 -7182 -9087 -6593
tri -9087 -7182 -8378 -6473 sw
tri -8378 -7182 -7669 -6473 ne
rect -7669 -7182 -6256 -6473
rect -10380 -7302 -8378 -7182
tri -8378 -7302 -8258 -7182 sw
tri -7669 -7302 -7549 -7182 ne
rect -7549 -7302 -6256 -7182
tri -6256 -7302 -5427 -6473 sw
tri 5427 -7302 6256 -6473 se
rect 6256 -6965 7886 -6473
tri 7886 -6965 8595 -6256 nw
tri 8595 -6965 9304 -6256 se
rect 9304 -6845 10837 -6256
tri 10837 -6845 11546 -6136 nw
tri 11546 -6845 12255 -6136 se
rect 12255 -6845 12375 -6136
rect 9304 -6965 10253 -6845
rect 6256 -7302 7549 -6965
tri 7549 -7302 7886 -6965 nw
tri 8258 -7302 8595 -6965 se
rect 8595 -7302 10253 -6965
tri -13211 -8131 -12382 -7302 ne
rect -12382 -8011 -11089 -7302
tri -11089 -8011 -10380 -7302 sw
tri -10380 -8011 -9671 -7302 ne
rect -9671 -7422 -8258 -7302
tri -8258 -7422 -8138 -7302 sw
tri -7549 -7422 -7429 -7302 ne
rect -7429 -7422 -5427 -7302
rect -9671 -8011 -8138 -7422
rect -12382 -8131 -10380 -8011
tri -10380 -8131 -10260 -8011 sw
tri -9671 -8131 -9551 -8011 ne
rect -9551 -8131 -8138 -8011
tri -8138 -8131 -7429 -7422 sw
tri -7429 -8131 -6720 -7422 ne
rect -6720 -8131 -5427 -7422
tri -5427 -8131 -4598 -7302 sw
tri 4598 -8131 5427 -7302 se
rect 5427 -7422 7429 -7302
tri 7429 -7422 7549 -7302 nw
tri 8138 -7422 8258 -7302 se
rect 8258 -7422 10253 -7302
rect 5427 -8131 6720 -7422
tri 6720 -8131 7429 -7422 nw
tri 7429 -8131 8138 -7422 se
rect 8138 -7429 10253 -7422
tri 10253 -7429 10837 -6845 nw
tri 10962 -7429 11546 -6845 se
rect 11546 -7429 12375 -6845
rect 8138 -8131 9551 -7429
tri 9551 -8131 10253 -7429 nw
tri 10260 -8131 10962 -7429 se
rect 10962 -8131 12375 -7429
tri -12382 -8138 -12375 -8131 ne
rect -12375 -8138 -10260 -8131
tri -10260 -8138 -10253 -8131 sw
tri -9551 -8138 -9544 -8131 ne
rect -9544 -8138 -7429 -8131
tri -7429 -8138 -7422 -8131 sw
tri -6720 -8138 -6713 -8131 ne
rect -6713 -8138 -4598 -8131
tri -4598 -8138 -4591 -8131 sw
tri 4591 -8138 4598 -8131 se
rect 4598 -8138 6713 -8131
tri 6713 -8138 6720 -8131 nw
tri 7422 -8138 7429 -8131 se
rect 7429 -8138 9544 -8131
tri 9544 -8138 9551 -8131 nw
tri 10253 -8138 10260 -8131 se
rect 10260 -8138 12375 -8131
tri 12375 -8138 14377 -6136 nw
tri -12375 -9424 -11089 -8138 ne
rect -11089 -8715 -10253 -8138
tri -10253 -8715 -9676 -8138 sw
tri -9544 -8715 -8967 -8138 ne
rect -8967 -8258 -7422 -8138
tri -7422 -8258 -7302 -8138 sw
tri -6713 -8258 -6593 -8138 ne
rect -6593 -8258 -4591 -8138
tri -4591 -8258 -4471 -8138 sw
tri 4471 -8258 4591 -8138 se
rect 4591 -8258 6593 -8138
tri 6593 -8258 6713 -8138 nw
tri 7302 -8258 7422 -8138 se
rect 7422 -8258 9424 -8138
tri 9424 -8258 9544 -8138 nw
tri 10133 -8258 10253 -8138 se
rect 10253 -8258 12255 -8138
tri 12255 -8258 12375 -8138 nw
rect -8967 -8595 -7302 -8258
tri -7302 -8595 -6965 -8258 sw
tri -6593 -8378 -6473 -8258 ne
rect -6473 -8378 -4471 -8258
tri -4471 -8378 -4351 -8258 sw
tri 4351 -8378 4471 -8258 se
rect 4471 -8378 6473 -8258
tri 6473 -8378 6593 -8258 nw
tri 7182 -8378 7302 -8258 se
rect 7302 -8378 8715 -8258
tri -6473 -8595 -6256 -8378 ne
rect -6256 -8595 -4351 -8378
tri -4351 -8595 -4134 -8378 sw
tri 4134 -8595 4351 -8378 se
rect 4351 -8595 5764 -8378
rect -8967 -8715 -6965 -8595
rect -11089 -9424 -9676 -8715
tri -9676 -9424 -8967 -8715 sw
tri -8967 -9424 -8258 -8715 ne
rect -8258 -9304 -6965 -8715
tri -6965 -9304 -6256 -8595 sw
tri -6256 -9304 -5547 -8595 ne
rect -5547 -9000 -4134 -8595
tri -4134 -9000 -3729 -8595 sw
tri 3729 -9000 4134 -8595 se
rect 4134 -9000 5764 -8595
rect -5547 -9087 5764 -9000
tri 5764 -9087 6473 -8378 nw
tri 6473 -9087 7182 -8378 se
rect 7182 -8967 8715 -8378
tri 8715 -8967 9424 -8258 nw
tri 9424 -8967 10133 -8258 se
rect 10133 -8967 10253 -8258
rect 7182 -9087 8131 -8967
rect -5547 -9304 5427 -9087
rect -8258 -9424 -6256 -9304
tri -6256 -9424 -6136 -9304 sw
tri -5547 -9424 -5427 -9304 ne
rect -5427 -9424 5427 -9304
tri 5427 -9424 5764 -9087 nw
tri 6136 -9424 6473 -9087 se
rect 6473 -9424 8131 -9087
tri -11089 -10253 -10260 -9424 ne
rect -10260 -10133 -8967 -9424
tri -8967 -10133 -8258 -9424 sw
tri -8258 -10133 -7549 -9424 ne
rect -7549 -9544 -6136 -9424
tri -6136 -9544 -6016 -9424 sw
tri -5427 -9544 -5307 -9424 ne
rect -5307 -9544 5307 -9424
tri 5307 -9544 5427 -9424 nw
tri 6016 -9544 6136 -9424 se
rect 6136 -9544 8131 -9424
rect -7549 -10133 -6016 -9544
rect -10260 -10253 -8258 -10133
tri -8258 -10253 -8138 -10133 sw
tri -7549 -10253 -7429 -10133 ne
rect -7429 -10253 -6016 -10133
tri -6016 -10253 -5307 -9544 sw
tri -5307 -10253 -4598 -9544 ne
rect -4598 -10253 4598 -9544
tri 4598 -10253 5307 -9544 nw
tri 5307 -10253 6016 -9544 se
rect 6016 -9551 8131 -9544
tri 8131 -9551 8715 -8967 nw
tri 8840 -9551 9424 -8967 se
rect 9424 -9551 10253 -8967
rect 6016 -10253 7429 -9551
tri 7429 -10253 8131 -9551 nw
tri 8138 -10253 8840 -9551 se
rect 8840 -10253 10253 -9551
tri -10260 -10260 -10253 -10253 ne
rect -10253 -10260 -8138 -10253
tri -8138 -10260 -8131 -10253 sw
tri -7429 -10260 -7422 -10253 ne
rect -7422 -10260 -5307 -10253
tri -5307 -10260 -5300 -10253 sw
tri -4598 -10260 -4591 -10253 ne
rect -4591 -10260 4591 -10253
tri 4591 -10260 4598 -10253 nw
tri 5300 -10260 5307 -10253 se
rect 5307 -10260 7422 -10253
tri 7422 -10260 7429 -10253 nw
tri 8131 -10260 8138 -10253 se
rect 8138 -10260 10253 -10253
tri 10253 -10260 12255 -8258 nw
tri -10253 -11004 -9509 -10260 ne
rect -9509 -10295 -8131 -10260
tri -8131 -10295 -8096 -10260 sw
tri -7422 -10295 -7387 -10260 ne
rect -7387 -10295 -5300 -10260
rect -9509 -11004 -8096 -10295
tri -8096 -11004 -7387 -10295 sw
tri -7387 -10380 -7302 -10295 ne
rect -7302 -10380 -5300 -10295
tri -5300 -10380 -5180 -10260 sw
tri -4591 -10380 -4471 -10260 ne
rect -4471 -10380 4471 -10260
tri 4471 -10380 4591 -10260 nw
tri 5180 -10380 5300 -10260 se
rect 5300 -10380 7302 -10260
tri 7302 -10380 7422 -10260 nw
tri 8011 -10380 8131 -10260 se
rect 8131 -10380 9509 -10260
tri -7302 -11004 -6678 -10380 ne
rect -6678 -10500 -5180 -10380
tri -5180 -10500 -5060 -10380 sw
tri -4471 -10500 -4351 -10380 ne
rect -4351 -10500 4351 -10380
tri 4351 -10500 4471 -10380 nw
tri 5060 -10500 5180 -10380 se
rect 5180 -10500 6678 -10380
rect -6678 -11004 -5060 -10500
tri -5060 -11004 -4556 -10500 sw
tri 4558 -11002 5060 -10500 se
rect 5060 -11002 6678 -10500
tri 1583 -11004 1585 -11002 se
rect 1585 -11004 6678 -11002
tri 6678 -11004 7302 -10380 nw
tri 7387 -11004 8011 -10380 se
rect 8011 -11004 9509 -10380
tri 9509 -11004 10253 -10260 nw
tri -9509 -11377 -9136 -11004 ne
rect -9136 -11377 -7387 -11004
tri -7387 -11377 -7014 -11004 sw
tri -6678 -11377 -6305 -11004 ne
rect -6305 -11377 -689 -11004
tri -689 -11377 -316 -11004 sw
tri 1311 -11276 1583 -11004 se
rect 1583 -11089 6593 -11004
tri 6593 -11089 6678 -11004 nw
tri 7302 -11089 7387 -11004 se
rect 7387 -11089 8131 -11004
rect 1583 -11276 6009 -11089
rect 1311 -11377 6009 -11276
tri -9136 -11546 -8967 -11377 ne
rect -8967 -11546 -7014 -11377
tri -7014 -11546 -6845 -11377 sw
tri -6305 -11546 -6136 -11377 ne
rect -6136 -11546 -316 -11377
tri -8967 -11633 -8880 -11546 ne
rect -8880 -11633 -6845 -11546
tri -6845 -11633 -6758 -11546 sw
tri -6136 -11633 -6049 -11546 ne
rect -6049 -11633 -316 -11546
tri -316 -11633 -60 -11377 sw
rect 1311 -11633 1410 -11377
rect 1666 -11633 1934 -11377
rect 2190 -11633 2488 -11377
rect 2744 -11633 3042 -11377
rect 3298 -11633 3566 -11377
rect 3822 -11633 6009 -11377
tri -8880 -11871 -8642 -11633 ne
rect -8642 -11871 -6758 -11633
tri -6758 -11871 -6520 -11633 sw
tri -6049 -11871 -5811 -11633 ne
rect -5811 -11871 -60 -11633
tri -60 -11871 178 -11633 sw
rect 1311 -11673 6009 -11633
tri 6009 -11673 6593 -11089 nw
tri 6718 -11673 7302 -11089 se
rect 7302 -11673 8131 -11089
rect 1311 -11871 5300 -11673
tri -8642 -12127 -8386 -11871 ne
rect -8386 -12127 -6520 -11871
tri -6520 -12127 -6264 -11871 sw
tri -5811 -12127 -5555 -11871 ne
rect -5555 -12127 178 -11871
tri 178 -12127 434 -11871 sw
rect 1311 -12127 1410 -11871
rect 1666 -12127 1934 -11871
rect 2190 -12127 2488 -11871
rect 2744 -12127 3042 -11871
rect 3298 -12127 3566 -11871
rect 3822 -12127 5300 -11871
tri -8386 -12375 -8138 -12127 ne
rect -8138 -12255 -6264 -12127
tri -6264 -12255 -6136 -12127 sw
tri -5555 -12255 -5427 -12127 ne
rect -5427 -12255 434 -12127
rect -8138 -12375 -6136 -12255
tri -6136 -12375 -6016 -12255 sw
tri -5427 -12375 -5307 -12255 ne
rect -5307 -12375 434 -12255
tri -8138 -12502 -8011 -12375 ne
rect -8011 -12502 -6016 -12375
tri -6016 -12502 -5889 -12375 sw
tri -5307 -12502 -5180 -12375 ne
rect -5180 -12502 434 -12375
tri 434 -12502 809 -12127 sw
rect 1311 -12228 5300 -12127
tri 1311 -12502 1585 -12228 ne
rect 1585 -12382 5300 -12228
tri 5300 -12382 6009 -11673 nw
tri 6009 -12382 6718 -11673 se
rect 6718 -12382 8131 -11673
tri 8131 -12382 9509 -11004 nw
rect 1585 -12502 5180 -12382
tri 5180 -12502 5300 -12382 nw
tri 5889 -12502 6009 -12382 se
rect 6009 -12502 8011 -12382
tri 8011 -12502 8131 -12382 nw
tri -8011 -13377 -7136 -12502 ne
rect -7136 -13004 -5889 -12502
tri -5889 -13004 -5387 -12502 sw
tri -1313 -13004 -811 -12502 ne
rect -811 -13004 809 -12502
tri 809 -13004 1311 -12502 sw
tri 5387 -13004 5889 -12502 se
rect 5889 -13004 7509 -12502
tri 7509 -13004 8011 -12502 nw
rect -7136 -13278 -1783 -13004
tri -1783 -13278 -1509 -13004 sw
rect -7136 -13377 -1509 -13278
tri -7136 -13633 -6880 -13377 ne
rect -6880 -13633 -4024 -13377
rect -3768 -13633 -3500 -13377
rect -3244 -13633 -2946 -13377
rect -2690 -13633 -2392 -13377
rect -2136 -13633 -1868 -13377
rect -1612 -13633 -1509 -13377
tri -6880 -13871 -6642 -13633 ne
rect -6642 -13871 -1509 -13633
tri -6642 -14127 -6386 -13871 ne
rect -6386 -14127 -4024 -13871
rect -3768 -14127 -3500 -13871
rect -3244 -14127 -2946 -13871
rect -2690 -14127 -2392 -13871
rect -2136 -14127 -1868 -13871
rect -1612 -14127 -1509 -13871
tri -6386 -14497 -6016 -14127 ne
rect -6016 -14230 -1509 -14127
rect -6016 -14497 -1776 -14230
tri -1776 -14497 -1509 -14230 nw
tri -811 -14497 682 -13004 ne
rect 682 -14497 6009 -13004
tri -6016 -14504 -6009 -14497 ne
rect -6009 -14504 -1783 -14497
tri -1783 -14504 -1776 -14497 nw
tri 682 -14504 689 -14497 ne
rect 689 -14504 6009 -14497
tri 6009 -14504 7509 -13004 nw
<< comment >>
tri -6009 6009 -2489 14504 ne
rect -2489 6009 2489 14504
tri 2489 6009 6009 14504 nw
tri -14504 2489 -6009 6009 sw
tri -2489 2489 -1031 6009 ne
rect -1031 2489 1031 6009
tri 1031 2490 2489 6009 nw
tri 6009 2490 14504 6009 se
rect -14504 427 -6009 2489
tri -6009 427 -1031 2489 sw
tri -1031 428 -177 2489 ne
rect -177 427 177 2489
tri 177 427 1031 2489 nw
tri 1031 427 6009 2489 se
rect 6009 427 14504 2490
rect -14504 73 -1031 427
tri -1031 73 -177 427 sw
tri -177 74 -31 427 ne
rect -31 73 30 427
tri 30 73 177 427 nw
tri 177 73 1031 427 se
rect 1031 73 14504 427
rect -14504 13 -177 73
tri -177 13 -31 73 sw
tri -31 13 -5 73 ne
rect -5 13 5 73
tri 5 13 30 73 nw
tri 30 13 177 73 se
rect 177 13 14504 73
rect -14504 2 -31 13
tri -31 2 -5 13 sw
tri -5 2 -1 13 ne
rect -1 2 1 13
tri 1 2 5 13 nw
tri 6 2 30 13 se
rect 30 2 14504 13
rect -14504 -2 -5 2
tri -5 0 -1 2 sw
tri -1 0 0 2 ne
tri 0 0 1 2 nw
tri 1 0 5 2 se
tri -5 -2 -1 0 nw
tri -1 -2 0 0 se
tri 0 -2 1 0 sw
tri 1 -2 5 0 ne
rect 5 -2 14504 2
rect -14504 -13 -30 -2
tri -30 -13 -5 -2 nw
tri -5 -13 -1 -2 se
rect -1 -12 1 -2
tri 1 -12 5 -2 sw
tri 5 -12 30 -2 ne
rect 30 -12 14504 -2
rect -1 -13 5 -12
rect -14504 -73 -177 -13
tri -177 -73 -30 -13 nw
tri -30 -73 -5 -13 se
rect -5 -73 5 -13
tri 5 -73 30 -12 sw
tri 30 -73 176 -12 ne
rect 176 -73 14504 -12
rect -14504 -427 -1031 -73
tri -1031 -427 -177 -73 nw
tri -177 -427 -30 -73 se
rect -30 -427 30 -73
tri 30 -427 177 -73 sw
tri 177 -427 1030 -73 ne
rect 1030 -427 14504 -73
rect -14504 -2489 -6009 -427
tri -6009 -2489 -1031 -427 nw
tri -1031 -2489 -177 -427 se
rect -177 -2489 177 -427
tri 177 -2489 1031 -427 sw
tri 1031 -2489 6008 -427 ne
rect 6008 -2489 14504 -427
tri -14504 -6009 -6009 -2489 nw
tri -2489 -6009 -1031 -2490 se
rect -1031 -6009 1031 -2489
tri 1031 -6009 2489 -2489 sw
tri 6009 -6009 14504 -2489 ne
tri -6009 -14504 -2489 -6009 se
rect -2489 -14504 2489 -6009
tri 2489 -14504 6009 -6009 sw
<< properties >>
string GDS_END 10489546
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10482838
string gencell sky130_fd_pr__rf_test_coil1
string library sky130
string parameter m=1
string path 343.850 -150.225 343.850 -43.750 
<< end >>
