magic
tech sky130B
magscale 12 1
timestamp 1598777186
<< metal5 >>
rect 10 70 35 75
rect 5 65 40 70
rect 0 55 45 65
rect 0 20 15 55
rect 30 20 45 55
rect 0 10 45 20
rect 5 5 45 10
rect 10 0 45 5
rect 30 -30 45 0
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
