magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 49 67 600 203
rect 49 21 503 67
rect 49 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 131 47 161 177
rect 215 47 245 177
rect 311 47 341 177
rect 395 47 425 177
rect 492 93 522 177
<< scpmoshvt >>
rect 131 297 161 497
rect 215 297 245 497
rect 311 297 341 497
rect 395 297 425 497
rect 492 336 522 420
<< ndiff >>
rect 75 89 131 177
rect 75 55 87 89
rect 121 55 131 89
rect 75 47 131 55
rect 161 116 215 177
rect 161 82 171 116
rect 205 82 215 116
rect 161 47 215 82
rect 245 95 311 177
rect 245 61 261 95
rect 295 61 311 95
rect 245 47 311 61
rect 341 116 395 177
rect 341 82 351 116
rect 385 82 395 116
rect 341 47 395 82
rect 425 163 492 177
rect 425 129 435 163
rect 469 129 492 163
rect 425 95 492 129
rect 425 61 435 95
rect 469 93 492 95
rect 522 149 574 177
rect 522 115 532 149
rect 566 115 574 149
rect 522 93 574 115
rect 469 61 477 93
rect 425 47 477 61
<< pdiff >>
rect 27 474 131 497
rect 27 440 35 474
rect 69 440 131 474
rect 27 406 131 440
rect 27 372 35 406
rect 69 372 131 406
rect 27 297 131 372
rect 161 297 215 497
rect 245 297 311 497
rect 341 297 395 497
rect 425 471 477 497
rect 425 437 435 471
rect 469 437 477 471
rect 425 420 477 437
rect 425 336 492 420
rect 522 397 574 420
rect 522 363 532 397
rect 566 363 574 397
rect 522 336 574 363
rect 425 297 477 336
<< ndiffc >>
rect 87 55 121 89
rect 171 82 205 116
rect 261 61 295 95
rect 351 82 385 116
rect 435 129 469 163
rect 435 61 469 95
rect 532 115 566 149
<< pdiffc >>
rect 35 440 69 474
rect 35 372 69 406
rect 435 437 469 471
rect 532 363 566 397
<< poly >>
rect 131 497 161 523
rect 215 497 245 523
rect 311 497 341 523
rect 395 497 425 523
rect 492 420 522 446
rect 131 265 161 297
rect 215 265 245 297
rect 311 265 341 297
rect 395 265 425 297
rect 492 265 522 336
rect 91 249 161 265
rect 91 215 107 249
rect 141 215 161 249
rect 91 199 161 215
rect 203 249 257 265
rect 203 215 213 249
rect 247 215 257 249
rect 203 199 257 215
rect 299 249 353 265
rect 299 215 309 249
rect 343 215 353 249
rect 299 199 353 215
rect 395 249 449 265
rect 395 215 405 249
rect 439 215 449 249
rect 395 199 449 215
rect 491 249 545 265
rect 491 215 501 249
rect 535 215 545 249
rect 491 199 545 215
rect 131 177 161 199
rect 215 177 245 199
rect 311 177 341 199
rect 395 177 425 199
rect 492 177 522 199
rect 492 67 522 93
rect 131 21 161 47
rect 215 21 245 47
rect 311 21 341 47
rect 395 21 425 47
<< polycont >>
rect 107 215 141 249
rect 213 215 247 249
rect 309 215 343 249
rect 405 215 439 249
rect 501 215 535 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 474 69 490
rect 17 440 35 474
rect 17 406 69 440
rect 419 471 485 527
rect 419 437 435 471
rect 469 437 485 471
rect 17 372 35 406
rect 17 165 69 372
rect 105 397 627 401
rect 105 363 532 397
rect 566 363 627 397
rect 105 359 627 363
rect 105 249 149 359
rect 105 215 107 249
rect 141 215 149 249
rect 105 199 149 215
rect 197 249 257 323
rect 197 215 213 249
rect 247 215 257 249
rect 197 199 257 215
rect 291 249 357 323
rect 291 215 309 249
rect 343 215 357 249
rect 291 199 357 215
rect 391 249 455 323
rect 391 215 405 249
rect 439 215 455 249
rect 391 199 455 215
rect 489 249 559 323
rect 489 215 501 249
rect 535 215 559 249
rect 489 199 559 215
rect 593 165 627 359
rect 17 131 385 165
rect 171 116 211 131
rect 71 89 137 96
rect 71 55 87 89
rect 121 55 137 89
rect 205 82 211 116
rect 345 116 385 131
rect 171 60 211 82
rect 245 95 311 97
rect 245 61 261 95
rect 295 61 311 95
rect 345 82 351 116
rect 345 62 385 82
rect 419 163 485 165
rect 419 129 435 163
rect 469 129 485 163
rect 419 95 485 129
rect 71 17 137 55
rect 245 17 311 61
rect 419 61 435 95
rect 469 61 485 95
rect 532 149 627 165
rect 566 131 627 149
rect 532 81 566 115
rect 419 17 485 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4b_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1176742
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1171536
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
