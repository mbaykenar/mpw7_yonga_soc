magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 99 157 623 203
rect 1 21 728 157
rect 29 -17 63 21
<< scnmos >>
rect 80 47 110 131
rect 252 47 282 177
rect 447 47 477 177
rect 619 47 649 131
<< scpmoshvt >>
rect 80 297 110 497
rect 252 333 282 497
rect 447 333 477 497
rect 619 297 649 497
<< ndiff >>
rect 125 131 252 177
rect 27 93 80 131
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 93 252 131
rect 110 59 132 93
rect 166 59 252 93
rect 110 47 252 59
rect 282 161 335 177
rect 282 127 293 161
rect 327 127 335 161
rect 282 93 335 127
rect 282 59 293 93
rect 327 59 335 93
rect 282 47 335 59
rect 394 93 447 177
rect 394 59 402 93
rect 436 59 447 93
rect 394 47 447 59
rect 477 131 597 177
rect 477 93 619 131
rect 477 59 558 93
rect 592 59 619 93
rect 477 47 619 59
rect 649 93 702 131
rect 649 59 660 93
rect 694 59 702 93
rect 649 47 702 59
<< pdiff >>
rect 27 478 80 497
rect 27 444 35 478
rect 69 444 80 478
rect 27 410 80 444
rect 27 376 35 410
rect 69 376 80 410
rect 27 297 80 376
rect 110 485 252 497
rect 110 451 135 485
rect 169 451 252 485
rect 110 417 252 451
rect 110 383 135 417
rect 169 383 252 417
rect 110 333 252 383
rect 282 485 335 497
rect 282 451 293 485
rect 327 451 335 485
rect 282 417 335 451
rect 282 383 293 417
rect 327 383 335 417
rect 282 333 335 383
rect 394 485 447 497
rect 394 451 402 485
rect 436 451 447 485
rect 394 417 447 451
rect 394 383 402 417
rect 436 383 447 417
rect 394 333 447 383
rect 477 485 619 497
rect 477 451 558 485
rect 592 451 619 485
rect 477 417 619 451
rect 477 383 558 417
rect 592 383 619 417
rect 477 333 619 383
rect 110 297 232 333
rect 509 297 619 333
rect 649 485 702 497
rect 649 451 660 485
rect 694 451 702 485
rect 649 417 702 451
rect 649 383 660 417
rect 694 383 702 417
rect 649 297 702 383
<< ndiffc >>
rect 35 59 69 93
rect 132 59 166 93
rect 293 127 327 161
rect 293 59 327 93
rect 402 59 436 93
rect 558 59 592 93
rect 660 59 694 93
<< pdiffc >>
rect 35 444 69 478
rect 35 376 69 410
rect 135 451 169 485
rect 135 383 169 417
rect 293 451 327 485
rect 293 383 327 417
rect 402 451 436 485
rect 402 383 436 417
rect 558 451 592 485
rect 558 383 592 417
rect 660 451 694 485
rect 660 383 694 417
<< poly >>
rect 80 497 110 523
rect 252 497 282 523
rect 447 497 477 523
rect 619 497 649 523
rect 80 265 110 297
rect 46 249 112 265
rect 252 259 282 333
rect 447 266 477 333
rect 619 266 649 297
rect 46 215 62 249
rect 96 215 112 249
rect 46 205 112 215
rect 154 249 282 259
rect 154 215 170 249
rect 204 215 282 249
rect 80 131 110 205
rect 154 199 282 215
rect 401 249 541 266
rect 401 215 417 249
rect 451 215 485 249
rect 519 215 541 249
rect 401 200 541 215
rect 583 249 649 266
rect 583 215 599 249
rect 633 215 649 249
rect 583 200 649 215
rect 252 177 282 199
rect 447 177 477 200
rect 619 131 649 200
rect 80 21 110 47
rect 252 21 282 47
rect 447 21 477 47
rect 619 21 649 47
<< polycont >>
rect 62 215 96 249
rect 170 215 204 249
rect 417 215 451 249
rect 485 215 519 249
rect 599 215 633 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 478 85 493
rect 17 444 35 478
rect 69 444 85 478
rect 17 410 85 444
rect 17 376 35 410
rect 69 376 85 410
rect 17 333 85 376
rect 119 485 185 527
rect 119 451 135 485
rect 169 451 185 485
rect 119 417 185 451
rect 119 383 135 417
rect 169 383 185 417
rect 119 367 185 383
rect 277 485 352 493
rect 277 451 293 485
rect 327 451 352 485
rect 277 417 352 451
rect 277 383 293 417
rect 327 383 352 417
rect 277 367 352 383
rect 17 299 243 333
rect 17 249 112 265
rect 17 215 62 249
rect 96 215 112 249
rect 17 211 112 215
rect 146 249 243 299
rect 146 215 170 249
rect 204 215 243 249
rect 146 177 243 215
rect 17 143 243 177
rect 318 250 352 367
rect 386 485 482 493
rect 386 451 402 485
rect 436 451 482 485
rect 386 417 482 451
rect 386 383 402 417
rect 436 383 482 417
rect 386 318 482 383
rect 528 485 608 527
rect 528 451 558 485
rect 592 451 608 485
rect 528 417 608 451
rect 528 383 558 417
rect 592 383 608 417
rect 528 352 608 383
rect 642 485 719 493
rect 642 451 660 485
rect 694 451 719 485
rect 642 417 719 451
rect 642 383 660 417
rect 694 383 719 417
rect 642 352 719 383
rect 386 284 639 318
rect 318 249 537 250
rect 318 215 417 249
rect 451 215 485 249
rect 519 215 537 249
rect 318 211 537 215
rect 571 249 639 284
rect 571 215 599 249
rect 633 215 639 249
rect 318 165 352 211
rect 571 177 639 215
rect 277 161 352 165
rect 17 93 85 143
rect 277 127 293 161
rect 327 127 352 161
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 119 93 182 109
rect 119 59 132 93
rect 166 59 182 93
rect 119 17 182 59
rect 277 93 352 127
rect 277 59 293 93
rect 327 59 352 93
rect 277 51 352 59
rect 386 143 639 177
rect 386 93 452 143
rect 673 109 719 352
rect 386 59 402 93
rect 436 59 452 93
rect 386 51 452 59
rect 542 93 608 109
rect 542 59 558 93
rect 592 59 608 93
rect 542 17 608 59
rect 642 93 719 109
rect 642 59 660 93
rect 694 59 719 93
rect 642 57 719 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 673 85 707 119 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 673 153 707 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 673 289 707 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 673 357 707 391 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 673 425 707 459 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 clkdlybuf4s15_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3188518
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3182366
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 18.400 13.600 
<< end >>
