magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfl1sd2__example_55959141808316  sky130_fd_pr__hvdfl1sd2__example_55959141808316_0
timestamp 1649977179
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_0
timestamp 1649977179
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808506  sky130_fd_pr__hvdftpl1s2__example_55959141808506_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 324 97 324 97 0 FreeSans 300 0 0 0 D
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 S
flabel comment s -130 97 -130 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 48476924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48475350
<< end >>
