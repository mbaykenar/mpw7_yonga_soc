magic
tech sky130A
timestamp 1649977179
<< properties >>
string GDS_END 11280140
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11273480
<< end >>
