magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 838 157 1195 203
rect 1 21 1195 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 355 47 385 131
rect 439 47 469 131
rect 547 47 577 119
rect 633 47 663 119
rect 728 47 758 131
rect 916 47 946 177
rect 1003 47 1033 177
rect 1087 47 1117 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 355 369 385 497
rect 439 369 469 497
rect 535 413 565 497
rect 656 413 686 497
rect 728 413 758 497
rect 916 297 946 497
rect 1003 297 1033 497
rect 1087 297 1117 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 303 119 355 131
rect 303 85 311 119
rect 345 85 355 119
rect 303 47 355 85
rect 385 89 439 131
rect 385 55 395 89
rect 429 55 439 89
rect 385 47 439 55
rect 469 119 519 131
rect 864 133 916 177
rect 678 119 728 131
rect 469 47 547 119
rect 577 107 633 119
rect 577 73 588 107
rect 622 73 633 107
rect 577 47 633 73
rect 663 47 728 119
rect 758 106 810 131
rect 758 72 768 106
rect 802 72 810 106
rect 758 47 810 72
rect 864 99 872 133
rect 906 99 916 133
rect 864 47 916 99
rect 946 127 1003 177
rect 946 93 959 127
rect 993 93 1003 127
rect 946 47 1003 93
rect 1033 133 1087 177
rect 1033 99 1043 133
rect 1077 99 1087 133
rect 1033 47 1087 99
rect 1117 93 1169 177
rect 1117 59 1127 93
rect 1161 59 1169 93
rect 1117 47 1169 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 303 483 355 497
rect 303 449 311 483
rect 345 449 355 483
rect 303 415 355 449
rect 303 381 311 415
rect 345 381 355 415
rect 303 369 355 381
rect 385 485 439 497
rect 385 451 395 485
rect 429 451 439 485
rect 385 417 439 451
rect 385 383 395 417
rect 429 383 439 417
rect 385 369 439 383
rect 469 413 535 497
rect 565 485 656 497
rect 565 451 600 485
rect 634 451 656 485
rect 565 413 656 451
rect 686 413 728 497
rect 758 477 810 497
rect 758 443 768 477
rect 802 443 810 477
rect 758 413 810 443
rect 864 471 916 497
rect 864 437 872 471
rect 906 437 916 471
rect 469 369 519 413
rect 864 368 916 437
rect 864 334 872 368
rect 906 334 916 368
rect 864 297 916 334
rect 946 484 1003 497
rect 946 450 959 484
rect 993 450 1003 484
rect 946 364 1003 450
rect 946 330 959 364
rect 993 330 1003 364
rect 946 297 1003 330
rect 1033 475 1087 497
rect 1033 441 1043 475
rect 1077 441 1087 475
rect 1033 384 1087 441
rect 1033 350 1043 384
rect 1077 350 1087 384
rect 1033 297 1087 350
rect 1117 485 1169 497
rect 1117 451 1127 485
rect 1161 451 1169 485
rect 1117 417 1169 451
rect 1117 383 1127 417
rect 1161 383 1169 417
rect 1117 297 1169 383
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 311 85 345 119
rect 395 55 429 89
rect 588 73 622 107
rect 768 72 802 106
rect 872 99 906 133
rect 959 93 993 127
rect 1043 99 1077 133
rect 1127 59 1161 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 311 449 345 483
rect 311 381 345 415
rect 395 451 429 485
rect 395 383 429 417
rect 600 451 634 485
rect 768 443 802 477
rect 872 437 906 471
rect 872 334 906 368
rect 959 450 993 484
rect 959 330 993 364
rect 1043 441 1077 475
rect 1043 350 1077 384
rect 1127 451 1161 485
rect 1127 383 1161 417
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 355 497 385 523
rect 439 497 469 523
rect 535 497 565 523
rect 656 497 686 523
rect 728 497 758 523
rect 916 497 946 523
rect 1003 497 1033 523
rect 1087 497 1117 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 355 241 385 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 302 225 385 241
rect 302 191 312 225
rect 346 191 385 225
rect 439 219 469 369
rect 535 337 565 413
rect 656 375 686 413
rect 511 321 565 337
rect 607 365 686 375
rect 607 331 623 365
rect 657 331 686 365
rect 607 321 686 331
rect 728 373 758 413
rect 728 357 816 373
rect 728 323 772 357
rect 806 323 816 357
rect 511 287 521 321
rect 555 287 565 321
rect 511 279 565 287
rect 728 307 816 323
rect 511 271 663 279
rect 535 249 663 271
rect 302 175 385 191
rect 355 131 385 175
rect 428 203 482 219
rect 428 169 438 203
rect 472 169 482 203
rect 428 153 482 169
rect 537 191 591 207
rect 537 157 547 191
rect 581 157 591 191
rect 439 131 469 153
rect 537 141 591 157
rect 547 119 577 141
rect 633 119 663 249
rect 728 131 758 307
rect 916 265 946 297
rect 1003 265 1033 297
rect 1087 265 1117 297
rect 800 249 946 265
rect 800 215 810 249
rect 844 215 946 249
rect 800 199 946 215
rect 988 249 1117 265
rect 988 215 998 249
rect 1032 215 1117 249
rect 988 199 1117 215
rect 916 177 946 199
rect 1003 177 1033 199
rect 1087 177 1117 199
rect 79 21 109 47
rect 163 21 193 47
rect 355 21 385 47
rect 439 21 469 47
rect 547 21 577 47
rect 633 21 663 47
rect 728 21 758 47
rect 916 21 946 47
rect 1003 21 1033 47
rect 1087 21 1117 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 312 191 346 225
rect 623 331 657 365
rect 772 323 806 357
rect 521 287 555 321
rect 438 169 472 203
rect 547 157 581 191
rect 810 215 844 249
rect 998 215 1032 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 395 485 458 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 295 449 311 483
rect 345 449 361 483
rect 295 415 361 449
rect 295 381 311 415
rect 345 381 361 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 295 333 361 381
rect 429 451 458 485
rect 584 451 600 485
rect 634 451 734 485
rect 395 417 458 451
rect 429 383 458 417
rect 395 367 458 383
rect 498 391 555 401
rect 532 357 555 391
rect 295 299 432 333
rect 296 225 362 265
rect 296 191 312 225
rect 346 191 362 225
rect 398 219 432 299
rect 498 321 555 357
rect 498 287 521 321
rect 498 271 555 287
rect 589 365 657 399
rect 589 331 623 365
rect 589 323 657 331
rect 589 289 590 323
rect 624 289 657 323
rect 589 283 657 289
rect 398 203 472 219
rect 589 207 623 283
rect 700 265 734 451
rect 768 477 828 527
rect 802 443 828 477
rect 768 427 828 443
rect 872 471 916 487
rect 906 437 916 471
rect 872 373 916 437
rect 772 368 916 373
rect 772 357 872 368
rect 806 334 872 357
rect 906 334 916 368
rect 806 323 916 334
rect 772 307 916 323
rect 882 265 916 307
rect 952 484 1009 527
rect 952 450 959 484
rect 993 450 1009 484
rect 952 364 1009 450
rect 952 330 959 364
rect 993 330 1009 364
rect 952 299 1009 330
rect 1043 475 1093 491
rect 1077 441 1093 475
rect 1043 384 1093 441
rect 1077 350 1093 384
rect 1127 485 1179 527
rect 1161 451 1179 485
rect 1127 417 1179 451
rect 1161 383 1179 417
rect 1127 351 1179 383
rect 1043 328 1093 350
rect 1043 299 1100 328
rect 1066 265 1100 299
rect 700 249 844 265
rect 700 233 810 249
rect 398 169 438 203
rect 398 157 472 169
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 311 153 472 157
rect 547 191 623 207
rect 581 157 623 191
rect 311 123 432 153
rect 547 141 623 157
rect 670 215 810 233
rect 670 199 844 215
rect 882 249 1032 265
rect 882 215 998 249
rect 882 199 1032 215
rect 1066 199 1179 265
rect 311 119 345 123
rect 670 107 704 199
rect 882 165 916 199
rect 1066 165 1100 199
rect 311 69 345 85
rect 103 17 169 59
rect 379 55 395 89
rect 429 55 445 89
rect 572 73 588 107
rect 622 73 704 107
rect 752 106 818 165
rect 379 17 445 55
rect 752 72 768 106
rect 802 72 818 106
rect 872 133 916 165
rect 906 99 916 133
rect 872 83 916 99
rect 952 127 1009 165
rect 952 93 959 127
rect 993 93 1009 127
rect 752 17 818 72
rect 952 17 1009 93
rect 1043 137 1100 165
rect 1043 133 1093 137
rect 1077 99 1093 133
rect 1043 83 1093 99
rect 1127 93 1179 110
rect 1161 59 1179 93
rect 1127 17 1179 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 498 357 532 391
rect 590 289 624 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 486 391 544 397
rect 486 388 498 391
rect 248 360 498 388
rect 248 357 260 360
rect 202 351 260 357
rect 486 357 498 360
rect 532 357 544 391
rect 486 351 544 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 578 323 636 329
rect 578 320 590 323
rect 156 292 590 320
rect 156 289 168 292
rect 110 283 168 289
rect 578 289 590 292
rect 624 289 636 323
rect 578 283 636 289
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 314 221 348 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1054 357 1088 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1054 425 1088 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1054 85 1088 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1139 221 1173 255 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 dlxtn_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 2854808
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2844736
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 29.900 13.600 
<< end >>
