magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect 172 3385 1880 3493
rect 172 3169 1895 3385
rect 172 2953 1102 3169
<< pwell >>
rect 399 1475 1369 1727
rect 399 639 1717 1291
rect 441 529 1651 639
<< mvnmos >>
rect 478 1501 578 1701
rect 754 1501 854 1701
rect 910 1501 1010 1701
rect 1190 1501 1290 1701
rect 478 665 578 1265
rect 634 665 734 1265
rect 790 665 890 1265
rect 946 665 1046 1265
rect 1102 665 1202 1265
rect 1258 665 1358 1265
rect 1538 665 1638 1265
<< mvpmos >>
rect 291 3019 391 3319
rect 447 3019 547 3319
rect 727 3019 827 3319
rect 883 3019 983 3319
rect 1320 3235 1520 3319
rect 1576 3235 1776 3319
<< mvndiff >>
rect 425 1689 478 1701
rect 425 1655 433 1689
rect 467 1655 478 1689
rect 425 1621 478 1655
rect 425 1587 433 1621
rect 467 1587 478 1621
rect 425 1553 478 1587
rect 425 1519 433 1553
rect 467 1519 478 1553
rect 425 1501 478 1519
rect 578 1689 631 1701
rect 578 1655 589 1689
rect 623 1655 631 1689
rect 578 1621 631 1655
rect 578 1587 589 1621
rect 623 1587 631 1621
rect 578 1553 631 1587
rect 578 1519 589 1553
rect 623 1519 631 1553
rect 578 1501 631 1519
rect 701 1683 754 1701
rect 701 1649 709 1683
rect 743 1649 754 1683
rect 701 1615 754 1649
rect 701 1581 709 1615
rect 743 1581 754 1615
rect 701 1547 754 1581
rect 701 1513 709 1547
rect 743 1513 754 1547
rect 701 1501 754 1513
rect 854 1683 910 1701
rect 854 1649 865 1683
rect 899 1649 910 1683
rect 854 1615 910 1649
rect 854 1581 865 1615
rect 899 1581 910 1615
rect 854 1547 910 1581
rect 854 1513 865 1547
rect 899 1513 910 1547
rect 854 1501 910 1513
rect 1010 1683 1063 1701
rect 1010 1649 1021 1683
rect 1055 1649 1063 1683
rect 1010 1615 1063 1649
rect 1010 1581 1021 1615
rect 1055 1581 1063 1615
rect 1010 1547 1063 1581
rect 1010 1513 1021 1547
rect 1055 1513 1063 1547
rect 1010 1501 1063 1513
rect 1137 1683 1190 1701
rect 1137 1649 1145 1683
rect 1179 1649 1190 1683
rect 1137 1615 1190 1649
rect 1137 1581 1145 1615
rect 1179 1581 1190 1615
rect 1137 1547 1190 1581
rect 1137 1513 1145 1547
rect 1179 1513 1190 1547
rect 1137 1501 1190 1513
rect 1290 1683 1343 1701
rect 1290 1649 1301 1683
rect 1335 1649 1343 1683
rect 1290 1615 1343 1649
rect 1290 1581 1301 1615
rect 1335 1581 1343 1615
rect 1290 1547 1343 1581
rect 1290 1513 1301 1547
rect 1335 1513 1343 1547
rect 1290 1501 1343 1513
rect 425 1187 478 1265
rect 425 1153 433 1187
rect 467 1153 478 1187
rect 425 1119 478 1153
rect 425 1085 433 1119
rect 467 1085 478 1119
rect 425 1051 478 1085
rect 425 1017 433 1051
rect 467 1017 478 1051
rect 425 983 478 1017
rect 425 949 433 983
rect 467 949 478 983
rect 425 915 478 949
rect 425 881 433 915
rect 467 881 478 915
rect 425 847 478 881
rect 425 813 433 847
rect 467 813 478 847
rect 425 779 478 813
rect 425 745 433 779
rect 467 745 478 779
rect 425 711 478 745
rect 425 677 433 711
rect 467 677 478 711
rect 425 665 478 677
rect 578 1187 634 1265
rect 578 1153 589 1187
rect 623 1153 634 1187
rect 578 1119 634 1153
rect 578 1085 589 1119
rect 623 1085 634 1119
rect 578 1051 634 1085
rect 578 1017 589 1051
rect 623 1017 634 1051
rect 578 983 634 1017
rect 578 949 589 983
rect 623 949 634 983
rect 578 915 634 949
rect 578 881 589 915
rect 623 881 634 915
rect 578 847 634 881
rect 578 813 589 847
rect 623 813 634 847
rect 578 779 634 813
rect 578 745 589 779
rect 623 745 634 779
rect 578 711 634 745
rect 578 677 589 711
rect 623 677 634 711
rect 578 665 634 677
rect 734 1187 790 1265
rect 734 1153 745 1187
rect 779 1153 790 1187
rect 734 1119 790 1153
rect 734 1085 745 1119
rect 779 1085 790 1119
rect 734 1051 790 1085
rect 734 1017 745 1051
rect 779 1017 790 1051
rect 734 983 790 1017
rect 734 949 745 983
rect 779 949 790 983
rect 734 915 790 949
rect 734 881 745 915
rect 779 881 790 915
rect 734 847 790 881
rect 734 813 745 847
rect 779 813 790 847
rect 734 779 790 813
rect 734 745 745 779
rect 779 745 790 779
rect 734 711 790 745
rect 734 677 745 711
rect 779 677 790 711
rect 734 665 790 677
rect 890 1187 946 1265
rect 890 1153 901 1187
rect 935 1153 946 1187
rect 890 1119 946 1153
rect 890 1085 901 1119
rect 935 1085 946 1119
rect 890 1051 946 1085
rect 890 1017 901 1051
rect 935 1017 946 1051
rect 890 983 946 1017
rect 890 949 901 983
rect 935 949 946 983
rect 890 915 946 949
rect 890 881 901 915
rect 935 881 946 915
rect 890 847 946 881
rect 890 813 901 847
rect 935 813 946 847
rect 890 779 946 813
rect 890 745 901 779
rect 935 745 946 779
rect 890 711 946 745
rect 890 677 901 711
rect 935 677 946 711
rect 890 665 946 677
rect 1046 1187 1102 1265
rect 1046 1153 1057 1187
rect 1091 1153 1102 1187
rect 1046 1119 1102 1153
rect 1046 1085 1057 1119
rect 1091 1085 1102 1119
rect 1046 1051 1102 1085
rect 1046 1017 1057 1051
rect 1091 1017 1102 1051
rect 1046 983 1102 1017
rect 1046 949 1057 983
rect 1091 949 1102 983
rect 1046 915 1102 949
rect 1046 881 1057 915
rect 1091 881 1102 915
rect 1046 847 1102 881
rect 1046 813 1057 847
rect 1091 813 1102 847
rect 1046 779 1102 813
rect 1046 745 1057 779
rect 1091 745 1102 779
rect 1046 711 1102 745
rect 1046 677 1057 711
rect 1091 677 1102 711
rect 1046 665 1102 677
rect 1202 1187 1258 1265
rect 1202 1153 1213 1187
rect 1247 1153 1258 1187
rect 1202 1119 1258 1153
rect 1202 1085 1213 1119
rect 1247 1085 1258 1119
rect 1202 1051 1258 1085
rect 1202 1017 1213 1051
rect 1247 1017 1258 1051
rect 1202 983 1258 1017
rect 1202 949 1213 983
rect 1247 949 1258 983
rect 1202 915 1258 949
rect 1202 881 1213 915
rect 1247 881 1258 915
rect 1202 847 1258 881
rect 1202 813 1213 847
rect 1247 813 1258 847
rect 1202 779 1258 813
rect 1202 745 1213 779
rect 1247 745 1258 779
rect 1202 711 1258 745
rect 1202 677 1213 711
rect 1247 677 1258 711
rect 1202 665 1258 677
rect 1358 1187 1411 1265
rect 1358 1153 1369 1187
rect 1403 1153 1411 1187
rect 1358 1119 1411 1153
rect 1358 1085 1369 1119
rect 1403 1085 1411 1119
rect 1358 1051 1411 1085
rect 1358 1017 1369 1051
rect 1403 1017 1411 1051
rect 1358 983 1411 1017
rect 1358 949 1369 983
rect 1403 949 1411 983
rect 1358 915 1411 949
rect 1358 881 1369 915
rect 1403 881 1411 915
rect 1358 847 1411 881
rect 1358 813 1369 847
rect 1403 813 1411 847
rect 1358 779 1411 813
rect 1358 745 1369 779
rect 1403 745 1411 779
rect 1358 711 1411 745
rect 1358 677 1369 711
rect 1403 677 1411 711
rect 1358 665 1411 677
rect 1485 1187 1538 1265
rect 1485 1153 1493 1187
rect 1527 1153 1538 1187
rect 1485 1119 1538 1153
rect 1485 1085 1493 1119
rect 1527 1085 1538 1119
rect 1485 1051 1538 1085
rect 1485 1017 1493 1051
rect 1527 1017 1538 1051
rect 1485 983 1538 1017
rect 1485 949 1493 983
rect 1527 949 1538 983
rect 1485 915 1538 949
rect 1485 881 1493 915
rect 1527 881 1538 915
rect 1485 847 1538 881
rect 1485 813 1493 847
rect 1527 813 1538 847
rect 1485 779 1538 813
rect 1485 745 1493 779
rect 1527 745 1538 779
rect 1485 711 1538 745
rect 1485 677 1493 711
rect 1527 677 1538 711
rect 1485 665 1538 677
rect 1638 1187 1691 1265
rect 1638 1153 1649 1187
rect 1683 1153 1691 1187
rect 1638 1119 1691 1153
rect 1638 1085 1649 1119
rect 1683 1085 1691 1119
rect 1638 1051 1691 1085
rect 1638 1017 1649 1051
rect 1683 1017 1691 1051
rect 1638 983 1691 1017
rect 1638 949 1649 983
rect 1683 949 1691 983
rect 1638 915 1691 949
rect 1638 881 1649 915
rect 1683 881 1691 915
rect 1638 847 1691 881
rect 1638 813 1649 847
rect 1683 813 1691 847
rect 1638 779 1691 813
rect 1638 745 1649 779
rect 1683 745 1691 779
rect 1638 711 1691 745
rect 1638 677 1649 711
rect 1683 677 1691 711
rect 1638 665 1691 677
<< mvpdiff >>
rect 238 3307 291 3319
rect 238 3273 246 3307
rect 280 3273 291 3307
rect 238 3239 291 3273
rect 238 3205 246 3239
rect 280 3205 291 3239
rect 238 3171 291 3205
rect 238 3137 246 3171
rect 280 3137 291 3171
rect 238 3103 291 3137
rect 238 3069 246 3103
rect 280 3069 291 3103
rect 238 3019 291 3069
rect 391 3307 447 3319
rect 391 3273 402 3307
rect 436 3273 447 3307
rect 391 3239 447 3273
rect 391 3205 402 3239
rect 436 3205 447 3239
rect 391 3171 447 3205
rect 391 3137 402 3171
rect 436 3137 447 3171
rect 391 3103 447 3137
rect 391 3069 402 3103
rect 436 3069 447 3103
rect 391 3019 447 3069
rect 547 3307 600 3319
rect 547 3273 558 3307
rect 592 3273 600 3307
rect 547 3239 600 3273
rect 547 3205 558 3239
rect 592 3205 600 3239
rect 547 3171 600 3205
rect 547 3137 558 3171
rect 592 3137 600 3171
rect 547 3103 600 3137
rect 547 3069 558 3103
rect 592 3069 600 3103
rect 547 3019 600 3069
rect 674 3269 727 3319
rect 674 3235 682 3269
rect 716 3235 727 3269
rect 674 3201 727 3235
rect 674 3167 682 3201
rect 716 3167 727 3201
rect 674 3133 727 3167
rect 674 3099 682 3133
rect 716 3099 727 3133
rect 674 3065 727 3099
rect 674 3031 682 3065
rect 716 3031 727 3065
rect 674 3019 727 3031
rect 827 3269 883 3319
rect 827 3235 838 3269
rect 872 3235 883 3269
rect 827 3201 883 3235
rect 827 3167 838 3201
rect 872 3167 883 3201
rect 827 3133 883 3167
rect 827 3099 838 3133
rect 872 3099 883 3133
rect 827 3065 883 3099
rect 827 3031 838 3065
rect 872 3031 883 3065
rect 827 3019 883 3031
rect 983 3269 1036 3319
rect 983 3235 994 3269
rect 1028 3235 1036 3269
rect 1267 3281 1320 3319
rect 1267 3247 1275 3281
rect 1309 3247 1320 3281
rect 1267 3235 1320 3247
rect 1520 3281 1576 3319
rect 1520 3247 1531 3281
rect 1565 3247 1576 3281
rect 1520 3235 1576 3247
rect 1776 3281 1829 3319
rect 1776 3247 1787 3281
rect 1821 3247 1829 3281
rect 1776 3235 1829 3247
rect 983 3201 1036 3235
rect 983 3167 994 3201
rect 1028 3167 1036 3201
rect 983 3133 1036 3167
rect 983 3099 994 3133
rect 1028 3099 1036 3133
rect 983 3065 1036 3099
rect 983 3031 994 3065
rect 1028 3031 1036 3065
rect 983 3019 1036 3031
<< mvndiffc >>
rect 433 1655 467 1689
rect 433 1587 467 1621
rect 433 1519 467 1553
rect 589 1655 623 1689
rect 589 1587 623 1621
rect 589 1519 623 1553
rect 709 1649 743 1683
rect 709 1581 743 1615
rect 709 1513 743 1547
rect 865 1649 899 1683
rect 865 1581 899 1615
rect 865 1513 899 1547
rect 1021 1649 1055 1683
rect 1021 1581 1055 1615
rect 1021 1513 1055 1547
rect 1145 1649 1179 1683
rect 1145 1581 1179 1615
rect 1145 1513 1179 1547
rect 1301 1649 1335 1683
rect 1301 1581 1335 1615
rect 1301 1513 1335 1547
rect 433 1153 467 1187
rect 433 1085 467 1119
rect 433 1017 467 1051
rect 433 949 467 983
rect 433 881 467 915
rect 433 813 467 847
rect 433 745 467 779
rect 433 677 467 711
rect 589 1153 623 1187
rect 589 1085 623 1119
rect 589 1017 623 1051
rect 589 949 623 983
rect 589 881 623 915
rect 589 813 623 847
rect 589 745 623 779
rect 589 677 623 711
rect 745 1153 779 1187
rect 745 1085 779 1119
rect 745 1017 779 1051
rect 745 949 779 983
rect 745 881 779 915
rect 745 813 779 847
rect 745 745 779 779
rect 745 677 779 711
rect 901 1153 935 1187
rect 901 1085 935 1119
rect 901 1017 935 1051
rect 901 949 935 983
rect 901 881 935 915
rect 901 813 935 847
rect 901 745 935 779
rect 901 677 935 711
rect 1057 1153 1091 1187
rect 1057 1085 1091 1119
rect 1057 1017 1091 1051
rect 1057 949 1091 983
rect 1057 881 1091 915
rect 1057 813 1091 847
rect 1057 745 1091 779
rect 1057 677 1091 711
rect 1213 1153 1247 1187
rect 1213 1085 1247 1119
rect 1213 1017 1247 1051
rect 1213 949 1247 983
rect 1213 881 1247 915
rect 1213 813 1247 847
rect 1213 745 1247 779
rect 1213 677 1247 711
rect 1369 1153 1403 1187
rect 1369 1085 1403 1119
rect 1369 1017 1403 1051
rect 1369 949 1403 983
rect 1369 881 1403 915
rect 1369 813 1403 847
rect 1369 745 1403 779
rect 1369 677 1403 711
rect 1493 1153 1527 1187
rect 1493 1085 1527 1119
rect 1493 1017 1527 1051
rect 1493 949 1527 983
rect 1493 881 1527 915
rect 1493 813 1527 847
rect 1493 745 1527 779
rect 1493 677 1527 711
rect 1649 1153 1683 1187
rect 1649 1085 1683 1119
rect 1649 1017 1683 1051
rect 1649 949 1683 983
rect 1649 881 1683 915
rect 1649 813 1683 847
rect 1649 745 1683 779
rect 1649 677 1683 711
<< mvpdiffc >>
rect 246 3273 280 3307
rect 246 3205 280 3239
rect 246 3137 280 3171
rect 246 3069 280 3103
rect 402 3273 436 3307
rect 402 3205 436 3239
rect 402 3137 436 3171
rect 402 3069 436 3103
rect 558 3273 592 3307
rect 558 3205 592 3239
rect 558 3137 592 3171
rect 558 3069 592 3103
rect 682 3235 716 3269
rect 682 3167 716 3201
rect 682 3099 716 3133
rect 682 3031 716 3065
rect 838 3235 872 3269
rect 838 3167 872 3201
rect 838 3099 872 3133
rect 838 3031 872 3065
rect 994 3235 1028 3269
rect 1275 3247 1309 3281
rect 1531 3247 1565 3281
rect 1787 3247 1821 3281
rect 994 3167 1028 3201
rect 994 3099 1028 3133
rect 994 3031 1028 3065
<< psubdiff >>
rect 467 555 491 589
rect 525 555 563 589
rect 597 555 635 589
rect 669 555 707 589
rect 741 555 779 589
rect 813 555 851 589
rect 885 555 923 589
rect 957 555 995 589
rect 1029 555 1067 589
rect 1101 555 1139 589
rect 1173 555 1211 589
rect 1245 555 1283 589
rect 1317 555 1354 589
rect 1388 555 1425 589
rect 1459 555 1496 589
rect 1530 555 1567 589
rect 1601 555 1625 589
<< mvnsubdiff >>
rect 238 3393 262 3427
rect 296 3393 334 3427
rect 368 3393 406 3427
rect 440 3393 478 3427
rect 512 3393 549 3427
rect 583 3393 620 3427
rect 654 3393 691 3427
rect 725 3393 762 3427
rect 796 3393 833 3427
rect 867 3393 904 3427
rect 938 3393 975 3427
rect 1009 3393 1046 3427
rect 1080 3393 1117 3427
rect 1151 3393 1188 3427
rect 1222 3393 1259 3427
rect 1293 3393 1330 3427
rect 1364 3393 1401 3427
rect 1435 3393 1472 3427
rect 1506 3393 1543 3427
rect 1577 3393 1614 3427
rect 1648 3393 1685 3427
rect 1719 3393 1756 3427
rect 1790 3393 1814 3427
<< psubdiffcont >>
rect 491 555 525 589
rect 563 555 597 589
rect 635 555 669 589
rect 707 555 741 589
rect 779 555 813 589
rect 851 555 885 589
rect 923 555 957 589
rect 995 555 1029 589
rect 1067 555 1101 589
rect 1139 555 1173 589
rect 1211 555 1245 589
rect 1283 555 1317 589
rect 1354 555 1388 589
rect 1425 555 1459 589
rect 1496 555 1530 589
rect 1567 555 1601 589
<< mvnsubdiffcont >>
rect 262 3393 296 3427
rect 334 3393 368 3427
rect 406 3393 440 3427
rect 478 3393 512 3427
rect 549 3393 583 3427
rect 620 3393 654 3427
rect 691 3393 725 3427
rect 762 3393 796 3427
rect 833 3393 867 3427
rect 904 3393 938 3427
rect 975 3393 1009 3427
rect 1046 3393 1080 3427
rect 1117 3393 1151 3427
rect 1188 3393 1222 3427
rect 1259 3393 1293 3427
rect 1330 3393 1364 3427
rect 1401 3393 1435 3427
rect 1472 3393 1506 3427
rect 1543 3393 1577 3427
rect 1614 3393 1648 3427
rect 1685 3393 1719 3427
rect 1756 3393 1790 3427
<< poly >>
rect 291 3319 391 3345
rect 447 3319 547 3345
rect 727 3319 827 3351
rect 883 3319 983 3351
rect 1320 3319 1520 3351
rect 1576 3319 1776 3351
rect 1320 3187 1520 3235
rect 1320 3153 1336 3187
rect 1370 3153 1470 3187
rect 1504 3153 1520 3187
rect 1320 3137 1520 3153
rect 1576 3187 1776 3235
rect 1576 3153 1592 3187
rect 1626 3153 1726 3187
rect 1760 3153 1776 3187
rect 1576 3137 1776 3153
rect 291 2987 391 3019
rect 447 2987 547 3019
rect 727 2987 827 3019
rect 291 2971 547 2987
rect 291 2937 307 2971
rect 341 2937 402 2971
rect 436 2937 497 2971
rect 531 2937 547 2971
rect 291 2921 547 2937
rect 693 2971 827 2987
rect 693 2937 709 2971
rect 743 2937 777 2971
rect 811 2937 827 2971
rect 693 2921 827 2937
rect 883 2984 983 3019
rect 883 2968 1017 2984
rect 883 2934 899 2968
rect 933 2934 967 2968
rect 1001 2934 1017 2968
rect 883 2918 1017 2934
rect 478 1701 578 1727
rect 754 1701 854 1727
rect 910 1701 1010 1727
rect 1190 1701 1290 1727
rect 478 1465 578 1501
rect 754 1476 854 1501
rect 464 1449 598 1465
rect 464 1415 480 1449
rect 514 1415 548 1449
rect 582 1415 598 1449
rect 464 1399 598 1415
rect 721 1460 855 1476
rect 910 1475 1010 1501
rect 1190 1475 1290 1501
rect 721 1426 737 1460
rect 771 1426 805 1460
rect 839 1426 855 1460
rect 721 1410 855 1426
rect 906 1459 1040 1475
rect 906 1425 922 1459
rect 956 1425 990 1459
rect 1024 1425 1040 1459
rect 906 1409 1040 1425
rect 1178 1459 1312 1475
rect 1178 1425 1194 1459
rect 1228 1425 1262 1459
rect 1296 1425 1312 1459
rect 1178 1409 1312 1425
rect 478 1341 890 1357
rect 478 1307 494 1341
rect 528 1307 564 1341
rect 598 1307 633 1341
rect 667 1307 702 1341
rect 736 1307 771 1341
rect 805 1307 840 1341
rect 874 1307 890 1341
rect 478 1291 890 1307
rect 478 1265 578 1291
rect 634 1265 734 1291
rect 790 1265 890 1291
rect 946 1341 1358 1357
rect 946 1307 962 1341
rect 996 1307 1031 1341
rect 1065 1307 1100 1341
rect 1134 1307 1169 1341
rect 1203 1307 1238 1341
rect 1272 1307 1308 1341
rect 1342 1307 1358 1341
rect 946 1291 1358 1307
rect 1534 1341 1676 1357
rect 1534 1307 1550 1341
rect 1584 1307 1626 1341
rect 1660 1307 1676 1341
rect 1534 1291 1676 1307
rect 946 1265 1046 1291
rect 1102 1265 1202 1291
rect 1258 1265 1358 1291
rect 1538 1265 1638 1291
rect 478 639 578 665
rect 634 639 734 665
rect 790 639 890 665
rect 946 639 1046 665
rect 1102 639 1202 665
rect 1258 639 1358 665
rect 1538 639 1638 665
<< polycont >>
rect 1336 3153 1370 3187
rect 1470 3153 1504 3187
rect 1592 3153 1626 3187
rect 1726 3153 1760 3187
rect 307 2937 341 2971
rect 402 2937 436 2971
rect 497 2937 531 2971
rect 709 2937 743 2971
rect 777 2937 811 2971
rect 899 2934 933 2968
rect 967 2934 1001 2968
rect 480 1415 514 1449
rect 548 1415 582 1449
rect 737 1426 771 1460
rect 805 1426 839 1460
rect 922 1425 956 1459
rect 990 1425 1024 1459
rect 1194 1425 1228 1459
rect 1262 1425 1296 1459
rect 494 1307 528 1341
rect 564 1307 598 1341
rect 633 1307 667 1341
rect 702 1307 736 1341
rect 771 1307 805 1341
rect 840 1307 874 1341
rect 962 1307 996 1341
rect 1031 1307 1065 1341
rect 1100 1307 1134 1341
rect 1169 1307 1203 1341
rect 1238 1307 1272 1341
rect 1308 1307 1342 1341
rect 1550 1307 1584 1341
rect 1626 1307 1660 1341
<< locali >>
rect 238 3393 252 3427
rect 296 3393 328 3427
rect 368 3393 404 3427
rect 440 3393 478 3427
rect 514 3393 549 3427
rect 590 3393 620 3427
rect 666 3393 691 3427
rect 742 3393 762 3427
rect 818 3393 833 3427
rect 894 3393 904 3427
rect 970 3393 975 3427
rect 1009 3393 1012 3427
rect 1080 3393 1088 3427
rect 1151 3393 1164 3427
rect 1222 3393 1240 3427
rect 1293 3393 1315 3427
rect 1364 3393 1390 3427
rect 1435 3393 1465 3427
rect 1506 3393 1540 3427
rect 1577 3393 1614 3427
rect 1648 3393 1685 3427
rect 1719 3393 1756 3427
rect 1790 3393 1814 3427
rect 246 3264 280 3273
rect 246 3171 280 3205
rect 246 3103 280 3137
rect 246 3053 280 3069
rect 402 3307 436 3323
rect 402 3239 436 3273
rect 402 3171 436 3205
rect 402 3103 436 3129
rect 402 3053 436 3057
rect 558 3264 592 3273
rect 558 3171 592 3205
rect 682 3269 716 3285
rect 682 3201 716 3235
rect 682 3139 716 3167
rect 558 3103 592 3137
rect 558 3053 592 3069
rect 715 3133 716 3139
rect 681 3099 682 3105
rect 681 3067 716 3099
rect 715 3065 716 3067
rect 838 3269 872 3302
rect 838 3201 872 3230
rect 838 3133 872 3167
rect 838 3065 872 3099
rect 682 3015 716 3031
rect 761 2982 795 3020
rect 994 3269 1028 3285
rect 994 3201 1028 3235
rect 994 3133 1028 3167
rect 994 3065 1028 3099
rect 838 3015 872 3031
rect 420 2971 458 2976
rect 291 2937 307 2971
rect 341 2942 386 2971
rect 436 2942 458 2971
rect 920 2982 954 3020
rect 1167 3281 1309 3297
rect 1167 3247 1275 3281
rect 1167 3231 1309 3247
rect 1531 3281 1565 3302
rect 1167 3110 1275 3231
rect 1787 3281 1926 3297
rect 1821 3247 1926 3281
rect 1787 3231 1926 3247
rect 1320 3153 1336 3187
rect 1370 3184 1470 3187
rect 1504 3184 1520 3187
rect 1370 3153 1401 3184
rect 1435 3153 1470 3184
rect 1507 3153 1520 3184
rect 1576 3153 1592 3187
rect 1626 3153 1726 3187
rect 1760 3153 1776 3187
rect 1435 3150 1473 3153
rect 1201 3076 1239 3110
rect 1273 3091 1275 3110
rect 1576 3091 1776 3153
rect 1820 3184 1926 3231
rect 1854 3150 1892 3184
rect 1273 3076 1776 3091
rect 994 3002 1006 3031
rect 1040 3002 1078 3036
rect 1167 3032 1776 3076
rect 492 2942 497 2971
rect 341 2937 402 2942
rect 436 2937 497 2942
rect 531 2937 547 2971
rect 693 2937 709 2971
rect 743 2948 761 2971
rect 743 2937 777 2948
rect 811 2937 827 2971
rect 883 2934 899 2968
rect 954 2948 967 2968
rect 933 2934 967 2948
rect 1001 2934 1017 2968
rect 1492 1978 1564 2012
rect 1598 1978 1639 2012
rect 1673 1978 1713 2012
rect 1747 1978 1787 2012
rect 1821 1978 1861 2012
rect 1895 1978 1935 2012
rect 1969 1978 2009 2012
rect 2043 1978 2083 2012
rect 2117 1978 2157 2012
rect 2191 1978 2231 2012
rect 2265 1978 2305 2012
rect 2339 1978 2379 2012
rect 2413 1978 2453 2012
rect 2487 1978 2527 2012
rect 2561 1978 2601 2012
rect 2635 1978 2675 2012
rect 2709 1978 2749 2012
rect 2783 1978 2823 2012
rect 2857 1978 2897 2012
rect 2931 1978 2971 2012
rect 3005 1978 3045 2012
rect 3079 1978 3119 2012
rect 3153 1978 3193 2012
rect 3227 1978 3267 2012
rect 3301 1978 3341 2012
rect 3375 1978 3415 2012
rect 3449 1978 3489 2012
rect 3523 1978 3563 2012
rect 3597 1978 3637 2012
rect 3671 1978 3711 2012
rect 3745 1978 3785 2012
rect 3819 1978 3859 2012
rect 3893 1978 3933 2012
rect 3967 1978 4007 2012
rect 1492 1958 4041 1978
rect 1156 1924 1196 1958
rect 1230 1924 1270 1958
rect 1304 1924 1344 1958
rect 1378 1924 1418 1958
rect 1452 1941 4041 1958
rect 1452 1924 1526 1941
rect 433 1689 467 1705
rect 589 1691 623 1705
rect 433 1621 467 1655
rect 433 1553 467 1587
rect 619 1689 623 1691
rect 585 1655 589 1657
rect 585 1621 623 1655
rect 585 1619 589 1621
rect 619 1585 623 1587
rect 589 1553 623 1585
rect 433 1503 467 1519
rect 589 1503 623 1519
rect 709 1683 743 1699
rect 709 1615 743 1624
rect 865 1683 899 1699
rect 865 1615 899 1649
rect 709 1547 743 1552
rect 709 1497 743 1513
rect 898 1567 899 1581
rect 864 1547 899 1567
rect 864 1529 865 1547
rect 898 1497 899 1513
rect 939 1687 973 1725
rect 507 1449 541 1486
rect 464 1415 480 1449
rect 514 1448 548 1449
rect 541 1415 548 1448
rect 582 1415 598 1449
rect 721 1448 737 1460
rect 771 1448 805 1460
rect 721 1426 727 1448
rect 771 1426 799 1448
rect 839 1426 855 1460
rect 939 1459 973 1653
rect 1021 1687 1055 1725
rect 1021 1615 1055 1649
rect 1021 1547 1055 1581
rect 1021 1497 1055 1513
rect 1145 1683 1179 1699
rect 1145 1615 1179 1649
rect 1145 1547 1179 1567
rect 1301 1683 1335 1699
rect 1301 1618 1335 1649
rect 1301 1547 1335 1581
rect 1301 1497 1335 1512
rect 761 1414 799 1426
rect 906 1425 922 1459
rect 956 1448 990 1459
rect 1024 1448 1040 1459
rect 963 1425 990 1448
rect 1035 1425 1040 1448
rect 1178 1425 1194 1459
rect 1228 1425 1262 1459
rect 1296 1453 1413 1459
rect 1296 1425 1307 1453
rect 963 1414 1001 1425
rect 1341 1419 1379 1453
rect 526 1341 564 1342
rect 478 1308 492 1341
rect 478 1307 494 1308
rect 528 1307 564 1341
rect 598 1307 633 1341
rect 667 1307 702 1341
rect 736 1307 771 1341
rect 805 1307 840 1341
rect 874 1307 890 1341
rect 946 1307 962 1341
rect 996 1307 1031 1341
rect 1065 1307 1100 1341
rect 1134 1307 1169 1341
rect 1203 1307 1238 1341
rect 1272 1307 1308 1341
rect 1347 1308 1385 1342
rect 1342 1307 1358 1308
rect 1534 1307 1550 1341
rect 1584 1340 1626 1341
rect 1660 1340 1676 1341
rect 1584 1307 1611 1340
rect 1660 1307 1683 1340
rect 1645 1306 1683 1307
rect 710 1239 986 1273
rect 1020 1239 1058 1273
rect 710 1237 1056 1239
rect 710 1203 816 1237
rect 415 1187 453 1203
rect 415 1169 433 1187
rect 589 1187 623 1203
rect 433 1119 467 1153
rect 433 1051 467 1085
rect 744 1187 782 1203
rect 744 1169 745 1187
rect 589 1119 623 1153
rect 589 1056 623 1085
rect 779 1169 782 1187
rect 901 1187 935 1203
rect 745 1119 779 1153
rect 587 1051 625 1056
rect 587 1022 589 1051
rect 433 983 467 1017
rect 433 915 467 949
rect 433 847 467 881
rect 433 779 467 813
rect 433 711 467 745
rect 433 661 467 677
rect 623 1022 625 1051
rect 745 1051 779 1085
rect 901 1119 935 1153
rect 1057 1187 1091 1203
rect 1057 1131 1091 1153
rect 1213 1187 1247 1203
rect 1055 1119 1093 1131
rect 1055 1097 1057 1119
rect 901 1056 935 1085
rect 1091 1097 1093 1119
rect 1213 1119 1247 1153
rect 1369 1187 1403 1203
rect 1369 1131 1403 1153
rect 1493 1187 1527 1203
rect 589 983 623 1017
rect 589 915 623 949
rect 589 847 623 881
rect 589 779 623 813
rect 589 711 623 745
rect 589 661 623 677
rect 897 1051 935 1056
rect 897 1022 901 1051
rect 745 983 779 1017
rect 745 915 779 949
rect 745 847 779 881
rect 745 779 779 813
rect 745 711 779 745
rect 745 661 779 677
rect 1057 1051 1091 1085
rect 1369 1119 1407 1131
rect 1213 1056 1247 1085
rect 1403 1097 1407 1119
rect 1493 1119 1527 1153
rect 901 983 935 1017
rect 901 915 935 949
rect 901 847 935 881
rect 901 779 935 813
rect 901 711 935 745
rect 901 661 935 677
rect 1207 1051 1245 1056
rect 1207 1022 1213 1051
rect 1369 1051 1403 1085
rect 1493 1056 1527 1085
rect 1649 1187 1683 1203
rect 1649 1119 1683 1153
rect 1057 983 1091 1017
rect 1057 915 1091 949
rect 1057 847 1091 881
rect 1057 779 1091 813
rect 1057 711 1091 745
rect 1057 661 1091 677
rect 1213 983 1247 1017
rect 1213 915 1247 949
rect 1213 847 1247 881
rect 1213 779 1247 813
rect 1213 711 1247 745
rect 1213 661 1247 677
rect 1491 1051 1529 1056
rect 1491 1022 1493 1051
rect 1369 983 1403 1017
rect 1369 915 1403 949
rect 1369 847 1403 881
rect 1369 779 1403 813
rect 1369 711 1403 745
rect 1369 661 1403 677
rect 1527 1022 1529 1051
rect 1649 1051 1683 1085
rect 1493 983 1527 1017
rect 1493 915 1527 949
rect 1493 847 1527 881
rect 1493 779 1527 813
rect 1493 711 1527 745
rect 1493 661 1527 677
rect 1649 983 1683 1017
rect 1649 915 1683 949
rect 1649 847 1683 881
rect 1649 779 1683 813
rect 1649 730 1683 745
rect 1649 711 1652 730
rect 1683 677 1686 696
rect 1649 661 1686 677
rect 1652 658 1686 661
rect 467 555 491 589
rect 525 555 563 589
rect 597 555 635 589
rect 669 555 707 589
rect 741 555 779 589
rect 813 555 851 589
rect 885 555 923 589
rect 957 587 995 589
rect 957 555 994 587
rect 1029 555 1067 589
rect 1101 587 1139 589
rect 1173 587 1211 589
rect 1245 587 1283 589
rect 1317 587 1354 589
rect 1388 587 1425 589
rect 1459 587 1496 589
rect 1530 587 1567 589
rect 1601 587 1625 589
rect 1102 555 1139 587
rect 1176 555 1211 587
rect 1250 555 1283 587
rect 1324 555 1354 587
rect 1398 555 1425 587
rect 1472 555 1496 587
rect 1546 555 1567 587
rect 1620 555 1625 587
rect 1028 553 1068 555
rect 1102 553 1142 555
rect 1176 553 1216 555
rect 1250 553 1290 555
rect 1324 553 1364 555
rect 1398 553 1438 555
rect 1472 553 1512 555
rect 1546 553 1586 555
<< viali >>
rect 252 3393 262 3427
rect 262 3393 286 3427
rect 328 3393 334 3427
rect 334 3393 362 3427
rect 404 3393 406 3427
rect 406 3393 438 3427
rect 480 3393 512 3427
rect 512 3393 514 3427
rect 556 3393 583 3427
rect 583 3393 590 3427
rect 632 3393 654 3427
rect 654 3393 666 3427
rect 708 3393 725 3427
rect 725 3393 742 3427
rect 784 3393 796 3427
rect 796 3393 818 3427
rect 860 3393 867 3427
rect 867 3393 894 3427
rect 936 3393 938 3427
rect 938 3393 970 3427
rect 1012 3393 1046 3427
rect 1088 3393 1117 3427
rect 1117 3393 1122 3427
rect 1164 3393 1188 3427
rect 1188 3393 1198 3427
rect 1240 3393 1259 3427
rect 1259 3393 1274 3427
rect 1315 3393 1330 3427
rect 1330 3393 1349 3427
rect 1390 3393 1401 3427
rect 1401 3393 1424 3427
rect 1465 3393 1472 3427
rect 1472 3393 1499 3427
rect 1540 3393 1543 3427
rect 1543 3393 1574 3427
rect 246 3307 280 3336
rect 246 3302 280 3307
rect 246 3239 280 3264
rect 246 3230 280 3239
rect 402 3137 436 3163
rect 402 3129 436 3137
rect 402 3069 436 3091
rect 402 3057 436 3069
rect 558 3307 592 3336
rect 558 3302 592 3307
rect 838 3302 872 3336
rect 558 3239 592 3264
rect 558 3230 592 3239
rect 681 3133 715 3139
rect 681 3105 682 3133
rect 682 3105 715 3133
rect 681 3065 715 3067
rect 681 3033 682 3065
rect 682 3033 715 3065
rect 1531 3302 1565 3336
rect 838 3235 872 3264
rect 838 3230 872 3235
rect 761 3020 795 3054
rect 920 3020 954 3054
rect 386 2971 420 2976
rect 386 2942 402 2971
rect 402 2942 420 2971
rect 458 2942 492 2976
rect 761 2971 795 2982
rect 1531 3247 1565 3264
rect 1531 3230 1565 3247
rect 1401 3150 1435 3184
rect 1473 3153 1504 3184
rect 1504 3153 1507 3184
rect 1473 3150 1507 3153
rect 1167 3076 1201 3110
rect 1239 3076 1273 3110
rect 1820 3150 1854 3184
rect 1892 3150 1926 3184
rect 1006 3031 1028 3036
rect 1028 3031 1040 3036
rect 1006 3002 1040 3031
rect 1078 3002 1112 3036
rect 761 2948 777 2971
rect 777 2948 795 2971
rect 920 2968 954 2982
rect 920 2948 933 2968
rect 933 2948 954 2968
rect 1564 1978 1598 2012
rect 1639 1978 1673 2012
rect 1713 1978 1747 2012
rect 1787 1978 1821 2012
rect 1861 1978 1895 2012
rect 1935 1978 1969 2012
rect 2009 1978 2043 2012
rect 2083 1978 2117 2012
rect 2157 1978 2191 2012
rect 2231 1978 2265 2012
rect 2305 1978 2339 2012
rect 2379 1978 2413 2012
rect 2453 1978 2487 2012
rect 2527 1978 2561 2012
rect 2601 1978 2635 2012
rect 2675 1978 2709 2012
rect 2749 1978 2783 2012
rect 2823 1978 2857 2012
rect 2897 1978 2931 2012
rect 2971 1978 3005 2012
rect 3045 1978 3079 2012
rect 3119 1978 3153 2012
rect 3193 1978 3227 2012
rect 3267 1978 3301 2012
rect 3341 1978 3375 2012
rect 3415 1978 3449 2012
rect 3489 1978 3523 2012
rect 3563 1978 3597 2012
rect 3637 1978 3671 2012
rect 3711 1978 3745 2012
rect 3785 1978 3819 2012
rect 3859 1978 3893 2012
rect 3933 1978 3967 2012
rect 4007 1978 4041 2012
rect 1122 1924 1156 1958
rect 1196 1924 1230 1958
rect 1270 1924 1304 1958
rect 1344 1924 1378 1958
rect 1418 1924 1452 1958
rect 939 1725 973 1759
rect 585 1689 619 1691
rect 585 1657 589 1689
rect 589 1657 619 1689
rect 585 1587 589 1619
rect 589 1587 619 1619
rect 585 1585 619 1587
rect 507 1486 541 1520
rect 709 1649 743 1658
rect 709 1624 743 1649
rect 709 1581 743 1586
rect 709 1552 743 1581
rect 864 1581 865 1601
rect 865 1581 898 1601
rect 864 1567 898 1581
rect 864 1513 865 1529
rect 865 1513 898 1529
rect 864 1495 898 1513
rect 939 1653 973 1687
rect 507 1415 514 1448
rect 514 1415 541 1448
rect 727 1426 737 1448
rect 737 1426 761 1448
rect 799 1426 805 1448
rect 805 1426 833 1448
rect 1021 1725 1055 1759
rect 1021 1683 1055 1687
rect 1021 1653 1055 1683
rect 1145 1581 1179 1601
rect 1145 1567 1179 1581
rect 1145 1513 1179 1529
rect 1145 1495 1179 1513
rect 1301 1615 1335 1618
rect 1301 1584 1335 1615
rect 1301 1513 1335 1546
rect 1301 1512 1335 1513
rect 507 1414 541 1415
rect 727 1414 761 1426
rect 799 1414 833 1426
rect 929 1425 956 1448
rect 956 1425 963 1448
rect 1001 1425 1024 1448
rect 1024 1425 1035 1448
rect 929 1414 963 1425
rect 1001 1414 1035 1425
rect 1307 1419 1341 1453
rect 1379 1419 1413 1453
rect 492 1341 526 1342
rect 564 1341 598 1342
rect 1313 1341 1347 1342
rect 492 1308 494 1341
rect 494 1308 526 1341
rect 564 1308 598 1341
rect 1313 1308 1342 1341
rect 1342 1308 1347 1341
rect 1385 1308 1419 1342
rect 1611 1307 1626 1340
rect 1626 1307 1645 1340
rect 1611 1306 1645 1307
rect 1683 1306 1717 1340
rect 986 1239 1020 1273
rect 1058 1239 1092 1273
rect 381 1169 415 1203
rect 453 1187 487 1203
rect 453 1169 467 1187
rect 467 1169 487 1187
rect 710 1169 744 1203
rect 782 1169 816 1203
rect 553 1022 587 1056
rect 625 1022 659 1056
rect 1021 1097 1055 1131
rect 1093 1097 1127 1131
rect 863 1022 897 1056
rect 935 1022 969 1056
rect 1335 1097 1369 1131
rect 1407 1097 1441 1131
rect 1173 1022 1207 1056
rect 1245 1051 1279 1056
rect 1245 1022 1247 1051
rect 1247 1022 1279 1051
rect 1457 1022 1491 1056
rect 1529 1022 1563 1056
rect 1652 711 1686 730
rect 1652 696 1683 711
rect 1683 696 1686 711
rect 1652 624 1686 658
rect 994 555 995 587
rect 995 555 1028 587
rect 1068 555 1101 587
rect 1101 555 1102 587
rect 1142 555 1173 587
rect 1173 555 1176 587
rect 1216 555 1245 587
rect 1245 555 1250 587
rect 1290 555 1317 587
rect 1317 555 1324 587
rect 1364 555 1388 587
rect 1388 555 1398 587
rect 1438 555 1459 587
rect 1459 555 1472 587
rect 1512 555 1530 587
rect 1530 555 1546 587
rect 1586 555 1601 587
rect 1601 555 1620 587
rect 994 553 1028 555
rect 1068 553 1102 555
rect 1142 553 1176 555
rect 1216 553 1250 555
rect 1290 553 1324 555
rect 1364 553 1398 555
rect 1438 553 1472 555
rect 1512 553 1546 555
rect 1586 553 1620 555
<< metal1 >>
rect 196 3427 1586 3433
rect 196 3393 252 3427
rect 286 3393 328 3427
rect 362 3393 404 3427
rect 438 3393 480 3427
rect 514 3393 556 3427
rect 590 3393 632 3427
rect 666 3393 708 3427
rect 742 3393 784 3427
rect 818 3393 860 3427
rect 894 3393 936 3427
rect 970 3393 1012 3427
rect 1046 3393 1088 3427
rect 1122 3393 1164 3427
rect 1198 3393 1240 3427
rect 1274 3393 1315 3427
rect 1349 3393 1390 3427
rect 1424 3393 1465 3427
rect 1499 3393 1540 3427
rect 1574 3393 1586 3427
rect 196 3336 1586 3393
rect 196 3302 246 3336
rect 280 3302 558 3336
rect 592 3302 838 3336
rect 872 3302 1531 3336
rect 1565 3302 1586 3336
rect 196 3264 1586 3302
rect 196 3230 246 3264
rect 280 3230 558 3264
rect 592 3230 838 3264
rect 872 3230 1531 3264
rect 1565 3230 1586 3264
rect 196 3218 1586 3230
rect 755 3184 1938 3190
rect 396 3163 442 3175
rect 396 3129 402 3163
rect 436 3139 442 3163
tri 442 3139 451 3148 sw
rect 675 3139 721 3151
rect 436 3129 451 3139
rect 396 3105 451 3129
tri 451 3105 485 3139 sw
rect 675 3105 681 3139
rect 715 3105 721 3139
rect 396 3091 485 3105
rect 396 3057 402 3091
rect 436 3088 485 3091
tri 485 3088 502 3105 sw
rect 436 3057 625 3088
rect 396 3045 625 3057
tri 545 3033 557 3045 ne
rect 557 3033 625 3045
tri 557 3020 570 3033 ne
rect 570 3020 625 3033
tri 570 3011 579 3020 ne
rect 374 2976 504 2982
rect 374 2942 386 2976
rect 420 2942 458 2976
rect 492 2942 504 2976
rect 374 2936 504 2942
tri 424 2902 458 2936 ne
rect 458 2629 504 2936
tri 504 2629 547 2672 sw
rect 458 2583 547 2629
tri 458 2540 501 2583 ne
tri 495 2413 501 2419 ne
rect 501 1520 547 2583
rect 579 1691 625 3020
rect 675 3067 721 3105
rect 675 3033 681 3067
rect 715 3033 721 3067
rect 675 2736 721 3033
rect 755 3150 1401 3184
rect 1435 3150 1473 3184
rect 1507 3150 1820 3184
rect 1854 3150 1892 3184
rect 1926 3150 1938 3184
rect 755 3144 1938 3150
rect 755 3054 801 3144
tri 801 3110 835 3144 nw
rect 914 3110 1285 3116
rect 755 3020 761 3054
rect 795 3020 801 3054
rect 755 2982 801 3020
rect 755 2948 761 2982
rect 795 2948 801 2982
rect 755 2864 801 2948
rect 914 3076 1167 3110
rect 1201 3076 1239 3110
rect 1273 3076 1285 3110
rect 914 3073 1285 3076
rect 914 3070 982 3073
tri 982 3070 985 3073 nw
tri 1152 3070 1155 3073 ne
rect 1155 3070 1285 3073
rect 914 3066 978 3070
tri 978 3066 982 3070 nw
rect 914 3054 960 3066
rect 914 3020 920 3054
rect 954 3020 960 3054
tri 960 3048 978 3066 nw
rect 914 2982 960 3020
rect 994 3036 1124 3042
rect 994 3002 1006 3036
rect 1040 3002 1078 3036
rect 1112 3002 1124 3036
rect 994 2996 1124 3002
tri 994 2992 998 2996 ne
rect 998 2992 1120 2996
tri 1120 2992 1124 2996 nw
rect 914 2948 920 2982
rect 954 2948 960 2982
tri 801 2864 827 2890 sw
rect 755 2818 827 2864
tri 755 2792 781 2818 ne
tri 721 2736 749 2764 sw
rect 675 2690 749 2736
tri 675 2662 703 2690 ne
tri 697 2602 703 2608 ne
tri 625 2375 631 2381 sw
tri 625 2241 631 2247 nw
rect 579 1657 585 1691
rect 619 1657 625 1691
rect 579 1619 625 1657
rect 579 1585 585 1619
rect 619 1585 625 1619
rect 579 1573 625 1585
rect 703 1658 749 2690
rect 703 1624 709 1658
rect 743 1624 749 1658
rect 703 1586 749 1624
rect 703 1552 709 1586
rect 743 1552 749 1586
rect 703 1540 749 1552
rect 501 1486 507 1520
rect 541 1486 547 1520
rect 501 1448 547 1486
rect 781 1454 827 2818
rect 914 1771 960 2948
rect 998 1884 1032 2992
tri 1032 2904 1120 2992 nw
rect 1486 2012 4053 2018
rect 1486 1978 1564 2012
rect 1598 1978 1639 2012
rect 1673 1978 1713 2012
rect 1747 1978 1787 2012
rect 1821 1978 1861 2012
rect 1895 1978 1935 2012
rect 1969 1978 2009 2012
rect 2043 1978 2083 2012
rect 2117 1978 2157 2012
rect 2191 1978 2231 2012
rect 2265 1978 2305 2012
rect 2339 1978 2379 2012
rect 2413 1978 2453 2012
rect 2487 1978 2527 2012
rect 2561 1978 2601 2012
rect 2635 1978 2675 2012
rect 2709 1978 2749 2012
rect 2783 1978 2823 2012
rect 2857 1978 2897 2012
rect 2931 1978 2971 2012
rect 3005 1978 3045 2012
rect 3079 1978 3119 2012
rect 3153 1978 3193 2012
rect 3227 1978 3267 2012
rect 3301 1978 3341 2012
rect 3375 1978 3415 2012
rect 3449 1978 3489 2012
rect 3523 1978 3563 2012
rect 3597 1978 3637 2012
rect 3671 1978 3711 2012
rect 3745 1978 3785 2012
rect 3819 1978 3859 2012
rect 3893 1978 3933 2012
rect 3967 1978 4007 2012
rect 4041 1978 4053 2012
rect 1486 1972 4053 1978
rect 1486 1964 1532 1972
rect 1110 1958 1532 1964
rect 1110 1924 1122 1958
rect 1156 1924 1196 1958
rect 1230 1924 1270 1958
rect 1304 1924 1344 1958
rect 1378 1924 1418 1958
rect 1452 1924 1532 1958
rect 1110 1918 1532 1924
tri 1032 1884 1056 1908 sw
rect 998 1856 1056 1884
tri 1056 1856 1084 1884 sw
rect 998 1850 1061 1856
tri 998 1833 1015 1850 ne
tri 960 1771 979 1790 sw
rect 914 1759 979 1771
rect 914 1725 939 1759
rect 973 1725 979 1759
rect 914 1687 979 1725
rect 914 1653 939 1687
rect 973 1653 979 1687
rect 914 1641 979 1653
rect 1015 1759 1061 1850
tri 1061 1777 1108 1824 nw
rect 1015 1725 1021 1759
rect 1055 1725 1061 1759
rect 1015 1687 1061 1725
rect 1015 1653 1021 1687
rect 1055 1653 1061 1687
rect 1015 1641 1061 1653
rect 1221 1618 1341 1630
rect 858 1601 1185 1613
rect 858 1567 864 1601
rect 898 1567 1145 1601
rect 1179 1567 1185 1601
rect 858 1529 1185 1567
rect 858 1495 864 1529
rect 898 1495 1145 1529
rect 1179 1495 1185 1529
rect 858 1483 1185 1495
rect 1221 1584 1301 1618
rect 1335 1584 1341 1618
rect 1221 1546 1341 1584
rect 1221 1512 1301 1546
rect 1335 1512 1341 1546
rect 1221 1500 1341 1512
rect 501 1414 507 1448
rect 541 1414 547 1448
rect 501 1402 547 1414
rect 715 1448 845 1454
rect 715 1414 727 1448
rect 761 1414 799 1448
rect 833 1414 845 1448
rect 715 1408 845 1414
rect 917 1448 1047 1454
rect 917 1414 929 1448
rect 963 1414 1001 1448
rect 1035 1414 1047 1448
rect 917 1408 1047 1414
rect 480 1342 610 1348
rect 480 1308 492 1342
rect 526 1308 564 1342
rect 598 1308 610 1342
rect 480 1302 610 1308
rect 773 1308 819 1408
tri 940 1374 974 1408 ne
tri 819 1308 850 1339 sw
rect 974 1308 1030 1408
tri 1030 1391 1047 1408 nw
tri 1030 1308 1035 1313 sw
rect 773 1306 850 1308
tri 850 1306 852 1308 sw
rect 974 1306 1035 1308
tri 1035 1306 1037 1308 sw
rect 773 1305 852 1306
tri 852 1305 853 1306 sw
rect 974 1305 1037 1306
tri 1037 1305 1038 1306 sw
rect 773 1259 937 1305
tri 857 1239 877 1259 ne
rect 877 1239 937 1259
tri 877 1225 891 1239 ne
rect 369 1203 835 1209
rect 369 1169 381 1203
rect 415 1169 453 1203
rect 487 1169 710 1203
rect 744 1169 782 1203
rect 816 1169 835 1203
rect 369 1163 835 1169
rect 891 1137 937 1239
rect 974 1279 1038 1305
tri 1038 1279 1064 1305 sw
rect 974 1273 1104 1279
rect 974 1239 986 1273
rect 1020 1239 1058 1273
rect 1092 1239 1104 1273
rect 974 1233 1104 1239
tri 937 1137 971 1171 sw
rect 1221 1137 1267 1500
rect 1295 1453 1425 1459
rect 1295 1419 1307 1453
rect 1341 1419 1379 1453
rect 1413 1419 1425 1453
rect 1295 1413 1425 1419
rect 1301 1342 1431 1348
rect 1301 1308 1313 1342
rect 1347 1308 1385 1342
rect 1419 1308 1431 1342
rect 1301 1302 1431 1308
rect 1599 1340 1729 1346
rect 1599 1306 1611 1340
rect 1645 1306 1683 1340
rect 1717 1306 1729 1340
rect 1599 1300 1729 1306
rect 891 1131 1453 1137
rect 891 1097 1021 1131
rect 1055 1097 1093 1131
rect 1127 1097 1335 1131
rect 1369 1097 1407 1131
rect 1441 1097 1453 1131
rect 891 1091 1453 1097
rect 541 1056 1575 1062
rect 541 1022 553 1056
rect 587 1022 625 1056
rect 659 1022 863 1056
rect 897 1022 935 1056
rect 969 1022 1173 1056
rect 1207 1022 1245 1056
rect 1279 1022 1457 1056
rect 1491 1022 1529 1056
rect 1563 1022 1575 1056
rect 541 1016 1575 1022
rect 1634 730 1704 742
rect 1634 696 1652 730
rect 1686 696 1704 730
rect 1634 658 1704 696
rect 1634 624 1652 658
rect 1686 624 1704 658
rect 1634 613 1704 624
rect 1646 612 1692 613
rect 982 587 1632 593
rect 982 553 994 587
rect 1028 553 1068 587
rect 1102 553 1142 587
rect 1176 553 1216 587
rect 1250 553 1290 587
rect 1324 553 1364 587
rect 1398 553 1438 587
rect 1472 553 1512 587
rect 1546 553 1586 587
rect 1620 553 1632 587
rect 982 547 1632 553
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808587  sky130_fd_pr__model__nfet_highvoltage__example_55959141808587_0
timestamp 1649977179
transform 1 0 478 0 -1 1701
box -28 0 128 97
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808588  sky130_fd_pr__model__pfet_highvoltage__example_55959141808588_0
timestamp 1649977179
transform 1 0 291 0 -1 3319
box -28 0 128 131
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808588  sky130_fd_pr__model__pfet_highvoltage__example_55959141808588_1
timestamp 1649977179
transform 1 0 447 0 -1 3319
box -28 0 128 131
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_0
timestamp 1649977179
transform 1 0 946 0 1 665
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_1
timestamp 1649977179
transform -1 0 890 0 1 665
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_0
timestamp 1649977179
transform 1 0 1190 0 1 1501
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_1
timestamp 1649977179
transform 1 0 910 0 1 1501
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_2
timestamp 1649977179
transform -1 0 854 0 1 1501
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808589  sky130_fd_pr__nfet_01v8__example_55959141808589_0
timestamp 1649977179
transform -1 0 1638 0 1 665
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_0
timestamp 1649977179
transform 1 0 883 0 1 3019
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_1
timestamp 1649977179
transform -1 0 827 0 1 3019
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1649977179
transform -1 0 1520 0 1 3235
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1649977179
transform 1 0 1576 0 1 3235
box -28 0 228 29
<< labels >>
flabel metal1 s 1340 1313 1368 1341 3 FreeSans 520 0 0 0 IN_B
port 1 nsew
flabel metal1 s 518 1314 546 1342 3 FreeSans 520 0 0 0 IN
port 2 nsew
flabel metal1 s 1338 1420 1366 1448 3 FreeSans 520 0 0 0 RST_H
port 3 nsew
flabel metal1 s 712 1584 740 1612 3 FreeSans 520 0 0 0 OUT_H_N
port 4 nsew
flabel metal1 s 1024 1667 1052 1695 3 FreeSans 520 0 0 0 OUT_H
port 5 nsew
flabel metal1 s 941 3275 969 3303 3 FreeSans 520 0 0 0 VPWR_HV
port 6 nsew
flabel metal1 s 1630 1310 1658 1338 3 FreeSans 520 0 0 0 HLD_H
port 7 nsew
flabel metal1 s 968 1534 996 1562 3 FreeSans 520 0 0 0 VGND
port 8 nsew
flabel metal1 s 1664 668 1692 696 3 FreeSans 520 0 0 0 VGND
port 8 nsew
<< properties >>
string GDS_END 8439222
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8412112
<< end >>
