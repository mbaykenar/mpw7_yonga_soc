magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 222 582
<< pwell >>
rect 3 38 181 195
<< psubdiff >>
rect 29 145 155 169
rect 63 111 121 145
rect 29 64 155 111
<< nsubdiff >>
rect 29 447 155 480
rect 63 413 121 447
rect 29 363 155 413
rect 63 329 121 363
rect 29 305 155 329
<< psubdiffcont >>
rect 29 111 63 145
rect 121 111 155 145
<< nsubdiffcont >>
rect 29 413 63 447
rect 121 413 155 447
rect 29 329 63 363
rect 121 329 155 363
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 17 447 167 491
rect 17 413 29 447
rect 63 413 121 447
rect 155 413 167 447
rect 17 363 167 413
rect 17 329 29 363
rect 63 329 121 363
rect 155 329 167 363
rect 17 294 167 329
rect 17 145 167 162
rect 17 111 29 145
rect 63 111 121 145
rect 155 111 167 145
rect 17 53 167 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 29 -17 63 17
rect 121 -17 155 17
<< metal1 >>
rect 0 561 184 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 0 496 184 527
rect 0 17 184 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
rect 0 -48 184 -17
<< labels >>
flabel metal1 s 19 -14 67 12 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 21 533 75 555 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
flabel locali s 35 431 60 456 0 FreeSans 250 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 120 92 155 122 0 FreeSans 250 0 0 0 VNB
port 2 nsew ground bidirectional
flabel locali s 128 425 150 454 0 FreeSans 250 0 0 0 VPB
port 3 nsew power bidirectional
rlabel comment s 0 0 0 0 4 tap_2
rlabel metal1 s 0 -48 184 48 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 496 184 592 1 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 184 544
string GDS_END 513316
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 511064
string LEFclass CORE WELLTAP
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 0.920 0.000 
<< end >>
