magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 17 21 707 203
rect 29 -17 63 21
<< scnmos >>
rect 95 47 125 177
rect 192 93 222 177
rect 418 47 448 177
rect 514 47 544 177
rect 598 47 628 177
<< scpmoshvt >>
rect 79 297 109 497
rect 192 297 222 381
rect 418 297 448 497
rect 514 297 544 497
rect 586 297 616 497
<< ndiff >>
rect 43 149 95 177
rect 43 115 51 149
rect 85 115 95 149
rect 43 47 95 115
rect 125 149 192 177
rect 125 115 142 149
rect 176 115 192 149
rect 125 93 192 115
rect 222 149 274 177
rect 222 115 232 149
rect 266 115 274 149
rect 222 93 274 115
rect 366 131 418 177
rect 366 97 374 131
rect 408 97 418 131
rect 125 47 177 93
rect 366 47 418 97
rect 448 163 514 177
rect 448 129 470 163
rect 504 129 514 163
rect 448 95 514 129
rect 448 61 470 95
rect 504 61 514 95
rect 448 47 514 61
rect 544 95 598 177
rect 544 61 554 95
rect 588 61 598 95
rect 544 47 598 61
rect 628 163 681 177
rect 628 129 638 163
rect 672 129 681 163
rect 628 95 681 129
rect 628 61 638 95
rect 672 61 681 95
rect 628 47 681 61
<< pdiff >>
rect 27 482 79 497
rect 27 448 35 482
rect 69 448 79 482
rect 27 414 79 448
rect 27 380 35 414
rect 69 380 79 414
rect 27 346 79 380
rect 27 312 35 346
rect 69 312 79 346
rect 27 297 79 312
rect 109 475 177 497
rect 109 441 135 475
rect 169 441 177 475
rect 109 381 177 441
rect 358 477 418 497
rect 358 443 366 477
rect 400 443 418 477
rect 109 297 192 381
rect 222 339 278 381
rect 222 305 232 339
rect 266 305 278 339
rect 222 297 278 305
rect 358 297 418 443
rect 448 477 514 497
rect 448 443 470 477
rect 504 443 514 477
rect 448 409 514 443
rect 448 375 470 409
rect 504 375 514 409
rect 448 341 514 375
rect 448 307 470 341
rect 504 307 514 341
rect 448 297 514 307
rect 544 297 586 497
rect 616 477 672 497
rect 616 443 626 477
rect 660 443 672 477
rect 616 409 672 443
rect 616 375 626 409
rect 660 375 672 409
rect 616 341 672 375
rect 616 307 626 341
rect 660 307 672 341
rect 616 297 672 307
<< ndiffc >>
rect 51 115 85 149
rect 142 115 176 149
rect 232 115 266 149
rect 374 97 408 131
rect 470 129 504 163
rect 470 61 504 95
rect 554 61 588 95
rect 638 129 672 163
rect 638 61 672 95
<< pdiffc >>
rect 35 448 69 482
rect 35 380 69 414
rect 35 312 69 346
rect 135 441 169 475
rect 366 443 400 477
rect 232 305 266 339
rect 470 443 504 477
rect 470 375 504 409
rect 470 307 504 341
rect 626 443 660 477
rect 626 375 660 409
rect 626 307 660 341
<< poly >>
rect 79 497 109 523
rect 418 497 448 523
rect 514 497 544 523
rect 586 497 616 523
rect 192 381 222 407
rect 79 265 109 297
rect 192 265 222 297
rect 418 265 448 297
rect 514 265 544 297
rect 79 249 146 265
rect 79 215 102 249
rect 136 215 146 249
rect 79 199 146 215
rect 192 249 254 265
rect 192 215 210 249
rect 244 215 254 249
rect 192 199 254 215
rect 296 249 448 265
rect 296 215 306 249
rect 340 215 448 249
rect 296 199 448 215
rect 490 249 544 265
rect 490 215 500 249
rect 534 215 544 249
rect 490 199 544 215
rect 586 265 616 297
rect 586 249 656 265
rect 586 215 606 249
rect 640 215 656 249
rect 586 199 656 215
rect 95 177 125 199
rect 192 177 222 199
rect 418 177 448 199
rect 514 177 544 199
rect 598 177 628 199
rect 192 67 222 93
rect 95 21 125 47
rect 418 21 448 47
rect 514 21 544 47
rect 598 21 628 47
<< polycont >>
rect 102 215 136 249
rect 210 215 244 249
rect 306 215 340 249
rect 500 215 534 249
rect 606 215 640 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 482 85 493
rect 17 448 35 482
rect 69 448 85 482
rect 17 414 85 448
rect 119 475 201 527
rect 119 441 135 475
rect 169 441 201 475
rect 350 477 416 527
rect 350 443 366 477
rect 400 443 416 477
rect 450 477 515 493
rect 450 443 470 477
rect 504 443 515 477
rect 17 380 35 414
rect 69 380 85 414
rect 450 409 515 443
rect 450 407 470 409
rect 17 346 85 380
rect 17 312 35 346
rect 69 312 85 346
rect 17 296 85 312
rect 119 375 470 407
rect 504 375 515 409
rect 119 373 515 375
rect 17 165 68 296
rect 119 265 172 373
rect 374 341 515 373
rect 215 305 232 339
rect 266 305 340 339
rect 102 249 172 265
rect 136 215 172 249
rect 102 199 172 215
rect 206 249 272 265
rect 206 215 210 249
rect 244 215 272 249
rect 206 199 272 215
rect 306 249 340 305
rect 306 165 340 215
rect 17 149 89 165
rect 17 115 51 149
rect 85 115 89 149
rect 17 90 89 115
rect 142 149 176 165
rect 142 17 176 115
rect 232 149 340 165
rect 266 131 340 149
rect 374 307 470 341
rect 504 307 515 341
rect 610 477 676 527
rect 610 443 626 477
rect 660 443 676 477
rect 610 409 676 443
rect 610 375 626 409
rect 660 375 676 409
rect 610 341 676 375
rect 610 307 626 341
rect 660 307 676 341
rect 374 291 515 307
rect 374 131 408 291
rect 442 249 556 257
rect 442 215 500 249
rect 534 215 556 249
rect 590 249 719 257
rect 590 215 606 249
rect 640 215 719 249
rect 232 90 266 115
rect 374 51 408 97
rect 454 163 688 181
rect 454 129 470 163
rect 504 147 638 163
rect 504 129 520 147
rect 454 95 520 129
rect 622 129 638 147
rect 672 129 688 163
rect 454 61 470 95
rect 504 61 520 95
rect 454 51 520 61
rect 554 95 588 111
rect 554 17 588 61
rect 622 95 688 129
rect 622 61 638 95
rect 672 61 688 95
rect 622 54 688 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 425 63 459 0 FreeSans 400 0 0 0 X
port 8 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o21ba_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1332384
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1326280
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.680 0.000 
<< end >>
