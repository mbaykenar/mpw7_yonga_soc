magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 5 21 735 203
rect 29 -17 63 21
rect 395 -13 429 21
<< scnmos >>
rect 179 47 209 177
rect 286 47 316 177
rect 390 47 420 177
rect 538 47 568 177
rect 620 47 650 177
<< scpmoshvt >>
rect 187 297 217 497
rect 286 297 316 497
rect 390 297 420 497
rect 536 297 566 497
rect 621 297 651 497
<< ndiff >>
rect 31 89 179 177
rect 31 55 79 89
rect 113 55 179 89
rect 31 47 179 55
rect 209 163 286 177
rect 209 129 224 163
rect 258 129 286 163
rect 209 95 286 129
rect 209 61 225 95
rect 259 61 286 95
rect 209 47 286 61
rect 316 91 390 177
rect 316 57 326 91
rect 360 57 390 91
rect 316 47 390 57
rect 420 163 538 177
rect 420 129 434 163
rect 468 129 538 163
rect 420 95 538 129
rect 420 61 434 95
rect 468 61 538 95
rect 420 47 538 61
rect 568 47 620 177
rect 650 112 709 177
rect 650 78 662 112
rect 696 78 709 112
rect 650 47 709 78
<< pdiff >>
rect 36 476 187 497
rect 36 442 72 476
rect 106 442 187 476
rect 36 408 187 442
rect 36 374 72 408
rect 106 374 187 408
rect 36 339 187 374
rect 36 305 72 339
rect 106 305 187 339
rect 36 297 187 305
rect 217 297 286 497
rect 316 297 390 497
rect 420 453 536 497
rect 420 419 491 453
rect 525 419 536 453
rect 420 385 536 419
rect 420 351 491 385
rect 525 351 536 385
rect 420 297 536 351
rect 566 486 621 497
rect 566 452 576 486
rect 610 452 621 486
rect 566 418 621 452
rect 566 384 576 418
rect 610 384 621 418
rect 566 297 621 384
rect 651 463 709 497
rect 651 429 662 463
rect 696 429 709 463
rect 651 395 709 429
rect 651 361 662 395
rect 696 361 709 395
rect 651 297 709 361
<< ndiffc >>
rect 79 55 113 89
rect 224 129 258 163
rect 225 61 259 95
rect 326 57 360 91
rect 434 129 468 163
rect 434 61 468 95
rect 662 78 696 112
<< pdiffc >>
rect 72 442 106 476
rect 72 374 106 408
rect 72 305 106 339
rect 491 419 525 453
rect 491 351 525 385
rect 576 452 610 486
rect 576 384 610 418
rect 662 429 696 463
rect 662 361 696 395
<< poly >>
rect 187 497 217 523
rect 286 497 316 523
rect 390 497 420 523
rect 536 497 566 523
rect 621 497 651 523
rect 187 265 217 297
rect 157 249 217 265
rect 157 215 173 249
rect 207 215 217 249
rect 157 199 217 215
rect 286 276 316 297
rect 286 249 348 276
rect 286 215 304 249
rect 338 215 348 249
rect 179 177 209 199
rect 286 194 348 215
rect 390 266 420 297
rect 390 249 449 266
rect 536 264 566 297
rect 621 265 651 297
rect 390 215 404 249
rect 438 215 449 249
rect 286 177 316 194
rect 390 192 449 215
rect 491 253 566 264
rect 491 249 568 253
rect 491 215 507 249
rect 541 215 568 249
rect 491 193 568 215
rect 390 177 420 192
rect 538 177 568 193
rect 620 249 688 265
rect 620 215 635 249
rect 669 215 688 249
rect 620 193 688 215
rect 620 177 650 193
rect 179 21 209 47
rect 286 21 316 47
rect 390 21 420 47
rect 538 21 568 47
rect 620 21 650 47
<< polycont >>
rect 173 215 207 249
rect 304 215 338 249
rect 404 215 438 249
rect 507 215 541 249
rect 635 215 669 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 29 476 106 492
rect 29 442 72 476
rect 29 408 106 442
rect 29 374 72 408
rect 29 339 106 374
rect 29 305 72 339
rect 29 176 106 305
rect 157 249 247 491
rect 157 215 173 249
rect 207 215 247 249
rect 157 210 247 215
rect 287 249 354 491
rect 287 215 304 249
rect 338 215 354 249
rect 287 210 354 215
rect 388 280 443 491
rect 479 453 525 492
rect 479 419 491 453
rect 479 385 525 419
rect 479 351 491 385
rect 560 486 626 527
rect 560 452 576 486
rect 610 452 626 486
rect 560 418 626 452
rect 560 384 576 418
rect 610 384 626 418
rect 662 463 701 492
rect 696 429 701 463
rect 662 395 701 429
rect 479 350 525 351
rect 696 361 701 395
rect 662 350 701 361
rect 479 316 701 350
rect 388 249 454 280
rect 388 215 404 249
rect 438 215 454 249
rect 388 210 454 215
rect 488 249 545 280
rect 488 215 507 249
rect 541 215 545 249
rect 488 199 545 215
rect 581 249 708 258
rect 581 215 635 249
rect 669 215 708 249
rect 581 204 708 215
rect 29 163 460 176
rect 29 140 224 163
rect 209 129 224 140
rect 258 141 434 163
rect 258 129 275 141
rect 63 89 126 105
rect 63 55 79 89
rect 113 55 126 89
rect 63 17 126 55
rect 209 95 275 129
rect 418 129 434 141
rect 468 129 484 163
rect 209 61 225 95
rect 259 61 275 95
rect 209 52 275 61
rect 310 91 376 107
rect 310 57 326 91
rect 360 57 376 91
rect 418 95 484 129
rect 418 61 434 95
rect 468 61 484 95
rect 581 70 618 204
rect 654 112 702 152
rect 654 78 662 112
rect 696 78 702 112
rect 310 17 376 57
rect 654 17 702 78
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 397 289 431 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 213 425 247 459 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 673 221 707 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 357 247 391 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 305 357 339 391 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 305 425 339 459 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 397 357 431 391 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 397 425 431 459 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 425 63 459 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 581 153 615 187 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 85 615 119 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel pwell s 395 -13 429 20 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111oi_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3791152
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3783370
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 18.400 13.600 
<< end >>
