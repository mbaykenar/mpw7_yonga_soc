magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< pwell >>
rect 15 163 655 817
<< nmoslvt >>
rect 171 189 201 791
rect 257 189 307 791
rect 363 189 413 791
rect 469 189 499 791
<< ndiff >>
rect 111 779 171 791
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 779 257 791
rect 201 513 212 779
rect 246 513 257 779
rect 201 467 257 513
rect 201 201 212 467
rect 246 201 257 467
rect 201 189 257 201
rect 307 779 363 791
rect 307 513 318 779
rect 352 513 363 779
rect 307 467 363 513
rect 307 201 318 467
rect 352 201 363 467
rect 307 189 363 201
rect 413 779 469 791
rect 413 513 424 779
rect 458 513 469 779
rect 413 467 469 513
rect 413 201 424 467
rect 458 201 469 467
rect 413 189 469 201
rect 499 779 559 791
rect 499 745 510 779
rect 544 745 559 779
rect 499 711 559 745
rect 499 677 510 711
rect 544 677 559 711
rect 499 643 559 677
rect 499 609 510 643
rect 544 609 559 643
rect 499 575 559 609
rect 499 541 510 575
rect 544 541 559 575
rect 499 507 559 541
rect 499 473 510 507
rect 544 473 559 507
rect 499 439 559 473
rect 499 405 510 439
rect 544 405 559 439
rect 499 371 559 405
rect 499 337 510 371
rect 544 337 559 371
rect 499 303 559 337
rect 499 269 510 303
rect 544 269 559 303
rect 499 235 559 269
rect 499 201 510 235
rect 544 201 559 235
rect 499 189 559 201
<< ndiffc >>
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 513 246 779
rect 212 201 246 467
rect 318 513 352 779
rect 318 201 352 467
rect 424 513 458 779
rect 424 201 458 467
rect 510 745 544 779
rect 510 677 544 711
rect 510 609 544 643
rect 510 541 544 575
rect 510 473 544 507
rect 510 405 544 439
rect 510 337 544 371
rect 510 269 544 303
rect 510 201 544 235
<< psubdiff >>
rect 41 779 111 791
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 559 779 629 791
rect 559 745 578 779
rect 612 745 629 779
rect 559 711 629 745
rect 559 677 578 711
rect 612 677 629 711
rect 559 643 629 677
rect 559 609 578 643
rect 612 609 629 643
rect 559 575 629 609
rect 559 541 578 575
rect 612 541 629 575
rect 559 507 629 541
rect 559 473 578 507
rect 612 473 629 507
rect 559 439 629 473
rect 559 405 578 439
rect 612 405 629 439
rect 559 371 629 405
rect 559 337 578 371
rect 612 337 629 371
rect 559 303 629 337
rect 559 269 578 303
rect 612 269 629 303
rect 559 235 629 269
rect 559 201 578 235
rect 612 201 629 235
rect 559 189 629 201
<< psubdiffcont >>
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 578 745 612 779
rect 578 677 612 711
rect 578 609 612 643
rect 578 541 612 575
rect 578 473 612 507
rect 578 405 612 439
rect 578 337 612 371
rect 578 269 612 303
rect 578 201 612 235
<< poly >>
rect 243 891 427 907
rect 120 867 201 883
rect 120 833 136 867
rect 170 833 201 867
rect 243 857 264 891
rect 406 857 427 891
rect 243 841 427 857
rect 469 867 550 883
rect 120 817 201 833
rect 171 791 201 817
rect 257 791 307 841
rect 363 791 413 841
rect 469 833 500 867
rect 534 833 550 867
rect 469 817 550 833
rect 469 791 499 817
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 307 189
rect 363 139 413 189
rect 469 163 499 189
rect 469 147 550 163
rect 120 97 201 113
rect 243 123 427 139
rect 243 89 264 123
rect 406 89 427 123
rect 469 113 500 147
rect 534 113 550 147
rect 469 97 550 113
rect 243 73 427 89
<< polycont >>
rect 136 833 170 867
rect 264 857 406 891
rect 500 833 534 867
rect 136 113 170 147
rect 264 89 406 123
rect 500 113 534 147
<< locali >>
rect 248 961 422 980
rect 248 927 276 961
rect 310 927 360 961
rect 394 927 422 961
rect 248 891 422 927
rect 120 867 186 883
rect 120 833 136 867
rect 170 833 186 867
rect 248 857 264 891
rect 406 857 422 891
rect 248 855 276 857
rect 310 855 360 857
rect 394 855 422 857
rect 248 841 422 855
rect 484 867 550 883
rect 120 817 186 833
rect 484 833 500 867
rect 534 833 550 867
rect 484 817 550 833
rect 120 795 160 817
rect 510 795 550 817
rect 41 779 160 795
rect 41 745 58 779
rect 92 759 126 779
rect 94 745 126 759
rect 41 725 60 745
rect 94 725 160 745
rect 41 711 160 725
rect 41 677 58 711
rect 92 687 126 711
rect 94 677 126 687
rect 41 653 60 677
rect 94 653 160 677
rect 41 643 160 653
rect 41 609 58 643
rect 92 615 126 643
rect 94 609 126 615
rect 41 581 60 609
rect 94 581 160 609
rect 41 575 160 581
rect 41 541 58 575
rect 92 543 126 575
rect 94 541 126 543
rect 41 509 60 541
rect 94 509 160 541
rect 41 507 160 509
rect 41 473 58 507
rect 92 473 126 507
rect 41 471 160 473
rect 41 439 60 471
rect 94 439 160 471
rect 41 405 58 439
rect 94 437 126 439
rect 92 405 126 437
rect 41 399 160 405
rect 41 371 60 399
rect 94 371 160 399
rect 41 337 58 371
rect 94 365 126 371
rect 92 337 126 365
rect 41 327 160 337
rect 41 303 60 327
rect 94 303 160 327
rect 41 269 58 303
rect 94 293 126 303
rect 92 269 126 293
rect 41 255 160 269
rect 41 235 60 255
rect 94 235 160 255
rect 41 201 58 235
rect 94 221 126 235
rect 92 201 126 221
rect 41 185 160 201
rect 212 779 246 795
rect 212 471 246 509
rect 212 185 246 201
rect 318 779 352 795
rect 318 471 352 509
rect 318 185 352 201
rect 424 779 458 795
rect 424 471 458 509
rect 424 185 458 201
rect 510 779 629 795
rect 544 759 578 779
rect 544 745 576 759
rect 612 745 629 779
rect 510 725 576 745
rect 610 725 629 745
rect 510 711 629 725
rect 544 687 578 711
rect 544 677 576 687
rect 612 677 629 711
rect 510 653 576 677
rect 610 653 629 677
rect 510 643 629 653
rect 544 615 578 643
rect 544 609 576 615
rect 612 609 629 643
rect 510 581 576 609
rect 610 581 629 609
rect 510 575 629 581
rect 544 543 578 575
rect 544 541 576 543
rect 612 541 629 575
rect 510 509 576 541
rect 610 509 629 541
rect 510 507 629 509
rect 544 473 578 507
rect 612 473 629 507
rect 510 471 629 473
rect 510 439 576 471
rect 610 439 629 471
rect 544 437 576 439
rect 544 405 578 437
rect 612 405 629 439
rect 510 399 629 405
rect 510 371 576 399
rect 610 371 629 399
rect 544 365 576 371
rect 544 337 578 365
rect 612 337 629 371
rect 510 327 629 337
rect 510 303 576 327
rect 610 303 629 327
rect 544 293 576 303
rect 544 269 578 293
rect 612 269 629 303
rect 510 255 629 269
rect 510 235 576 255
rect 610 235 629 255
rect 544 221 576 235
rect 544 201 578 221
rect 612 201 629 235
rect 510 185 629 201
rect 120 163 160 185
rect 510 163 550 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 484 147 550 163
rect 120 97 186 113
rect 248 125 422 139
rect 248 123 276 125
rect 310 123 360 125
rect 394 123 422 125
rect 248 89 264 123
rect 406 89 422 123
rect 484 113 500 147
rect 534 113 550 147
rect 484 97 550 113
rect 248 53 422 89
rect 248 19 276 53
rect 310 19 360 53
rect 394 19 422 53
rect 248 0 422 19
<< viali >>
rect 276 927 310 961
rect 360 927 394 961
rect 276 857 310 889
rect 360 857 394 889
rect 276 855 310 857
rect 360 855 394 857
rect 60 745 92 759
rect 92 745 94 759
rect 60 725 94 745
rect 60 677 92 687
rect 92 677 94 687
rect 60 653 94 677
rect 60 609 92 615
rect 92 609 94 615
rect 60 581 94 609
rect 60 541 92 543
rect 92 541 94 543
rect 60 509 94 541
rect 60 439 94 471
rect 60 437 92 439
rect 92 437 94 439
rect 60 371 94 399
rect 60 365 92 371
rect 92 365 94 371
rect 60 303 94 327
rect 60 293 92 303
rect 92 293 94 303
rect 60 235 94 255
rect 60 221 92 235
rect 92 221 94 235
rect 212 725 246 759
rect 212 653 246 687
rect 212 581 246 615
rect 212 513 246 543
rect 212 509 246 513
rect 212 467 246 471
rect 212 437 246 467
rect 212 365 246 399
rect 212 293 246 327
rect 212 221 246 255
rect 318 725 352 759
rect 318 653 352 687
rect 318 581 352 615
rect 318 513 352 543
rect 318 509 352 513
rect 318 467 352 471
rect 318 437 352 467
rect 318 365 352 399
rect 318 293 352 327
rect 318 221 352 255
rect 424 725 458 759
rect 424 653 458 687
rect 424 581 458 615
rect 424 513 458 543
rect 424 509 458 513
rect 424 467 458 471
rect 424 437 458 467
rect 424 365 458 399
rect 424 293 458 327
rect 424 221 458 255
rect 576 745 578 759
rect 578 745 610 759
rect 576 725 610 745
rect 576 677 578 687
rect 578 677 610 687
rect 576 653 610 677
rect 576 609 578 615
rect 578 609 610 615
rect 576 581 610 609
rect 576 541 578 543
rect 578 541 610 543
rect 576 509 610 541
rect 576 439 610 471
rect 576 437 578 439
rect 578 437 610 439
rect 576 371 610 399
rect 576 365 578 371
rect 578 365 610 371
rect 576 303 610 327
rect 576 293 578 303
rect 578 293 610 303
rect 576 235 610 255
rect 576 221 578 235
rect 578 221 610 235
rect 276 123 310 125
rect 360 123 394 125
rect 276 91 310 123
rect 360 91 394 123
rect 276 19 310 53
rect 360 19 394 53
<< metal1 >>
rect 250 961 420 980
rect 250 927 276 961
rect 310 927 360 961
rect 394 927 420 961
rect 250 889 420 927
rect 250 855 276 889
rect 310 855 360 889
rect 394 855 420 889
rect 250 843 420 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 203 759 255 771
rect 203 725 212 759
rect 246 725 255 759
rect 203 687 255 725
rect 203 653 212 687
rect 246 653 255 687
rect 203 615 255 653
rect 203 581 212 615
rect 246 581 255 615
rect 203 543 255 581
rect 203 509 212 543
rect 246 509 255 543
rect 203 471 255 509
rect 203 459 212 471
rect 246 459 255 471
rect 203 399 255 407
rect 203 395 212 399
rect 246 395 255 399
rect 203 331 255 343
rect 203 267 255 279
rect 203 209 255 215
rect 309 765 361 771
rect 309 701 361 713
rect 309 637 361 649
rect 309 581 318 585
rect 352 581 361 585
rect 309 573 361 581
rect 309 509 318 521
rect 352 509 361 521
rect 309 471 361 509
rect 309 437 318 471
rect 352 437 361 471
rect 309 399 361 437
rect 309 365 318 399
rect 352 365 361 399
rect 309 327 361 365
rect 309 293 318 327
rect 352 293 361 327
rect 309 255 361 293
rect 309 221 318 255
rect 352 221 361 255
rect 309 209 361 221
rect 415 759 467 771
rect 415 725 424 759
rect 458 725 467 759
rect 415 687 467 725
rect 415 653 424 687
rect 458 653 467 687
rect 415 615 467 653
rect 415 581 424 615
rect 458 581 467 615
rect 415 543 467 581
rect 415 509 424 543
rect 458 509 467 543
rect 415 471 467 509
rect 415 459 424 471
rect 458 459 467 471
rect 415 399 467 407
rect 415 395 424 399
rect 458 395 467 399
rect 415 331 467 343
rect 415 267 467 279
rect 415 209 467 215
rect 570 759 629 771
rect 570 725 576 759
rect 610 725 629 759
rect 570 687 629 725
rect 570 653 576 687
rect 610 653 629 687
rect 570 615 629 653
rect 570 581 576 615
rect 610 581 629 615
rect 570 543 629 581
rect 570 509 576 543
rect 610 509 629 543
rect 570 471 629 509
rect 570 437 576 471
rect 610 437 629 471
rect 570 399 629 437
rect 570 365 576 399
rect 610 365 629 399
rect 570 327 629 365
rect 570 293 576 327
rect 610 293 629 327
rect 570 255 629 293
rect 570 221 576 255
rect 610 221 629 255
rect 570 209 629 221
rect 250 125 420 137
rect 250 91 276 125
rect 310 91 360 125
rect 394 91 420 125
rect 250 53 420 91
rect 250 19 276 53
rect 310 19 360 53
rect 394 19 420 53
rect 250 0 420 19
<< via1 >>
rect 203 437 212 459
rect 212 437 246 459
rect 246 437 255 459
rect 203 407 255 437
rect 203 365 212 395
rect 212 365 246 395
rect 246 365 255 395
rect 203 343 255 365
rect 203 327 255 331
rect 203 293 212 327
rect 212 293 246 327
rect 246 293 255 327
rect 203 279 255 293
rect 203 255 255 267
rect 203 221 212 255
rect 212 221 246 255
rect 246 221 255 255
rect 203 215 255 221
rect 309 759 361 765
rect 309 725 318 759
rect 318 725 352 759
rect 352 725 361 759
rect 309 713 361 725
rect 309 687 361 701
rect 309 653 318 687
rect 318 653 352 687
rect 352 653 361 687
rect 309 649 361 653
rect 309 615 361 637
rect 309 585 318 615
rect 318 585 352 615
rect 352 585 361 615
rect 309 543 361 573
rect 309 521 318 543
rect 318 521 352 543
rect 352 521 361 543
rect 415 437 424 459
rect 424 437 458 459
rect 458 437 467 459
rect 415 407 467 437
rect 415 365 424 395
rect 424 365 458 395
rect 458 365 467 395
rect 415 343 467 365
rect 415 327 467 331
rect 415 293 424 327
rect 424 293 458 327
rect 458 293 467 327
rect 415 279 467 293
rect 415 255 467 267
rect 415 221 424 255
rect 424 221 458 255
rect 458 221 467 255
rect 415 215 467 221
<< metal2 >>
rect 14 765 656 771
rect 14 713 309 765
rect 361 713 656 765
rect 14 701 656 713
rect 14 649 309 701
rect 361 649 656 701
rect 14 637 656 649
rect 14 585 309 637
rect 361 585 656 637
rect 14 573 656 585
rect 14 521 309 573
rect 361 521 656 573
rect 14 515 656 521
rect 14 459 656 465
rect 14 407 203 459
rect 255 407 415 459
rect 467 407 656 459
rect 14 395 656 407
rect 14 343 203 395
rect 255 343 415 395
rect 467 343 656 395
rect 14 331 656 343
rect 14 279 203 331
rect 255 279 415 331
rect 467 279 656 331
rect 14 267 656 279
rect 14 215 203 267
rect 255 215 415 267
rect 467 215 656 267
rect 14 209 656 215
<< labels >>
flabel comment s 182 506 182 506 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 482 499 482 499 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 44 414 95 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 255 880 414 931 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 570 469 629 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 14 280 35 408 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 589 35 717 7 FreeSans 300 180 0 0 DRAIN
port 4 nsew
<< properties >>
string GDS_END 6686672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6673808
<< end >>
