magic
tech sky130B
magscale 12 1
timestamp 1598786254
<< metal5 >>
rect 0 75 30 105
rect 15 60 30 75
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
