VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO peripherals
  CLASS BLOCK ;
  FOREIGN peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 2200.000 ;
  PIN axi_spi_master_ar_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 2196.000 621.830 2200.000 ;
    END
  END axi_spi_master_ar_addr[0]
  PIN axi_spi_master_ar_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END axi_spi_master_ar_addr[10]
  PIN axi_spi_master_ar_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END axi_spi_master_ar_addr[11]
  PIN axi_spi_master_ar_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 180.240 700.000 180.840 ;
    END
  END axi_spi_master_ar_addr[12]
  PIN axi_spi_master_ar_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 989.440 700.000 990.040 ;
    END
  END axi_spi_master_ar_addr[13]
  PIN axi_spi_master_ar_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END axi_spi_master_ar_addr[14]
  PIN axi_spi_master_ar_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END axi_spi_master_ar_addr[15]
  PIN axi_spi_master_ar_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END axi_spi_master_ar_addr[16]
  PIN axi_spi_master_ar_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2053.640 700.000 2054.240 ;
    END
  END axi_spi_master_ar_addr[17]
  PIN axi_spi_master_ar_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END axi_spi_master_ar_addr[18]
  PIN axi_spi_master_ar_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1706.840 4.000 1707.440 ;
    END
  END axi_spi_master_ar_addr[19]
  PIN axi_spi_master_ar_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END axi_spi_master_ar_addr[1]
  PIN axi_spi_master_ar_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 2196.000 695.890 2200.000 ;
    END
  END axi_spi_master_ar_addr[20]
  PIN axi_spi_master_ar_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.240 4.000 1914.840 ;
    END
  END axi_spi_master_ar_addr[21]
  PIN axi_spi_master_ar_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1638.840 700.000 1639.440 ;
    END
  END axi_spi_master_ar_addr[22]
  PIN axi_spi_master_ar_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 112.240 700.000 112.840 ;
    END
  END axi_spi_master_ar_addr[23]
  PIN axi_spi_master_ar_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 707.240 700.000 707.840 ;
    END
  END axi_spi_master_ar_addr[24]
  PIN axi_spi_master_ar_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END axi_spi_master_ar_addr[25]
  PIN axi_spi_master_ar_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 2196.000 512.350 2200.000 ;
    END
  END axi_spi_master_ar_addr[26]
  PIN axi_spi_master_ar_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 289.040 700.000 289.640 ;
    END
  END axi_spi_master_ar_addr[27]
  PIN axi_spi_master_ar_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 2196.000 351.350 2200.000 ;
    END
  END axi_spi_master_ar_addr[28]
  PIN axi_spi_master_ar_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1774.840 4.000 1775.440 ;
    END
  END axi_spi_master_ar_addr[29]
  PIN axi_spi_master_ar_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END axi_spi_master_ar_addr[2]
  PIN axi_spi_master_ar_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 567.840 700.000 568.440 ;
    END
  END axi_spi_master_ar_addr[30]
  PIN axi_spi_master_ar_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 2196.000 576.750 2200.000 ;
    END
  END axi_spi_master_ar_addr[31]
  PIN axi_spi_master_ar_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END axi_spi_master_ar_addr[3]
  PIN axi_spi_master_ar_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 2196.000 245.090 2200.000 ;
    END
  END axi_spi_master_ar_addr[4]
  PIN axi_spi_master_ar_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 2196.000 425.410 2200.000 ;
    END
  END axi_spi_master_ar_addr[5]
  PIN axi_spi_master_ar_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END axi_spi_master_ar_addr[6]
  PIN axi_spi_master_ar_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1880.240 700.000 1880.840 ;
    END
  END axi_spi_master_ar_addr[7]
  PIN axi_spi_master_ar_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 2196.000 676.570 2200.000 ;
    END
  END axi_spi_master_ar_addr[8]
  PIN axi_spi_master_ar_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 646.040 700.000 646.640 ;
    END
  END axi_spi_master_ar_addr[9]
  PIN axi_spi_master_ar_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END axi_spi_master_ar_burst[0]
  PIN axi_spi_master_ar_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 2196.000 602.510 2200.000 ;
    END
  END axi_spi_master_ar_burst[1]
  PIN axi_spi_master_ar_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END axi_spi_master_ar_cache[0]
  PIN axi_spi_master_ar_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END axi_spi_master_ar_cache[1]
  PIN axi_spi_master_ar_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2189.640 700.000 2190.240 ;
    END
  END axi_spi_master_ar_cache[2]
  PIN axi_spi_master_ar_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1938.040 4.000 1938.640 ;
    END
  END axi_spi_master_ar_cache[3]
  PIN axi_spi_master_ar_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2094.440 700.000 2095.040 ;
    END
  END axi_spi_master_ar_id[0]
  PIN axi_spi_master_ar_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 452.240 700.000 452.840 ;
    END
  END axi_spi_master_ar_id[1]
  PIN axi_spi_master_ar_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 459.040 700.000 459.640 ;
    END
  END axi_spi_master_ar_id[2]
  PIN axi_spi_master_ar_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 523.640 700.000 524.240 ;
    END
  END axi_spi_master_ar_id[3]
  PIN axi_spi_master_ar_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1247.840 700.000 1248.440 ;
    END
  END axi_spi_master_ar_id[4]
  PIN axi_spi_master_ar_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 4.000 1850.240 ;
    END
  END axi_spi_master_ar_id[5]
  PIN axi_spi_master_ar_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END axi_spi_master_ar_len[0]
  PIN axi_spi_master_ar_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 37.440 700.000 38.040 ;
    END
  END axi_spi_master_ar_len[1]
  PIN axi_spi_master_ar_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END axi_spi_master_ar_len[2]
  PIN axi_spi_master_ar_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END axi_spi_master_ar_len[3]
  PIN axi_spi_master_ar_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 132.640 700.000 133.240 ;
    END
  END axi_spi_master_ar_len[4]
  PIN axi_spi_master_ar_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END axi_spi_master_ar_len[5]
  PIN axi_spi_master_ar_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END axi_spi_master_ar_len[6]
  PIN axi_spi_master_ar_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END axi_spi_master_ar_len[7]
  PIN axi_spi_master_ar_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END axi_spi_master_ar_lock
  PIN axi_spi_master_ar_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 153.040 700.000 153.640 ;
    END
  END axi_spi_master_ar_prot[0]
  PIN axi_spi_master_ar_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2029.840 700.000 2030.440 ;
    END
  END axi_spi_master_ar_prot[1]
  PIN axi_spi_master_ar_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END axi_spi_master_ar_prot[2]
  PIN axi_spi_master_ar_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2063.840 4.000 2064.440 ;
    END
  END axi_spi_master_ar_qos[0]
  PIN axi_spi_master_ar_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1050.640 700.000 1051.240 ;
    END
  END axi_spi_master_ar_qos[1]
  PIN axi_spi_master_ar_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END axi_spi_master_ar_qos[2]
  PIN axi_spi_master_ar_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2193.040 700.000 2193.640 ;
    END
  END axi_spi_master_ar_qos[3]
  PIN axi_spi_master_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 2196.000 373.890 2200.000 ;
    END
  END axi_spi_master_ar_ready
  PIN axi_spi_master_ar_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END axi_spi_master_ar_region[0]
  PIN axi_spi_master_ar_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1149.240 700.000 1149.840 ;
    END
  END axi_spi_master_ar_region[1]
  PIN axi_spi_master_ar_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 632.440 700.000 633.040 ;
    END
  END axi_spi_master_ar_region[2]
  PIN axi_spi_master_ar_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END axi_spi_master_ar_region[3]
  PIN axi_spi_master_ar_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1812.240 700.000 1812.840 ;
    END
  END axi_spi_master_ar_size[0]
  PIN axi_spi_master_ar_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2084.240 700.000 2084.840 ;
    END
  END axi_spi_master_ar_size[1]
  PIN axi_spi_master_ar_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 901.040 700.000 901.640 ;
    END
  END axi_spi_master_ar_size[2]
  PIN axi_spi_master_ar_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END axi_spi_master_ar_user[0]
  PIN axi_spi_master_ar_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END axi_spi_master_ar_user[1]
  PIN axi_spi_master_ar_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1876.840 700.000 1877.440 ;
    END
  END axi_spi_master_ar_user[2]
  PIN axi_spi_master_ar_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END axi_spi_master_ar_user[3]
  PIN axi_spi_master_ar_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END axi_spi_master_ar_user[4]
  PIN axi_spi_master_ar_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END axi_spi_master_ar_user[5]
  PIN axi_spi_master_ar_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1958.440 700.000 1959.040 ;
    END
  END axi_spi_master_ar_valid
  PIN axi_spi_master_aw_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END axi_spi_master_aw_addr[0]
  PIN axi_spi_master_aw_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 431.840 700.000 432.440 ;
    END
  END axi_spi_master_aw_addr[10]
  PIN axi_spi_master_aw_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END axi_spi_master_aw_addr[11]
  PIN axi_spi_master_aw_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 2196.000 431.850 2200.000 ;
    END
  END axi_spi_master_aw_addr[12]
  PIN axi_spi_master_aw_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 2196.000 615.390 2200.000 ;
    END
  END axi_spi_master_aw_addr[13]
  PIN axi_spi_master_aw_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 2196.000 679.790 2200.000 ;
    END
  END axi_spi_master_aw_addr[14]
  PIN axi_spi_master_aw_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END axi_spi_master_aw_addr[15]
  PIN axi_spi_master_aw_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1499.440 700.000 1500.040 ;
    END
  END axi_spi_master_aw_addr[16]
  PIN axi_spi_master_aw_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END axi_spi_master_aw_addr[17]
  PIN axi_spi_master_aw_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END axi_spi_master_aw_addr[18]
  PIN axi_spi_master_aw_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 591.640 700.000 592.240 ;
    END
  END axi_spi_master_aw_addr[19]
  PIN axi_spi_master_aw_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 2196.000 283.730 2200.000 ;
    END
  END axi_spi_master_aw_addr[1]
  PIN axi_spi_master_aw_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1873.440 700.000 1874.040 ;
    END
  END axi_spi_master_aw_addr[20]
  PIN axi_spi_master_aw_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END axi_spi_master_aw_addr[21]
  PIN axi_spi_master_aw_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 2196.000 625.050 2200.000 ;
    END
  END axi_spi_master_aw_addr[22]
  PIN axi_spi_master_aw_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1836.040 4.000 1836.640 ;
    END
  END axi_spi_master_aw_addr[23]
  PIN axi_spi_master_aw_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END axi_spi_master_aw_addr[24]
  PIN axi_spi_master_aw_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END axi_spi_master_aw_addr[25]
  PIN axi_spi_master_aw_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END axi_spi_master_aw_addr[26]
  PIN axi_spi_master_aw_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END axi_spi_master_aw_addr[27]
  PIN axi_spi_master_aw_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1795.240 4.000 1795.840 ;
    END
  END axi_spi_master_aw_addr[28]
  PIN axi_spi_master_aw_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 2196.000 225.770 2200.000 ;
    END
  END axi_spi_master_aw_addr[29]
  PIN axi_spi_master_aw_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1625.240 700.000 1625.840 ;
    END
  END axi_spi_master_aw_addr[2]
  PIN axi_spi_master_aw_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1856.440 4.000 1857.040 ;
    END
  END axi_spi_master_aw_addr[30]
  PIN axi_spi_master_aw_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END axi_spi_master_aw_addr[31]
  PIN axi_spi_master_aw_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1176.440 700.000 1177.040 ;
    END
  END axi_spi_master_aw_addr[3]
  PIN axi_spi_master_aw_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END axi_spi_master_aw_addr[4]
  PIN axi_spi_master_aw_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1757.840 700.000 1758.440 ;
    END
  END axi_spi_master_aw_addr[5]
  PIN axi_spi_master_aw_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END axi_spi_master_aw_addr[6]
  PIN axi_spi_master_aw_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1968.640 4.000 1969.240 ;
    END
  END axi_spi_master_aw_addr[7]
  PIN axi_spi_master_aw_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END axi_spi_master_aw_addr[8]
  PIN axi_spi_master_aw_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END axi_spi_master_aw_addr[9]
  PIN axi_spi_master_aw_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 2196.000 544.550 2200.000 ;
    END
  END axi_spi_master_aw_burst[0]
  PIN axi_spi_master_aw_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END axi_spi_master_aw_burst[1]
  PIN axi_spi_master_aw_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END axi_spi_master_aw_cache[0]
  PIN axi_spi_master_aw_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1519.840 700.000 1520.440 ;
    END
  END axi_spi_master_aw_cache[1]
  PIN axi_spi_master_aw_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1805.440 4.000 1806.040 ;
    END
  END axi_spi_master_aw_cache[2]
  PIN axi_spi_master_aw_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1098.240 700.000 1098.840 ;
    END
  END axi_spi_master_aw_cache[3]
  PIN axi_spi_master_aw_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1387.240 700.000 1387.840 ;
    END
  END axi_spi_master_aw_id[0]
  PIN axi_spi_master_aw_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1880.240 4.000 1880.840 ;
    END
  END axi_spi_master_aw_id[1]
  PIN axi_spi_master_aw_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1883.640 700.000 1884.240 ;
    END
  END axi_spi_master_aw_id[2]
  PIN axi_spi_master_aw_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 897.640 700.000 898.240 ;
    END
  END axi_spi_master_aw_id[3]
  PIN axi_spi_master_aw_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2036.640 700.000 2037.240 ;
    END
  END axi_spi_master_aw_id[4]
  PIN axi_spi_master_aw_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1217.240 700.000 1217.840 ;
    END
  END axi_spi_master_aw_id[5]
  PIN axi_spi_master_aw_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1043.840 700.000 1044.440 ;
    END
  END axi_spi_master_aw_len[0]
  PIN axi_spi_master_aw_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1822.440 4.000 1823.040 ;
    END
  END axi_spi_master_aw_len[1]
  PIN axi_spi_master_aw_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END axi_spi_master_aw_len[2]
  PIN axi_spi_master_aw_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2006.040 700.000 2006.640 ;
    END
  END axi_spi_master_aw_len[3]
  PIN axi_spi_master_aw_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END axi_spi_master_aw_len[4]
  PIN axi_spi_master_aw_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 741.240 700.000 741.840 ;
    END
  END axi_spi_master_aw_len[5]
  PIN axi_spi_master_aw_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 142.840 700.000 143.440 ;
    END
  END axi_spi_master_aw_len[6]
  PIN axi_spi_master_aw_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END axi_spi_master_aw_len[7]
  PIN axi_spi_master_aw_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1455.240 700.000 1455.840 ;
    END
  END axi_spi_master_aw_lock
  PIN axi_spi_master_aw_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END axi_spi_master_aw_prot[0]
  PIN axi_spi_master_aw_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2043.440 700.000 2044.040 ;
    END
  END axi_spi_master_aw_prot[1]
  PIN axi_spi_master_aw_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END axi_spi_master_aw_prot[2]
  PIN axi_spi_master_aw_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 2196.000 303.050 2200.000 ;
    END
  END axi_spi_master_aw_qos[0]
  PIN axi_spi_master_aw_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1989.040 4.000 1989.640 ;
    END
  END axi_spi_master_aw_qos[1]
  PIN axi_spi_master_aw_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 2196.000 151.710 2200.000 ;
    END
  END axi_spi_master_aw_qos[2]
  PIN axi_spi_master_aw_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END axi_spi_master_aw_qos[3]
  PIN axi_spi_master_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END axi_spi_master_aw_ready
  PIN axi_spi_master_aw_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END axi_spi_master_aw_region[0]
  PIN axi_spi_master_aw_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END axi_spi_master_aw_region[1]
  PIN axi_spi_master_aw_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1162.840 700.000 1163.440 ;
    END
  END axi_spi_master_aw_region[2]
  PIN axi_spi_master_aw_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END axi_spi_master_aw_region[3]
  PIN axi_spi_master_aw_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END axi_spi_master_aw_size[0]
  PIN axi_spi_master_aw_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END axi_spi_master_aw_size[1]
  PIN axi_spi_master_aw_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 571.240 700.000 571.840 ;
    END
  END axi_spi_master_aw_size[2]
  PIN axi_spi_master_aw_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 2196.000 531.670 2200.000 ;
    END
  END axi_spi_master_aw_user[0]
  PIN axi_spi_master_aw_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1751.040 700.000 1751.640 ;
    END
  END axi_spi_master_aw_user[1]
  PIN axi_spi_master_aw_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END axi_spi_master_aw_user[2]
  PIN axi_spi_master_aw_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END axi_spi_master_aw_user[3]
  PIN axi_spi_master_aw_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 2196.000 666.910 2200.000 ;
    END
  END axi_spi_master_aw_user[4]
  PIN axi_spi_master_aw_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 221.040 700.000 221.640 ;
    END
  END axi_spi_master_aw_user[5]
  PIN axi_spi_master_aw_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 2196.000 264.410 2200.000 ;
    END
  END axi_spi_master_aw_valid
  PIN axi_spi_master_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1768.040 700.000 1768.640 ;
    END
  END axi_spi_master_b_id[0]
  PIN axi_spi_master_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1108.440 700.000 1109.040 ;
    END
  END axi_spi_master_b_id[1]
  PIN axi_spi_master_b_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 146.240 700.000 146.840 ;
    END
  END axi_spi_master_b_id[2]
  PIN axi_spi_master_b_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 2196.000 483.370 2200.000 ;
    END
  END axi_spi_master_b_id[3]
  PIN axi_spi_master_b_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END axi_spi_master_b_id[4]
  PIN axi_spi_master_b_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END axi_spi_master_b_id[5]
  PIN axi_spi_master_b_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.840 4.000 1469.440 ;
    END
  END axi_spi_master_b_ready
  PIN axi_spi_master_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END axi_spi_master_b_resp[0]
  PIN axi_spi_master_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1394.040 700.000 1394.640 ;
    END
  END axi_spi_master_b_resp[1]
  PIN axi_spi_master_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 2196.000 193.570 2200.000 ;
    END
  END axi_spi_master_b_user[0]
  PIN axi_spi_master_b_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END axi_spi_master_b_user[1]
  PIN axi_spi_master_b_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 496.440 700.000 497.040 ;
    END
  END axi_spi_master_b_user[2]
  PIN axi_spi_master_b_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END axi_spi_master_b_user[3]
  PIN axi_spi_master_b_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1203.640 4.000 1204.240 ;
    END
  END axi_spi_master_b_user[4]
  PIN axi_spi_master_b_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 2196.000 418.970 2200.000 ;
    END
  END axi_spi_master_b_user[5]
  PIN axi_spi_master_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END axi_spi_master_b_valid
  PIN axi_spi_master_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END axi_spi_master_r_data[0]
  PIN axi_spi_master_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1037.040 700.000 1037.640 ;
    END
  END axi_spi_master_r_data[10]
  PIN axi_spi_master_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 159.840 700.000 160.440 ;
    END
  END axi_spi_master_r_data[11]
  PIN axi_spi_master_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 421.640 700.000 422.240 ;
    END
  END axi_spi_master_r_data[12]
  PIN axi_spi_master_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1717.040 700.000 1717.640 ;
    END
  END axi_spi_master_r_data[13]
  PIN axi_spi_master_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2193.040 4.000 2193.640 ;
    END
  END axi_spi_master_r_data[14]
  PIN axi_spi_master_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END axi_spi_master_r_data[15]
  PIN axi_spi_master_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2114.840 4.000 2115.440 ;
    END
  END axi_spi_master_r_data[16]
  PIN axi_spi_master_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2121.640 700.000 2122.240 ;
    END
  END axi_spi_master_r_data[17]
  PIN axi_spi_master_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END axi_spi_master_r_data[18]
  PIN axi_spi_master_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 2196.000 344.910 2200.000 ;
    END
  END axi_spi_master_r_data[19]
  PIN axi_spi_master_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END axi_spi_master_r_data[1]
  PIN axi_spi_master_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1356.640 700.000 1357.240 ;
    END
  END axi_spi_master_r_data[20]
  PIN axi_spi_master_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 2196.000 58.330 2200.000 ;
    END
  END axi_spi_master_r_data[21]
  PIN axi_spi_master_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 884.040 700.000 884.640 ;
    END
  END axi_spi_master_r_data[22]
  PIN axi_spi_master_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END axi_spi_master_r_data[23]
  PIN axi_spi_master_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 2196.000 663.690 2200.000 ;
    END
  END axi_spi_master_r_data[24]
  PIN axi_spi_master_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END axi_spi_master_r_data[25]
  PIN axi_spi_master_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 442.040 700.000 442.640 ;
    END
  END axi_spi_master_r_data[26]
  PIN axi_spi_master_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1859.840 4.000 1860.440 ;
    END
  END axi_spi_master_r_data[27]
  PIN axi_spi_master_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1540.240 4.000 1540.840 ;
    END
  END axi_spi_master_r_data[28]
  PIN axi_spi_master_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END axi_spi_master_r_data[29]
  PIN axi_spi_master_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 394.440 700.000 395.040 ;
    END
  END axi_spi_master_r_data[2]
  PIN axi_spi_master_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 224.440 700.000 225.040 ;
    END
  END axi_spi_master_r_data[30]
  PIN axi_spi_master_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END axi_spi_master_r_data[31]
  PIN axi_spi_master_r_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1747.640 700.000 1748.240 ;
    END
  END axi_spi_master_r_data[32]
  PIN axi_spi_master_r_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 673.240 700.000 673.840 ;
    END
  END axi_spi_master_r_data[33]
  PIN axi_spi_master_r_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 887.440 700.000 888.040 ;
    END
  END axi_spi_master_r_data[34]
  PIN axi_spi_master_r_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 2196.000 171.030 2200.000 ;
    END
  END axi_spi_master_r_data[35]
  PIN axi_spi_master_r_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 540.640 700.000 541.240 ;
    END
  END axi_spi_master_r_data[36]
  PIN axi_spi_master_r_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.040 4.000 1496.640 ;
    END
  END axi_spi_master_r_data[37]
  PIN axi_spi_master_r_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1635.440 4.000 1636.040 ;
    END
  END axi_spi_master_r_data[38]
  PIN axi_spi_master_r_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1363.440 700.000 1364.040 ;
    END
  END axi_spi_master_r_data[39]
  PIN axi_spi_master_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1237.640 700.000 1238.240 ;
    END
  END axi_spi_master_r_data[3]
  PIN axi_spi_master_r_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END axi_spi_master_r_data[40]
  PIN axi_spi_master_r_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END axi_spi_master_r_data[41]
  PIN axi_spi_master_r_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END axi_spi_master_r_data[42]
  PIN axi_spi_master_r_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.840 700.000 296.440 ;
    END
  END axi_spi_master_r_data[43]
  PIN axi_spi_master_r_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1288.640 700.000 1289.240 ;
    END
  END axi_spi_master_r_data[44]
  PIN axi_spi_master_r_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1948.240 4.000 1948.840 ;
    END
  END axi_spi_master_r_data[45]
  PIN axi_spi_master_r_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1999.240 4.000 1999.840 ;
    END
  END axi_spi_master_r_data[46]
  PIN axi_spi_master_r_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 2196.000 422.190 2200.000 ;
    END
  END axi_spi_master_r_data[47]
  PIN axi_spi_master_r_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2002.640 4.000 2003.240 ;
    END
  END axi_spi_master_r_data[48]
  PIN axi_spi_master_r_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END axi_spi_master_r_data[49]
  PIN axi_spi_master_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1618.440 700.000 1619.040 ;
    END
  END axi_spi_master_r_data[4]
  PIN axi_spi_master_r_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1965.240 4.000 1965.840 ;
    END
  END axi_spi_master_r_data[50]
  PIN axi_spi_master_r_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END axi_spi_master_r_data[51]
  PIN axi_spi_master_r_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2172.640 4.000 2173.240 ;
    END
  END axi_spi_master_r_data[52]
  PIN axi_spi_master_r_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1890.440 4.000 1891.040 ;
    END
  END axi_spi_master_r_data[53]
  PIN axi_spi_master_r_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1944.840 700.000 1945.440 ;
    END
  END axi_spi_master_r_data[54]
  PIN axi_spi_master_r_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END axi_spi_master_r_data[55]
  PIN axi_spi_master_r_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2182.840 4.000 2183.440 ;
    END
  END axi_spi_master_r_data[56]
  PIN axi_spi_master_r_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1985.640 700.000 1986.240 ;
    END
  END axi_spi_master_r_data[57]
  PIN axi_spi_master_r_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END axi_spi_master_r_data[58]
  PIN axi_spi_master_r_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2029.840 4.000 2030.440 ;
    END
  END axi_spi_master_r_data[59]
  PIN axi_spi_master_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1832.640 4.000 1833.240 ;
    END
  END axi_spi_master_r_data[5]
  PIN axi_spi_master_r_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END axi_spi_master_r_data[60]
  PIN axi_spi_master_r_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 2196.000 338.470 2200.000 ;
    END
  END axi_spi_master_r_data[61]
  PIN axi_spi_master_r_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1370.240 700.000 1370.840 ;
    END
  END axi_spi_master_r_data[62]
  PIN axi_spi_master_r_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 2196.000 135.610 2200.000 ;
    END
  END axi_spi_master_r_data[63]
  PIN axi_spi_master_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1737.440 4.000 1738.040 ;
    END
  END axi_spi_master_r_data[6]
  PIN axi_spi_master_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END axi_spi_master_r_data[7]
  PIN axi_spi_master_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 792.240 700.000 792.840 ;
    END
  END axi_spi_master_r_data[8]
  PIN axi_spi_master_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END axi_spi_master_r_data[9]
  PIN axi_spi_master_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1917.640 700.000 1918.240 ;
    END
  END axi_spi_master_r_id[0]
  PIN axi_spi_master_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END axi_spi_master_r_id[1]
  PIN axi_spi_master_r_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1832.640 700.000 1833.240 ;
    END
  END axi_spi_master_r_id[2]
  PIN axi_spi_master_r_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 2196.000 518.790 2200.000 ;
    END
  END axi_spi_master_r_id[3]
  PIN axi_spi_master_r_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END axi_spi_master_r_id[4]
  PIN axi_spi_master_r_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.240 4.000 1608.840 ;
    END
  END axi_spi_master_r_id[5]
  PIN axi_spi_master_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END axi_spi_master_r_last
  PIN axi_spi_master_r_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 652.840 700.000 653.440 ;
    END
  END axi_spi_master_r_ready
  PIN axi_spi_master_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2026.440 700.000 2027.040 ;
    END
  END axi_spi_master_r_resp[0]
  PIN axi_spi_master_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END axi_spi_master_r_resp[1]
  PIN axi_spi_master_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 292.440 700.000 293.040 ;
    END
  END axi_spi_master_r_user[0]
  PIN axi_spi_master_r_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1366.840 700.000 1367.440 ;
    END
  END axi_spi_master_r_user[1]
  PIN axi_spi_master_r_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END axi_spi_master_r_user[2]
  PIN axi_spi_master_r_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END axi_spi_master_r_user[3]
  PIN axi_spi_master_r_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 856.840 700.000 857.440 ;
    END
  END axi_spi_master_r_user[4]
  PIN axi_spi_master_r_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 312.840 700.000 313.440 ;
    END
  END axi_spi_master_r_user[5]
  PIN axi_spi_master_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2026.440 4.000 2027.040 ;
    END
  END axi_spi_master_r_valid
  PIN axi_spi_master_w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 2196.000 415.750 2200.000 ;
    END
  END axi_spi_master_w_data[0]
  PIN axi_spi_master_w_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1904.040 700.000 1904.640 ;
    END
  END axi_spi_master_w_data[10]
  PIN axi_spi_master_w_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1982.240 4.000 1982.840 ;
    END
  END axi_spi_master_w_data[11]
  PIN axi_spi_master_w_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END axi_spi_master_w_data[12]
  PIN axi_spi_master_w_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END axi_spi_master_w_data[13]
  PIN axi_spi_master_w_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 2196.000 251.530 2200.000 ;
    END
  END axi_spi_master_w_data[14]
  PIN axi_spi_master_w_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END axi_spi_master_w_data[15]
  PIN axi_spi_master_w_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END axi_spi_master_w_data[16]
  PIN axi_spi_master_w_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1771.440 700.000 1772.040 ;
    END
  END axi_spi_master_w_data[17]
  PIN axi_spi_master_w_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 2196.000 42.230 2200.000 ;
    END
  END axi_spi_master_w_data[18]
  PIN axi_spi_master_w_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 928.240 700.000 928.840 ;
    END
  END axi_spi_master_w_data[19]
  PIN axi_spi_master_w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END axi_spi_master_w_data[1]
  PIN axi_spi_master_w_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 282.240 700.000 282.840 ;
    END
  END axi_spi_master_w_data[20]
  PIN axi_spi_master_w_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 2196.000 39.010 2200.000 ;
    END
  END axi_spi_master_w_data[21]
  PIN axi_spi_master_w_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 833.040 700.000 833.640 ;
    END
  END axi_spi_master_w_data[22]
  PIN axi_spi_master_w_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1560.640 4.000 1561.240 ;
    END
  END axi_spi_master_w_data[23]
  PIN axi_spi_master_w_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 2196.000 380.330 2200.000 ;
    END
  END axi_spi_master_w_data[24]
  PIN axi_spi_master_w_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2077.440 700.000 2078.040 ;
    END
  END axi_spi_master_w_data[25]
  PIN axi_spi_master_w_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1978.840 700.000 1979.440 ;
    END
  END axi_spi_master_w_data[26]
  PIN axi_spi_master_w_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END axi_spi_master_w_data[27]
  PIN axi_spi_master_w_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END axi_spi_master_w_data[28]
  PIN axi_spi_master_w_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1118.640 700.000 1119.240 ;
    END
  END axi_spi_master_w_data[29]
  PIN axi_spi_master_w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 771.840 700.000 772.440 ;
    END
  END axi_spi_master_w_data[2]
  PIN axi_spi_master_w_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1516.440 700.000 1517.040 ;
    END
  END axi_spi_master_w_data[30]
  PIN axi_spi_master_w_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END axi_spi_master_w_data[31]
  PIN axi_spi_master_w_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END axi_spi_master_w_data[32]
  PIN axi_spi_master_w_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 527.040 700.000 527.640 ;
    END
  END axi_spi_master_w_data[33]
  PIN axi_spi_master_w_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END axi_spi_master_w_data[34]
  PIN axi_spi_master_w_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1023.440 700.000 1024.040 ;
    END
  END axi_spi_master_w_data[35]
  PIN axi_spi_master_w_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 809.240 700.000 809.840 ;
    END
  END axi_spi_master_w_data[36]
  PIN axi_spi_master_w_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 2196.000 261.190 2200.000 ;
    END
  END axi_spi_master_w_data[37]
  PIN axi_spi_master_w_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1492.640 700.000 1493.240 ;
    END
  END axi_spi_master_w_data[38]
  PIN axi_spi_master_w_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END axi_spi_master_w_data[39]
  PIN axi_spi_master_w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1955.040 4.000 1955.640 ;
    END
  END axi_spi_master_w_data[3]
  PIN axi_spi_master_w_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END axi_spi_master_w_data[40]
  PIN axi_spi_master_w_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1897.240 700.000 1897.840 ;
    END
  END axi_spi_master_w_data[41]
  PIN axi_spi_master_w_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END axi_spi_master_w_data[42]
  PIN axi_spi_master_w_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 799.040 700.000 799.640 ;
    END
  END axi_spi_master_w_data[43]
  PIN axi_spi_master_w_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1628.640 700.000 1629.240 ;
    END
  END axi_spi_master_w_data[44]
  PIN axi_spi_master_w_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END axi_spi_master_w_data[45]
  PIN axi_spi_master_w_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END axi_spi_master_w_data[46]
  PIN axi_spi_master_w_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 622.240 700.000 622.840 ;
    END
  END axi_spi_master_w_data[47]
  PIN axi_spi_master_w_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 996.240 700.000 996.840 ;
    END
  END axi_spi_master_w_data[48]
  PIN axi_spi_master_w_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 2196.000 232.210 2200.000 ;
    END
  END axi_spi_master_w_data[49]
  PIN axi_spi_master_w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END axi_spi_master_w_data[4]
  PIN axi_spi_master_w_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END axi_spi_master_w_data[50]
  PIN axi_spi_master_w_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END axi_spi_master_w_data[51]
  PIN axi_spi_master_w_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1397.440 4.000 1398.040 ;
    END
  END axi_spi_master_w_data[52]
  PIN axi_spi_master_w_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END axi_spi_master_w_data[53]
  PIN axi_spi_master_w_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END axi_spi_master_w_data[54]
  PIN axi_spi_master_w_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END axi_spi_master_w_data[55]
  PIN axi_spi_master_w_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1513.040 4.000 1513.640 ;
    END
  END axi_spi_master_w_data[56]
  PIN axi_spi_master_w_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1448.440 700.000 1449.040 ;
    END
  END axi_spi_master_w_data[57]
  PIN axi_spi_master_w_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END axi_spi_master_w_data[58]
  PIN axi_spi_master_w_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 2196.000 325.590 2200.000 ;
    END
  END axi_spi_master_w_data[59]
  PIN axi_spi_master_w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1999.240 700.000 1999.840 ;
    END
  END axi_spi_master_w_data[5]
  PIN axi_spi_master_w_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.240 4.000 1438.840 ;
    END
  END axi_spi_master_w_data[60]
  PIN axi_spi_master_w_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 2196.000 341.690 2200.000 ;
    END
  END axi_spi_master_w_data[61]
  PIN axi_spi_master_w_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END axi_spi_master_w_data[62]
  PIN axi_spi_master_w_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 561.040 700.000 561.640 ;
    END
  END axi_spi_master_w_data[63]
  PIN axi_spi_master_w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 782.040 700.000 782.640 ;
    END
  END axi_spi_master_w_data[6]
  PIN axi_spi_master_w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END axi_spi_master_w_data[7]
  PIN axi_spi_master_w_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END axi_spi_master_w_data[8]
  PIN axi_spi_master_w_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 2196.000 493.030 2200.000 ;
    END
  END axi_spi_master_w_data[9]
  PIN axi_spi_master_w_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END axi_spi_master_w_last
  PIN axi_spi_master_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2060.440 4.000 2061.040 ;
    END
  END axi_spi_master_w_ready
  PIN axi_spi_master_w_strb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END axi_spi_master_w_strb[0]
  PIN axi_spi_master_w_strb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END axi_spi_master_w_strb[1]
  PIN axi_spi_master_w_strb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 183.640 700.000 184.240 ;
    END
  END axi_spi_master_w_strb[2]
  PIN axi_spi_master_w_strb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 414.840 700.000 415.440 ;
    END
  END axi_spi_master_w_strb[3]
  PIN axi_spi_master_w_strb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END axi_spi_master_w_strb[4]
  PIN axi_spi_master_w_strb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END axi_spi_master_w_strb[5]
  PIN axi_spi_master_w_strb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END axi_spi_master_w_strb[6]
  PIN axi_spi_master_w_strb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2077.440 4.000 2078.040 ;
    END
  END axi_spi_master_w_strb[7]
  PIN axi_spi_master_w_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 81.640 700.000 82.240 ;
    END
  END axi_spi_master_w_user[0]
  PIN axi_spi_master_w_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 27.240 700.000 27.840 ;
    END
  END axi_spi_master_w_user[1]
  PIN axi_spi_master_w_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 2196.000 583.190 2200.000 ;
    END
  END axi_spi_master_w_user[2]
  PIN axi_spi_master_w_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END axi_spi_master_w_user[3]
  PIN axi_spi_master_w_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1839.440 4.000 1840.040 ;
    END
  END axi_spi_master_w_user[4]
  PIN axi_spi_master_w_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END axi_spi_master_w_user[5]
  PIN axi_spi_master_w_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END axi_spi_master_w_valid
  PIN boot_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1893.840 4.000 1894.440 ;
    END
  END boot_addr_o[0]
  PIN boot_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2145.440 4.000 2146.040 ;
    END
  END boot_addr_o[10]
  PIN boot_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END boot_addr_o[11]
  PIN boot_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1451.840 700.000 1452.440 ;
    END
  END boot_addr_o[12]
  PIN boot_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END boot_addr_o[13]
  PIN boot_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 119.040 700.000 119.640 ;
    END
  END boot_addr_o[14]
  PIN boot_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 95.240 700.000 95.840 ;
    END
  END boot_addr_o[15]
  PIN boot_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END boot_addr_o[16]
  PIN boot_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2046.840 4.000 2047.440 ;
    END
  END boot_addr_o[17]
  PIN boot_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END boot_addr_o[18]
  PIN boot_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1662.640 4.000 1663.240 ;
    END
  END boot_addr_o[19]
  PIN boot_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1744.240 700.000 1744.840 ;
    END
  END boot_addr_o[1]
  PIN boot_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END boot_addr_o[20]
  PIN boot_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END boot_addr_o[21]
  PIN boot_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1094.840 700.000 1095.440 ;
    END
  END boot_addr_o[22]
  PIN boot_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 2196.000 10.030 2200.000 ;
    END
  END boot_addr_o[23]
  PIN boot_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 479.440 700.000 480.040 ;
    END
  END boot_addr_o[24]
  PIN boot_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1428.040 700.000 1428.640 ;
    END
  END boot_addr_o[25]
  PIN boot_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 40.840 700.000 41.440 ;
    END
  END boot_addr_o[26]
  PIN boot_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 618.840 700.000 619.440 ;
    END
  END boot_addr_o[27]
  PIN boot_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2009.440 700.000 2010.040 ;
    END
  END boot_addr_o[28]
  PIN boot_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2009.440 4.000 2010.040 ;
    END
  END boot_addr_o[29]
  PIN boot_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 469.240 700.000 469.840 ;
    END
  END boot_addr_o[2]
  PIN boot_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END boot_addr_o[30]
  PIN boot_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END boot_addr_o[31]
  PIN boot_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2108.040 4.000 2108.640 ;
    END
  END boot_addr_o[3]
  PIN boot_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END boot_addr_o[4]
  PIN boot_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 2196.000 138.830 2200.000 ;
    END
  END boot_addr_o[5]
  PIN boot_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END boot_addr_o[6]
  PIN boot_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END boot_addr_o[7]
  PIN boot_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END boot_addr_o[8]
  PIN boot_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END boot_addr_o[9]
  PIN clk_gate_core_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END clk_gate_core_o
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END clk_i
  PIN clk_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1152.640 700.000 1153.240 ;
    END
  END clk_i_pll
  PIN clk_o_pll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END clk_o_pll
  PIN clk_sel_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END clk_sel_i_pll
  PIN clk_standalone_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 377.440 700.000 378.040 ;
    END
  END clk_standalone_i_pll
  PIN core_busy_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END core_busy_i
  PIN debug_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 2196.000 525.230 2200.000 ;
    END
  END debug_addr[0]
  PIN debug_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 2196.000 238.650 2200.000 ;
    END
  END debug_addr[10]
  PIN debug_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2138.640 4.000 2139.240 ;
    END
  END debug_addr[11]
  PIN debug_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END debug_addr[12]
  PIN debug_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END debug_addr[13]
  PIN debug_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 2196.000 399.650 2200.000 ;
    END
  END debug_addr[14]
  PIN debug_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1863.240 4.000 1863.840 ;
    END
  END debug_addr[1]
  PIN debug_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 2196.000 257.970 2200.000 ;
    END
  END debug_addr[2]
  PIN debug_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END debug_addr[3]
  PIN debug_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END debug_addr[4]
  PIN debug_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 2196.000 473.710 2200.000 ;
    END
  END debug_addr[5]
  PIN debug_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.040 4.000 1734.640 ;
    END
  END debug_addr[6]
  PIN debug_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END debug_addr[7]
  PIN debug_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END debug_addr[8]
  PIN debug_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 2196.000 109.850 2200.000 ;
    END
  END debug_addr[9]
  PIN debug_gnt
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END debug_gnt
  PIN debug_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 380.840 700.000 381.440 ;
    END
  END debug_rdata[0]
  PIN debug_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END debug_rdata[10]
  PIN debug_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END debug_rdata[11]
  PIN debug_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 122.440 700.000 123.040 ;
    END
  END debug_rdata[12]
  PIN debug_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 690.240 700.000 690.840 ;
    END
  END debug_rdata[13]
  PIN debug_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1479.040 700.000 1479.640 ;
    END
  END debug_rdata[14]
  PIN debug_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END debug_rdata[15]
  PIN debug_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 836.440 700.000 837.040 ;
    END
  END debug_rdata[16]
  PIN debug_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1373.640 700.000 1374.240 ;
    END
  END debug_rdata[17]
  PIN debug_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 547.440 700.000 548.040 ;
    END
  END debug_rdata[18]
  PIN debug_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 357.040 700.000 357.640 ;
    END
  END debug_rdata[19]
  PIN debug_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1883.640 4.000 1884.240 ;
    END
  END debug_rdata[1]
  PIN debug_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END debug_rdata[20]
  PIN debug_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END debug_rdata[21]
  PIN debug_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END debug_rdata[22]
  PIN debug_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END debug_rdata[23]
  PIN debug_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END debug_rdata[24]
  PIN debug_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END debug_rdata[25]
  PIN debug_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1944.840 4.000 1945.440 ;
    END
  END debug_rdata[26]
  PIN debug_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 17.040 700.000 17.640 ;
    END
  END debug_rdata[27]
  PIN debug_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END debug_rdata[28]
  PIN debug_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 948.640 700.000 949.240 ;
    END
  END debug_rdata[29]
  PIN debug_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 193.840 700.000 194.440 ;
    END
  END debug_rdata[2]
  PIN debug_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 2196.000 190.350 2200.000 ;
    END
  END debug_rdata[30]
  PIN debug_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END debug_rdata[31]
  PIN debug_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2196.440 700.000 2197.040 ;
    END
  END debug_rdata[3]
  PIN debug_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END debug_rdata[4]
  PIN debug_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END debug_rdata[5]
  PIN debug_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2111.440 4.000 2112.040 ;
    END
  END debug_rdata[6]
  PIN debug_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 248.240 700.000 248.840 ;
    END
  END debug_rdata[7]
  PIN debug_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END debug_rdata[8]
  PIN debug_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END debug_rdata[9]
  PIN debug_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1533.440 700.000 1534.040 ;
    END
  END debug_req
  PIN debug_rvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1679.640 700.000 1680.240 ;
    END
  END debug_rvalid
  PIN debug_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 68.040 700.000 68.640 ;
    END
  END debug_wdata[0]
  PIN debug_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 629.040 700.000 629.640 ;
    END
  END debug_wdata[10]
  PIN debug_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1798.640 700.000 1799.240 ;
    END
  END debug_wdata[11]
  PIN debug_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END debug_wdata[12]
  PIN debug_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END debug_wdata[13]
  PIN debug_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2043.440 4.000 2044.040 ;
    END
  END debug_wdata[14]
  PIN debug_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END debug_wdata[15]
  PIN debug_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 2196.000 647.590 2200.000 ;
    END
  END debug_wdata[16]
  PIN debug_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 204.040 700.000 204.640 ;
    END
  END debug_wdata[17]
  PIN debug_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 751.440 700.000 752.040 ;
    END
  END debug_wdata[18]
  PIN debug_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 775.240 700.000 775.840 ;
    END
  END debug_wdata[19]
  PIN debug_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END debug_wdata[1]
  PIN debug_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.040 4.000 1649.640 ;
    END
  END debug_wdata[20]
  PIN debug_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1132.240 700.000 1132.840 ;
    END
  END debug_wdata[21]
  PIN debug_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END debug_wdata[22]
  PIN debug_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 2196.000 270.850 2200.000 ;
    END
  END debug_wdata[23]
  PIN debug_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1829.240 700.000 1829.840 ;
    END
  END debug_wdata[24]
  PIN debug_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1700.040 4.000 1700.640 ;
    END
  END debug_wdata[25]
  PIN debug_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2070.640 700.000 2071.240 ;
    END
  END debug_wdata[26]
  PIN debug_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END debug_wdata[27]
  PIN debug_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END debug_wdata[28]
  PIN debug_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 2196.000 293.390 2200.000 ;
    END
  END debug_wdata[29]
  PIN debug_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END debug_wdata[2]
  PIN debug_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 880.640 700.000 881.240 ;
    END
  END debug_wdata[30]
  PIN debug_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END debug_wdata[31]
  PIN debug_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 2196.000 476.930 2200.000 ;
    END
  END debug_wdata[3]
  PIN debug_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END debug_wdata[4]
  PIN debug_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END debug_wdata[5]
  PIN debug_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END debug_wdata[6]
  PIN debug_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END debug_wdata[7]
  PIN debug_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 3.440 700.000 4.040 ;
    END
  END debug_wdata[8]
  PIN debug_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END debug_wdata[9]
  PIN debug_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 2196.000 454.390 2200.000 ;
    END
  END debug_we
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 231.240 700.000 231.840 ;
    END
  END fetch_enable_i
  PIN fetch_enable_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1978.840 4.000 1979.440 ;
    END
  END fetch_enable_o
  PIN fll1_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 537.240 700.000 537.840 ;
    END
  END fll1_ack_i
  PIN fll1_add_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END fll1_add_o[0]
  PIN fll1_add_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1071.040 700.000 1071.640 ;
    END
  END fll1_add_o[1]
  PIN fll1_lock_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END fll1_lock_i
  PIN fll1_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1057.440 700.000 1058.040 ;
    END
  END fll1_rdata_i[0]
  PIN fll1_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 2196.000 222.550 2200.000 ;
    END
  END fll1_rdata_i[10]
  PIN fll1_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END fll1_rdata_i[11]
  PIN fll1_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END fll1_rdata_i[12]
  PIN fll1_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END fll1_rdata_i[13]
  PIN fll1_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1669.440 4.000 1670.040 ;
    END
  END fll1_rdata_i[14]
  PIN fll1_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END fll1_rdata_i[15]
  PIN fll1_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1462.040 700.000 1462.640 ;
    END
  END fll1_rdata_i[16]
  PIN fll1_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END fll1_rdata_i[17]
  PIN fll1_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 2196.000 74.430 2200.000 ;
    END
  END fll1_rdata_i[18]
  PIN fll1_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END fll1_rdata_i[19]
  PIN fll1_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END fll1_rdata_i[1]
  PIN fll1_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2125.040 4.000 2125.640 ;
    END
  END fll1_rdata_i[20]
  PIN fll1_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2012.840 700.000 2013.440 ;
    END
  END fll1_rdata_i[21]
  PIN fll1_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 438.640 700.000 439.240 ;
    END
  END fll1_rdata_i[22]
  PIN fll1_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2108.040 700.000 2108.640 ;
    END
  END fll1_rdata_i[23]
  PIN fll1_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 125.840 700.000 126.440 ;
    END
  END fll1_rdata_i[24]
  PIN fll1_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 13.640 700.000 14.240 ;
    END
  END fll1_rdata_i[25]
  PIN fll1_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 2196.000 132.390 2200.000 ;
    END
  END fll1_rdata_i[26]
  PIN fll1_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2128.440 700.000 2129.040 ;
    END
  END fll1_rdata_i[27]
  PIN fll1_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 2196.000 567.090 2200.000 ;
    END
  END fll1_rdata_i[28]
  PIN fll1_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 2196.000 235.430 2200.000 ;
    END
  END fll1_rdata_i[29]
  PIN fll1_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END fll1_rdata_i[2]
  PIN fll1_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1033.640 700.000 1034.240 ;
    END
  END fll1_rdata_i[30]
  PIN fll1_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1377.040 700.000 1377.640 ;
    END
  END fll1_rdata_i[31]
  PIN fll1_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END fll1_rdata_i[3]
  PIN fll1_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1016.640 700.000 1017.240 ;
    END
  END fll1_rdata_i[4]
  PIN fll1_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END fll1_rdata_i[5]
  PIN fll1_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2162.440 700.000 2163.040 ;
    END
  END fll1_rdata_i[6]
  PIN fll1_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 625.640 700.000 626.240 ;
    END
  END fll1_rdata_i[7]
  PIN fll1_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 493.040 700.000 493.640 ;
    END
  END fll1_rdata_i[8]
  PIN fll1_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END fll1_rdata_i[9]
  PIN fll1_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 156.440 700.000 157.040 ;
    END
  END fll1_req_o
  PIN fll1_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END fll1_wdata_o[0]
  PIN fll1_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 639.240 700.000 639.840 ;
    END
  END fll1_wdata_o[10]
  PIN fll1_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 4.000 1415.040 ;
    END
  END fll1_wdata_o[11]
  PIN fll1_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 513.440 700.000 514.040 ;
    END
  END fll1_wdata_o[12]
  PIN fll1_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END fll1_wdata_o[13]
  PIN fll1_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END fll1_wdata_o[14]
  PIN fll1_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 2196.000 438.290 2200.000 ;
    END
  END fll1_wdata_o[15]
  PIN fll1_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2050.240 700.000 2050.840 ;
    END
  END fll1_wdata_o[16]
  PIN fll1_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 656.240 700.000 656.840 ;
    END
  END fll1_wdata_o[17]
  PIN fll1_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END fll1_wdata_o[18]
  PIN fll1_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END fll1_wdata_o[19]
  PIN fll1_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 2196.000 560.650 2200.000 ;
    END
  END fll1_wdata_o[1]
  PIN fll1_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 2196.000 599.290 2200.000 ;
    END
  END fll1_wdata_o[20]
  PIN fll1_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1278.440 700.000 1279.040 ;
    END
  END fll1_wdata_o[21]
  PIN fll1_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1142.440 700.000 1143.040 ;
    END
  END fll1_wdata_o[22]
  PIN fll1_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END fll1_wdata_o[23]
  PIN fll1_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1621.840 4.000 1622.440 ;
    END
  END fll1_wdata_o[24]
  PIN fll1_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1081.240 700.000 1081.840 ;
    END
  END fll1_wdata_o[25]
  PIN fll1_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END fll1_wdata_o[26]
  PIN fll1_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 2196.000 200.010 2200.000 ;
    END
  END fll1_wdata_o[27]
  PIN fll1_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1771.440 4.000 1772.040 ;
    END
  END fll1_wdata_o[28]
  PIN fll1_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1468.840 700.000 1469.440 ;
    END
  END fll1_wdata_o[29]
  PIN fll1_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1281.840 700.000 1282.440 ;
    END
  END fll1_wdata_o[2]
  PIN fll1_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1441.640 700.000 1442.240 ;
    END
  END fll1_wdata_o[30]
  PIN fll1_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END fll1_wdata_o[31]
  PIN fll1_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1264.840 700.000 1265.440 ;
    END
  END fll1_wdata_o[3]
  PIN fll1_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END fll1_wdata_o[4]
  PIN fll1_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END fll1_wdata_o[5]
  PIN fll1_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2135.240 4.000 2135.840 ;
    END
  END fll1_wdata_o[6]
  PIN fll1_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END fll1_wdata_o[7]
  PIN fll1_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END fll1_wdata_o[8]
  PIN fll1_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END fll1_wdata_o[9]
  PIN fll1_wrn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1812.240 4.000 1812.840 ;
    END
  END fll1_wrn_o
  PIN fll_ack_o_pll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END fll_ack_o_pll
  PIN fll_add_i_pll[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.840 4.000 1520.440 ;
    END
  END fll_add_i_pll[0]
  PIN fll_add_i_pll[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1302.240 700.000 1302.840 ;
    END
  END fll_add_i_pll[1]
  PIN fll_data_i_pll[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END fll_data_i_pll[0]
  PIN fll_data_i_pll[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1431.440 700.000 1432.040 ;
    END
  END fll_data_i_pll[10]
  PIN fll_data_i_pll[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END fll_data_i_pll[11]
  PIN fll_data_i_pll[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1397.440 700.000 1398.040 ;
    END
  END fll_data_i_pll[12]
  PIN fll_data_i_pll[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1781.640 700.000 1782.240 ;
    END
  END fll_data_i_pll[13]
  PIN fll_data_i_pll[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2172.640 700.000 2173.240 ;
    END
  END fll_data_i_pll[14]
  PIN fll_data_i_pll[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END fll_data_i_pll[15]
  PIN fll_data_i_pll[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END fll_data_i_pll[16]
  PIN fll_data_i_pll[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 911.240 700.000 911.840 ;
    END
  END fll_data_i_pll[17]
  PIN fll_data_i_pll[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END fll_data_i_pll[18]
  PIN fll_data_i_pll[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 863.640 700.000 864.240 ;
    END
  END fll_data_i_pll[19]
  PIN fll_data_i_pll[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END fll_data_i_pll[1]
  PIN fll_data_i_pll[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1482.440 700.000 1483.040 ;
    END
  END fll_data_i_pll[20]
  PIN fll_data_i_pll[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END fll_data_i_pll[21]
  PIN fll_data_i_pll[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 2196.000 145.270 2200.000 ;
    END
  END fll_data_i_pll[22]
  PIN fll_data_i_pll[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1876.840 4.000 1877.440 ;
    END
  END fll_data_i_pll[23]
  PIN fll_data_i_pll[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END fll_data_i_pll[24]
  PIN fll_data_i_pll[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 336.640 700.000 337.240 ;
    END
  END fll_data_i_pll[25]
  PIN fll_data_i_pll[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 210.840 700.000 211.440 ;
    END
  END fll_data_i_pll[26]
  PIN fll_data_i_pll[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END fll_data_i_pll[27]
  PIN fll_data_i_pll[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1730.640 4.000 1731.240 ;
    END
  END fll_data_i_pll[28]
  PIN fll_data_i_pll[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1261.440 700.000 1262.040 ;
    END
  END fll_data_i_pll[29]
  PIN fll_data_i_pll[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END fll_data_i_pll[2]
  PIN fll_data_i_pll[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 197.240 700.000 197.840 ;
    END
  END fll_data_i_pll[30]
  PIN fll_data_i_pll[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END fll_data_i_pll[31]
  PIN fll_data_i_pll[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 499.840 700.000 500.440 ;
    END
  END fll_data_i_pll[3]
  PIN fll_data_i_pll[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 2196.000 306.270 2200.000 ;
    END
  END fll_data_i_pll[4]
  PIN fll_data_i_pll[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 992.840 700.000 993.440 ;
    END
  END fll_data_i_pll[5]
  PIN fll_data_i_pll[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END fll_data_i_pll[6]
  PIN fll_data_i_pll[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END fll_data_i_pll[7]
  PIN fll_data_i_pll[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END fll_data_i_pll[8]
  PIN fll_data_i_pll[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1669.440 700.000 1670.040 ;
    END
  END fll_data_i_pll[9]
  PIN fll_lock_o_pll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2067.240 700.000 2067.840 ;
    END
  END fll_lock_o_pll
  PIN fll_r_data_o_pll[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 962.240 700.000 962.840 ;
    END
  END fll_r_data_o_pll[0]
  PIN fll_r_data_o_pll[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END fll_r_data_o_pll[10]
  PIN fll_r_data_o_pll[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1496.040 700.000 1496.640 ;
    END
  END fll_r_data_o_pll[11]
  PIN fll_r_data_o_pll[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1322.640 700.000 1323.240 ;
    END
  END fll_r_data_o_pll[12]
  PIN fll_r_data_o_pll[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 2196.000 203.230 2200.000 ;
    END
  END fll_r_data_o_pll[13]
  PIN fll_r_data_o_pll[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1567.440 700.000 1568.040 ;
    END
  END fll_r_data_o_pll[14]
  PIN fll_r_data_o_pll[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 2196.000 628.270 2200.000 ;
    END
  END fll_r_data_o_pll[15]
  PIN fll_r_data_o_pll[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1873.440 4.000 1874.040 ;
    END
  END fll_r_data_o_pll[16]
  PIN fll_r_data_o_pll[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 108.840 700.000 109.440 ;
    END
  END fll_r_data_o_pll[17]
  PIN fll_r_data_o_pll[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END fll_r_data_o_pll[18]
  PIN fll_r_data_o_pll[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 115.640 700.000 116.240 ;
    END
  END fll_r_data_o_pll[19]
  PIN fll_r_data_o_pll[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2033.240 700.000 2033.840 ;
    END
  END fll_r_data_o_pll[1]
  PIN fll_r_data_o_pll[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1536.840 700.000 1537.440 ;
    END
  END fll_r_data_o_pll[20]
  PIN fll_r_data_o_pll[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END fll_r_data_o_pll[21]
  PIN fll_r_data_o_pll[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END fll_r_data_o_pll[22]
  PIN fll_r_data_o_pll[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1689.840 4.000 1690.440 ;
    END
  END fll_r_data_o_pll[23]
  PIN fll_r_data_o_pll[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END fll_r_data_o_pll[24]
  PIN fll_r_data_o_pll[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END fll_r_data_o_pll[25]
  PIN fll_r_data_o_pll[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END fll_r_data_o_pll[26]
  PIN fll_r_data_o_pll[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END fll_r_data_o_pll[27]
  PIN fll_r_data_o_pll[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END fll_r_data_o_pll[28]
  PIN fll_r_data_o_pll[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END fll_r_data_o_pll[29]
  PIN fll_r_data_o_pll[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END fll_r_data_o_pll[2]
  PIN fll_r_data_o_pll[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END fll_r_data_o_pll[30]
  PIN fll_r_data_o_pll[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 907.840 700.000 908.440 ;
    END
  END fll_r_data_o_pll[31]
  PIN fll_r_data_o_pll[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 2196.000 496.250 2200.000 ;
    END
  END fll_r_data_o_pll[3]
  PIN fll_r_data_o_pll[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END fll_r_data_o_pll[4]
  PIN fll_r_data_o_pll[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1972.040 700.000 1972.640 ;
    END
  END fll_r_data_o_pll[5]
  PIN fll_r_data_o_pll[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END fll_r_data_o_pll[6]
  PIN fll_r_data_o_pll[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END fll_r_data_o_pll[7]
  PIN fll_r_data_o_pll[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END fll_r_data_o_pll[8]
  PIN fll_r_data_o_pll[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1914.240 700.000 1914.840 ;
    END
  END fll_r_data_o_pll[9]
  PIN fll_req_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 2196.000 122.730 2200.000 ;
    END
  END fll_req_i_pll
  PIN fll_wrn_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 904.440 700.000 905.040 ;
    END
  END fll_wrn_i_pll
  PIN gpio_dir[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END gpio_dir[0]
  PIN gpio_dir[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1856.440 700.000 1857.040 ;
    END
  END gpio_dir[10]
  PIN gpio_dir[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END gpio_dir[11]
  PIN gpio_dir[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END gpio_dir[12]
  PIN gpio_dir[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 102.040 700.000 102.640 ;
    END
  END gpio_dir[13]
  PIN gpio_dir[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 578.040 700.000 578.640 ;
    END
  END gpio_dir[14]
  PIN gpio_dir[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1407.640 700.000 1408.240 ;
    END
  END gpio_dir[15]
  PIN gpio_dir[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1047.240 700.000 1047.840 ;
    END
  END gpio_dir[16]
  PIN gpio_dir[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END gpio_dir[17]
  PIN gpio_dir[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 2196.000 154.930 2200.000 ;
    END
  END gpio_dir[18]
  PIN gpio_dir[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END gpio_dir[19]
  PIN gpio_dir[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1689.840 700.000 1690.440 ;
    END
  END gpio_dir[1]
  PIN gpio_dir[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1842.840 700.000 1843.440 ;
    END
  END gpio_dir[20]
  PIN gpio_dir[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 2196.000 699.110 2200.000 ;
    END
  END gpio_dir[21]
  PIN gpio_dir[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END gpio_dir[22]
  PIN gpio_dir[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 2196.000 32.570 2200.000 ;
    END
  END gpio_dir[23]
  PIN gpio_dir[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END gpio_dir[24]
  PIN gpio_dir[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END gpio_dir[25]
  PIN gpio_dir[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END gpio_dir[26]
  PIN gpio_dir[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1193.440 700.000 1194.040 ;
    END
  END gpio_dir[27]
  PIN gpio_dir[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END gpio_dir[28]
  PIN gpio_dir[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1604.840 700.000 1605.440 ;
    END
  END gpio_dir[29]
  PIN gpio_dir[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 2196.000 19.690 2200.000 ;
    END
  END gpio_dir[2]
  PIN gpio_dir[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END gpio_dir[30]
  PIN gpio_dir[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 931.640 700.000 932.240 ;
    END
  END gpio_dir[31]
  PIN gpio_dir[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 642.640 700.000 643.240 ;
    END
  END gpio_dir[3]
  PIN gpio_dir[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2019.640 4.000 2020.240 ;
    END
  END gpio_dir[4]
  PIN gpio_dir[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1764.640 4.000 1765.240 ;
    END
  END gpio_dir[5]
  PIN gpio_dir[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END gpio_dir[6]
  PIN gpio_dir[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END gpio_dir[7]
  PIN gpio_dir[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END gpio_dir[8]
  PIN gpio_dir[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END gpio_dir[9]
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 853.440 700.000 854.040 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 503.240 700.000 503.840 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 2196.000 71.210 2200.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1703.440 700.000 1704.040 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 74.840 700.000 75.440 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 2196.000 396.430 2200.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1587.840 700.000 1588.440 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1730.640 700.000 1731.240 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 2196.000 579.970 2200.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 265.240 700.000 265.840 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1941.440 700.000 1942.040 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 30.640 700.000 31.240 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 91.840 700.000 92.440 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 2196.000 125.950 2200.000 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 2196.000 386.770 2200.000 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1210.440 4.000 1211.040 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END gpio_in[31]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1632.040 700.000 1632.640 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 251.640 700.000 252.240 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1258.040 700.000 1258.640 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1842.840 4.000 1843.440 ;
    END
  END gpio_in[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 2196.000 354.570 2200.000 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1067.640 700.000 1068.240 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 2196.000 451.170 2200.000 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2070.640 4.000 2071.240 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1754.440 700.000 1755.040 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1584.440 700.000 1585.040 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 2196.000 290.170 2200.000 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 819.440 700.000 820.040 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1349.840 700.000 1350.440 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1244.440 700.000 1245.040 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1785.040 4.000 1785.640 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 2196.000 93.750 2200.000 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1312.440 700.000 1313.040 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 418.240 700.000 418.840 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1897.240 4.000 1897.840 ;
    END
  END gpio_out[31]
  PIN gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 2196.000 502.690 2200.000 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 411.440 700.000 412.040 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1292.040 700.000 1292.640 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2012.840 4.000 2013.440 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1863.240 700.000 1863.840 ;
    END
  END gpio_out[9]
  PIN gpio_padcfg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1009.840 700.000 1010.440 ;
    END
  END gpio_padcfg[0]
  PIN gpio_padcfg[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 227.840 700.000 228.440 ;
    END
  END gpio_padcfg[100]
  PIN gpio_padcfg[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1203.640 700.000 1204.240 ;
    END
  END gpio_padcfg[101]
  PIN gpio_padcfg[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END gpio_padcfg[102]
  PIN gpio_padcfg[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END gpio_padcfg[103]
  PIN gpio_padcfg[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 649.440 700.000 650.040 ;
    END
  END gpio_padcfg[104]
  PIN gpio_padcfg[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 2196.000 370.670 2200.000 ;
    END
  END gpio_padcfg[105]
  PIN gpio_padcfg[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END gpio_padcfg[106]
  PIN gpio_padcfg[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END gpio_padcfg[107]
  PIN gpio_padcfg[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2111.440 700.000 2112.040 ;
    END
  END gpio_padcfg[108]
  PIN gpio_padcfg[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END gpio_padcfg[109]
  PIN gpio_padcfg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END gpio_padcfg[10]
  PIN gpio_padcfg[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2176.040 700.000 2176.640 ;
    END
  END gpio_padcfg[110]
  PIN gpio_padcfg[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 2196.000 274.070 2200.000 ;
    END
  END gpio_padcfg[111]
  PIN gpio_padcfg[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 163.240 700.000 163.840 ;
    END
  END gpio_padcfg[112]
  PIN gpio_padcfg[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1713.640 4.000 1714.240 ;
    END
  END gpio_padcfg[113]
  PIN gpio_padcfg[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END gpio_padcfg[114]
  PIN gpio_padcfg[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END gpio_padcfg[115]
  PIN gpio_padcfg[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1207.040 700.000 1207.640 ;
    END
  END gpio_padcfg[116]
  PIN gpio_padcfg[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END gpio_padcfg[117]
  PIN gpio_padcfg[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 2196.000 322.370 2200.000 ;
    END
  END gpio_padcfg[118]
  PIN gpio_padcfg[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END gpio_padcfg[119]
  PIN gpio_padcfg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END gpio_padcfg[11]
  PIN gpio_padcfg[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2179.440 4.000 2180.040 ;
    END
  END gpio_padcfg[120]
  PIN gpio_padcfg[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END gpio_padcfg[121]
  PIN gpio_padcfg[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END gpio_padcfg[122]
  PIN gpio_padcfg[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END gpio_padcfg[123]
  PIN gpio_padcfg[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 2196.000 64.770 2200.000 ;
    END
  END gpio_padcfg[124]
  PIN gpio_padcfg[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END gpio_padcfg[125]
  PIN gpio_padcfg[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 2196.000 383.550 2200.000 ;
    END
  END gpio_padcfg[126]
  PIN gpio_padcfg[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2169.240 4.000 2169.840 ;
    END
  END gpio_padcfg[127]
  PIN gpio_padcfg[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 2196.000 660.470 2200.000 ;
    END
  END gpio_padcfg[128]
  PIN gpio_padcfg[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2063.840 700.000 2064.440 ;
    END
  END gpio_padcfg[129]
  PIN gpio_padcfg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END gpio_padcfg[12]
  PIN gpio_padcfg[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END gpio_padcfg[130]
  PIN gpio_padcfg[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1091.440 700.000 1092.040 ;
    END
  END gpio_padcfg[131]
  PIN gpio_padcfg[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2019.640 700.000 2020.240 ;
    END
  END gpio_padcfg[132]
  PIN gpio_padcfg[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1666.040 700.000 1666.640 ;
    END
  END gpio_padcfg[133]
  PIN gpio_padcfg[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 860.240 700.000 860.840 ;
    END
  END gpio_padcfg[134]
  PIN gpio_padcfg[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 2196.000 522.010 2200.000 ;
    END
  END gpio_padcfg[135]
  PIN gpio_padcfg[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END gpio_padcfg[136]
  PIN gpio_padcfg[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END gpio_padcfg[137]
  PIN gpio_padcfg[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1159.440 700.000 1160.040 ;
    END
  END gpio_padcfg[138]
  PIN gpio_padcfg[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 952.040 700.000 952.640 ;
    END
  END gpio_padcfg[139]
  PIN gpio_padcfg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 408.040 700.000 408.640 ;
    END
  END gpio_padcfg[13]
  PIN gpio_padcfg[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 2196.000 554.210 2200.000 ;
    END
  END gpio_padcfg[140]
  PIN gpio_padcfg[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 965.640 700.000 966.240 ;
    END
  END gpio_padcfg[141]
  PIN gpio_padcfg[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END gpio_padcfg[142]
  PIN gpio_padcfg[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2057.040 700.000 2057.640 ;
    END
  END gpio_padcfg[143]
  PIN gpio_padcfg[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 2196.000 563.870 2200.000 ;
    END
  END gpio_padcfg[144]
  PIN gpio_padcfg[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END gpio_padcfg[145]
  PIN gpio_padcfg[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2155.640 4.000 2156.240 ;
    END
  END gpio_padcfg[146]
  PIN gpio_padcfg[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END gpio_padcfg[147]
  PIN gpio_padcfg[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2091.040 700.000 2091.640 ;
    END
  END gpio_padcfg[148]
  PIN gpio_padcfg[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1186.640 700.000 1187.240 ;
    END
  END gpio_padcfg[149]
  PIN gpio_padcfg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END gpio_padcfg[14]
  PIN gpio_padcfg[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END gpio_padcfg[150]
  PIN gpio_padcfg[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2053.640 4.000 2054.240 ;
    END
  END gpio_padcfg[151]
  PIN gpio_padcfg[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END gpio_padcfg[152]
  PIN gpio_padcfg[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 2196.000 96.970 2200.000 ;
    END
  END gpio_padcfg[153]
  PIN gpio_padcfg[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1251.240 700.000 1251.840 ;
    END
  END gpio_padcfg[154]
  PIN gpio_padcfg[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 894.240 700.000 894.840 ;
    END
  END gpio_padcfg[155]
  PIN gpio_padcfg[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END gpio_padcfg[156]
  PIN gpio_padcfg[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 778.640 700.000 779.240 ;
    END
  END gpio_padcfg[157]
  PIN gpio_padcfg[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 788.840 700.000 789.440 ;
    END
  END gpio_padcfg[158]
  PIN gpio_padcfg[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2104.640 700.000 2105.240 ;
    END
  END gpio_padcfg[159]
  PIN gpio_padcfg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1166.240 700.000 1166.840 ;
    END
  END gpio_padcfg[15]
  PIN gpio_padcfg[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 2196.000 3.590 2200.000 ;
    END
  END gpio_padcfg[160]
  PIN gpio_padcfg[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END gpio_padcfg[161]
  PIN gpio_padcfg[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 54.440 700.000 55.040 ;
    END
  END gpio_padcfg[162]
  PIN gpio_padcfg[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 2196.000 277.290 2200.000 ;
    END
  END gpio_padcfg[163]
  PIN gpio_padcfg[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1982.240 700.000 1982.840 ;
    END
  END gpio_padcfg[164]
  PIN gpio_padcfg[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1213.840 700.000 1214.440 ;
    END
  END gpio_padcfg[165]
  PIN gpio_padcfg[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2182.840 700.000 2183.440 ;
    END
  END gpio_padcfg[166]
  PIN gpio_padcfg[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1156.040 700.000 1156.640 ;
    END
  END gpio_padcfg[167]
  PIN gpio_padcfg[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 2196.000 480.150 2200.000 ;
    END
  END gpio_padcfg[168]
  PIN gpio_padcfg[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 486.240 700.000 486.840 ;
    END
  END gpio_padcfg[169]
  PIN gpio_padcfg[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END gpio_padcfg[16]
  PIN gpio_padcfg[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END gpio_padcfg[170]
  PIN gpio_padcfg[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 697.040 700.000 697.640 ;
    END
  END gpio_padcfg[171]
  PIN gpio_padcfg[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END gpio_padcfg[172]
  PIN gpio_padcfg[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1815.640 4.000 1816.240 ;
    END
  END gpio_padcfg[173]
  PIN gpio_padcfg[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 2196.000 296.610 2200.000 ;
    END
  END gpio_padcfg[174]
  PIN gpio_padcfg[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1774.840 700.000 1775.440 ;
    END
  END gpio_padcfg[175]
  PIN gpio_padcfg[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 795.640 700.000 796.240 ;
    END
  END gpio_padcfg[176]
  PIN gpio_padcfg[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1645.640 700.000 1646.240 ;
    END
  END gpio_padcfg[177]
  PIN gpio_padcfg[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END gpio_padcfg[178]
  PIN gpio_padcfg[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END gpio_padcfg[179]
  PIN gpio_padcfg[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 748.040 700.000 748.640 ;
    END
  END gpio_padcfg[17]
  PIN gpio_padcfg[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 2196.000 116.290 2200.000 ;
    END
  END gpio_padcfg[180]
  PIN gpio_padcfg[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END gpio_padcfg[181]
  PIN gpio_padcfg[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END gpio_padcfg[182]
  PIN gpio_padcfg[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1961.840 700.000 1962.440 ;
    END
  END gpio_padcfg[183]
  PIN gpio_padcfg[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 241.440 700.000 242.040 ;
    END
  END gpio_padcfg[184]
  PIN gpio_padcfg[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 2196.000 103.410 2200.000 ;
    END
  END gpio_padcfg[185]
  PIN gpio_padcfg[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END gpio_padcfg[186]
  PIN gpio_padcfg[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END gpio_padcfg[187]
  PIN gpio_padcfg[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 2196.000 212.890 2200.000 ;
    END
  END gpio_padcfg[188]
  PIN gpio_padcfg[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END gpio_padcfg[189]
  PIN gpio_padcfg[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 346.840 700.000 347.440 ;
    END
  END gpio_padcfg[18]
  PIN gpio_padcfg[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio_padcfg[190]
  PIN gpio_padcfg[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1798.640 4.000 1799.240 ;
    END
  END gpio_padcfg[191]
  PIN gpio_padcfg[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END gpio_padcfg[19]
  PIN gpio_padcfg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END gpio_padcfg[1]
  PIN gpio_padcfg[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END gpio_padcfg[20]
  PIN gpio_padcfg[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END gpio_padcfg[21]
  PIN gpio_padcfg[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END gpio_padcfg[22]
  PIN gpio_padcfg[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END gpio_padcfg[23]
  PIN gpio_padcfg[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 608.640 700.000 609.240 ;
    END
  END gpio_padcfg[24]
  PIN gpio_padcfg[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END gpio_padcfg[25]
  PIN gpio_padcfg[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1234.240 700.000 1234.840 ;
    END
  END gpio_padcfg[26]
  PIN gpio_padcfg[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 666.440 700.000 667.040 ;
    END
  END gpio_padcfg[27]
  PIN gpio_padcfg[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1054.040 700.000 1054.640 ;
    END
  END gpio_padcfg[28]
  PIN gpio_padcfg[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1390.640 700.000 1391.240 ;
    END
  END gpio_padcfg[29]
  PIN gpio_padcfg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1652.440 700.000 1653.040 ;
    END
  END gpio_padcfg[2]
  PIN gpio_padcfg[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 938.440 700.000 939.040 ;
    END
  END gpio_padcfg[30]
  PIN gpio_padcfg[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 2196.000 541.330 2200.000 ;
    END
  END gpio_padcfg[31]
  PIN gpio_padcfg[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 2196.000 84.090 2200.000 ;
    END
  END gpio_padcfg[32]
  PIN gpio_padcfg[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gpio_padcfg[33]
  PIN gpio_padcfg[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END gpio_padcfg[34]
  PIN gpio_padcfg[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END gpio_padcfg[35]
  PIN gpio_padcfg[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END gpio_padcfg[36]
  PIN gpio_padcfg[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END gpio_padcfg[37]
  PIN gpio_padcfg[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END gpio_padcfg[38]
  PIN gpio_padcfg[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1064.240 700.000 1064.840 ;
    END
  END gpio_padcfg[39]
  PIN gpio_padcfg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END gpio_padcfg[3]
  PIN gpio_padcfg[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 78.240 700.000 78.840 ;
    END
  END gpio_padcfg[40]
  PIN gpio_padcfg[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 714.040 700.000 714.640 ;
    END
  END gpio_padcfg[41]
  PIN gpio_padcfg[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END gpio_padcfg[42]
  PIN gpio_padcfg[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 2196.000 618.610 2200.000 ;
    END
  END gpio_padcfg[43]
  PIN gpio_padcfg[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END gpio_padcfg[44]
  PIN gpio_padcfg[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END gpio_padcfg[45]
  PIN gpio_padcfg[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 612.040 700.000 612.640 ;
    END
  END gpio_padcfg[46]
  PIN gpio_padcfg[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1543.640 700.000 1544.240 ;
    END
  END gpio_padcfg[47]
  PIN gpio_padcfg[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1574.240 700.000 1574.840 ;
    END
  END gpio_padcfg[48]
  PIN gpio_padcfg[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 683.440 700.000 684.040 ;
    END
  END gpio_padcfg[49]
  PIN gpio_padcfg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1679.640 4.000 1680.240 ;
    END
  END gpio_padcfg[4]
  PIN gpio_padcfg[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END gpio_padcfg[50]
  PIN gpio_padcfg[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END gpio_padcfg[51]
  PIN gpio_padcfg[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END gpio_padcfg[52]
  PIN gpio_padcfg[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gpio_padcfg[53]
  PIN gpio_padcfg[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END gpio_padcfg[54]
  PIN gpio_padcfg[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1618.440 4.000 1619.040 ;
    END
  END gpio_padcfg[55]
  PIN gpio_padcfg[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1764.640 700.000 1765.240 ;
    END
  END gpio_padcfg[56]
  PIN gpio_padcfg[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END gpio_padcfg[57]
  PIN gpio_padcfg[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.240 4.000 1574.840 ;
    END
  END gpio_padcfg[58]
  PIN gpio_padcfg[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1900.640 4.000 1901.240 ;
    END
  END gpio_padcfg[59]
  PIN gpio_padcfg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 2196.000 80.870 2200.000 ;
    END
  END gpio_padcfg[5]
  PIN gpio_padcfg[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1948.240 700.000 1948.840 ;
    END
  END gpio_padcfg[60]
  PIN gpio_padcfg[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END gpio_padcfg[61]
  PIN gpio_padcfg[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.840 4.000 1282.440 ;
    END
  END gpio_padcfg[62]
  PIN gpio_padcfg[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1686.440 700.000 1687.040 ;
    END
  END gpio_padcfg[63]
  PIN gpio_padcfg[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END gpio_padcfg[64]
  PIN gpio_padcfg[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 2196.000 357.790 2200.000 ;
    END
  END gpio_padcfg[65]
  PIN gpio_padcfg[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1615.040 4.000 1615.640 ;
    END
  END gpio_padcfg[66]
  PIN gpio_padcfg[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END gpio_padcfg[67]
  PIN gpio_padcfg[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1737.440 700.000 1738.040 ;
    END
  END gpio_padcfg[68]
  PIN gpio_padcfg[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END gpio_padcfg[69]
  PIN gpio_padcfg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1438.240 700.000 1438.840 ;
    END
  END gpio_padcfg[6]
  PIN gpio_padcfg[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1659.240 700.000 1659.840 ;
    END
  END gpio_padcfg[70]
  PIN gpio_padcfg[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1111.840 700.000 1112.440 ;
    END
  END gpio_padcfg[71]
  PIN gpio_padcfg[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 669.840 700.000 670.440 ;
    END
  END gpio_padcfg[72]
  PIN gpio_padcfg[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END gpio_padcfg[73]
  PIN gpio_padcfg[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END gpio_padcfg[74]
  PIN gpio_padcfg[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpio_padcfg[75]
  PIN gpio_padcfg[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 2196.000 35.790 2200.000 ;
    END
  END gpio_padcfg[76]
  PIN gpio_padcfg[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END gpio_padcfg[77]
  PIN gpio_padcfg[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END gpio_padcfg[78]
  PIN gpio_padcfg[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1414.440 700.000 1415.040 ;
    END
  END gpio_padcfg[79]
  PIN gpio_padcfg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END gpio_padcfg[7]
  PIN gpio_padcfg[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 6.840 700.000 7.440 ;
    END
  END gpio_padcfg[80]
  PIN gpio_padcfg[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 2196.000 0.370 2200.000 ;
    END
  END gpio_padcfg[81]
  PIN gpio_padcfg[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1938.040 700.000 1938.640 ;
    END
  END gpio_padcfg[82]
  PIN gpio_padcfg[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END gpio_padcfg[83]
  PIN gpio_padcfg[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1077.840 700.000 1078.440 ;
    END
  END gpio_padcfg[84]
  PIN gpio_padcfg[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END gpio_padcfg[85]
  PIN gpio_padcfg[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END gpio_padcfg[86]
  PIN gpio_padcfg[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1139.040 700.000 1139.640 ;
    END
  END gpio_padcfg[87]
  PIN gpio_padcfg[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 520.240 700.000 520.840 ;
    END
  END gpio_padcfg[88]
  PIN gpio_padcfg[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 323.040 700.000 323.640 ;
    END
  END gpio_padcfg[89]
  PIN gpio_padcfg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END gpio_padcfg[8]
  PIN gpio_padcfg[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END gpio_padcfg[90]
  PIN gpio_padcfg[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END gpio_padcfg[91]
  PIN gpio_padcfg[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 139.440 700.000 140.040 ;
    END
  END gpio_padcfg[92]
  PIN gpio_padcfg[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END gpio_padcfg[93]
  PIN gpio_padcfg[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.840 4.000 1673.440 ;
    END
  END gpio_padcfg[94]
  PIN gpio_padcfg[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1346.440 700.000 1347.040 ;
    END
  END gpio_padcfg[95]
  PIN gpio_padcfg[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 2196.000 673.350 2200.000 ;
    END
  END gpio_padcfg[96]
  PIN gpio_padcfg[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END gpio_padcfg[97]
  PIN gpio_padcfg[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 2196.000 180.690 2200.000 ;
    END
  END gpio_padcfg[98]
  PIN gpio_padcfg[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END gpio_padcfg[99]
  PIN gpio_padcfg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END gpio_padcfg[9]
  PIN io_oeb_pll[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 918.040 700.000 918.640 ;
    END
  END io_oeb_pll[0]
  PIN io_oeb_pll[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END io_oeb_pll[10]
  PIN io_oeb_pll[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_oeb_pll[11]
  PIN io_oeb_pll[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END io_oeb_pll[12]
  PIN io_oeb_pll[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1326.040 700.000 1326.640 ;
    END
  END io_oeb_pll[13]
  PIN io_oeb_pll[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 826.240 700.000 826.840 ;
    END
  END io_oeb_pll[14]
  PIN io_oeb_pll[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_oeb_pll[15]
  PIN io_oeb_pll[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1336.240 700.000 1336.840 ;
    END
  END io_oeb_pll[16]
  PIN io_oeb_pll[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 4.000 2118.840 ;
    END
  END io_oeb_pll[17]
  PIN io_oeb_pll[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END io_oeb_pll[18]
  PIN io_oeb_pll[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 476.040 700.000 476.640 ;
    END
  END io_oeb_pll[19]
  PIN io_oeb_pll[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 2196.000 457.610 2200.000 ;
    END
  END io_oeb_pll[1]
  PIN io_oeb_pll[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 2196.000 441.510 2200.000 ;
    END
  END io_oeb_pll[20]
  PIN io_oeb_pll[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END io_oeb_pll[21]
  PIN io_oeb_pll[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END io_oeb_pll[22]
  PIN io_oeb_pll[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 693.640 700.000 694.240 ;
    END
  END io_oeb_pll[23]
  PIN io_oeb_pll[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1802.040 700.000 1802.640 ;
    END
  END io_oeb_pll[24]
  PIN io_oeb_pll[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END io_oeb_pll[25]
  PIN io_oeb_pll[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1621.840 700.000 1622.440 ;
    END
  END io_oeb_pll[26]
  PIN io_oeb_pll[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END io_oeb_pll[27]
  PIN io_oeb_pll[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_oeb_pll[28]
  PIN io_oeb_pll[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_oeb_pll[29]
  PIN io_oeb_pll[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1088.040 700.000 1088.640 ;
    END
  END io_oeb_pll[2]
  PIN io_oeb_pll[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_oeb_pll[30]
  PIN io_oeb_pll[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1128.840 700.000 1129.440 ;
    END
  END io_oeb_pll[31]
  PIN io_oeb_pll[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END io_oeb_pll[32]
  PIN io_oeb_pll[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END io_oeb_pll[33]
  PIN io_oeb_pll[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1502.840 700.000 1503.440 ;
    END
  END io_oeb_pll[34]
  PIN io_oeb_pll[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 2196.000 464.050 2200.000 ;
    END
  END io_oeb_pll[35]
  PIN io_oeb_pll[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 200.640 700.000 201.240 ;
    END
  END io_oeb_pll[36]
  PIN io_oeb_pll[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2189.640 4.000 2190.240 ;
    END
  END io_oeb_pll[37]
  PIN io_oeb_pll[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END io_oeb_pll[3]
  PIN io_oeb_pll[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 2196.000 657.250 2200.000 ;
    END
  END io_oeb_pll[4]
  PIN io_oeb_pll[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1958.440 4.000 1959.040 ;
    END
  END io_oeb_pll[5]
  PIN io_oeb_pll[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 343.440 700.000 344.040 ;
    END
  END io_oeb_pll[6]
  PIN io_oeb_pll[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1305.640 700.000 1306.240 ;
    END
  END io_oeb_pll[7]
  PIN io_oeb_pll[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 588.240 700.000 588.840 ;
    END
  END io_oeb_pll[8]
  PIN io_oeb_pll[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1887.040 700.000 1887.640 ;
    END
  END io_oeb_pll[9]
  PIN io_out_pll[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1866.640 700.000 1867.240 ;
    END
  END io_out_pll[0]
  PIN io_out_pll[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END io_out_pll[10]
  PIN io_out_pll[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1853.040 700.000 1853.640 ;
    END
  END io_out_pll[11]
  PIN io_out_pll[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END io_out_pll[12]
  PIN io_out_pll[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2023.040 700.000 2023.640 ;
    END
  END io_out_pll[13]
  PIN io_out_pll[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END io_out_pll[14]
  PIN io_out_pll[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 2196.000 377.110 2200.000 ;
    END
  END io_out_pll[15]
  PIN io_out_pll[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 363.840 700.000 364.440 ;
    END
  END io_out_pll[16]
  PIN io_out_pll[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1200.240 700.000 1200.840 ;
    END
  END io_out_pll[17]
  PIN io_out_pll[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 207.440 700.000 208.040 ;
    END
  END io_out_pll[18]
  PIN io_out_pll[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END io_out_pll[19]
  PIN io_out_pll[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 605.240 700.000 605.840 ;
    END
  END io_out_pll[1]
  PIN io_out_pll[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2152.240 4.000 2152.840 ;
    END
  END io_out_pll[20]
  PIN io_out_pll[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1788.440 700.000 1789.040 ;
    END
  END io_out_pll[21]
  PIN io_out_pll[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1577.640 700.000 1578.240 ;
    END
  END io_out_pll[22]
  PIN io_out_pll[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 47.640 700.000 48.240 ;
    END
  END io_out_pll[23]
  PIN io_out_pll[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END io_out_pll[24]
  PIN io_out_pll[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_out_pll[25]
  PIN io_out_pll[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_out_pll[2]
  PIN io_out_pll[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 2196.000 142.050 2200.000 ;
    END
  END io_out_pll[3]
  PIN io_out_pll[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1900.640 700.000 1901.240 ;
    END
  END io_out_pll[4]
  PIN io_out_pll[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 2196.000 444.730 2200.000 ;
    END
  END io_out_pll[5]
  PIN io_out_pll[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 2196.000 113.070 2200.000 ;
    END
  END io_out_pll[6]
  PIN io_out_pll[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1581.040 4.000 1581.640 ;
    END
  END io_out_pll[7]
  PIN io_out_pll[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1383.840 700.000 1384.440 ;
    END
  END io_out_pll[8]
  PIN io_out_pll[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END io_out_pll[9]
  PIN irq_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END irq_o[0]
  PIN irq_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1115.240 700.000 1115.840 ;
    END
  END irq_o[10]
  PIN irq_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 472.640 700.000 473.240 ;
    END
  END irq_o[11]
  PIN irq_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 285.640 700.000 286.240 ;
    END
  END irq_o[12]
  PIN irq_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 2196.000 393.210 2200.000 ;
    END
  END irq_o[13]
  PIN irq_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END irq_o[14]
  PIN irq_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 737.840 700.000 738.440 ;
    END
  END irq_o[15]
  PIN irq_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 435.240 700.000 435.840 ;
    END
  END irq_o[16]
  PIN irq_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.040 4.000 1530.640 ;
    END
  END irq_o[17]
  PIN irq_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END irq_o[18]
  PIN irq_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END irq_o[19]
  PIN irq_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1604.840 4.000 1605.440 ;
    END
  END irq_o[1]
  PIN irq_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END irq_o[20]
  PIN irq_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1475.640 700.000 1476.240 ;
    END
  END irq_o[21]
  PIN irq_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END irq_o[22]
  PIN irq_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1404.240 700.000 1404.840 ;
    END
  END irq_o[23]
  PIN irq_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END irq_o[24]
  PIN irq_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END irq_o[25]
  PIN irq_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 2196.000 61.550 2200.000 ;
    END
  END irq_o[26]
  PIN irq_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END irq_o[27]
  PIN irq_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END irq_o[28]
  PIN irq_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2179.440 700.000 2180.040 ;
    END
  END irq_o[29]
  PIN irq_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END irq_o[2]
  PIN irq_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END irq_o[30]
  PIN irq_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 2196.000 90.530 2200.000 ;
    END
  END irq_o[31]
  PIN irq_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 353.640 700.000 354.240 ;
    END
  END irq_o[3]
  PIN irq_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2131.840 4.000 2132.440 ;
    END
  END irq_o[4]
  PIN irq_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1101.640 700.000 1102.240 ;
    END
  END irq_o[5]
  PIN irq_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END irq_o[6]
  PIN irq_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1961.840 4.000 1962.440 ;
    END
  END irq_o[7]
  PIN irq_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END irq_o[8]
  PIN irq_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END irq_o[9]
  PIN la_data_out_pll[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1808.840 700.000 1809.440 ;
    END
  END la_data_out_pll[0]
  PIN la_data_out_pll[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 2196.000 605.730 2200.000 ;
    END
  END la_data_out_pll[10]
  PIN la_data_out_pll[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END la_data_out_pll[11]
  PIN la_data_out_pll[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1523.240 700.000 1523.840 ;
    END
  END la_data_out_pll[12]
  PIN la_data_out_pll[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END la_data_out_pll[13]
  PIN la_data_out_pll[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1241.040 700.000 1241.640 ;
    END
  END la_data_out_pll[14]
  PIN la_data_out_pll[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2131.840 700.000 2132.440 ;
    END
  END la_data_out_pll[15]
  PIN la_data_out_pll[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 173.440 700.000 174.040 ;
    END
  END la_data_out_pll[16]
  PIN la_data_out_pll[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.840 4.000 1418.440 ;
    END
  END la_data_out_pll[17]
  PIN la_data_out_pll[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 2196.000 219.330 2200.000 ;
    END
  END la_data_out_pll[18]
  PIN la_data_out_pll[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1224.040 700.000 1224.640 ;
    END
  END la_data_out_pll[19]
  PIN la_data_out_pll[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END la_data_out_pll[1]
  PIN la_data_out_pll[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END la_data_out_pll[20]
  PIN la_data_out_pll[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1839.440 700.000 1840.040 ;
    END
  END la_data_out_pll[21]
  PIN la_data_out_pll[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1271.640 700.000 1272.240 ;
    END
  END la_data_out_pll[22]
  PIN la_data_out_pll[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 663.040 700.000 663.640 ;
    END
  END la_data_out_pll[23]
  PIN la_data_out_pll[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END la_data_out_pll[24]
  PIN la_data_out_pll[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END la_data_out_pll[25]
  PIN la_data_out_pll[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1795.240 700.000 1795.840 ;
    END
  END la_data_out_pll[26]
  PIN la_data_out_pll[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 2196.000 29.350 2200.000 ;
    END
  END la_data_out_pll[27]
  PIN la_data_out_pll[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 2196.000 77.650 2200.000 ;
    END
  END la_data_out_pll[28]
  PIN la_data_out_pll[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1220.640 700.000 1221.240 ;
    END
  END la_data_out_pll[29]
  PIN la_data_out_pll[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END la_data_out_pll[2]
  PIN la_data_out_pll[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1921.040 4.000 1921.640 ;
    END
  END la_data_out_pll[30]
  PIN la_data_out_pll[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1941.440 4.000 1942.040 ;
    END
  END la_data_out_pll[31]
  PIN la_data_out_pll[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1649.040 700.000 1649.640 ;
    END
  END la_data_out_pll[32]
  PIN la_data_out_pll[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_data_out_pll[33]
  PIN la_data_out_pll[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END la_data_out_pll[34]
  PIN la_data_out_pll[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END la_data_out_pll[35]
  PIN la_data_out_pll[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END la_data_out_pll[36]
  PIN la_data_out_pll[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 754.840 700.000 755.440 ;
    END
  END la_data_out_pll[37]
  PIN la_data_out_pll[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1329.440 700.000 1330.040 ;
    END
  END la_data_out_pll[38]
  PIN la_data_out_pll[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_out_pll[39]
  PIN la_data_out_pll[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1472.240 700.000 1472.840 ;
    END
  END la_data_out_pll[3]
  PIN la_data_out_pll[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1581.040 700.000 1581.640 ;
    END
  END la_data_out_pll[40]
  PIN la_data_out_pll[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 516.840 700.000 517.440 ;
    END
  END la_data_out_pll[41]
  PIN la_data_out_pll[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1951.640 700.000 1952.240 ;
    END
  END la_data_out_pll[42]
  PIN la_data_out_pll[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 2196.000 683.010 2200.000 ;
    END
  END la_data_out_pll[43]
  PIN la_data_out_pll[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 2196.000 183.910 2200.000 ;
    END
  END la_data_out_pll[44]
  PIN la_data_out_pll[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END la_data_out_pll[45]
  PIN la_data_out_pll[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1927.840 700.000 1928.440 ;
    END
  END la_data_out_pll[46]
  PIN la_data_out_pll[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 768.440 700.000 769.040 ;
    END
  END la_data_out_pll[47]
  PIN la_data_out_pll[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END la_data_out_pll[48]
  PIN la_data_out_pll[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_data_out_pll[49]
  PIN la_data_out_pll[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 601.840 700.000 602.440 ;
    END
  END la_data_out_pll[4]
  PIN la_data_out_pll[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1298.840 700.000 1299.440 ;
    END
  END la_data_out_pll[50]
  PIN la_data_out_pll[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 238.040 700.000 238.640 ;
    END
  END la_data_out_pll[51]
  PIN la_data_out_pll[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END la_data_out_pll[52]
  PIN la_data_out_pll[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 2196.000 692.670 2200.000 ;
    END
  END la_data_out_pll[53]
  PIN la_data_out_pll[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_data_out_pll[54]
  PIN la_data_out_pll[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 187.040 700.000 187.640 ;
    END
  END la_data_out_pll[55]
  PIN la_data_out_pll[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1744.240 4.000 1744.840 ;
    END
  END la_data_out_pll[56]
  PIN la_data_out_pll[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1968.640 700.000 1969.240 ;
    END
  END la_data_out_pll[57]
  PIN la_data_out_pll[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1122.040 700.000 1122.640 ;
    END
  END la_data_out_pll[58]
  PIN la_data_out_pll[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2142.040 700.000 2142.640 ;
    END
  END la_data_out_pll[59]
  PIN la_data_out_pll[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1285.240 700.000 1285.840 ;
    END
  END la_data_out_pll[5]
  PIN la_data_out_pll[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1547.040 700.000 1547.640 ;
    END
  END la_data_out_pll[60]
  PIN la_data_out_pll[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 533.840 700.000 534.440 ;
    END
  END la_data_out_pll[61]
  PIN la_data_out_pll[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END la_data_out_pll[62]
  PIN la_data_out_pll[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END la_data_out_pll[63]
  PIN la_data_out_pll[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_out_pll[6]
  PIN la_data_out_pll[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END la_data_out_pll[7]
  PIN la_data_out_pll[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2046.840 700.000 2047.440 ;
    END
  END la_data_out_pll[8]
  PIN la_data_out_pll[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END la_data_out_pll[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END rst_n
  PIN rstn_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 822.840 700.000 823.440 ;
    END
  END rstn_i_pll
  PIN rstn_o_pll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END rstn_o_pll
  PIN scan_en_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1710.240 700.000 1710.840 ;
    END
  END scan_en_i_pll
  PIN scan_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1819.040 700.000 1819.640 ;
    END
  END scan_i_pll
  PIN scan_o_pll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2087.640 700.000 2088.240 ;
    END
  END scan_o_pll
  PIN scl_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2074.040 4.000 2074.640 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END scl_pad_o
  PIN scl_padoen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END scl_padoen_o
  PIN sda_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END sda_padoen_o
  PIN slave_ar_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END slave_ar_addr[0]
  PIN slave_ar_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2094.440 4.000 2095.040 ;
    END
  END slave_ar_addr[10]
  PIN slave_ar_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 2196.000 335.250 2200.000 ;
    END
  END slave_ar_addr[11]
  PIN slave_ar_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END slave_ar_addr[12]
  PIN slave_ar_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2087.640 4.000 2088.240 ;
    END
  END slave_ar_addr[13]
  PIN slave_ar_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 2196.000 16.470 2200.000 ;
    END
  END slave_ar_addr[14]
  PIN slave_ar_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END slave_ar_addr[15]
  PIN slave_ar_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END slave_ar_addr[16]
  PIN slave_ar_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 2196.000 534.890 2200.000 ;
    END
  END slave_ar_addr[17]
  PIN slave_ar_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 2196.000 637.930 2200.000 ;
    END
  END slave_ar_addr[18]
  PIN slave_ar_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 758.240 700.000 758.840 ;
    END
  END slave_ar_addr[19]
  PIN slave_ar_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 455.640 700.000 456.240 ;
    END
  END slave_ar_addr[1]
  PIN slave_ar_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END slave_ar_addr[20]
  PIN slave_ar_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 71.440 700.000 72.040 ;
    END
  END slave_ar_addr[21]
  PIN slave_ar_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1989.040 700.000 1989.640 ;
    END
  END slave_ar_addr[22]
  PIN slave_ar_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END slave_ar_addr[23]
  PIN slave_ar_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1985.640 4.000 1986.240 ;
    END
  END slave_ar_addr[24]
  PIN slave_ar_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1672.840 700.000 1673.440 ;
    END
  END slave_ar_addr[25]
  PIN slave_ar_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1992.440 4.000 1993.040 ;
    END
  END slave_ar_addr[26]
  PIN slave_ar_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END slave_ar_addr[27]
  PIN slave_ar_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END slave_ar_addr[28]
  PIN slave_ar_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END slave_ar_addr[29]
  PIN slave_ar_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END slave_ar_addr[2]
  PIN slave_ar_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 391.040 700.000 391.640 ;
    END
  END slave_ar_addr[30]
  PIN slave_ar_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1564.040 700.000 1564.640 ;
    END
  END slave_ar_addr[31]
  PIN slave_ar_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END slave_ar_addr[3]
  PIN slave_ar_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1683.040 700.000 1683.640 ;
    END
  END slave_ar_addr[4]
  PIN slave_ar_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END slave_ar_addr[5]
  PIN slave_ar_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 2196.000 100.190 2200.000 ;
    END
  END slave_ar_addr[6]
  PIN slave_ar_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 23.840 700.000 24.440 ;
    END
  END slave_ar_addr[7]
  PIN slave_ar_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2148.840 700.000 2149.440 ;
    END
  END slave_ar_addr[8]
  PIN slave_ar_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 258.440 700.000 259.040 ;
    END
  END slave_ar_addr[9]
  PIN slave_ar_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END slave_ar_burst[0]
  PIN slave_ar_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 2196.000 592.850 2200.000 ;
    END
  END slave_ar_burst[1]
  PIN slave_ar_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2023.040 4.000 2023.640 ;
    END
  END slave_ar_cache[0]
  PIN slave_ar_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1642.240 700.000 1642.840 ;
    END
  END slave_ar_cache[1]
  PIN slave_ar_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END slave_ar_cache[2]
  PIN slave_ar_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END slave_ar_cache[3]
  PIN slave_ar_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END slave_ar_id[0]
  PIN slave_ar_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 2196.000 412.530 2200.000 ;
    END
  END slave_ar_id[1]
  PIN slave_ar_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END slave_ar_id[2]
  PIN slave_ar_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END slave_ar_id[3]
  PIN slave_ar_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END slave_ar_id[4]
  PIN slave_ar_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2162.440 4.000 2163.040 ;
    END
  END slave_ar_id[5]
  PIN slave_ar_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.840 4.000 1724.440 ;
    END
  END slave_ar_len[0]
  PIN slave_ar_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1557.240 700.000 1557.840 ;
    END
  END slave_ar_len[1]
  PIN slave_ar_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 979.240 700.000 979.840 ;
    END
  END slave_ar_len[2]
  PIN slave_ar_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1026.840 700.000 1027.440 ;
    END
  END slave_ar_len[3]
  PIN slave_ar_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 2196.000 573.530 2200.000 ;
    END
  END slave_ar_len[4]
  PIN slave_ar_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END slave_ar_len[5]
  PIN slave_ar_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 34.040 700.000 34.640 ;
    END
  END slave_ar_len[6]
  PIN slave_ar_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END slave_ar_len[7]
  PIN slave_ar_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2138.640 700.000 2139.240 ;
    END
  END slave_ar_lock
  PIN slave_ar_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 816.040 700.000 816.640 ;
    END
  END slave_ar_prot[0]
  PIN slave_ar_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END slave_ar_prot[1]
  PIN slave_ar_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 2196.000 51.890 2200.000 ;
    END
  END slave_ar_prot[2]
  PIN slave_ar_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1553.840 700.000 1554.440 ;
    END
  END slave_ar_qos[0]
  PIN slave_ar_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 2196.000 460.830 2200.000 ;
    END
  END slave_ar_qos[1]
  PIN slave_ar_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END slave_ar_qos[2]
  PIN slave_ar_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 244.840 700.000 245.440 ;
    END
  END slave_ar_qos[3]
  PIN slave_ar_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 2196.000 596.070 2200.000 ;
    END
  END slave_ar_ready
  PIN slave_ar_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 727.640 700.000 728.240 ;
    END
  END slave_ar_region[0]
  PIN slave_ar_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END slave_ar_region[1]
  PIN slave_ar_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2006.040 4.000 2006.640 ;
    END
  END slave_ar_region[2]
  PIN slave_ar_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END slave_ar_region[3]
  PIN slave_ar_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 2196.000 505.910 2200.000 ;
    END
  END slave_ar_size[0]
  PIN slave_ar_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 98.640 700.000 99.240 ;
    END
  END slave_ar_size[1]
  PIN slave_ar_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1560.640 700.000 1561.240 ;
    END
  END slave_ar_size[2]
  PIN slave_ar_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 710.640 700.000 711.240 ;
    END
  END slave_ar_user[0]
  PIN slave_ar_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END slave_ar_user[1]
  PIN slave_ar_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END slave_ar_user[2]
  PIN slave_ar_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 2196.000 45.450 2200.000 ;
    END
  END slave_ar_user[3]
  PIN slave_ar_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END slave_ar_user[4]
  PIN slave_ar_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2159.040 4.000 2159.640 ;
    END
  END slave_ar_user[5]
  PIN slave_ar_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1696.640 700.000 1697.240 ;
    END
  END slave_ar_valid
  PIN slave_aw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1074.440 700.000 1075.040 ;
    END
  END slave_aw_addr[0]
  PIN slave_aw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END slave_aw_addr[10]
  PIN slave_aw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END slave_aw_addr[11]
  PIN slave_aw_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2152.240 700.000 2152.840 ;
    END
  END slave_aw_addr[12]
  PIN slave_aw_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END slave_aw_addr[13]
  PIN slave_aw_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 941.840 700.000 942.440 ;
    END
  END slave_aw_addr[14]
  PIN slave_aw_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2196.440 4.000 2197.040 ;
    END
  END slave_aw_addr[15]
  PIN slave_aw_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 2196.000 319.150 2200.000 ;
    END
  END slave_aw_addr[16]
  PIN slave_aw_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END slave_aw_addr[17]
  PIN slave_aw_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 350.240 700.000 350.840 ;
    END
  END slave_aw_addr[18]
  PIN slave_aw_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END slave_aw_addr[19]
  PIN slave_aw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 2196.000 161.370 2200.000 ;
    END
  END slave_aw_addr[1]
  PIN slave_aw_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END slave_aw_addr[20]
  PIN slave_aw_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END slave_aw_addr[21]
  PIN slave_aw_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1992.440 700.000 1993.040 ;
    END
  END slave_aw_addr[22]
  PIN slave_aw_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 374.040 700.000 374.640 ;
    END
  END slave_aw_addr[23]
  PIN slave_aw_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1815.640 700.000 1816.240 ;
    END
  END slave_aw_addr[24]
  PIN slave_aw_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END slave_aw_addr[25]
  PIN slave_aw_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END slave_aw_addr[26]
  PIN slave_aw_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1526.640 700.000 1527.240 ;
    END
  END slave_aw_addr[27]
  PIN slave_aw_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1723.840 700.000 1724.440 ;
    END
  END slave_aw_addr[28]
  PIN slave_aw_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END slave_aw_addr[29]
  PIN slave_aw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 2196.000 486.590 2200.000 ;
    END
  END slave_aw_addr[2]
  PIN slave_aw_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 370.640 700.000 371.240 ;
    END
  END slave_aw_addr[30]
  PIN slave_aw_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 2196.000 686.230 2200.000 ;
    END
  END slave_aw_addr[31]
  PIN slave_aw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END slave_aw_addr[3]
  PIN slave_aw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 867.040 700.000 867.640 ;
    END
  END slave_aw_addr[4]
  PIN slave_aw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 557.640 700.000 558.240 ;
    END
  END slave_aw_addr[5]
  PIN slave_aw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END slave_aw_addr[6]
  PIN slave_aw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END slave_aw_addr[7]
  PIN slave_aw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END slave_aw_addr[8]
  PIN slave_aw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1611.640 700.000 1612.240 ;
    END
  END slave_aw_addr[9]
  PIN slave_aw_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END slave_aw_burst[0]
  PIN slave_aw_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2118.240 700.000 2118.840 ;
    END
  END slave_aw_burst[1]
  PIN slave_aw_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END slave_aw_cache[0]
  PIN slave_aw_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END slave_aw_cache[1]
  PIN slave_aw_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END slave_aw_cache[2]
  PIN slave_aw_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END slave_aw_cache[3]
  PIN slave_aw_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END slave_aw_id[0]
  PIN slave_aw_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END slave_aw_id[1]
  PIN slave_aw_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 2196.000 299.830 2200.000 ;
    END
  END slave_aw_id[2]
  PIN slave_aw_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1608.240 700.000 1608.840 ;
    END
  END slave_aw_id[3]
  PIN slave_aw_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 2196.000 364.230 2200.000 ;
    END
  END slave_aw_id[4]
  PIN slave_aw_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 448.840 700.000 449.440 ;
    END
  END slave_aw_id[5]
  PIN slave_aw_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END slave_aw_len[0]
  PIN slave_aw_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END slave_aw_len[1]
  PIN slave_aw_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END slave_aw_len[2]
  PIN slave_aw_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END slave_aw_len[3]
  PIN slave_aw_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END slave_aw_len[4]
  PIN slave_aw_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 986.040 700.000 986.640 ;
    END
  END slave_aw_len[5]
  PIN slave_aw_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1179.840 700.000 1180.440 ;
    END
  END slave_aw_len[6]
  PIN slave_aw_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 2196.000 312.710 2200.000 ;
    END
  END slave_aw_len[7]
  PIN slave_aw_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1921.040 700.000 1921.640 ;
    END
  END slave_aw_lock
  PIN slave_aw_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END slave_aw_prot[0]
  PIN slave_aw_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 302.640 700.000 303.240 ;
    END
  END slave_aw_prot[1]
  PIN slave_aw_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 802.440 700.000 803.040 ;
    END
  END slave_aw_prot[2]
  PIN slave_aw_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 61.240 700.000 61.840 ;
    END
  END slave_aw_qos[0]
  PIN slave_aw_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END slave_aw_qos[1]
  PIN slave_aw_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 428.440 700.000 429.040 ;
    END
  END slave_aw_qos[2]
  PIN slave_aw_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 877.240 700.000 877.840 ;
    END
  END slave_aw_qos[3]
  PIN slave_aw_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 554.240 700.000 554.840 ;
    END
  END slave_aw_ready
  PIN slave_aw_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END slave_aw_region[0]
  PIN slave_aw_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 2196.000 332.030 2200.000 ;
    END
  END slave_aw_region[1]
  PIN slave_aw_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 326.440 700.000 327.040 ;
    END
  END slave_aw_region[2]
  PIN slave_aw_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1591.240 700.000 1591.840 ;
    END
  END slave_aw_region[3]
  PIN slave_aw_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1268.240 700.000 1268.840 ;
    END
  END slave_aw_size[0]
  PIN slave_aw_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1836.040 700.000 1836.640 ;
    END
  END slave_aw_size[1]
  PIN slave_aw_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1727.240 700.000 1727.840 ;
    END
  END slave_aw_size[2]
  PIN slave_aw_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END slave_aw_user[0]
  PIN slave_aw_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END slave_aw_user[1]
  PIN slave_aw_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 734.440 700.000 735.040 ;
    END
  END slave_aw_user[2]
  PIN slave_aw_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END slave_aw_user[3]
  PIN slave_aw_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 969.040 700.000 969.640 ;
    END
  END slave_aw_user[4]
  PIN slave_aw_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1904.040 4.000 1904.640 ;
    END
  END slave_aw_user[5]
  PIN slave_aw_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END slave_aw_valid
  PIN slave_b_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1332.840 700.000 1333.440 ;
    END
  END slave_b_id[0]
  PIN slave_b_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END slave_b_id[1]
  PIN slave_b_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 367.240 700.000 367.840 ;
    END
  END slave_b_id[2]
  PIN slave_b_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 584.840 700.000 585.440 ;
    END
  END slave_b_id[3]
  PIN slave_b_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END slave_b_id[4]
  PIN slave_b_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END slave_b_id[5]
  PIN slave_b_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END slave_b_ready
  PIN slave_b_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1003.040 700.000 1003.640 ;
    END
  END slave_b_resp[0]
  PIN slave_b_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END slave_b_resp[1]
  PIN slave_b_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END slave_b_user[0]
  PIN slave_b_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1917.640 4.000 1918.240 ;
    END
  END slave_b_user[1]
  PIN slave_b_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 846.640 700.000 847.240 ;
    END
  END slave_b_user[2]
  PIN slave_b_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1907.440 700.000 1908.040 ;
    END
  END slave_b_user[3]
  PIN slave_b_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1533.440 4.000 1534.040 ;
    END
  END slave_b_user[4]
  PIN slave_b_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END slave_b_user[5]
  PIN slave_b_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1309.040 700.000 1309.640 ;
    END
  END slave_b_valid
  PIN slave_r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 176.840 700.000 177.440 ;
    END
  END slave_r_data[0]
  PIN slave_r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 333.240 700.000 333.840 ;
    END
  END slave_r_data[10]
  PIN slave_r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1907.440 4.000 1908.040 ;
    END
  END slave_r_data[11]
  PIN slave_r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1513.040 700.000 1513.640 ;
    END
  END slave_r_data[12]
  PIN slave_r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END slave_r_data[13]
  PIN slave_r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END slave_r_data[14]
  PIN slave_r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 2196.000 515.570 2200.000 ;
    END
  END slave_r_data[15]
  PIN slave_r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 724.240 700.000 724.840 ;
    END
  END slave_r_data[16]
  PIN slave_r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1870.040 4.000 1870.640 ;
    END
  END slave_r_data[17]
  PIN slave_r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 2196.000 547.770 2200.000 ;
    END
  END slave_r_data[18]
  PIN slave_r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END slave_r_data[19]
  PIN slave_r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1499.440 4.000 1500.040 ;
    END
  END slave_r_data[1]
  PIN slave_r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 57.840 700.000 58.440 ;
    END
  END slave_r_data[20]
  PIN slave_r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 2196.000 209.670 2200.000 ;
    END
  END slave_r_data[21]
  PIN slave_r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 703.840 700.000 704.440 ;
    END
  END slave_r_data[22]
  PIN slave_r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 2196.000 654.030 2200.000 ;
    END
  END slave_r_data[23]
  PIN slave_r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END slave_r_data[24]
  PIN slave_r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END slave_r_data[25]
  PIN slave_r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 401.240 700.000 401.840 ;
    END
  END slave_r_data[26]
  PIN slave_r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 272.040 700.000 272.640 ;
    END
  END slave_r_data[27]
  PIN slave_r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2091.040 4.000 2091.640 ;
    END
  END slave_r_data[28]
  PIN slave_r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1965.240 700.000 1965.840 ;
    END
  END slave_r_data[29]
  PIN slave_r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1319.240 700.000 1319.840 ;
    END
  END slave_r_data[2]
  PIN slave_r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 2196.000 612.170 2200.000 ;
    END
  END slave_r_data[30]
  PIN slave_r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 506.640 700.000 507.240 ;
    END
  END slave_r_data[31]
  PIN slave_r_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END slave_r_data[32]
  PIN slave_r_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END slave_r_data[33]
  PIN slave_r_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END slave_r_data[34]
  PIN slave_r_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1822.440 700.000 1823.040 ;
    END
  END slave_r_data[35]
  PIN slave_r_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2097.840 700.000 2098.440 ;
    END
  END slave_r_data[36]
  PIN slave_r_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 843.240 700.000 843.840 ;
    END
  END slave_r_data[37]
  PIN slave_r_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1662.640 700.000 1663.240 ;
    END
  END slave_r_data[38]
  PIN slave_r_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 2196.000 435.070 2200.000 ;
    END
  END slave_r_data[39]
  PIN slave_r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END slave_r_data[3]
  PIN slave_r_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END slave_r_data[40]
  PIN slave_r_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 278.840 700.000 279.440 ;
    END
  END slave_r_data[41]
  PIN slave_r_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END slave_r_data[42]
  PIN slave_r_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1489.240 700.000 1489.840 ;
    END
  END slave_r_data[43]
  PIN slave_r_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END slave_r_data[44]
  PIN slave_r_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END slave_r_data[45]
  PIN slave_r_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1434.840 700.000 1435.440 ;
    END
  END slave_r_data[46]
  PIN slave_r_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 2196.000 55.110 2200.000 ;
    END
  END slave_r_data[47]
  PIN slave_r_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1924.440 700.000 1925.040 ;
    END
  END slave_r_data[48]
  PIN slave_r_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END slave_r_data[49]
  PIN slave_r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1778.240 700.000 1778.840 ;
    END
  END slave_r_data[4]
  PIN slave_r_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 564.440 700.000 565.040 ;
    END
  END slave_r_data[50]
  PIN slave_r_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1934.640 4.000 1935.240 ;
    END
  END slave_r_data[51]
  PIN slave_r_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 462.440 700.000 463.040 ;
    END
  END slave_r_data[52]
  PIN slave_r_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2135.240 700.000 2135.840 ;
    END
  END slave_r_data[53]
  PIN slave_r_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2176.040 4.000 2176.640 ;
    END
  END slave_r_data[54]
  PIN slave_r_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1975.440 4.000 1976.040 ;
    END
  END slave_r_data[55]
  PIN slave_r_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END slave_r_data[56]
  PIN slave_r_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 2196.000 13.250 2200.000 ;
    END
  END slave_r_data[57]
  PIN slave_r_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END slave_r_data[58]
  PIN slave_r_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END slave_r_data[59]
  PIN slave_r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1227.440 700.000 1228.040 ;
    END
  END slave_r_data[5]
  PIN slave_r_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1693.240 700.000 1693.840 ;
    END
  END slave_r_data[60]
  PIN slave_r_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2155.640 700.000 2156.240 ;
    END
  END slave_r_data[61]
  PIN slave_r_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END slave_r_data[62]
  PIN slave_r_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 676.640 700.000 677.240 ;
    END
  END slave_r_data[63]
  PIN slave_r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 2196.000 361.010 2200.000 ;
    END
  END slave_r_data[6]
  PIN slave_r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 2196.000 586.410 2200.000 ;
    END
  END slave_r_data[7]
  PIN slave_r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2097.840 4.000 2098.440 ;
    END
  END slave_r_data[8]
  PIN slave_r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 2196.000 216.110 2200.000 ;
    END
  END slave_r_data[9]
  PIN slave_r_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 945.240 700.000 945.840 ;
    END
  END slave_r_id[0]
  PIN slave_r_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 2196.000 196.790 2200.000 ;
    END
  END slave_r_id[1]
  PIN slave_r_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 873.840 700.000 874.440 ;
    END
  END slave_r_id[2]
  PIN slave_r_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1183.240 700.000 1183.840 ;
    END
  END slave_r_id[3]
  PIN slave_r_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END slave_r_id[4]
  PIN slave_r_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END slave_r_id[5]
  PIN slave_r_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 982.640 700.000 983.240 ;
    END
  END slave_r_last
  PIN slave_r_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1601.440 700.000 1602.040 ;
    END
  END slave_r_ready
  PIN slave_r_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END slave_r_resp[0]
  PIN slave_r_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END slave_r_resp[1]
  PIN slave_r_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END slave_r_user[0]
  PIN slave_r_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END slave_r_user[1]
  PIN slave_r_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END slave_r_user[2]
  PIN slave_r_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 2196.000 254.750 2200.000 ;
    END
  END slave_r_user[3]
  PIN slave_r_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1135.640 700.000 1136.240 ;
    END
  END slave_r_user[4]
  PIN slave_r_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END slave_r_user[5]
  PIN slave_r_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END slave_r_valid
  PIN slave_w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 2196.000 467.270 2200.000 ;
    END
  END slave_w_data[0]
  PIN slave_w_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1819.040 4.000 1819.640 ;
    END
  END slave_w_data[10]
  PIN slave_w_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END slave_w_data[11]
  PIN slave_w_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2040.040 4.000 2040.640 ;
    END
  END slave_w_data[12]
  PIN slave_w_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2128.440 4.000 2129.040 ;
    END
  END slave_w_data[13]
  PIN slave_w_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2148.840 4.000 2149.440 ;
    END
  END slave_w_data[14]
  PIN slave_w_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END slave_w_data[15]
  PIN slave_w_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END slave_w_data[16]
  PIN slave_w_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END slave_w_data[17]
  PIN slave_w_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END slave_w_data[18]
  PIN slave_w_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 812.640 700.000 813.240 ;
    END
  END slave_w_data[19]
  PIN slave_w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END slave_w_data[1]
  PIN slave_w_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END slave_w_data[20]
  PIN slave_w_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1778.240 4.000 1778.840 ;
    END
  END slave_w_data[21]
  PIN slave_w_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1506.240 700.000 1506.840 ;
    END
  END slave_w_data[22]
  PIN slave_w_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END slave_w_data[23]
  PIN slave_w_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END slave_w_data[24]
  PIN slave_w_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END slave_w_data[25]
  PIN slave_w_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 136.040 700.000 136.640 ;
    END
  END slave_w_data[26]
  PIN slave_w_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END slave_w_data[27]
  PIN slave_w_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 839.840 700.000 840.440 ;
    END
  END slave_w_data[28]
  PIN slave_w_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 10.240 700.000 10.840 ;
    END
  END slave_w_data[29]
  PIN slave_w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 731.040 700.000 731.640 ;
    END
  END slave_w_data[2]
  PIN slave_w_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END slave_w_data[30]
  PIN slave_w_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 2196.000 406.090 2200.000 ;
    END
  END slave_w_data[31]
  PIN slave_w_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 761.640 700.000 762.240 ;
    END
  END slave_w_data[32]
  PIN slave_w_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END slave_w_data[33]
  PIN slave_w_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1173.040 700.000 1173.640 ;
    END
  END slave_w_data[34]
  PIN slave_w_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END slave_w_data[35]
  PIN slave_w_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END slave_w_data[36]
  PIN slave_w_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2159.040 700.000 2159.640 ;
    END
  END slave_w_data[37]
  PIN slave_w_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 717.440 700.000 718.040 ;
    END
  END slave_w_data[38]
  PIN slave_w_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1853.040 4.000 1853.640 ;
    END
  END slave_w_data[39]
  PIN slave_w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1353.240 700.000 1353.840 ;
    END
  END slave_w_data[3]
  PIN slave_w_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1322.640 4.000 1323.240 ;
    END
  END slave_w_data[40]
  PIN slave_w_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1013.240 700.000 1013.840 ;
    END
  END slave_w_data[41]
  PIN slave_w_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END slave_w_data[42]
  PIN slave_w_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END slave_w_data[43]
  PIN slave_w_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2074.040 700.000 2074.640 ;
    END
  END slave_w_data[44]
  PIN slave_w_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 316.240 700.000 316.840 ;
    END
  END slave_w_data[45]
  PIN slave_w_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 2196.000 557.430 2200.000 ;
    END
  END slave_w_data[46]
  PIN slave_w_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END slave_w_data[47]
  PIN slave_w_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1030.240 700.000 1030.840 ;
    END
  END slave_w_data[48]
  PIN slave_w_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END slave_w_data[49]
  PIN slave_w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1924.440 4.000 1925.040 ;
    END
  END slave_w_data[4]
  PIN slave_w_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 2196.000 402.870 2200.000 ;
    END
  END slave_w_data[50]
  PIN slave_w_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END slave_w_data[51]
  PIN slave_w_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END slave_w_data[52]
  PIN slave_w_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END slave_w_data[53]
  PIN slave_w_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END slave_w_data[54]
  PIN slave_w_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1713.640 700.000 1714.240 ;
    END
  END slave_w_data[55]
  PIN slave_w_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1642.240 4.000 1642.840 ;
    END
  END slave_w_data[56]
  PIN slave_w_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END slave_w_data[57]
  PIN slave_w_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END slave_w_data[58]
  PIN slave_w_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END slave_w_data[59]
  PIN slave_w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 268.640 700.000 269.240 ;
    END
  END slave_w_data[5]
  PIN slave_w_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 2196.000 538.110 2200.000 ;
    END
  END slave_w_data[60]
  PIN slave_w_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 2196.000 644.370 2200.000 ;
    END
  END slave_w_data[61]
  PIN slave_w_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 397.840 700.000 398.440 ;
    END
  END slave_w_data[62]
  PIN slave_w_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2114.840 700.000 2115.440 ;
    END
  END slave_w_data[63]
  PIN slave_w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1598.040 700.000 1598.640 ;
    END
  END slave_w_data[6]
  PIN slave_w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 972.440 700.000 973.040 ;
    END
  END slave_w_data[7]
  PIN slave_w_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1720.440 4.000 1721.040 ;
    END
  END slave_w_data[8]
  PIN slave_w_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 2196.000 22.910 2200.000 ;
    END
  END slave_w_data[9]
  PIN slave_w_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 261.840 700.000 262.440 ;
    END
  END slave_w_last
  PIN slave_w_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 686.840 700.000 687.440 ;
    END
  END slave_w_ready
  PIN slave_w_strb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1417.840 700.000 1418.440 ;
    END
  END slave_w_strb[0]
  PIN slave_w_strb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END slave_w_strb[1]
  PIN slave_w_strb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END slave_w_strb[2]
  PIN slave_w_strb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END slave_w_strb[3]
  PIN slave_w_strb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END slave_w_strb[4]
  PIN slave_w_strb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2002.640 700.000 2003.240 ;
    END
  END slave_w_strb[5]
  PIN slave_w_strb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 2196.000 280.510 2200.000 ;
    END
  END slave_w_strb[6]
  PIN slave_w_strb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END slave_w_strb[7]
  PIN slave_w_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2084.240 4.000 2084.840 ;
    END
  END slave_w_user[0]
  PIN slave_w_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1706.840 700.000 1707.440 ;
    END
  END slave_w_user[1]
  PIN slave_w_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 598.440 700.000 599.040 ;
    END
  END slave_w_user[2]
  PIN slave_w_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2067.240 4.000 2067.840 ;
    END
  END slave_w_user[3]
  PIN slave_w_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 544.040 700.000 544.640 ;
    END
  END slave_w_user[4]
  PIN slave_w_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END slave_w_user[5]
  PIN slave_w_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END slave_w_valid
  PIN spi_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 958.840 700.000 959.440 ;
    END
  END spi_clk_i
  PIN spi_cs_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1411.040 700.000 1411.640 ;
    END
  END spi_cs_i
  PIN spi_master_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END spi_master_clk
  PIN spi_master_csn0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 2196.000 499.470 2200.000 ;
    END
  END spi_master_csn0
  PIN spi_master_csn1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END spi_master_csn1
  PIN spi_master_csn2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END spi_master_csn2
  PIN spi_master_csn3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END spi_master_csn3
  PIN spi_master_mode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END spi_master_mode[0]
  PIN spi_master_mode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END spi_master_mode[1]
  PIN spi_master_sdi0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1791.840 700.000 1792.440 ;
    END
  END spi_master_sdi0
  PIN spi_master_sdi1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 217.640 700.000 218.240 ;
    END
  END spi_master_sdi1
  PIN spi_master_sdi2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2050.240 4.000 2050.840 ;
    END
  END spi_master_sdi2
  PIN spi_master_sdi3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 2196.000 241.870 2200.000 ;
    END
  END spi_master_sdi3
  PIN spi_master_sdo0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END spi_master_sdo0
  PIN spi_master_sdo1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END spi_master_sdo1
  PIN spi_master_sdo2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1893.840 700.000 1894.440 ;
    END
  END spi_master_sdo2
  PIN spi_master_sdo3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 2196.000 315.930 2200.000 ;
    END
  END spi_master_sdo3
  PIN spi_mode_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END spi_mode_o[0]
  PIN spi_mode_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2169.240 700.000 2169.840 ;
    END
  END spi_mode_o[1]
  PIN spi_sdi0_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1421.240 700.000 1421.840 ;
    END
  END spi_sdi0_i
  PIN spi_sdi1_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 387.640 700.000 388.240 ;
    END
  END spi_sdi1_i
  PIN spi_sdi2_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END spi_sdi2_i
  PIN spi_sdi3_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1424.640 4.000 1425.240 ;
    END
  END spi_sdi3_i
  PIN spi_sdo0_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END spi_sdo0_o
  PIN spi_sdo1_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1849.640 700.000 1850.240 ;
    END
  END spi_sdo1_o
  PIN spi_sdo2_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 581.440 700.000 582.040 ;
    END
  END spi_sdo2_o
  PIN spi_sdo3_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1343.040 700.000 1343.640 ;
    END
  END spi_sdo3_o
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END testmode_i
  PIN testmode_i_pll
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 921.440 700.000 922.040 ;
    END
  END testmode_i_pll
  PIN uart_cts
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END uart_cts
  PIN uart_dsr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 51.040 700.000 51.640 ;
    END
  END uart_dsr
  PIN uart_dtr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1540.240 700.000 1540.840 ;
    END
  END uart_dtr
  PIN uart_rts
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 2196.000 174.250 2200.000 ;
    END
  END uart_rts
  PIN uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 2196.000 641.150 2200.000 ;
    END
  END uart_rx
  PIN uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 924.840 700.000 925.440 ;
    END
  END uart_tx
  PIN user_irq_pll[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END user_irq_pll[0]
  PIN user_irq_pll[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1734.040 700.000 1734.640 ;
    END
  END user_irq_pll[1]
  PIN user_irq_pll[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END user_irq_pll[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 2196.000 634.710 2200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2187.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 2196.000 158.150 2200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2187.120 ;
    END
  END vssd1
  PIN wbs_ack_o_pll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1006.440 700.000 1007.040 ;
    END
  END wbs_ack_o_pll
  PIN wbs_dat_o_pll[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 2196.000 119.510 2200.000 ;
    END
  END wbs_dat_o_pll[0]
  PIN wbs_dat_o_pll[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 309.440 700.000 310.040 ;
    END
  END wbs_dat_o_pll[10]
  PIN wbs_dat_o_pll[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wbs_dat_o_pll[11]
  PIN wbs_dat_o_pll[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 306.040 700.000 306.640 ;
    END
  END wbs_dat_o_pll[12]
  PIN wbs_dat_o_pll[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wbs_dat_o_pll[13]
  PIN wbs_dat_o_pll[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 482.840 700.000 483.440 ;
    END
  END wbs_dat_o_pll[14]
  PIN wbs_dat_o_pll[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END wbs_dat_o_pll[15]
  PIN wbs_dat_o_pll[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END wbs_dat_o_pll[16]
  PIN wbs_dat_o_pll[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1703.440 4.000 1704.040 ;
    END
  END wbs_dat_o_pll[17]
  PIN wbs_dat_o_pll[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wbs_dat_o_pll[18]
  PIN wbs_dat_o_pll[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_dat_o_pll[19]
  PIN wbs_dat_o_pll[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_dat_o_pll[1]
  PIN wbs_dat_o_pll[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2104.640 4.000 2105.240 ;
    END
  END wbs_dat_o_pll[20]
  PIN wbs_dat_o_pll[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END wbs_dat_o_pll[21]
  PIN wbs_dat_o_pll[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 88.440 700.000 89.040 ;
    END
  END wbs_dat_o_pll[22]
  PIN wbs_dat_o_pll[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_dat_o_pll[23]
  PIN wbs_dat_o_pll[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1196.840 700.000 1197.440 ;
    END
  END wbs_dat_o_pll[24]
  PIN wbs_dat_o_pll[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END wbs_dat_o_pll[25]
  PIN wbs_dat_o_pll[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1934.640 700.000 1935.240 ;
    END
  END wbs_dat_o_pll[26]
  PIN wbs_dat_o_pll[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END wbs_dat_o_pll[27]
  PIN wbs_dat_o_pll[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END wbs_dat_o_pll[28]
  PIN wbs_dat_o_pll[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_dat_o_pll[29]
  PIN wbs_dat_o_pll[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1859.840 700.000 1860.440 ;
    END
  END wbs_dat_o_pll[2]
  PIN wbs_dat_o_pll[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 166.640 700.000 167.240 ;
    END
  END wbs_dat_o_pll[30]
  PIN wbs_dat_o_pll[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 2196.000 177.470 2200.000 ;
    END
  END wbs_dat_o_pll[31]
  PIN wbs_dat_o_pll[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 2196.000 164.590 2200.000 ;
    END
  END wbs_dat_o_pll[3]
  PIN wbs_dat_o_pll[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END wbs_dat_o_pll[4]
  PIN wbs_dat_o_pll[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1587.840 4.000 1588.440 ;
    END
  END wbs_dat_o_pll[5]
  PIN wbs_dat_o_pll[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 329.840 700.000 330.440 ;
    END
  END wbs_dat_o_pll[6]
  PIN wbs_dat_o_pll[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wbs_dat_o_pll[7]
  PIN wbs_dat_o_pll[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END wbs_dat_o_pll[8]
  PIN wbs_dat_o_pll[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 1458.640 700.000 1459.240 ;
    END
  END wbs_dat_o_pll[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 2186.965 ;
      LAYER met1 ;
        RECT 0.070 6.840 699.960 2187.120 ;
      LAYER met2 ;
        RECT 0.650 2195.720 3.030 2196.925 ;
        RECT 3.870 2195.720 9.470 2196.925 ;
        RECT 10.310 2195.720 12.690 2196.925 ;
        RECT 13.530 2195.720 15.910 2196.925 ;
        RECT 16.750 2195.720 19.130 2196.925 ;
        RECT 19.970 2195.720 22.350 2196.925 ;
        RECT 23.190 2195.720 28.790 2196.925 ;
        RECT 29.630 2195.720 32.010 2196.925 ;
        RECT 32.850 2195.720 35.230 2196.925 ;
        RECT 36.070 2195.720 38.450 2196.925 ;
        RECT 39.290 2195.720 41.670 2196.925 ;
        RECT 42.510 2195.720 44.890 2196.925 ;
        RECT 45.730 2195.720 51.330 2196.925 ;
        RECT 52.170 2195.720 54.550 2196.925 ;
        RECT 55.390 2195.720 57.770 2196.925 ;
        RECT 58.610 2195.720 60.990 2196.925 ;
        RECT 61.830 2195.720 64.210 2196.925 ;
        RECT 65.050 2195.720 70.650 2196.925 ;
        RECT 71.490 2195.720 73.870 2196.925 ;
        RECT 74.710 2195.720 77.090 2196.925 ;
        RECT 77.930 2195.720 80.310 2196.925 ;
        RECT 81.150 2195.720 83.530 2196.925 ;
        RECT 84.370 2195.720 89.970 2196.925 ;
        RECT 90.810 2195.720 93.190 2196.925 ;
        RECT 94.030 2195.720 96.410 2196.925 ;
        RECT 97.250 2195.720 99.630 2196.925 ;
        RECT 100.470 2195.720 102.850 2196.925 ;
        RECT 103.690 2195.720 109.290 2196.925 ;
        RECT 110.130 2195.720 112.510 2196.925 ;
        RECT 113.350 2195.720 115.730 2196.925 ;
        RECT 116.570 2195.720 118.950 2196.925 ;
        RECT 119.790 2195.720 122.170 2196.925 ;
        RECT 123.010 2195.720 125.390 2196.925 ;
        RECT 126.230 2195.720 131.830 2196.925 ;
        RECT 132.670 2195.720 135.050 2196.925 ;
        RECT 135.890 2195.720 138.270 2196.925 ;
        RECT 139.110 2195.720 141.490 2196.925 ;
        RECT 142.330 2195.720 144.710 2196.925 ;
        RECT 145.550 2195.720 151.150 2196.925 ;
        RECT 151.990 2195.720 154.370 2196.925 ;
        RECT 155.210 2195.720 157.590 2196.925 ;
        RECT 158.430 2195.720 160.810 2196.925 ;
        RECT 161.650 2195.720 164.030 2196.925 ;
        RECT 164.870 2195.720 170.470 2196.925 ;
        RECT 171.310 2195.720 173.690 2196.925 ;
        RECT 174.530 2195.720 176.910 2196.925 ;
        RECT 177.750 2195.720 180.130 2196.925 ;
        RECT 180.970 2195.720 183.350 2196.925 ;
        RECT 184.190 2195.720 189.790 2196.925 ;
        RECT 190.630 2195.720 193.010 2196.925 ;
        RECT 193.850 2195.720 196.230 2196.925 ;
        RECT 197.070 2195.720 199.450 2196.925 ;
        RECT 200.290 2195.720 202.670 2196.925 ;
        RECT 203.510 2195.720 209.110 2196.925 ;
        RECT 209.950 2195.720 212.330 2196.925 ;
        RECT 213.170 2195.720 215.550 2196.925 ;
        RECT 216.390 2195.720 218.770 2196.925 ;
        RECT 219.610 2195.720 221.990 2196.925 ;
        RECT 222.830 2195.720 225.210 2196.925 ;
        RECT 226.050 2195.720 231.650 2196.925 ;
        RECT 232.490 2195.720 234.870 2196.925 ;
        RECT 235.710 2195.720 238.090 2196.925 ;
        RECT 238.930 2195.720 241.310 2196.925 ;
        RECT 242.150 2195.720 244.530 2196.925 ;
        RECT 245.370 2195.720 250.970 2196.925 ;
        RECT 251.810 2195.720 254.190 2196.925 ;
        RECT 255.030 2195.720 257.410 2196.925 ;
        RECT 258.250 2195.720 260.630 2196.925 ;
        RECT 261.470 2195.720 263.850 2196.925 ;
        RECT 264.690 2195.720 270.290 2196.925 ;
        RECT 271.130 2195.720 273.510 2196.925 ;
        RECT 274.350 2195.720 276.730 2196.925 ;
        RECT 277.570 2195.720 279.950 2196.925 ;
        RECT 280.790 2195.720 283.170 2196.925 ;
        RECT 284.010 2195.720 289.610 2196.925 ;
        RECT 290.450 2195.720 292.830 2196.925 ;
        RECT 293.670 2195.720 296.050 2196.925 ;
        RECT 296.890 2195.720 299.270 2196.925 ;
        RECT 300.110 2195.720 302.490 2196.925 ;
        RECT 303.330 2195.720 305.710 2196.925 ;
        RECT 306.550 2195.720 312.150 2196.925 ;
        RECT 312.990 2195.720 315.370 2196.925 ;
        RECT 316.210 2195.720 318.590 2196.925 ;
        RECT 319.430 2195.720 321.810 2196.925 ;
        RECT 322.650 2195.720 325.030 2196.925 ;
        RECT 325.870 2195.720 331.470 2196.925 ;
        RECT 332.310 2195.720 334.690 2196.925 ;
        RECT 335.530 2195.720 337.910 2196.925 ;
        RECT 338.750 2195.720 341.130 2196.925 ;
        RECT 341.970 2195.720 344.350 2196.925 ;
        RECT 345.190 2195.720 350.790 2196.925 ;
        RECT 351.630 2195.720 354.010 2196.925 ;
        RECT 354.850 2195.720 357.230 2196.925 ;
        RECT 358.070 2195.720 360.450 2196.925 ;
        RECT 361.290 2195.720 363.670 2196.925 ;
        RECT 364.510 2195.720 370.110 2196.925 ;
        RECT 370.950 2195.720 373.330 2196.925 ;
        RECT 374.170 2195.720 376.550 2196.925 ;
        RECT 377.390 2195.720 379.770 2196.925 ;
        RECT 380.610 2195.720 382.990 2196.925 ;
        RECT 383.830 2195.720 386.210 2196.925 ;
        RECT 387.050 2195.720 392.650 2196.925 ;
        RECT 393.490 2195.720 395.870 2196.925 ;
        RECT 396.710 2195.720 399.090 2196.925 ;
        RECT 399.930 2195.720 402.310 2196.925 ;
        RECT 403.150 2195.720 405.530 2196.925 ;
        RECT 406.370 2195.720 411.970 2196.925 ;
        RECT 412.810 2195.720 415.190 2196.925 ;
        RECT 416.030 2195.720 418.410 2196.925 ;
        RECT 419.250 2195.720 421.630 2196.925 ;
        RECT 422.470 2195.720 424.850 2196.925 ;
        RECT 425.690 2195.720 431.290 2196.925 ;
        RECT 432.130 2195.720 434.510 2196.925 ;
        RECT 435.350 2195.720 437.730 2196.925 ;
        RECT 438.570 2195.720 440.950 2196.925 ;
        RECT 441.790 2195.720 444.170 2196.925 ;
        RECT 445.010 2195.720 450.610 2196.925 ;
        RECT 451.450 2195.720 453.830 2196.925 ;
        RECT 454.670 2195.720 457.050 2196.925 ;
        RECT 457.890 2195.720 460.270 2196.925 ;
        RECT 461.110 2195.720 463.490 2196.925 ;
        RECT 464.330 2195.720 466.710 2196.925 ;
        RECT 467.550 2195.720 473.150 2196.925 ;
        RECT 473.990 2195.720 476.370 2196.925 ;
        RECT 477.210 2195.720 479.590 2196.925 ;
        RECT 480.430 2195.720 482.810 2196.925 ;
        RECT 483.650 2195.720 486.030 2196.925 ;
        RECT 486.870 2195.720 492.470 2196.925 ;
        RECT 493.310 2195.720 495.690 2196.925 ;
        RECT 496.530 2195.720 498.910 2196.925 ;
        RECT 499.750 2195.720 502.130 2196.925 ;
        RECT 502.970 2195.720 505.350 2196.925 ;
        RECT 506.190 2195.720 511.790 2196.925 ;
        RECT 512.630 2195.720 515.010 2196.925 ;
        RECT 515.850 2195.720 518.230 2196.925 ;
        RECT 519.070 2195.720 521.450 2196.925 ;
        RECT 522.290 2195.720 524.670 2196.925 ;
        RECT 525.510 2195.720 531.110 2196.925 ;
        RECT 531.950 2195.720 534.330 2196.925 ;
        RECT 535.170 2195.720 537.550 2196.925 ;
        RECT 538.390 2195.720 540.770 2196.925 ;
        RECT 541.610 2195.720 543.990 2196.925 ;
        RECT 544.830 2195.720 547.210 2196.925 ;
        RECT 548.050 2195.720 553.650 2196.925 ;
        RECT 554.490 2195.720 556.870 2196.925 ;
        RECT 557.710 2195.720 560.090 2196.925 ;
        RECT 560.930 2195.720 563.310 2196.925 ;
        RECT 564.150 2195.720 566.530 2196.925 ;
        RECT 567.370 2195.720 572.970 2196.925 ;
        RECT 573.810 2195.720 576.190 2196.925 ;
        RECT 577.030 2195.720 579.410 2196.925 ;
        RECT 580.250 2195.720 582.630 2196.925 ;
        RECT 583.470 2195.720 585.850 2196.925 ;
        RECT 586.690 2195.720 592.290 2196.925 ;
        RECT 593.130 2195.720 595.510 2196.925 ;
        RECT 596.350 2195.720 598.730 2196.925 ;
        RECT 599.570 2195.720 601.950 2196.925 ;
        RECT 602.790 2195.720 605.170 2196.925 ;
        RECT 606.010 2195.720 611.610 2196.925 ;
        RECT 612.450 2195.720 614.830 2196.925 ;
        RECT 615.670 2195.720 618.050 2196.925 ;
        RECT 618.890 2195.720 621.270 2196.925 ;
        RECT 622.110 2195.720 624.490 2196.925 ;
        RECT 625.330 2195.720 627.710 2196.925 ;
        RECT 628.550 2195.720 634.150 2196.925 ;
        RECT 634.990 2195.720 637.370 2196.925 ;
        RECT 638.210 2195.720 640.590 2196.925 ;
        RECT 641.430 2195.720 643.810 2196.925 ;
        RECT 644.650 2195.720 647.030 2196.925 ;
        RECT 647.870 2195.720 653.470 2196.925 ;
        RECT 654.310 2195.720 656.690 2196.925 ;
        RECT 657.530 2195.720 659.910 2196.925 ;
        RECT 660.750 2195.720 663.130 2196.925 ;
        RECT 663.970 2195.720 666.350 2196.925 ;
        RECT 667.190 2195.720 672.790 2196.925 ;
        RECT 673.630 2195.720 676.010 2196.925 ;
        RECT 676.850 2195.720 679.230 2196.925 ;
        RECT 680.070 2195.720 682.450 2196.925 ;
        RECT 683.290 2195.720 685.670 2196.925 ;
        RECT 686.510 2195.720 692.110 2196.925 ;
        RECT 692.950 2195.720 695.330 2196.925 ;
        RECT 696.170 2195.720 698.550 2196.925 ;
        RECT 699.390 2195.720 699.960 2196.925 ;
        RECT 0.100 4.280 699.960 2195.720 ;
        RECT 0.650 3.555 3.030 4.280 ;
        RECT 3.870 3.555 6.250 4.280 ;
        RECT 7.090 3.555 9.470 4.280 ;
        RECT 10.310 3.555 12.690 4.280 ;
        RECT 13.530 3.555 15.910 4.280 ;
        RECT 16.750 3.555 22.350 4.280 ;
        RECT 23.190 3.555 25.570 4.280 ;
        RECT 26.410 3.555 28.790 4.280 ;
        RECT 29.630 3.555 32.010 4.280 ;
        RECT 32.850 3.555 35.230 4.280 ;
        RECT 36.070 3.555 41.670 4.280 ;
        RECT 42.510 3.555 44.890 4.280 ;
        RECT 45.730 3.555 48.110 4.280 ;
        RECT 48.950 3.555 51.330 4.280 ;
        RECT 52.170 3.555 54.550 4.280 ;
        RECT 55.390 3.555 60.990 4.280 ;
        RECT 61.830 3.555 64.210 4.280 ;
        RECT 65.050 3.555 67.430 4.280 ;
        RECT 68.270 3.555 70.650 4.280 ;
        RECT 71.490 3.555 73.870 4.280 ;
        RECT 74.710 3.555 80.310 4.280 ;
        RECT 81.150 3.555 83.530 4.280 ;
        RECT 84.370 3.555 86.750 4.280 ;
        RECT 87.590 3.555 89.970 4.280 ;
        RECT 90.810 3.555 93.190 4.280 ;
        RECT 94.030 3.555 96.410 4.280 ;
        RECT 97.250 3.555 102.850 4.280 ;
        RECT 103.690 3.555 106.070 4.280 ;
        RECT 106.910 3.555 109.290 4.280 ;
        RECT 110.130 3.555 112.510 4.280 ;
        RECT 113.350 3.555 115.730 4.280 ;
        RECT 116.570 3.555 122.170 4.280 ;
        RECT 123.010 3.555 125.390 4.280 ;
        RECT 126.230 3.555 128.610 4.280 ;
        RECT 129.450 3.555 131.830 4.280 ;
        RECT 132.670 3.555 135.050 4.280 ;
        RECT 135.890 3.555 141.490 4.280 ;
        RECT 142.330 3.555 144.710 4.280 ;
        RECT 145.550 3.555 147.930 4.280 ;
        RECT 148.770 3.555 151.150 4.280 ;
        RECT 151.990 3.555 154.370 4.280 ;
        RECT 155.210 3.555 160.810 4.280 ;
        RECT 161.650 3.555 164.030 4.280 ;
        RECT 164.870 3.555 167.250 4.280 ;
        RECT 168.090 3.555 170.470 4.280 ;
        RECT 171.310 3.555 173.690 4.280 ;
        RECT 174.530 3.555 176.910 4.280 ;
        RECT 177.750 3.555 183.350 4.280 ;
        RECT 184.190 3.555 186.570 4.280 ;
        RECT 187.410 3.555 189.790 4.280 ;
        RECT 190.630 3.555 193.010 4.280 ;
        RECT 193.850 3.555 196.230 4.280 ;
        RECT 197.070 3.555 202.670 4.280 ;
        RECT 203.510 3.555 205.890 4.280 ;
        RECT 206.730 3.555 209.110 4.280 ;
        RECT 209.950 3.555 212.330 4.280 ;
        RECT 213.170 3.555 215.550 4.280 ;
        RECT 216.390 3.555 221.990 4.280 ;
        RECT 222.830 3.555 225.210 4.280 ;
        RECT 226.050 3.555 228.430 4.280 ;
        RECT 229.270 3.555 231.650 4.280 ;
        RECT 232.490 3.555 234.870 4.280 ;
        RECT 235.710 3.555 241.310 4.280 ;
        RECT 242.150 3.555 244.530 4.280 ;
        RECT 245.370 3.555 247.750 4.280 ;
        RECT 248.590 3.555 250.970 4.280 ;
        RECT 251.810 3.555 254.190 4.280 ;
        RECT 255.030 3.555 257.410 4.280 ;
        RECT 258.250 3.555 263.850 4.280 ;
        RECT 264.690 3.555 267.070 4.280 ;
        RECT 267.910 3.555 270.290 4.280 ;
        RECT 271.130 3.555 273.510 4.280 ;
        RECT 274.350 3.555 276.730 4.280 ;
        RECT 277.570 3.555 283.170 4.280 ;
        RECT 284.010 3.555 286.390 4.280 ;
        RECT 287.230 3.555 289.610 4.280 ;
        RECT 290.450 3.555 292.830 4.280 ;
        RECT 293.670 3.555 296.050 4.280 ;
        RECT 296.890 3.555 302.490 4.280 ;
        RECT 303.330 3.555 305.710 4.280 ;
        RECT 306.550 3.555 308.930 4.280 ;
        RECT 309.770 3.555 312.150 4.280 ;
        RECT 312.990 3.555 315.370 4.280 ;
        RECT 316.210 3.555 321.810 4.280 ;
        RECT 322.650 3.555 325.030 4.280 ;
        RECT 325.870 3.555 328.250 4.280 ;
        RECT 329.090 3.555 331.470 4.280 ;
        RECT 332.310 3.555 334.690 4.280 ;
        RECT 335.530 3.555 337.910 4.280 ;
        RECT 338.750 3.555 344.350 4.280 ;
        RECT 345.190 3.555 347.570 4.280 ;
        RECT 348.410 3.555 350.790 4.280 ;
        RECT 351.630 3.555 354.010 4.280 ;
        RECT 354.850 3.555 357.230 4.280 ;
        RECT 358.070 3.555 363.670 4.280 ;
        RECT 364.510 3.555 366.890 4.280 ;
        RECT 367.730 3.555 370.110 4.280 ;
        RECT 370.950 3.555 373.330 4.280 ;
        RECT 374.170 3.555 376.550 4.280 ;
        RECT 377.390 3.555 382.990 4.280 ;
        RECT 383.830 3.555 386.210 4.280 ;
        RECT 387.050 3.555 389.430 4.280 ;
        RECT 390.270 3.555 392.650 4.280 ;
        RECT 393.490 3.555 395.870 4.280 ;
        RECT 396.710 3.555 402.310 4.280 ;
        RECT 403.150 3.555 405.530 4.280 ;
        RECT 406.370 3.555 408.750 4.280 ;
        RECT 409.590 3.555 411.970 4.280 ;
        RECT 412.810 3.555 415.190 4.280 ;
        RECT 416.030 3.555 418.410 4.280 ;
        RECT 419.250 3.555 424.850 4.280 ;
        RECT 425.690 3.555 428.070 4.280 ;
        RECT 428.910 3.555 431.290 4.280 ;
        RECT 432.130 3.555 434.510 4.280 ;
        RECT 435.350 3.555 437.730 4.280 ;
        RECT 438.570 3.555 444.170 4.280 ;
        RECT 445.010 3.555 447.390 4.280 ;
        RECT 448.230 3.555 450.610 4.280 ;
        RECT 451.450 3.555 453.830 4.280 ;
        RECT 454.670 3.555 457.050 4.280 ;
        RECT 457.890 3.555 463.490 4.280 ;
        RECT 464.330 3.555 466.710 4.280 ;
        RECT 467.550 3.555 469.930 4.280 ;
        RECT 470.770 3.555 473.150 4.280 ;
        RECT 473.990 3.555 476.370 4.280 ;
        RECT 477.210 3.555 482.810 4.280 ;
        RECT 483.650 3.555 486.030 4.280 ;
        RECT 486.870 3.555 489.250 4.280 ;
        RECT 490.090 3.555 492.470 4.280 ;
        RECT 493.310 3.555 495.690 4.280 ;
        RECT 496.530 3.555 498.910 4.280 ;
        RECT 499.750 3.555 505.350 4.280 ;
        RECT 506.190 3.555 508.570 4.280 ;
        RECT 509.410 3.555 511.790 4.280 ;
        RECT 512.630 3.555 515.010 4.280 ;
        RECT 515.850 3.555 518.230 4.280 ;
        RECT 519.070 3.555 524.670 4.280 ;
        RECT 525.510 3.555 527.890 4.280 ;
        RECT 528.730 3.555 531.110 4.280 ;
        RECT 531.950 3.555 534.330 4.280 ;
        RECT 535.170 3.555 537.550 4.280 ;
        RECT 538.390 3.555 543.990 4.280 ;
        RECT 544.830 3.555 547.210 4.280 ;
        RECT 548.050 3.555 550.430 4.280 ;
        RECT 551.270 3.555 553.650 4.280 ;
        RECT 554.490 3.555 556.870 4.280 ;
        RECT 557.710 3.555 563.310 4.280 ;
        RECT 564.150 3.555 566.530 4.280 ;
        RECT 567.370 3.555 569.750 4.280 ;
        RECT 570.590 3.555 572.970 4.280 ;
        RECT 573.810 3.555 576.190 4.280 ;
        RECT 577.030 3.555 579.410 4.280 ;
        RECT 580.250 3.555 585.850 4.280 ;
        RECT 586.690 3.555 589.070 4.280 ;
        RECT 589.910 3.555 592.290 4.280 ;
        RECT 593.130 3.555 595.510 4.280 ;
        RECT 596.350 3.555 598.730 4.280 ;
        RECT 599.570 3.555 605.170 4.280 ;
        RECT 606.010 3.555 608.390 4.280 ;
        RECT 609.230 3.555 611.610 4.280 ;
        RECT 612.450 3.555 614.830 4.280 ;
        RECT 615.670 3.555 618.050 4.280 ;
        RECT 618.890 3.555 624.490 4.280 ;
        RECT 625.330 3.555 627.710 4.280 ;
        RECT 628.550 3.555 630.930 4.280 ;
        RECT 631.770 3.555 634.150 4.280 ;
        RECT 634.990 3.555 637.370 4.280 ;
        RECT 638.210 3.555 643.810 4.280 ;
        RECT 644.650 3.555 647.030 4.280 ;
        RECT 647.870 3.555 650.250 4.280 ;
        RECT 651.090 3.555 653.470 4.280 ;
        RECT 654.310 3.555 656.690 4.280 ;
        RECT 657.530 3.555 659.910 4.280 ;
        RECT 660.750 3.555 666.350 4.280 ;
        RECT 667.190 3.555 669.570 4.280 ;
        RECT 670.410 3.555 672.790 4.280 ;
        RECT 673.630 3.555 676.010 4.280 ;
        RECT 676.850 3.555 679.230 4.280 ;
        RECT 680.070 3.555 685.670 4.280 ;
        RECT 686.510 3.555 688.890 4.280 ;
        RECT 689.730 3.555 692.110 4.280 ;
        RECT 692.950 3.555 695.330 4.280 ;
        RECT 696.170 3.555 698.550 4.280 ;
        RECT 699.390 3.555 699.960 4.280 ;
      LAYER met3 ;
        RECT 4.400 2196.040 695.600 2196.905 ;
        RECT 0.985 2194.040 699.850 2196.040 ;
        RECT 4.400 2192.640 695.600 2194.040 ;
        RECT 0.985 2190.640 699.850 2192.640 ;
        RECT 4.400 2189.240 695.600 2190.640 ;
        RECT 0.985 2183.840 699.850 2189.240 ;
        RECT 4.400 2182.440 695.600 2183.840 ;
        RECT 0.985 2180.440 699.850 2182.440 ;
        RECT 4.400 2179.040 695.600 2180.440 ;
        RECT 0.985 2177.040 699.850 2179.040 ;
        RECT 4.400 2175.640 695.600 2177.040 ;
        RECT 0.985 2173.640 699.850 2175.640 ;
        RECT 4.400 2172.240 695.600 2173.640 ;
        RECT 0.985 2170.240 699.850 2172.240 ;
        RECT 4.400 2168.840 695.600 2170.240 ;
        RECT 0.985 2163.440 699.850 2168.840 ;
        RECT 4.400 2162.040 695.600 2163.440 ;
        RECT 0.985 2160.040 699.850 2162.040 ;
        RECT 4.400 2158.640 695.600 2160.040 ;
        RECT 0.985 2156.640 699.850 2158.640 ;
        RECT 4.400 2155.240 695.600 2156.640 ;
        RECT 0.985 2153.240 699.850 2155.240 ;
        RECT 4.400 2151.840 695.600 2153.240 ;
        RECT 0.985 2149.840 699.850 2151.840 ;
        RECT 4.400 2148.440 695.600 2149.840 ;
        RECT 0.985 2146.440 699.850 2148.440 ;
        RECT 4.400 2145.040 699.850 2146.440 ;
        RECT 0.985 2143.040 699.850 2145.040 ;
        RECT 0.985 2141.640 695.600 2143.040 ;
        RECT 0.985 2139.640 699.850 2141.640 ;
        RECT 4.400 2138.240 695.600 2139.640 ;
        RECT 0.985 2136.240 699.850 2138.240 ;
        RECT 4.400 2134.840 695.600 2136.240 ;
        RECT 0.985 2132.840 699.850 2134.840 ;
        RECT 4.400 2131.440 695.600 2132.840 ;
        RECT 0.985 2129.440 699.850 2131.440 ;
        RECT 4.400 2128.040 695.600 2129.440 ;
        RECT 0.985 2126.040 699.850 2128.040 ;
        RECT 4.400 2124.640 699.850 2126.040 ;
        RECT 0.985 2122.640 699.850 2124.640 ;
        RECT 0.985 2121.240 695.600 2122.640 ;
        RECT 0.985 2119.240 699.850 2121.240 ;
        RECT 4.400 2117.840 695.600 2119.240 ;
        RECT 0.985 2115.840 699.850 2117.840 ;
        RECT 4.400 2114.440 695.600 2115.840 ;
        RECT 0.985 2112.440 699.850 2114.440 ;
        RECT 4.400 2111.040 695.600 2112.440 ;
        RECT 0.985 2109.040 699.850 2111.040 ;
        RECT 4.400 2107.640 695.600 2109.040 ;
        RECT 0.985 2105.640 699.850 2107.640 ;
        RECT 4.400 2104.240 695.600 2105.640 ;
        RECT 0.985 2098.840 699.850 2104.240 ;
        RECT 4.400 2097.440 695.600 2098.840 ;
        RECT 0.985 2095.440 699.850 2097.440 ;
        RECT 4.400 2094.040 695.600 2095.440 ;
        RECT 0.985 2092.040 699.850 2094.040 ;
        RECT 4.400 2090.640 695.600 2092.040 ;
        RECT 0.985 2088.640 699.850 2090.640 ;
        RECT 4.400 2087.240 695.600 2088.640 ;
        RECT 0.985 2085.240 699.850 2087.240 ;
        RECT 4.400 2083.840 695.600 2085.240 ;
        RECT 0.985 2078.440 699.850 2083.840 ;
        RECT 4.400 2077.040 695.600 2078.440 ;
        RECT 0.985 2075.040 699.850 2077.040 ;
        RECT 4.400 2073.640 695.600 2075.040 ;
        RECT 0.985 2071.640 699.850 2073.640 ;
        RECT 4.400 2070.240 695.600 2071.640 ;
        RECT 0.985 2068.240 699.850 2070.240 ;
        RECT 4.400 2066.840 695.600 2068.240 ;
        RECT 0.985 2064.840 699.850 2066.840 ;
        RECT 4.400 2063.440 695.600 2064.840 ;
        RECT 0.985 2061.440 699.850 2063.440 ;
        RECT 4.400 2060.040 699.850 2061.440 ;
        RECT 0.985 2058.040 699.850 2060.040 ;
        RECT 0.985 2056.640 695.600 2058.040 ;
        RECT 0.985 2054.640 699.850 2056.640 ;
        RECT 4.400 2053.240 695.600 2054.640 ;
        RECT 0.985 2051.240 699.850 2053.240 ;
        RECT 4.400 2049.840 695.600 2051.240 ;
        RECT 0.985 2047.840 699.850 2049.840 ;
        RECT 4.400 2046.440 695.600 2047.840 ;
        RECT 0.985 2044.440 699.850 2046.440 ;
        RECT 4.400 2043.040 695.600 2044.440 ;
        RECT 0.985 2041.040 699.850 2043.040 ;
        RECT 4.400 2039.640 699.850 2041.040 ;
        RECT 0.985 2037.640 699.850 2039.640 ;
        RECT 0.985 2036.240 695.600 2037.640 ;
        RECT 0.985 2034.240 699.850 2036.240 ;
        RECT 4.400 2032.840 695.600 2034.240 ;
        RECT 0.985 2030.840 699.850 2032.840 ;
        RECT 4.400 2029.440 695.600 2030.840 ;
        RECT 0.985 2027.440 699.850 2029.440 ;
        RECT 4.400 2026.040 695.600 2027.440 ;
        RECT 0.985 2024.040 699.850 2026.040 ;
        RECT 4.400 2022.640 695.600 2024.040 ;
        RECT 0.985 2020.640 699.850 2022.640 ;
        RECT 4.400 2019.240 695.600 2020.640 ;
        RECT 0.985 2013.840 699.850 2019.240 ;
        RECT 4.400 2012.440 695.600 2013.840 ;
        RECT 0.985 2010.440 699.850 2012.440 ;
        RECT 4.400 2009.040 695.600 2010.440 ;
        RECT 0.985 2007.040 699.850 2009.040 ;
        RECT 4.400 2005.640 695.600 2007.040 ;
        RECT 0.985 2003.640 699.850 2005.640 ;
        RECT 4.400 2002.240 695.600 2003.640 ;
        RECT 0.985 2000.240 699.850 2002.240 ;
        RECT 4.400 1998.840 695.600 2000.240 ;
        RECT 0.985 1993.440 699.850 1998.840 ;
        RECT 4.400 1992.040 695.600 1993.440 ;
        RECT 0.985 1990.040 699.850 1992.040 ;
        RECT 4.400 1988.640 695.600 1990.040 ;
        RECT 0.985 1986.640 699.850 1988.640 ;
        RECT 4.400 1985.240 695.600 1986.640 ;
        RECT 0.985 1983.240 699.850 1985.240 ;
        RECT 4.400 1981.840 695.600 1983.240 ;
        RECT 0.985 1979.840 699.850 1981.840 ;
        RECT 4.400 1978.440 695.600 1979.840 ;
        RECT 0.985 1976.440 699.850 1978.440 ;
        RECT 4.400 1975.040 699.850 1976.440 ;
        RECT 0.985 1973.040 699.850 1975.040 ;
        RECT 0.985 1971.640 695.600 1973.040 ;
        RECT 0.985 1969.640 699.850 1971.640 ;
        RECT 4.400 1968.240 695.600 1969.640 ;
        RECT 0.985 1966.240 699.850 1968.240 ;
        RECT 4.400 1964.840 695.600 1966.240 ;
        RECT 0.985 1962.840 699.850 1964.840 ;
        RECT 4.400 1961.440 695.600 1962.840 ;
        RECT 0.985 1959.440 699.850 1961.440 ;
        RECT 4.400 1958.040 695.600 1959.440 ;
        RECT 0.985 1956.040 699.850 1958.040 ;
        RECT 4.400 1954.640 699.850 1956.040 ;
        RECT 0.985 1952.640 699.850 1954.640 ;
        RECT 0.985 1951.240 695.600 1952.640 ;
        RECT 0.985 1949.240 699.850 1951.240 ;
        RECT 4.400 1947.840 695.600 1949.240 ;
        RECT 0.985 1945.840 699.850 1947.840 ;
        RECT 4.400 1944.440 695.600 1945.840 ;
        RECT 0.985 1942.440 699.850 1944.440 ;
        RECT 4.400 1941.040 695.600 1942.440 ;
        RECT 0.985 1939.040 699.850 1941.040 ;
        RECT 4.400 1937.640 695.600 1939.040 ;
        RECT 0.985 1935.640 699.850 1937.640 ;
        RECT 4.400 1934.240 695.600 1935.640 ;
        RECT 0.985 1928.840 699.850 1934.240 ;
        RECT 4.400 1927.440 695.600 1928.840 ;
        RECT 0.985 1925.440 699.850 1927.440 ;
        RECT 4.400 1924.040 695.600 1925.440 ;
        RECT 0.985 1922.040 699.850 1924.040 ;
        RECT 4.400 1920.640 695.600 1922.040 ;
        RECT 0.985 1918.640 699.850 1920.640 ;
        RECT 4.400 1917.240 695.600 1918.640 ;
        RECT 0.985 1915.240 699.850 1917.240 ;
        RECT 4.400 1913.840 695.600 1915.240 ;
        RECT 0.985 1908.440 699.850 1913.840 ;
        RECT 4.400 1907.040 695.600 1908.440 ;
        RECT 0.985 1905.040 699.850 1907.040 ;
        RECT 4.400 1903.640 695.600 1905.040 ;
        RECT 0.985 1901.640 699.850 1903.640 ;
        RECT 4.400 1900.240 695.600 1901.640 ;
        RECT 0.985 1898.240 699.850 1900.240 ;
        RECT 4.400 1896.840 695.600 1898.240 ;
        RECT 0.985 1894.840 699.850 1896.840 ;
        RECT 4.400 1893.440 695.600 1894.840 ;
        RECT 0.985 1891.440 699.850 1893.440 ;
        RECT 4.400 1890.040 699.850 1891.440 ;
        RECT 0.985 1888.040 699.850 1890.040 ;
        RECT 0.985 1886.640 695.600 1888.040 ;
        RECT 0.985 1884.640 699.850 1886.640 ;
        RECT 4.400 1883.240 695.600 1884.640 ;
        RECT 0.985 1881.240 699.850 1883.240 ;
        RECT 4.400 1879.840 695.600 1881.240 ;
        RECT 0.985 1877.840 699.850 1879.840 ;
        RECT 4.400 1876.440 695.600 1877.840 ;
        RECT 0.985 1874.440 699.850 1876.440 ;
        RECT 4.400 1873.040 695.600 1874.440 ;
        RECT 0.985 1871.040 699.850 1873.040 ;
        RECT 4.400 1869.640 699.850 1871.040 ;
        RECT 0.985 1867.640 699.850 1869.640 ;
        RECT 0.985 1866.240 695.600 1867.640 ;
        RECT 0.985 1864.240 699.850 1866.240 ;
        RECT 4.400 1862.840 695.600 1864.240 ;
        RECT 0.985 1860.840 699.850 1862.840 ;
        RECT 4.400 1859.440 695.600 1860.840 ;
        RECT 0.985 1857.440 699.850 1859.440 ;
        RECT 4.400 1856.040 695.600 1857.440 ;
        RECT 0.985 1854.040 699.850 1856.040 ;
        RECT 4.400 1852.640 695.600 1854.040 ;
        RECT 0.985 1850.640 699.850 1852.640 ;
        RECT 4.400 1849.240 695.600 1850.640 ;
        RECT 0.985 1843.840 699.850 1849.240 ;
        RECT 4.400 1842.440 695.600 1843.840 ;
        RECT 0.985 1840.440 699.850 1842.440 ;
        RECT 4.400 1839.040 695.600 1840.440 ;
        RECT 0.985 1837.040 699.850 1839.040 ;
        RECT 4.400 1835.640 695.600 1837.040 ;
        RECT 0.985 1833.640 699.850 1835.640 ;
        RECT 4.400 1832.240 695.600 1833.640 ;
        RECT 0.985 1830.240 699.850 1832.240 ;
        RECT 4.400 1828.840 695.600 1830.240 ;
        RECT 0.985 1823.440 699.850 1828.840 ;
        RECT 4.400 1822.040 695.600 1823.440 ;
        RECT 0.985 1820.040 699.850 1822.040 ;
        RECT 4.400 1818.640 695.600 1820.040 ;
        RECT 0.985 1816.640 699.850 1818.640 ;
        RECT 4.400 1815.240 695.600 1816.640 ;
        RECT 0.985 1813.240 699.850 1815.240 ;
        RECT 4.400 1811.840 695.600 1813.240 ;
        RECT 0.985 1809.840 699.850 1811.840 ;
        RECT 4.400 1808.440 695.600 1809.840 ;
        RECT 0.985 1806.440 699.850 1808.440 ;
        RECT 4.400 1805.040 699.850 1806.440 ;
        RECT 0.985 1803.040 699.850 1805.040 ;
        RECT 0.985 1801.640 695.600 1803.040 ;
        RECT 0.985 1799.640 699.850 1801.640 ;
        RECT 4.400 1798.240 695.600 1799.640 ;
        RECT 0.985 1796.240 699.850 1798.240 ;
        RECT 4.400 1794.840 695.600 1796.240 ;
        RECT 0.985 1792.840 699.850 1794.840 ;
        RECT 4.400 1791.440 695.600 1792.840 ;
        RECT 0.985 1789.440 699.850 1791.440 ;
        RECT 4.400 1788.040 695.600 1789.440 ;
        RECT 0.985 1786.040 699.850 1788.040 ;
        RECT 4.400 1784.640 699.850 1786.040 ;
        RECT 0.985 1782.640 699.850 1784.640 ;
        RECT 0.985 1781.240 695.600 1782.640 ;
        RECT 0.985 1779.240 699.850 1781.240 ;
        RECT 4.400 1777.840 695.600 1779.240 ;
        RECT 0.985 1775.840 699.850 1777.840 ;
        RECT 4.400 1774.440 695.600 1775.840 ;
        RECT 0.985 1772.440 699.850 1774.440 ;
        RECT 4.400 1771.040 695.600 1772.440 ;
        RECT 0.985 1769.040 699.850 1771.040 ;
        RECT 4.400 1767.640 695.600 1769.040 ;
        RECT 0.985 1765.640 699.850 1767.640 ;
        RECT 4.400 1764.240 695.600 1765.640 ;
        RECT 0.985 1758.840 699.850 1764.240 ;
        RECT 4.400 1757.440 695.600 1758.840 ;
        RECT 0.985 1755.440 699.850 1757.440 ;
        RECT 4.400 1754.040 695.600 1755.440 ;
        RECT 0.985 1752.040 699.850 1754.040 ;
        RECT 4.400 1750.640 695.600 1752.040 ;
        RECT 0.985 1748.640 699.850 1750.640 ;
        RECT 4.400 1747.240 695.600 1748.640 ;
        RECT 0.985 1745.240 699.850 1747.240 ;
        RECT 4.400 1743.840 695.600 1745.240 ;
        RECT 0.985 1738.440 699.850 1743.840 ;
        RECT 4.400 1737.040 695.600 1738.440 ;
        RECT 0.985 1735.040 699.850 1737.040 ;
        RECT 4.400 1733.640 695.600 1735.040 ;
        RECT 0.985 1731.640 699.850 1733.640 ;
        RECT 4.400 1730.240 695.600 1731.640 ;
        RECT 0.985 1728.240 699.850 1730.240 ;
        RECT 4.400 1726.840 695.600 1728.240 ;
        RECT 0.985 1724.840 699.850 1726.840 ;
        RECT 4.400 1723.440 695.600 1724.840 ;
        RECT 0.985 1721.440 699.850 1723.440 ;
        RECT 4.400 1720.040 699.850 1721.440 ;
        RECT 0.985 1718.040 699.850 1720.040 ;
        RECT 0.985 1716.640 695.600 1718.040 ;
        RECT 0.985 1714.640 699.850 1716.640 ;
        RECT 4.400 1713.240 695.600 1714.640 ;
        RECT 0.985 1711.240 699.850 1713.240 ;
        RECT 4.400 1709.840 695.600 1711.240 ;
        RECT 0.985 1707.840 699.850 1709.840 ;
        RECT 4.400 1706.440 695.600 1707.840 ;
        RECT 0.985 1704.440 699.850 1706.440 ;
        RECT 4.400 1703.040 695.600 1704.440 ;
        RECT 0.985 1701.040 699.850 1703.040 ;
        RECT 4.400 1699.640 699.850 1701.040 ;
        RECT 0.985 1697.640 699.850 1699.640 ;
        RECT 0.985 1696.240 695.600 1697.640 ;
        RECT 0.985 1694.240 699.850 1696.240 ;
        RECT 4.400 1692.840 695.600 1694.240 ;
        RECT 0.985 1690.840 699.850 1692.840 ;
        RECT 4.400 1689.440 695.600 1690.840 ;
        RECT 0.985 1687.440 699.850 1689.440 ;
        RECT 4.400 1686.040 695.600 1687.440 ;
        RECT 0.985 1684.040 699.850 1686.040 ;
        RECT 4.400 1682.640 695.600 1684.040 ;
        RECT 0.985 1680.640 699.850 1682.640 ;
        RECT 4.400 1679.240 695.600 1680.640 ;
        RECT 0.985 1673.840 699.850 1679.240 ;
        RECT 4.400 1672.440 695.600 1673.840 ;
        RECT 0.985 1670.440 699.850 1672.440 ;
        RECT 4.400 1669.040 695.600 1670.440 ;
        RECT 0.985 1667.040 699.850 1669.040 ;
        RECT 4.400 1665.640 695.600 1667.040 ;
        RECT 0.985 1663.640 699.850 1665.640 ;
        RECT 4.400 1662.240 695.600 1663.640 ;
        RECT 0.985 1660.240 699.850 1662.240 ;
        RECT 4.400 1658.840 695.600 1660.240 ;
        RECT 0.985 1653.440 699.850 1658.840 ;
        RECT 4.400 1652.040 695.600 1653.440 ;
        RECT 0.985 1650.040 699.850 1652.040 ;
        RECT 4.400 1648.640 695.600 1650.040 ;
        RECT 0.985 1646.640 699.850 1648.640 ;
        RECT 4.400 1645.240 695.600 1646.640 ;
        RECT 0.985 1643.240 699.850 1645.240 ;
        RECT 4.400 1641.840 695.600 1643.240 ;
        RECT 0.985 1639.840 699.850 1641.840 ;
        RECT 4.400 1638.440 695.600 1639.840 ;
        RECT 0.985 1636.440 699.850 1638.440 ;
        RECT 4.400 1635.040 699.850 1636.440 ;
        RECT 0.985 1633.040 699.850 1635.040 ;
        RECT 0.985 1631.640 695.600 1633.040 ;
        RECT 0.985 1629.640 699.850 1631.640 ;
        RECT 4.400 1628.240 695.600 1629.640 ;
        RECT 0.985 1626.240 699.850 1628.240 ;
        RECT 4.400 1624.840 695.600 1626.240 ;
        RECT 0.985 1622.840 699.850 1624.840 ;
        RECT 4.400 1621.440 695.600 1622.840 ;
        RECT 0.985 1619.440 699.850 1621.440 ;
        RECT 4.400 1618.040 695.600 1619.440 ;
        RECT 0.985 1616.040 699.850 1618.040 ;
        RECT 4.400 1614.640 699.850 1616.040 ;
        RECT 0.985 1612.640 699.850 1614.640 ;
        RECT 0.985 1611.240 695.600 1612.640 ;
        RECT 0.985 1609.240 699.850 1611.240 ;
        RECT 4.400 1607.840 695.600 1609.240 ;
        RECT 0.985 1605.840 699.850 1607.840 ;
        RECT 4.400 1604.440 695.600 1605.840 ;
        RECT 0.985 1602.440 699.850 1604.440 ;
        RECT 4.400 1601.040 695.600 1602.440 ;
        RECT 0.985 1599.040 699.850 1601.040 ;
        RECT 4.400 1597.640 695.600 1599.040 ;
        RECT 0.985 1595.640 699.850 1597.640 ;
        RECT 4.400 1594.240 699.850 1595.640 ;
        RECT 0.985 1592.240 699.850 1594.240 ;
        RECT 0.985 1590.840 695.600 1592.240 ;
        RECT 0.985 1588.840 699.850 1590.840 ;
        RECT 4.400 1587.440 695.600 1588.840 ;
        RECT 0.985 1585.440 699.850 1587.440 ;
        RECT 4.400 1584.040 695.600 1585.440 ;
        RECT 0.985 1582.040 699.850 1584.040 ;
        RECT 4.400 1580.640 695.600 1582.040 ;
        RECT 0.985 1578.640 699.850 1580.640 ;
        RECT 4.400 1577.240 695.600 1578.640 ;
        RECT 0.985 1575.240 699.850 1577.240 ;
        RECT 4.400 1573.840 695.600 1575.240 ;
        RECT 0.985 1568.440 699.850 1573.840 ;
        RECT 4.400 1567.040 695.600 1568.440 ;
        RECT 0.985 1565.040 699.850 1567.040 ;
        RECT 4.400 1563.640 695.600 1565.040 ;
        RECT 0.985 1561.640 699.850 1563.640 ;
        RECT 4.400 1560.240 695.600 1561.640 ;
        RECT 0.985 1558.240 699.850 1560.240 ;
        RECT 4.400 1556.840 695.600 1558.240 ;
        RECT 0.985 1554.840 699.850 1556.840 ;
        RECT 4.400 1553.440 695.600 1554.840 ;
        RECT 0.985 1551.440 699.850 1553.440 ;
        RECT 4.400 1550.040 699.850 1551.440 ;
        RECT 0.985 1548.040 699.850 1550.040 ;
        RECT 0.985 1546.640 695.600 1548.040 ;
        RECT 0.985 1544.640 699.850 1546.640 ;
        RECT 4.400 1543.240 695.600 1544.640 ;
        RECT 0.985 1541.240 699.850 1543.240 ;
        RECT 4.400 1539.840 695.600 1541.240 ;
        RECT 0.985 1537.840 699.850 1539.840 ;
        RECT 4.400 1536.440 695.600 1537.840 ;
        RECT 0.985 1534.440 699.850 1536.440 ;
        RECT 4.400 1533.040 695.600 1534.440 ;
        RECT 0.985 1531.040 699.850 1533.040 ;
        RECT 4.400 1529.640 699.850 1531.040 ;
        RECT 0.985 1527.640 699.850 1529.640 ;
        RECT 0.985 1526.240 695.600 1527.640 ;
        RECT 0.985 1524.240 699.850 1526.240 ;
        RECT 4.400 1522.840 695.600 1524.240 ;
        RECT 0.985 1520.840 699.850 1522.840 ;
        RECT 4.400 1519.440 695.600 1520.840 ;
        RECT 0.985 1517.440 699.850 1519.440 ;
        RECT 4.400 1516.040 695.600 1517.440 ;
        RECT 0.985 1514.040 699.850 1516.040 ;
        RECT 4.400 1512.640 695.600 1514.040 ;
        RECT 0.985 1510.640 699.850 1512.640 ;
        RECT 4.400 1509.240 699.850 1510.640 ;
        RECT 0.985 1507.240 699.850 1509.240 ;
        RECT 0.985 1505.840 695.600 1507.240 ;
        RECT 0.985 1503.840 699.850 1505.840 ;
        RECT 4.400 1502.440 695.600 1503.840 ;
        RECT 0.985 1500.440 699.850 1502.440 ;
        RECT 4.400 1499.040 695.600 1500.440 ;
        RECT 0.985 1497.040 699.850 1499.040 ;
        RECT 4.400 1495.640 695.600 1497.040 ;
        RECT 0.985 1493.640 699.850 1495.640 ;
        RECT 4.400 1492.240 695.600 1493.640 ;
        RECT 0.985 1490.240 699.850 1492.240 ;
        RECT 4.400 1488.840 695.600 1490.240 ;
        RECT 0.985 1483.440 699.850 1488.840 ;
        RECT 4.400 1482.040 695.600 1483.440 ;
        RECT 0.985 1480.040 699.850 1482.040 ;
        RECT 4.400 1478.640 695.600 1480.040 ;
        RECT 0.985 1476.640 699.850 1478.640 ;
        RECT 4.400 1475.240 695.600 1476.640 ;
        RECT 0.985 1473.240 699.850 1475.240 ;
        RECT 4.400 1471.840 695.600 1473.240 ;
        RECT 0.985 1469.840 699.850 1471.840 ;
        RECT 4.400 1468.440 695.600 1469.840 ;
        RECT 0.985 1466.440 699.850 1468.440 ;
        RECT 4.400 1465.040 699.850 1466.440 ;
        RECT 0.985 1463.040 699.850 1465.040 ;
        RECT 0.985 1461.640 695.600 1463.040 ;
        RECT 0.985 1459.640 699.850 1461.640 ;
        RECT 4.400 1458.240 695.600 1459.640 ;
        RECT 0.985 1456.240 699.850 1458.240 ;
        RECT 4.400 1454.840 695.600 1456.240 ;
        RECT 0.985 1452.840 699.850 1454.840 ;
        RECT 4.400 1451.440 695.600 1452.840 ;
        RECT 0.985 1449.440 699.850 1451.440 ;
        RECT 4.400 1448.040 695.600 1449.440 ;
        RECT 0.985 1446.040 699.850 1448.040 ;
        RECT 4.400 1444.640 699.850 1446.040 ;
        RECT 0.985 1442.640 699.850 1444.640 ;
        RECT 0.985 1441.240 695.600 1442.640 ;
        RECT 0.985 1439.240 699.850 1441.240 ;
        RECT 4.400 1437.840 695.600 1439.240 ;
        RECT 0.985 1435.840 699.850 1437.840 ;
        RECT 4.400 1434.440 695.600 1435.840 ;
        RECT 0.985 1432.440 699.850 1434.440 ;
        RECT 4.400 1431.040 695.600 1432.440 ;
        RECT 0.985 1429.040 699.850 1431.040 ;
        RECT 4.400 1427.640 695.600 1429.040 ;
        RECT 0.985 1425.640 699.850 1427.640 ;
        RECT 4.400 1424.240 699.850 1425.640 ;
        RECT 0.985 1422.240 699.850 1424.240 ;
        RECT 0.985 1420.840 695.600 1422.240 ;
        RECT 0.985 1418.840 699.850 1420.840 ;
        RECT 4.400 1417.440 695.600 1418.840 ;
        RECT 0.985 1415.440 699.850 1417.440 ;
        RECT 4.400 1414.040 695.600 1415.440 ;
        RECT 0.985 1412.040 699.850 1414.040 ;
        RECT 4.400 1410.640 695.600 1412.040 ;
        RECT 0.985 1408.640 699.850 1410.640 ;
        RECT 4.400 1407.240 695.600 1408.640 ;
        RECT 0.985 1405.240 699.850 1407.240 ;
        RECT 4.400 1403.840 695.600 1405.240 ;
        RECT 0.985 1398.440 699.850 1403.840 ;
        RECT 4.400 1397.040 695.600 1398.440 ;
        RECT 0.985 1395.040 699.850 1397.040 ;
        RECT 4.400 1393.640 695.600 1395.040 ;
        RECT 0.985 1391.640 699.850 1393.640 ;
        RECT 4.400 1390.240 695.600 1391.640 ;
        RECT 0.985 1388.240 699.850 1390.240 ;
        RECT 4.400 1386.840 695.600 1388.240 ;
        RECT 0.985 1384.840 699.850 1386.840 ;
        RECT 4.400 1383.440 695.600 1384.840 ;
        RECT 0.985 1381.440 699.850 1383.440 ;
        RECT 4.400 1380.040 699.850 1381.440 ;
        RECT 0.985 1378.040 699.850 1380.040 ;
        RECT 0.985 1376.640 695.600 1378.040 ;
        RECT 0.985 1374.640 699.850 1376.640 ;
        RECT 4.400 1373.240 695.600 1374.640 ;
        RECT 0.985 1371.240 699.850 1373.240 ;
        RECT 4.400 1369.840 695.600 1371.240 ;
        RECT 0.985 1367.840 699.850 1369.840 ;
        RECT 4.400 1366.440 695.600 1367.840 ;
        RECT 0.985 1364.440 699.850 1366.440 ;
        RECT 4.400 1363.040 695.600 1364.440 ;
        RECT 0.985 1361.040 699.850 1363.040 ;
        RECT 4.400 1359.640 699.850 1361.040 ;
        RECT 0.985 1357.640 699.850 1359.640 ;
        RECT 0.985 1356.240 695.600 1357.640 ;
        RECT 0.985 1354.240 699.850 1356.240 ;
        RECT 4.400 1352.840 695.600 1354.240 ;
        RECT 0.985 1350.840 699.850 1352.840 ;
        RECT 4.400 1349.440 695.600 1350.840 ;
        RECT 0.985 1347.440 699.850 1349.440 ;
        RECT 4.400 1346.040 695.600 1347.440 ;
        RECT 0.985 1344.040 699.850 1346.040 ;
        RECT 4.400 1342.640 695.600 1344.040 ;
        RECT 0.985 1340.640 699.850 1342.640 ;
        RECT 4.400 1339.240 699.850 1340.640 ;
        RECT 0.985 1337.240 699.850 1339.240 ;
        RECT 0.985 1335.840 695.600 1337.240 ;
        RECT 0.985 1333.840 699.850 1335.840 ;
        RECT 4.400 1332.440 695.600 1333.840 ;
        RECT 0.985 1330.440 699.850 1332.440 ;
        RECT 4.400 1329.040 695.600 1330.440 ;
        RECT 0.985 1327.040 699.850 1329.040 ;
        RECT 4.400 1325.640 695.600 1327.040 ;
        RECT 0.985 1323.640 699.850 1325.640 ;
        RECT 4.400 1322.240 695.600 1323.640 ;
        RECT 0.985 1320.240 699.850 1322.240 ;
        RECT 4.400 1318.840 695.600 1320.240 ;
        RECT 0.985 1313.440 699.850 1318.840 ;
        RECT 4.400 1312.040 695.600 1313.440 ;
        RECT 0.985 1310.040 699.850 1312.040 ;
        RECT 4.400 1308.640 695.600 1310.040 ;
        RECT 0.985 1306.640 699.850 1308.640 ;
        RECT 4.400 1305.240 695.600 1306.640 ;
        RECT 0.985 1303.240 699.850 1305.240 ;
        RECT 4.400 1301.840 695.600 1303.240 ;
        RECT 0.985 1299.840 699.850 1301.840 ;
        RECT 4.400 1298.440 695.600 1299.840 ;
        RECT 0.985 1296.440 699.850 1298.440 ;
        RECT 4.400 1295.040 699.850 1296.440 ;
        RECT 0.985 1293.040 699.850 1295.040 ;
        RECT 0.985 1291.640 695.600 1293.040 ;
        RECT 0.985 1289.640 699.850 1291.640 ;
        RECT 4.400 1288.240 695.600 1289.640 ;
        RECT 0.985 1286.240 699.850 1288.240 ;
        RECT 4.400 1284.840 695.600 1286.240 ;
        RECT 0.985 1282.840 699.850 1284.840 ;
        RECT 4.400 1281.440 695.600 1282.840 ;
        RECT 0.985 1279.440 699.850 1281.440 ;
        RECT 4.400 1278.040 695.600 1279.440 ;
        RECT 0.985 1276.040 699.850 1278.040 ;
        RECT 4.400 1274.640 699.850 1276.040 ;
        RECT 0.985 1272.640 699.850 1274.640 ;
        RECT 0.985 1271.240 695.600 1272.640 ;
        RECT 0.985 1269.240 699.850 1271.240 ;
        RECT 4.400 1267.840 695.600 1269.240 ;
        RECT 0.985 1265.840 699.850 1267.840 ;
        RECT 4.400 1264.440 695.600 1265.840 ;
        RECT 0.985 1262.440 699.850 1264.440 ;
        RECT 4.400 1261.040 695.600 1262.440 ;
        RECT 0.985 1259.040 699.850 1261.040 ;
        RECT 4.400 1257.640 695.600 1259.040 ;
        RECT 0.985 1255.640 699.850 1257.640 ;
        RECT 4.400 1254.240 699.850 1255.640 ;
        RECT 0.985 1252.240 699.850 1254.240 ;
        RECT 0.985 1250.840 695.600 1252.240 ;
        RECT 0.985 1248.840 699.850 1250.840 ;
        RECT 4.400 1247.440 695.600 1248.840 ;
        RECT 0.985 1245.440 699.850 1247.440 ;
        RECT 4.400 1244.040 695.600 1245.440 ;
        RECT 0.985 1242.040 699.850 1244.040 ;
        RECT 4.400 1240.640 695.600 1242.040 ;
        RECT 0.985 1238.640 699.850 1240.640 ;
        RECT 4.400 1237.240 695.600 1238.640 ;
        RECT 0.985 1235.240 699.850 1237.240 ;
        RECT 4.400 1233.840 695.600 1235.240 ;
        RECT 0.985 1228.440 699.850 1233.840 ;
        RECT 4.400 1227.040 695.600 1228.440 ;
        RECT 0.985 1225.040 699.850 1227.040 ;
        RECT 4.400 1223.640 695.600 1225.040 ;
        RECT 0.985 1221.640 699.850 1223.640 ;
        RECT 4.400 1220.240 695.600 1221.640 ;
        RECT 0.985 1218.240 699.850 1220.240 ;
        RECT 4.400 1216.840 695.600 1218.240 ;
        RECT 0.985 1214.840 699.850 1216.840 ;
        RECT 4.400 1213.440 695.600 1214.840 ;
        RECT 0.985 1211.440 699.850 1213.440 ;
        RECT 4.400 1210.040 699.850 1211.440 ;
        RECT 0.985 1208.040 699.850 1210.040 ;
        RECT 0.985 1206.640 695.600 1208.040 ;
        RECT 0.985 1204.640 699.850 1206.640 ;
        RECT 4.400 1203.240 695.600 1204.640 ;
        RECT 0.985 1201.240 699.850 1203.240 ;
        RECT 4.400 1199.840 695.600 1201.240 ;
        RECT 0.985 1197.840 699.850 1199.840 ;
        RECT 4.400 1196.440 695.600 1197.840 ;
        RECT 0.985 1194.440 699.850 1196.440 ;
        RECT 4.400 1193.040 695.600 1194.440 ;
        RECT 0.985 1191.040 699.850 1193.040 ;
        RECT 4.400 1189.640 699.850 1191.040 ;
        RECT 0.985 1187.640 699.850 1189.640 ;
        RECT 0.985 1186.240 695.600 1187.640 ;
        RECT 0.985 1184.240 699.850 1186.240 ;
        RECT 4.400 1182.840 695.600 1184.240 ;
        RECT 0.985 1180.840 699.850 1182.840 ;
        RECT 4.400 1179.440 695.600 1180.840 ;
        RECT 0.985 1177.440 699.850 1179.440 ;
        RECT 4.400 1176.040 695.600 1177.440 ;
        RECT 0.985 1174.040 699.850 1176.040 ;
        RECT 4.400 1172.640 695.600 1174.040 ;
        RECT 0.985 1170.640 699.850 1172.640 ;
        RECT 4.400 1169.240 699.850 1170.640 ;
        RECT 0.985 1167.240 699.850 1169.240 ;
        RECT 0.985 1165.840 695.600 1167.240 ;
        RECT 0.985 1163.840 699.850 1165.840 ;
        RECT 4.400 1162.440 695.600 1163.840 ;
        RECT 0.985 1160.440 699.850 1162.440 ;
        RECT 4.400 1159.040 695.600 1160.440 ;
        RECT 0.985 1157.040 699.850 1159.040 ;
        RECT 4.400 1155.640 695.600 1157.040 ;
        RECT 0.985 1153.640 699.850 1155.640 ;
        RECT 4.400 1152.240 695.600 1153.640 ;
        RECT 0.985 1150.240 699.850 1152.240 ;
        RECT 4.400 1148.840 695.600 1150.240 ;
        RECT 0.985 1143.440 699.850 1148.840 ;
        RECT 4.400 1142.040 695.600 1143.440 ;
        RECT 0.985 1140.040 699.850 1142.040 ;
        RECT 4.400 1138.640 695.600 1140.040 ;
        RECT 0.985 1136.640 699.850 1138.640 ;
        RECT 4.400 1135.240 695.600 1136.640 ;
        RECT 0.985 1133.240 699.850 1135.240 ;
        RECT 4.400 1131.840 695.600 1133.240 ;
        RECT 0.985 1129.840 699.850 1131.840 ;
        RECT 4.400 1128.440 695.600 1129.840 ;
        RECT 0.985 1123.040 699.850 1128.440 ;
        RECT 4.400 1121.640 695.600 1123.040 ;
        RECT 0.985 1119.640 699.850 1121.640 ;
        RECT 4.400 1118.240 695.600 1119.640 ;
        RECT 0.985 1116.240 699.850 1118.240 ;
        RECT 4.400 1114.840 695.600 1116.240 ;
        RECT 0.985 1112.840 699.850 1114.840 ;
        RECT 4.400 1111.440 695.600 1112.840 ;
        RECT 0.985 1109.440 699.850 1111.440 ;
        RECT 4.400 1108.040 695.600 1109.440 ;
        RECT 0.985 1106.040 699.850 1108.040 ;
        RECT 4.400 1104.640 699.850 1106.040 ;
        RECT 0.985 1102.640 699.850 1104.640 ;
        RECT 0.985 1101.240 695.600 1102.640 ;
        RECT 0.985 1099.240 699.850 1101.240 ;
        RECT 4.400 1097.840 695.600 1099.240 ;
        RECT 0.985 1095.840 699.850 1097.840 ;
        RECT 4.400 1094.440 695.600 1095.840 ;
        RECT 0.985 1092.440 699.850 1094.440 ;
        RECT 4.400 1091.040 695.600 1092.440 ;
        RECT 0.985 1089.040 699.850 1091.040 ;
        RECT 4.400 1087.640 695.600 1089.040 ;
        RECT 0.985 1085.640 699.850 1087.640 ;
        RECT 4.400 1084.240 699.850 1085.640 ;
        RECT 0.985 1082.240 699.850 1084.240 ;
        RECT 0.985 1080.840 695.600 1082.240 ;
        RECT 0.985 1078.840 699.850 1080.840 ;
        RECT 4.400 1077.440 695.600 1078.840 ;
        RECT 0.985 1075.440 699.850 1077.440 ;
        RECT 4.400 1074.040 695.600 1075.440 ;
        RECT 0.985 1072.040 699.850 1074.040 ;
        RECT 4.400 1070.640 695.600 1072.040 ;
        RECT 0.985 1068.640 699.850 1070.640 ;
        RECT 4.400 1067.240 695.600 1068.640 ;
        RECT 0.985 1065.240 699.850 1067.240 ;
        RECT 4.400 1063.840 695.600 1065.240 ;
        RECT 0.985 1058.440 699.850 1063.840 ;
        RECT 4.400 1057.040 695.600 1058.440 ;
        RECT 0.985 1055.040 699.850 1057.040 ;
        RECT 4.400 1053.640 695.600 1055.040 ;
        RECT 0.985 1051.640 699.850 1053.640 ;
        RECT 4.400 1050.240 695.600 1051.640 ;
        RECT 0.985 1048.240 699.850 1050.240 ;
        RECT 4.400 1046.840 695.600 1048.240 ;
        RECT 0.985 1044.840 699.850 1046.840 ;
        RECT 4.400 1043.440 695.600 1044.840 ;
        RECT 0.985 1038.040 699.850 1043.440 ;
        RECT 4.400 1036.640 695.600 1038.040 ;
        RECT 0.985 1034.640 699.850 1036.640 ;
        RECT 4.400 1033.240 695.600 1034.640 ;
        RECT 0.985 1031.240 699.850 1033.240 ;
        RECT 4.400 1029.840 695.600 1031.240 ;
        RECT 0.985 1027.840 699.850 1029.840 ;
        RECT 4.400 1026.440 695.600 1027.840 ;
        RECT 0.985 1024.440 699.850 1026.440 ;
        RECT 4.400 1023.040 695.600 1024.440 ;
        RECT 0.985 1021.040 699.850 1023.040 ;
        RECT 4.400 1019.640 699.850 1021.040 ;
        RECT 0.985 1017.640 699.850 1019.640 ;
        RECT 0.985 1016.240 695.600 1017.640 ;
        RECT 0.985 1014.240 699.850 1016.240 ;
        RECT 4.400 1012.840 695.600 1014.240 ;
        RECT 0.985 1010.840 699.850 1012.840 ;
        RECT 4.400 1009.440 695.600 1010.840 ;
        RECT 0.985 1007.440 699.850 1009.440 ;
        RECT 4.400 1006.040 695.600 1007.440 ;
        RECT 0.985 1004.040 699.850 1006.040 ;
        RECT 4.400 1002.640 695.600 1004.040 ;
        RECT 0.985 1000.640 699.850 1002.640 ;
        RECT 4.400 999.240 699.850 1000.640 ;
        RECT 0.985 997.240 699.850 999.240 ;
        RECT 0.985 995.840 695.600 997.240 ;
        RECT 0.985 993.840 699.850 995.840 ;
        RECT 4.400 992.440 695.600 993.840 ;
        RECT 0.985 990.440 699.850 992.440 ;
        RECT 4.400 989.040 695.600 990.440 ;
        RECT 0.985 987.040 699.850 989.040 ;
        RECT 4.400 985.640 695.600 987.040 ;
        RECT 0.985 983.640 699.850 985.640 ;
        RECT 4.400 982.240 695.600 983.640 ;
        RECT 0.985 980.240 699.850 982.240 ;
        RECT 4.400 978.840 695.600 980.240 ;
        RECT 0.985 973.440 699.850 978.840 ;
        RECT 4.400 972.040 695.600 973.440 ;
        RECT 0.985 970.040 699.850 972.040 ;
        RECT 4.400 968.640 695.600 970.040 ;
        RECT 0.985 966.640 699.850 968.640 ;
        RECT 4.400 965.240 695.600 966.640 ;
        RECT 0.985 963.240 699.850 965.240 ;
        RECT 4.400 961.840 695.600 963.240 ;
        RECT 0.985 959.840 699.850 961.840 ;
        RECT 4.400 958.440 695.600 959.840 ;
        RECT 0.985 953.040 699.850 958.440 ;
        RECT 4.400 951.640 695.600 953.040 ;
        RECT 0.985 949.640 699.850 951.640 ;
        RECT 4.400 948.240 695.600 949.640 ;
        RECT 0.985 946.240 699.850 948.240 ;
        RECT 4.400 944.840 695.600 946.240 ;
        RECT 0.985 942.840 699.850 944.840 ;
        RECT 4.400 941.440 695.600 942.840 ;
        RECT 0.985 939.440 699.850 941.440 ;
        RECT 4.400 938.040 695.600 939.440 ;
        RECT 0.985 936.040 699.850 938.040 ;
        RECT 4.400 934.640 699.850 936.040 ;
        RECT 0.985 932.640 699.850 934.640 ;
        RECT 0.985 931.240 695.600 932.640 ;
        RECT 0.985 929.240 699.850 931.240 ;
        RECT 4.400 927.840 695.600 929.240 ;
        RECT 0.985 925.840 699.850 927.840 ;
        RECT 4.400 924.440 695.600 925.840 ;
        RECT 0.985 922.440 699.850 924.440 ;
        RECT 4.400 921.040 695.600 922.440 ;
        RECT 0.985 919.040 699.850 921.040 ;
        RECT 4.400 917.640 695.600 919.040 ;
        RECT 0.985 915.640 699.850 917.640 ;
        RECT 4.400 914.240 699.850 915.640 ;
        RECT 0.985 912.240 699.850 914.240 ;
        RECT 0.985 910.840 695.600 912.240 ;
        RECT 0.985 908.840 699.850 910.840 ;
        RECT 4.400 907.440 695.600 908.840 ;
        RECT 0.985 905.440 699.850 907.440 ;
        RECT 4.400 904.040 695.600 905.440 ;
        RECT 0.985 902.040 699.850 904.040 ;
        RECT 4.400 900.640 695.600 902.040 ;
        RECT 0.985 898.640 699.850 900.640 ;
        RECT 4.400 897.240 695.600 898.640 ;
        RECT 0.985 895.240 699.850 897.240 ;
        RECT 4.400 893.840 695.600 895.240 ;
        RECT 0.985 888.440 699.850 893.840 ;
        RECT 4.400 887.040 695.600 888.440 ;
        RECT 0.985 885.040 699.850 887.040 ;
        RECT 4.400 883.640 695.600 885.040 ;
        RECT 0.985 881.640 699.850 883.640 ;
        RECT 4.400 880.240 695.600 881.640 ;
        RECT 0.985 878.240 699.850 880.240 ;
        RECT 4.400 876.840 695.600 878.240 ;
        RECT 0.985 874.840 699.850 876.840 ;
        RECT 4.400 873.440 695.600 874.840 ;
        RECT 0.985 868.040 699.850 873.440 ;
        RECT 4.400 866.640 695.600 868.040 ;
        RECT 0.985 864.640 699.850 866.640 ;
        RECT 4.400 863.240 695.600 864.640 ;
        RECT 0.985 861.240 699.850 863.240 ;
        RECT 4.400 859.840 695.600 861.240 ;
        RECT 0.985 857.840 699.850 859.840 ;
        RECT 4.400 856.440 695.600 857.840 ;
        RECT 0.985 854.440 699.850 856.440 ;
        RECT 4.400 853.040 695.600 854.440 ;
        RECT 0.985 851.040 699.850 853.040 ;
        RECT 4.400 849.640 699.850 851.040 ;
        RECT 0.985 847.640 699.850 849.640 ;
        RECT 0.985 846.240 695.600 847.640 ;
        RECT 0.985 844.240 699.850 846.240 ;
        RECT 4.400 842.840 695.600 844.240 ;
        RECT 0.985 840.840 699.850 842.840 ;
        RECT 4.400 839.440 695.600 840.840 ;
        RECT 0.985 837.440 699.850 839.440 ;
        RECT 4.400 836.040 695.600 837.440 ;
        RECT 0.985 834.040 699.850 836.040 ;
        RECT 4.400 832.640 695.600 834.040 ;
        RECT 0.985 830.640 699.850 832.640 ;
        RECT 4.400 829.240 699.850 830.640 ;
        RECT 0.985 827.240 699.850 829.240 ;
        RECT 0.985 825.840 695.600 827.240 ;
        RECT 0.985 823.840 699.850 825.840 ;
        RECT 4.400 822.440 695.600 823.840 ;
        RECT 0.985 820.440 699.850 822.440 ;
        RECT 4.400 819.040 695.600 820.440 ;
        RECT 0.985 817.040 699.850 819.040 ;
        RECT 4.400 815.640 695.600 817.040 ;
        RECT 0.985 813.640 699.850 815.640 ;
        RECT 4.400 812.240 695.600 813.640 ;
        RECT 0.985 810.240 699.850 812.240 ;
        RECT 4.400 808.840 695.600 810.240 ;
        RECT 0.985 803.440 699.850 808.840 ;
        RECT 4.400 802.040 695.600 803.440 ;
        RECT 0.985 800.040 699.850 802.040 ;
        RECT 4.400 798.640 695.600 800.040 ;
        RECT 0.985 796.640 699.850 798.640 ;
        RECT 4.400 795.240 695.600 796.640 ;
        RECT 0.985 793.240 699.850 795.240 ;
        RECT 4.400 791.840 695.600 793.240 ;
        RECT 0.985 789.840 699.850 791.840 ;
        RECT 4.400 788.440 695.600 789.840 ;
        RECT 0.985 783.040 699.850 788.440 ;
        RECT 4.400 781.640 695.600 783.040 ;
        RECT 0.985 779.640 699.850 781.640 ;
        RECT 4.400 778.240 695.600 779.640 ;
        RECT 0.985 776.240 699.850 778.240 ;
        RECT 4.400 774.840 695.600 776.240 ;
        RECT 0.985 772.840 699.850 774.840 ;
        RECT 4.400 771.440 695.600 772.840 ;
        RECT 0.985 769.440 699.850 771.440 ;
        RECT 4.400 768.040 695.600 769.440 ;
        RECT 0.985 766.040 699.850 768.040 ;
        RECT 4.400 764.640 699.850 766.040 ;
        RECT 0.985 762.640 699.850 764.640 ;
        RECT 0.985 761.240 695.600 762.640 ;
        RECT 0.985 759.240 699.850 761.240 ;
        RECT 4.400 757.840 695.600 759.240 ;
        RECT 0.985 755.840 699.850 757.840 ;
        RECT 4.400 754.440 695.600 755.840 ;
        RECT 0.985 752.440 699.850 754.440 ;
        RECT 4.400 751.040 695.600 752.440 ;
        RECT 0.985 749.040 699.850 751.040 ;
        RECT 4.400 747.640 695.600 749.040 ;
        RECT 0.985 745.640 699.850 747.640 ;
        RECT 4.400 744.240 699.850 745.640 ;
        RECT 0.985 742.240 699.850 744.240 ;
        RECT 0.985 740.840 695.600 742.240 ;
        RECT 0.985 738.840 699.850 740.840 ;
        RECT 4.400 737.440 695.600 738.840 ;
        RECT 0.985 735.440 699.850 737.440 ;
        RECT 4.400 734.040 695.600 735.440 ;
        RECT 0.985 732.040 699.850 734.040 ;
        RECT 4.400 730.640 695.600 732.040 ;
        RECT 0.985 728.640 699.850 730.640 ;
        RECT 4.400 727.240 695.600 728.640 ;
        RECT 0.985 725.240 699.850 727.240 ;
        RECT 4.400 723.840 695.600 725.240 ;
        RECT 0.985 718.440 699.850 723.840 ;
        RECT 4.400 717.040 695.600 718.440 ;
        RECT 0.985 715.040 699.850 717.040 ;
        RECT 4.400 713.640 695.600 715.040 ;
        RECT 0.985 711.640 699.850 713.640 ;
        RECT 4.400 710.240 695.600 711.640 ;
        RECT 0.985 708.240 699.850 710.240 ;
        RECT 4.400 706.840 695.600 708.240 ;
        RECT 0.985 704.840 699.850 706.840 ;
        RECT 4.400 703.440 695.600 704.840 ;
        RECT 0.985 698.040 699.850 703.440 ;
        RECT 4.400 696.640 695.600 698.040 ;
        RECT 0.985 694.640 699.850 696.640 ;
        RECT 4.400 693.240 695.600 694.640 ;
        RECT 0.985 691.240 699.850 693.240 ;
        RECT 4.400 689.840 695.600 691.240 ;
        RECT 0.985 687.840 699.850 689.840 ;
        RECT 4.400 686.440 695.600 687.840 ;
        RECT 0.985 684.440 699.850 686.440 ;
        RECT 4.400 683.040 695.600 684.440 ;
        RECT 0.985 681.040 699.850 683.040 ;
        RECT 4.400 679.640 699.850 681.040 ;
        RECT 0.985 677.640 699.850 679.640 ;
        RECT 0.985 676.240 695.600 677.640 ;
        RECT 0.985 674.240 699.850 676.240 ;
        RECT 4.400 672.840 695.600 674.240 ;
        RECT 0.985 670.840 699.850 672.840 ;
        RECT 4.400 669.440 695.600 670.840 ;
        RECT 0.985 667.440 699.850 669.440 ;
        RECT 4.400 666.040 695.600 667.440 ;
        RECT 0.985 664.040 699.850 666.040 ;
        RECT 4.400 662.640 695.600 664.040 ;
        RECT 0.985 660.640 699.850 662.640 ;
        RECT 4.400 659.240 699.850 660.640 ;
        RECT 0.985 657.240 699.850 659.240 ;
        RECT 0.985 655.840 695.600 657.240 ;
        RECT 0.985 653.840 699.850 655.840 ;
        RECT 4.400 652.440 695.600 653.840 ;
        RECT 0.985 650.440 699.850 652.440 ;
        RECT 4.400 649.040 695.600 650.440 ;
        RECT 0.985 647.040 699.850 649.040 ;
        RECT 4.400 645.640 695.600 647.040 ;
        RECT 0.985 643.640 699.850 645.640 ;
        RECT 4.400 642.240 695.600 643.640 ;
        RECT 0.985 640.240 699.850 642.240 ;
        RECT 4.400 638.840 695.600 640.240 ;
        RECT 0.985 633.440 699.850 638.840 ;
        RECT 4.400 632.040 695.600 633.440 ;
        RECT 0.985 630.040 699.850 632.040 ;
        RECT 4.400 628.640 695.600 630.040 ;
        RECT 0.985 626.640 699.850 628.640 ;
        RECT 4.400 625.240 695.600 626.640 ;
        RECT 0.985 623.240 699.850 625.240 ;
        RECT 4.400 621.840 695.600 623.240 ;
        RECT 0.985 619.840 699.850 621.840 ;
        RECT 4.400 618.440 695.600 619.840 ;
        RECT 0.985 613.040 699.850 618.440 ;
        RECT 4.400 611.640 695.600 613.040 ;
        RECT 0.985 609.640 699.850 611.640 ;
        RECT 4.400 608.240 695.600 609.640 ;
        RECT 0.985 606.240 699.850 608.240 ;
        RECT 4.400 604.840 695.600 606.240 ;
        RECT 0.985 602.840 699.850 604.840 ;
        RECT 4.400 601.440 695.600 602.840 ;
        RECT 0.985 599.440 699.850 601.440 ;
        RECT 4.400 598.040 695.600 599.440 ;
        RECT 0.985 596.040 699.850 598.040 ;
        RECT 4.400 594.640 699.850 596.040 ;
        RECT 0.985 592.640 699.850 594.640 ;
        RECT 0.985 591.240 695.600 592.640 ;
        RECT 0.985 589.240 699.850 591.240 ;
        RECT 4.400 587.840 695.600 589.240 ;
        RECT 0.985 585.840 699.850 587.840 ;
        RECT 4.400 584.440 695.600 585.840 ;
        RECT 0.985 582.440 699.850 584.440 ;
        RECT 4.400 581.040 695.600 582.440 ;
        RECT 0.985 579.040 699.850 581.040 ;
        RECT 4.400 577.640 695.600 579.040 ;
        RECT 0.985 575.640 699.850 577.640 ;
        RECT 4.400 574.240 699.850 575.640 ;
        RECT 0.985 572.240 699.850 574.240 ;
        RECT 0.985 570.840 695.600 572.240 ;
        RECT 0.985 568.840 699.850 570.840 ;
        RECT 4.400 567.440 695.600 568.840 ;
        RECT 0.985 565.440 699.850 567.440 ;
        RECT 4.400 564.040 695.600 565.440 ;
        RECT 0.985 562.040 699.850 564.040 ;
        RECT 4.400 560.640 695.600 562.040 ;
        RECT 0.985 558.640 699.850 560.640 ;
        RECT 4.400 557.240 695.600 558.640 ;
        RECT 0.985 555.240 699.850 557.240 ;
        RECT 4.400 553.840 695.600 555.240 ;
        RECT 0.985 548.440 699.850 553.840 ;
        RECT 4.400 547.040 695.600 548.440 ;
        RECT 0.985 545.040 699.850 547.040 ;
        RECT 4.400 543.640 695.600 545.040 ;
        RECT 0.985 541.640 699.850 543.640 ;
        RECT 4.400 540.240 695.600 541.640 ;
        RECT 0.985 538.240 699.850 540.240 ;
        RECT 4.400 536.840 695.600 538.240 ;
        RECT 0.985 534.840 699.850 536.840 ;
        RECT 4.400 533.440 695.600 534.840 ;
        RECT 0.985 528.040 699.850 533.440 ;
        RECT 4.400 526.640 695.600 528.040 ;
        RECT 0.985 524.640 699.850 526.640 ;
        RECT 4.400 523.240 695.600 524.640 ;
        RECT 0.985 521.240 699.850 523.240 ;
        RECT 4.400 519.840 695.600 521.240 ;
        RECT 0.985 517.840 699.850 519.840 ;
        RECT 4.400 516.440 695.600 517.840 ;
        RECT 0.985 514.440 699.850 516.440 ;
        RECT 4.400 513.040 695.600 514.440 ;
        RECT 0.985 511.040 699.850 513.040 ;
        RECT 4.400 509.640 699.850 511.040 ;
        RECT 0.985 507.640 699.850 509.640 ;
        RECT 0.985 506.240 695.600 507.640 ;
        RECT 0.985 504.240 699.850 506.240 ;
        RECT 4.400 502.840 695.600 504.240 ;
        RECT 0.985 500.840 699.850 502.840 ;
        RECT 4.400 499.440 695.600 500.840 ;
        RECT 0.985 497.440 699.850 499.440 ;
        RECT 4.400 496.040 695.600 497.440 ;
        RECT 0.985 494.040 699.850 496.040 ;
        RECT 4.400 492.640 695.600 494.040 ;
        RECT 0.985 490.640 699.850 492.640 ;
        RECT 4.400 489.240 699.850 490.640 ;
        RECT 0.985 487.240 699.850 489.240 ;
        RECT 0.985 485.840 695.600 487.240 ;
        RECT 0.985 483.840 699.850 485.840 ;
        RECT 4.400 482.440 695.600 483.840 ;
        RECT 0.985 480.440 699.850 482.440 ;
        RECT 4.400 479.040 695.600 480.440 ;
        RECT 0.985 477.040 699.850 479.040 ;
        RECT 4.400 475.640 695.600 477.040 ;
        RECT 0.985 473.640 699.850 475.640 ;
        RECT 4.400 472.240 695.600 473.640 ;
        RECT 0.985 470.240 699.850 472.240 ;
        RECT 4.400 468.840 695.600 470.240 ;
        RECT 0.985 463.440 699.850 468.840 ;
        RECT 4.400 462.040 695.600 463.440 ;
        RECT 0.985 460.040 699.850 462.040 ;
        RECT 4.400 458.640 695.600 460.040 ;
        RECT 0.985 456.640 699.850 458.640 ;
        RECT 4.400 455.240 695.600 456.640 ;
        RECT 0.985 453.240 699.850 455.240 ;
        RECT 4.400 451.840 695.600 453.240 ;
        RECT 0.985 449.840 699.850 451.840 ;
        RECT 4.400 448.440 695.600 449.840 ;
        RECT 0.985 443.040 699.850 448.440 ;
        RECT 4.400 441.640 695.600 443.040 ;
        RECT 0.985 439.640 699.850 441.640 ;
        RECT 4.400 438.240 695.600 439.640 ;
        RECT 0.985 436.240 699.850 438.240 ;
        RECT 4.400 434.840 695.600 436.240 ;
        RECT 0.985 432.840 699.850 434.840 ;
        RECT 4.400 431.440 695.600 432.840 ;
        RECT 0.985 429.440 699.850 431.440 ;
        RECT 4.400 428.040 695.600 429.440 ;
        RECT 0.985 426.040 699.850 428.040 ;
        RECT 4.400 424.640 699.850 426.040 ;
        RECT 0.985 422.640 699.850 424.640 ;
        RECT 0.985 421.240 695.600 422.640 ;
        RECT 0.985 419.240 699.850 421.240 ;
        RECT 4.400 417.840 695.600 419.240 ;
        RECT 0.985 415.840 699.850 417.840 ;
        RECT 4.400 414.440 695.600 415.840 ;
        RECT 0.985 412.440 699.850 414.440 ;
        RECT 4.400 411.040 695.600 412.440 ;
        RECT 0.985 409.040 699.850 411.040 ;
        RECT 4.400 407.640 695.600 409.040 ;
        RECT 0.985 405.640 699.850 407.640 ;
        RECT 4.400 404.240 699.850 405.640 ;
        RECT 0.985 402.240 699.850 404.240 ;
        RECT 0.985 400.840 695.600 402.240 ;
        RECT 0.985 398.840 699.850 400.840 ;
        RECT 4.400 397.440 695.600 398.840 ;
        RECT 0.985 395.440 699.850 397.440 ;
        RECT 4.400 394.040 695.600 395.440 ;
        RECT 0.985 392.040 699.850 394.040 ;
        RECT 4.400 390.640 695.600 392.040 ;
        RECT 0.985 388.640 699.850 390.640 ;
        RECT 4.400 387.240 695.600 388.640 ;
        RECT 0.985 385.240 699.850 387.240 ;
        RECT 4.400 383.840 699.850 385.240 ;
        RECT 0.985 381.840 699.850 383.840 ;
        RECT 0.985 380.440 695.600 381.840 ;
        RECT 0.985 378.440 699.850 380.440 ;
        RECT 4.400 377.040 695.600 378.440 ;
        RECT 0.985 375.040 699.850 377.040 ;
        RECT 4.400 373.640 695.600 375.040 ;
        RECT 0.985 371.640 699.850 373.640 ;
        RECT 4.400 370.240 695.600 371.640 ;
        RECT 0.985 368.240 699.850 370.240 ;
        RECT 4.400 366.840 695.600 368.240 ;
        RECT 0.985 364.840 699.850 366.840 ;
        RECT 4.400 363.440 695.600 364.840 ;
        RECT 0.985 358.040 699.850 363.440 ;
        RECT 4.400 356.640 695.600 358.040 ;
        RECT 0.985 354.640 699.850 356.640 ;
        RECT 4.400 353.240 695.600 354.640 ;
        RECT 0.985 351.240 699.850 353.240 ;
        RECT 4.400 349.840 695.600 351.240 ;
        RECT 0.985 347.840 699.850 349.840 ;
        RECT 4.400 346.440 695.600 347.840 ;
        RECT 0.985 344.440 699.850 346.440 ;
        RECT 4.400 343.040 695.600 344.440 ;
        RECT 0.985 341.040 699.850 343.040 ;
        RECT 4.400 339.640 699.850 341.040 ;
        RECT 0.985 337.640 699.850 339.640 ;
        RECT 0.985 336.240 695.600 337.640 ;
        RECT 0.985 334.240 699.850 336.240 ;
        RECT 4.400 332.840 695.600 334.240 ;
        RECT 0.985 330.840 699.850 332.840 ;
        RECT 4.400 329.440 695.600 330.840 ;
        RECT 0.985 327.440 699.850 329.440 ;
        RECT 4.400 326.040 695.600 327.440 ;
        RECT 0.985 324.040 699.850 326.040 ;
        RECT 4.400 322.640 695.600 324.040 ;
        RECT 0.985 320.640 699.850 322.640 ;
        RECT 4.400 319.240 699.850 320.640 ;
        RECT 0.985 317.240 699.850 319.240 ;
        RECT 0.985 315.840 695.600 317.240 ;
        RECT 0.985 313.840 699.850 315.840 ;
        RECT 4.400 312.440 695.600 313.840 ;
        RECT 0.985 310.440 699.850 312.440 ;
        RECT 4.400 309.040 695.600 310.440 ;
        RECT 0.985 307.040 699.850 309.040 ;
        RECT 4.400 305.640 695.600 307.040 ;
        RECT 0.985 303.640 699.850 305.640 ;
        RECT 4.400 302.240 695.600 303.640 ;
        RECT 0.985 300.240 699.850 302.240 ;
        RECT 4.400 298.840 699.850 300.240 ;
        RECT 0.985 296.840 699.850 298.840 ;
        RECT 0.985 295.440 695.600 296.840 ;
        RECT 0.985 293.440 699.850 295.440 ;
        RECT 4.400 292.040 695.600 293.440 ;
        RECT 0.985 290.040 699.850 292.040 ;
        RECT 4.400 288.640 695.600 290.040 ;
        RECT 0.985 286.640 699.850 288.640 ;
        RECT 4.400 285.240 695.600 286.640 ;
        RECT 0.985 283.240 699.850 285.240 ;
        RECT 4.400 281.840 695.600 283.240 ;
        RECT 0.985 279.840 699.850 281.840 ;
        RECT 4.400 278.440 695.600 279.840 ;
        RECT 0.985 273.040 699.850 278.440 ;
        RECT 4.400 271.640 695.600 273.040 ;
        RECT 0.985 269.640 699.850 271.640 ;
        RECT 4.400 268.240 695.600 269.640 ;
        RECT 0.985 266.240 699.850 268.240 ;
        RECT 4.400 264.840 695.600 266.240 ;
        RECT 0.985 262.840 699.850 264.840 ;
        RECT 4.400 261.440 695.600 262.840 ;
        RECT 0.985 259.440 699.850 261.440 ;
        RECT 4.400 258.040 695.600 259.440 ;
        RECT 0.985 256.040 699.850 258.040 ;
        RECT 4.400 254.640 699.850 256.040 ;
        RECT 0.985 252.640 699.850 254.640 ;
        RECT 0.985 251.240 695.600 252.640 ;
        RECT 0.985 249.240 699.850 251.240 ;
        RECT 4.400 247.840 695.600 249.240 ;
        RECT 0.985 245.840 699.850 247.840 ;
        RECT 4.400 244.440 695.600 245.840 ;
        RECT 0.985 242.440 699.850 244.440 ;
        RECT 4.400 241.040 695.600 242.440 ;
        RECT 0.985 239.040 699.850 241.040 ;
        RECT 4.400 237.640 695.600 239.040 ;
        RECT 0.985 235.640 699.850 237.640 ;
        RECT 4.400 234.240 699.850 235.640 ;
        RECT 0.985 232.240 699.850 234.240 ;
        RECT 0.985 230.840 695.600 232.240 ;
        RECT 0.985 228.840 699.850 230.840 ;
        RECT 4.400 227.440 695.600 228.840 ;
        RECT 0.985 225.440 699.850 227.440 ;
        RECT 4.400 224.040 695.600 225.440 ;
        RECT 0.985 222.040 699.850 224.040 ;
        RECT 4.400 220.640 695.600 222.040 ;
        RECT 0.985 218.640 699.850 220.640 ;
        RECT 4.400 217.240 695.600 218.640 ;
        RECT 0.985 215.240 699.850 217.240 ;
        RECT 4.400 213.840 699.850 215.240 ;
        RECT 0.985 211.840 699.850 213.840 ;
        RECT 0.985 210.440 695.600 211.840 ;
        RECT 0.985 208.440 699.850 210.440 ;
        RECT 4.400 207.040 695.600 208.440 ;
        RECT 0.985 205.040 699.850 207.040 ;
        RECT 4.400 203.640 695.600 205.040 ;
        RECT 0.985 201.640 699.850 203.640 ;
        RECT 4.400 200.240 695.600 201.640 ;
        RECT 0.985 198.240 699.850 200.240 ;
        RECT 4.400 196.840 695.600 198.240 ;
        RECT 0.985 194.840 699.850 196.840 ;
        RECT 4.400 193.440 695.600 194.840 ;
        RECT 0.985 188.040 699.850 193.440 ;
        RECT 4.400 186.640 695.600 188.040 ;
        RECT 0.985 184.640 699.850 186.640 ;
        RECT 4.400 183.240 695.600 184.640 ;
        RECT 0.985 181.240 699.850 183.240 ;
        RECT 4.400 179.840 695.600 181.240 ;
        RECT 0.985 177.840 699.850 179.840 ;
        RECT 4.400 176.440 695.600 177.840 ;
        RECT 0.985 174.440 699.850 176.440 ;
        RECT 4.400 173.040 695.600 174.440 ;
        RECT 0.985 171.040 699.850 173.040 ;
        RECT 4.400 169.640 699.850 171.040 ;
        RECT 0.985 167.640 699.850 169.640 ;
        RECT 0.985 166.240 695.600 167.640 ;
        RECT 0.985 164.240 699.850 166.240 ;
        RECT 4.400 162.840 695.600 164.240 ;
        RECT 0.985 160.840 699.850 162.840 ;
        RECT 4.400 159.440 695.600 160.840 ;
        RECT 0.985 157.440 699.850 159.440 ;
        RECT 4.400 156.040 695.600 157.440 ;
        RECT 0.985 154.040 699.850 156.040 ;
        RECT 4.400 152.640 695.600 154.040 ;
        RECT 0.985 150.640 699.850 152.640 ;
        RECT 4.400 149.240 699.850 150.640 ;
        RECT 0.985 147.240 699.850 149.240 ;
        RECT 0.985 145.840 695.600 147.240 ;
        RECT 0.985 143.840 699.850 145.840 ;
        RECT 4.400 142.440 695.600 143.840 ;
        RECT 0.985 140.440 699.850 142.440 ;
        RECT 4.400 139.040 695.600 140.440 ;
        RECT 0.985 137.040 699.850 139.040 ;
        RECT 4.400 135.640 695.600 137.040 ;
        RECT 0.985 133.640 699.850 135.640 ;
        RECT 4.400 132.240 695.600 133.640 ;
        RECT 0.985 130.240 699.850 132.240 ;
        RECT 4.400 128.840 699.850 130.240 ;
        RECT 0.985 126.840 699.850 128.840 ;
        RECT 0.985 125.440 695.600 126.840 ;
        RECT 0.985 123.440 699.850 125.440 ;
        RECT 4.400 122.040 695.600 123.440 ;
        RECT 0.985 120.040 699.850 122.040 ;
        RECT 4.400 118.640 695.600 120.040 ;
        RECT 0.985 116.640 699.850 118.640 ;
        RECT 4.400 115.240 695.600 116.640 ;
        RECT 0.985 113.240 699.850 115.240 ;
        RECT 4.400 111.840 695.600 113.240 ;
        RECT 0.985 109.840 699.850 111.840 ;
        RECT 4.400 108.440 695.600 109.840 ;
        RECT 0.985 103.040 699.850 108.440 ;
        RECT 4.400 101.640 695.600 103.040 ;
        RECT 0.985 99.640 699.850 101.640 ;
        RECT 4.400 98.240 695.600 99.640 ;
        RECT 0.985 96.240 699.850 98.240 ;
        RECT 4.400 94.840 695.600 96.240 ;
        RECT 0.985 92.840 699.850 94.840 ;
        RECT 4.400 91.440 695.600 92.840 ;
        RECT 0.985 89.440 699.850 91.440 ;
        RECT 4.400 88.040 695.600 89.440 ;
        RECT 0.985 86.040 699.850 88.040 ;
        RECT 4.400 84.640 699.850 86.040 ;
        RECT 0.985 82.640 699.850 84.640 ;
        RECT 0.985 81.240 695.600 82.640 ;
        RECT 0.985 79.240 699.850 81.240 ;
        RECT 4.400 77.840 695.600 79.240 ;
        RECT 0.985 75.840 699.850 77.840 ;
        RECT 4.400 74.440 695.600 75.840 ;
        RECT 0.985 72.440 699.850 74.440 ;
        RECT 4.400 71.040 695.600 72.440 ;
        RECT 0.985 69.040 699.850 71.040 ;
        RECT 4.400 67.640 695.600 69.040 ;
        RECT 0.985 65.640 699.850 67.640 ;
        RECT 4.400 64.240 699.850 65.640 ;
        RECT 0.985 62.240 699.850 64.240 ;
        RECT 0.985 60.840 695.600 62.240 ;
        RECT 0.985 58.840 699.850 60.840 ;
        RECT 4.400 57.440 695.600 58.840 ;
        RECT 0.985 55.440 699.850 57.440 ;
        RECT 4.400 54.040 695.600 55.440 ;
        RECT 0.985 52.040 699.850 54.040 ;
        RECT 4.400 50.640 695.600 52.040 ;
        RECT 0.985 48.640 699.850 50.640 ;
        RECT 4.400 47.240 695.600 48.640 ;
        RECT 0.985 45.240 699.850 47.240 ;
        RECT 4.400 43.840 699.850 45.240 ;
        RECT 0.985 41.840 699.850 43.840 ;
        RECT 0.985 40.440 695.600 41.840 ;
        RECT 0.985 38.440 699.850 40.440 ;
        RECT 4.400 37.040 695.600 38.440 ;
        RECT 0.985 35.040 699.850 37.040 ;
        RECT 4.400 33.640 695.600 35.040 ;
        RECT 0.985 31.640 699.850 33.640 ;
        RECT 4.400 30.240 695.600 31.640 ;
        RECT 0.985 28.240 699.850 30.240 ;
        RECT 4.400 26.840 695.600 28.240 ;
        RECT 0.985 24.840 699.850 26.840 ;
        RECT 4.400 23.440 695.600 24.840 ;
        RECT 0.985 18.040 699.850 23.440 ;
        RECT 4.400 16.640 695.600 18.040 ;
        RECT 0.985 14.640 699.850 16.640 ;
        RECT 4.400 13.240 695.600 14.640 ;
        RECT 0.985 11.240 699.850 13.240 ;
        RECT 4.400 9.840 695.600 11.240 ;
        RECT 0.985 7.840 699.850 9.840 ;
        RECT 4.400 6.440 695.600 7.840 ;
        RECT 0.985 4.440 699.850 6.440 ;
        RECT 4.400 3.575 695.600 4.440 ;
      LAYER met4 ;
        RECT 2.135 10.240 20.640 2186.025 ;
        RECT 23.040 10.240 97.440 2186.025 ;
        RECT 99.840 10.240 174.240 2186.025 ;
        RECT 176.640 10.240 251.040 2186.025 ;
        RECT 253.440 10.240 327.840 2186.025 ;
        RECT 330.240 10.240 404.640 2186.025 ;
        RECT 407.040 10.240 481.440 2186.025 ;
        RECT 483.840 10.240 558.240 2186.025 ;
        RECT 560.640 10.240 635.040 2186.025 ;
        RECT 637.440 10.240 699.825 2186.025 ;
        RECT 2.135 8.335 699.825 10.240 ;
  END
END peripherals
END LIBRARY

