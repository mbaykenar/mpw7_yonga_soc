magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 5 13 731 203
rect 26 -24 70 13
<< ndiff >>
rect 31 39 705 177
<< pdiff >>
rect 31 305 705 505
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel metal1 s 35 -20 67 10 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 29 523 67 555 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel nwell s 20 522 77 553 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel pwell s 26 -24 70 10 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 fill_8
rlabel metal1 s 0 -48 736 48 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3952840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3950588
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
