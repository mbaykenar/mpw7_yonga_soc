magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 183
rect 29 -17 63 21
<< scnmos >>
rect 79 47 1025 157
<< scpmoshvt >>
rect 79 323 1025 497
<< ndiff >>
rect 27 112 79 157
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 1025 112 1077 157
rect 1025 78 1035 112
rect 1069 78 1077 112
rect 1025 47 1077 78
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 383 79 451
rect 27 349 35 383
rect 69 349 79 383
rect 27 323 79 349
rect 1025 485 1077 497
rect 1025 451 1035 485
rect 1069 451 1077 485
rect 1025 383 1077 451
rect 1025 349 1035 383
rect 1069 349 1077 383
rect 1025 323 1077 349
<< ndiffc >>
rect 35 78 69 112
rect 1035 78 1069 112
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 1035 451 1069 485
rect 1035 349 1069 383
<< poly >>
rect 79 497 1025 523
rect 79 297 1025 323
rect 79 275 529 297
rect 79 241 95 275
rect 129 241 223 275
rect 257 241 351 275
rect 385 241 479 275
rect 513 241 529 275
rect 79 225 529 241
rect 571 239 1025 255
rect 571 205 587 239
rect 621 205 715 239
rect 749 205 843 239
rect 877 205 971 239
rect 1005 205 1025 239
rect 571 183 1025 205
rect 79 157 1025 183
rect 79 21 1025 47
<< polycont >>
rect 95 241 129 275
rect 223 241 257 275
rect 351 241 385 275
rect 479 241 513 275
rect 587 205 621 239
rect 715 205 749 239
rect 843 205 877 239
rect 971 205 1005 239
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 485 1086 493
rect 17 459 35 485
rect 69 459 1035 485
rect 1069 459 1086 485
rect 17 425 29 459
rect 69 451 121 459
rect 63 425 121 451
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 397 459
rect 431 425 489 459
rect 523 425 581 459
rect 615 425 673 459
rect 707 425 765 459
rect 799 425 857 459
rect 891 425 949 459
rect 983 451 1035 459
rect 983 425 1041 451
rect 1075 425 1086 459
rect 17 383 1086 425
rect 17 349 35 383
rect 69 349 1035 383
rect 1069 349 1086 383
rect 17 309 1086 349
rect 17 241 95 275
rect 129 241 223 275
rect 257 241 351 275
rect 385 241 479 275
rect 513 241 533 275
rect 17 171 533 241
rect 567 239 1086 309
rect 567 205 587 239
rect 621 205 715 239
rect 749 205 843 239
rect 877 205 971 239
rect 1005 205 1086 239
rect 17 112 1086 171
rect 17 78 35 112
rect 69 78 1035 112
rect 1069 78 1086 112
rect 17 17 1086 78
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 451 35 459
rect 35 451 63 459
rect 29 425 63 451
rect 121 425 155 459
rect 213 425 247 459
rect 305 425 339 459
rect 397 425 431 459
rect 489 425 523 459
rect 581 425 615 459
rect 673 425 707 459
rect 765 425 799 459
rect 857 425 891 459
rect 949 425 983 459
rect 1041 451 1069 459
rect 1069 451 1075 459
rect 1041 425 1075 451
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 14 459 1090 468
rect 14 428 29 459
rect 17 425 29 428
rect 63 425 121 459
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 397 459
rect 431 425 489 459
rect 523 425 581 459
rect 615 425 673 459
rect 707 425 765 459
rect 799 425 857 459
rect 891 425 949 459
rect 983 425 1041 459
rect 1075 428 1090 459
rect 1075 425 1087 428
rect 17 416 1087 425
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 33 429 68 460 0 FreeSans 200 0 0 0 KAPWR
port 1 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 lpflow_decapkapwr_12
rlabel metal1 s 17 416 1087 428 1 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 1090 468 1 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1104 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 2344016
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2338900
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 27.600 0.000 
<< end >>
