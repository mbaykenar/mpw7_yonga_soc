magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 821 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 175 47 205 177
rect 247 47 277 177
rect 435 47 465 177
rect 531 47 561 177
rect 624 47 654 177
rect 708 47 738 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 435 297 465 497
rect 531 297 561 497
rect 624 297 654 497
rect 708 297 738 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 105 175 177
rect 109 71 119 105
rect 153 71 175 105
rect 109 47 175 71
rect 205 47 247 177
rect 277 101 329 177
rect 277 67 287 101
rect 321 67 329 101
rect 277 47 329 67
rect 383 101 435 177
rect 383 67 391 101
rect 425 67 435 101
rect 383 47 435 67
rect 465 47 531 177
rect 561 97 624 177
rect 561 63 571 97
rect 605 63 624 97
rect 561 47 624 63
rect 654 101 708 177
rect 654 67 664 101
rect 698 67 708 101
rect 654 47 708 67
rect 738 169 795 177
rect 738 135 749 169
rect 783 135 795 169
rect 738 101 795 135
rect 738 67 749 101
rect 783 67 795 101
rect 738 47 795 67
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 347 79 443
rect 27 313 35 347
rect 69 313 79 347
rect 27 297 79 313
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 409 247 497
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 485 329 497
rect 277 451 287 485
rect 321 451 329 485
rect 277 297 329 451
rect 383 477 435 497
rect 383 443 391 477
rect 425 443 435 477
rect 383 297 435 443
rect 465 477 531 497
rect 465 443 480 477
rect 514 443 531 477
rect 465 407 531 443
rect 465 373 480 407
rect 514 373 531 407
rect 465 297 531 373
rect 561 477 624 497
rect 561 443 580 477
rect 614 443 624 477
rect 561 409 624 443
rect 561 375 580 409
rect 614 375 624 409
rect 561 297 624 375
rect 654 477 708 497
rect 654 443 664 477
rect 698 443 708 477
rect 654 409 708 443
rect 654 375 664 409
rect 698 375 708 409
rect 654 297 708 375
rect 738 477 795 497
rect 738 443 749 477
rect 783 443 795 477
rect 738 409 795 443
rect 738 375 749 409
rect 783 375 795 409
rect 738 341 795 375
rect 738 307 749 341
rect 783 307 795 341
rect 738 297 795 307
<< ndiffc >>
rect 35 95 69 129
rect 119 71 153 105
rect 287 67 321 101
rect 391 67 425 101
rect 571 63 605 97
rect 664 67 698 101
rect 749 135 783 169
rect 749 67 783 101
<< pdiffc >>
rect 35 443 69 477
rect 35 313 69 347
rect 119 443 153 477
rect 119 375 153 409
rect 203 375 237 409
rect 287 451 321 485
rect 391 443 425 477
rect 480 443 514 477
rect 480 373 514 407
rect 580 443 614 477
rect 580 375 614 409
rect 664 443 698 477
rect 664 375 698 409
rect 749 443 783 477
rect 749 375 783 409
rect 749 307 783 341
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 435 497 465 523
rect 531 497 561 523
rect 624 497 654 523
rect 708 497 738 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 435 265 465 297
rect 531 265 561 297
rect 624 265 654 297
rect 708 265 738 297
rect 28 249 109 265
rect 28 215 38 249
rect 72 215 109 249
rect 28 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 79 177 109 199
rect 175 177 205 199
rect 247 249 305 265
rect 247 215 261 249
rect 295 215 305 249
rect 247 199 305 215
rect 400 249 465 265
rect 400 215 410 249
rect 444 215 465 249
rect 400 199 465 215
rect 507 249 561 265
rect 507 215 517 249
rect 551 215 561 249
rect 507 199 561 215
rect 603 249 738 265
rect 603 215 613 249
rect 647 215 738 249
rect 603 199 738 215
rect 247 177 277 199
rect 435 177 465 199
rect 531 177 561 199
rect 624 177 654 199
rect 708 177 738 199
rect 79 21 109 47
rect 175 21 205 47
rect 247 21 277 47
rect 435 21 465 47
rect 531 21 561 47
rect 624 21 654 47
rect 708 21 738 47
<< polycont >>
rect 38 215 72 249
rect 161 215 195 249
rect 261 215 295 249
rect 410 215 444 249
rect 517 215 551 249
rect 613 215 647 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 35 477 69 493
rect 35 347 69 443
rect 103 485 337 493
rect 103 477 287 485
rect 103 443 119 477
rect 153 459 287 477
rect 153 443 169 459
rect 271 451 287 459
rect 321 451 337 485
rect 375 477 446 527
rect 375 443 391 477
rect 425 443 446 477
rect 480 477 530 493
rect 514 443 530 477
rect 103 409 169 443
rect 103 375 119 409
rect 153 375 169 409
rect 103 359 169 375
rect 203 409 249 425
rect 237 407 249 409
rect 480 407 530 443
rect 237 375 480 407
rect 203 373 480 375
rect 514 373 530 407
rect 564 477 630 527
rect 564 443 580 477
rect 614 443 630 477
rect 564 409 630 443
rect 564 375 580 409
rect 614 375 630 409
rect 664 477 715 493
rect 698 443 715 477
rect 664 409 715 443
rect 698 375 715 409
rect 203 359 530 373
rect 664 359 715 375
rect 69 313 647 325
rect 35 291 647 313
rect 17 249 88 257
rect 17 215 38 249
rect 72 215 88 249
rect 122 249 211 255
rect 122 215 161 249
rect 195 215 211 249
rect 245 249 340 255
rect 245 215 261 249
rect 295 215 340 249
rect 35 147 248 181
rect 35 129 69 147
rect 35 51 69 95
rect 103 105 169 113
rect 103 71 119 105
rect 153 71 169 105
rect 103 17 169 71
rect 214 101 248 147
rect 284 135 340 215
rect 394 249 460 255
rect 394 215 410 249
rect 444 215 460 249
rect 494 249 567 255
rect 494 215 517 249
rect 551 215 567 249
rect 613 249 647 291
rect 394 135 451 215
rect 613 181 647 215
rect 487 147 647 181
rect 487 101 521 147
rect 681 133 715 359
rect 749 477 783 527
rect 749 409 783 443
rect 749 341 783 375
rect 749 289 783 307
rect 678 117 715 133
rect 214 67 287 101
rect 321 67 391 101
rect 425 67 521 101
rect 214 51 521 67
rect 555 97 621 113
rect 555 63 571 97
rect 605 63 621 97
rect 555 17 621 63
rect 664 101 715 117
rect 698 67 715 101
rect 664 51 715 67
rect 749 169 783 196
rect 749 101 783 135
rect 749 17 783 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 678 85 712 119 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 306 153 340 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 402 153 436 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 678 425 712 459 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 494 221 528 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 122 -17 156 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel locali s 122 527 156 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a221o_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3579030
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3571354
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 20.700 13.600 
<< end >>
