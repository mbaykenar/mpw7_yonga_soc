magic
tech sky130B
magscale 1 2
timestamp 1662725136
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 484394 700680 484400 700732
rect 484452 700720 484458 700732
rect 543458 700720 543464 700732
rect 484452 700692 543464 700720
rect 484452 700680 484458 700692
rect 543458 700680 543464 700692
rect 543516 700680 543522 700732
rect 332502 700612 332508 700664
rect 332560 700652 332566 700664
rect 398190 700652 398196 700664
rect 332560 700624 398196 700652
rect 332560 700612 332566 700624
rect 398190 700612 398196 700624
rect 398248 700612 398254 700664
rect 402882 700612 402888 700664
rect 402940 700652 402946 700664
rect 527174 700652 527180 700664
rect 402940 700624 527180 700652
rect 402940 700612 402946 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 283834 700544 283840 700596
rect 283892 700584 283898 700596
rect 399478 700584 399484 700596
rect 283892 700556 399484 700584
rect 283892 700544 283898 700556
rect 399478 700544 399484 700556
rect 399536 700544 399542 700596
rect 404998 700544 405004 700596
rect 405056 700584 405062 700596
rect 559650 700584 559656 700596
rect 405056 700556 559656 700584
rect 405056 700544 405062 700556
rect 559650 700544 559656 700556
rect 559708 700544 559714 700596
rect 364978 700476 364984 700528
rect 365036 700516 365042 700528
rect 551370 700516 551376 700528
rect 365036 700488 551376 700516
rect 365036 700476 365042 700488
rect 551370 700476 551376 700488
rect 551428 700476 551434 700528
rect 218974 700408 218980 700460
rect 219032 700448 219038 700460
rect 342990 700448 342996 700460
rect 219032 700420 342996 700448
rect 219032 700408 219038 700420
rect 342990 700408 342996 700420
rect 343048 700408 343054 700460
rect 348786 700408 348792 700460
rect 348844 700448 348850 700460
rect 565998 700448 566004 700460
rect 348844 700420 566004 700448
rect 348844 700408 348850 700420
rect 565998 700408 566004 700420
rect 566056 700408 566062 700460
rect 300118 700340 300124 700392
rect 300176 700380 300182 700392
rect 551462 700380 551468 700392
rect 300176 700352 551468 700380
rect 300176 700340 300182 700352
rect 551462 700340 551468 700352
rect 551520 700340 551526 700392
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 566182 700312 566188 700324
rect 267700 700284 566188 700312
rect 267700 700272 267706 700284
rect 566182 700272 566188 700284
rect 566240 700272 566246 700324
rect 105446 698912 105452 698964
rect 105504 698952 105510 698964
rect 399386 698952 399392 698964
rect 105504 698924 399392 698952
rect 105504 698912 105510 698924
rect 399386 698912 399392 698924
rect 399444 698912 399450 698964
rect 429838 698912 429844 698964
rect 429896 698952 429902 698964
rect 550266 698952 550272 698964
rect 429896 698924 550272 698952
rect 429896 698912 429902 698924
rect 550266 698912 550272 698924
rect 550324 698912 550330 698964
rect 137830 697552 137836 697604
rect 137888 697592 137894 697604
rect 389910 697592 389916 697604
rect 137888 697564 389916 697592
rect 137888 697552 137894 697564
rect 389910 697552 389916 697564
rect 389968 697552 389974 697604
rect 413646 697552 413652 697604
rect 413704 697592 413710 697604
rect 552198 697592 552204 697604
rect 413704 697564 552204 697592
rect 413704 697552 413710 697564
rect 552198 697552 552204 697564
rect 552256 697552 552262 697604
rect 154114 696192 154120 696244
rect 154172 696232 154178 696244
rect 552842 696232 552848 696244
rect 154172 696204 552848 696232
rect 154172 696192 154178 696204
rect 552842 696192 552848 696204
rect 552900 696192 552906 696244
rect 201494 694764 201500 694816
rect 201552 694804 201558 694816
rect 498194 694804 498200 694816
rect 201552 694776 498200 694804
rect 201552 694764 201558 694776
rect 498194 694764 498200 694776
rect 498252 694764 498258 694816
rect 88334 693404 88340 693456
rect 88392 693444 88398 693456
rect 551094 693444 551100 693456
rect 88392 693416 551100 693444
rect 88392 693404 88398 693416
rect 551094 693404 551100 693416
rect 551152 693404 551158 693456
rect 6914 692044 6920 692096
rect 6972 692084 6978 692096
rect 550082 692084 550088 692096
rect 6972 692056 550088 692084
rect 6972 692044 6978 692056
rect 550082 692044 550088 692056
rect 550140 692044 550146 692096
rect 71774 690616 71780 690668
rect 71832 690656 71838 690668
rect 383010 690656 383016 690668
rect 71832 690628 383016 690656
rect 71832 690616 71838 690628
rect 383010 690616 383016 690628
rect 383068 690616 383074 690668
rect 234614 687964 234620 688016
rect 234672 688004 234678 688016
rect 538214 688004 538220 688016
rect 234672 687976 538220 688004
rect 234672 687964 234678 687976
rect 538214 687964 538220 687976
rect 538272 687964 538278 688016
rect 40034 687896 40040 687948
rect 40092 687936 40098 687948
rect 373626 687936 373632 687948
rect 40092 687908 373632 687936
rect 40092 687896 40098 687908
rect 373626 687896 373632 687908
rect 373684 687896 373690 687948
rect 462314 687896 462320 687948
rect 462372 687936 462378 687948
rect 550634 687936 550640 687948
rect 462372 687908 550640 687936
rect 462372 687896 462378 687908
rect 550634 687896 550640 687908
rect 550692 687896 550698 687948
rect 405090 687284 405096 687336
rect 405148 687324 405154 687336
rect 457346 687324 457352 687336
rect 405148 687296 457352 687324
rect 405148 687284 405154 687296
rect 457346 687284 457352 687296
rect 457404 687284 457410 687336
rect 399754 687216 399760 687268
rect 399812 687256 399818 687268
rect 554866 687256 554872 687268
rect 399812 687228 554872 687256
rect 399812 687216 399818 687228
rect 554866 687216 554872 687228
rect 554924 687216 554930 687268
rect 367738 686060 367744 686112
rect 367796 686100 367802 686112
rect 476574 686100 476580 686112
rect 367796 686072 476580 686100
rect 367796 686060 367802 686072
rect 476574 686060 476580 686072
rect 476632 686060 476638 686112
rect 407758 685992 407764 686044
rect 407816 686032 407822 686044
rect 554958 686032 554964 686044
rect 407816 686004 554964 686032
rect 407816 685992 407822 686004
rect 554958 685992 554964 686004
rect 555016 685992 555022 686044
rect 378778 685924 378784 685976
rect 378836 685964 378842 685976
rect 528830 685964 528836 685976
rect 378836 685936 528836 685964
rect 378836 685924 378842 685936
rect 528830 685924 528836 685936
rect 528888 685924 528894 685976
rect 405182 685856 405188 685908
rect 405240 685896 405246 685908
rect 580902 685896 580908 685908
rect 405240 685868 580908 685896
rect 405240 685856 405246 685868
rect 580902 685856 580908 685868
rect 580960 685856 580966 685908
rect 409138 685312 409144 685364
rect 409196 685352 409202 685364
rect 470870 685352 470876 685364
rect 409196 685324 470876 685352
rect 409196 685312 409202 685324
rect 470870 685312 470876 685324
rect 470928 685312 470934 685364
rect 409046 685244 409052 685296
rect 409104 685284 409110 685296
rect 454218 685284 454224 685296
rect 409104 685256 454224 685284
rect 409104 685244 409110 685256
rect 454218 685244 454224 685256
rect 454276 685244 454282 685296
rect 408402 685176 408408 685228
rect 408460 685216 408466 685228
rect 436094 685216 436100 685228
rect 408460 685188 436100 685216
rect 408460 685176 408466 685188
rect 436094 685176 436100 685188
rect 436152 685176 436158 685228
rect 409690 685108 409696 685160
rect 409748 685148 409754 685160
rect 450262 685148 450268 685160
rect 409748 685120 450268 685148
rect 409748 685108 409754 685120
rect 450262 685108 450268 685120
rect 450320 685108 450326 685160
rect 402422 685040 402428 685092
rect 402480 685080 402486 685092
rect 490006 685080 490012 685092
rect 402480 685052 490012 685080
rect 402480 685040 402486 685052
rect 490006 685040 490012 685052
rect 490064 685040 490070 685092
rect 510522 685040 510528 685092
rect 510580 685080 510586 685092
rect 580994 685080 581000 685092
rect 510580 685052 581000 685080
rect 510580 685040 510586 685052
rect 580994 685040 581000 685052
rect 581052 685040 581058 685092
rect 407942 684972 407948 685024
rect 408000 685012 408006 685024
rect 456886 685012 456892 685024
rect 408000 684984 456892 685012
rect 408000 684972 408006 684984
rect 456886 684972 456892 684984
rect 456944 684972 456950 685024
rect 472802 684972 472808 685024
rect 472860 685012 472866 685024
rect 582374 685012 582380 685024
rect 472860 684984 582380 685012
rect 472860 684972 472866 684984
rect 582374 684972 582380 684984
rect 582432 684972 582438 685024
rect 409230 684904 409236 684956
rect 409288 684944 409294 684956
rect 523034 684944 523040 684956
rect 409288 684916 523040 684944
rect 409288 684904 409294 684916
rect 523034 684904 523040 684916
rect 523092 684904 523098 684956
rect 467006 684836 467012 684888
rect 467064 684876 467070 684888
rect 582466 684876 582472 684888
rect 467064 684848 582472 684876
rect 467064 684836 467070 684848
rect 582466 684836 582472 684848
rect 582524 684836 582530 684888
rect 398742 684768 398748 684820
rect 398800 684808 398806 684820
rect 521838 684808 521844 684820
rect 398800 684780 521844 684808
rect 398800 684768 398806 684780
rect 521838 684768 521844 684780
rect 521896 684768 521902 684820
rect 409506 684700 409512 684752
rect 409564 684740 409570 684752
rect 535454 684740 535460 684752
rect 409564 684712 535460 684740
rect 409564 684700 409570 684712
rect 535454 684700 535460 684712
rect 535512 684700 535518 684752
rect 396810 684632 396816 684684
rect 396868 684672 396874 684684
rect 539134 684672 539140 684684
rect 396868 684644 539140 684672
rect 396868 684632 396874 684644
rect 539134 684632 539140 684644
rect 539192 684632 539198 684684
rect 435450 684564 435456 684616
rect 435508 684604 435514 684616
rect 576854 684604 576860 684616
rect 435508 684576 576860 684604
rect 435508 684564 435514 684576
rect 576854 684564 576860 684576
rect 576912 684564 576918 684616
rect 408034 684496 408040 684548
rect 408092 684536 408098 684548
rect 555142 684536 555148 684548
rect 408092 684508 555148 684536
rect 408092 684496 408098 684508
rect 555142 684496 555148 684508
rect 555200 684496 555206 684548
rect 393958 684088 393964 684140
rect 394016 684128 394022 684140
rect 470686 684128 470692 684140
rect 394016 684100 470692 684128
rect 394016 684088 394022 684100
rect 470686 684088 470692 684100
rect 470744 684088 470750 684140
rect 409782 684020 409788 684072
rect 409840 684060 409846 684072
rect 449894 684060 449900 684072
rect 409840 684032 449900 684060
rect 409840 684020 409846 684032
rect 449894 684020 449900 684032
rect 449952 684020 449958 684072
rect 399846 683952 399852 684004
rect 399904 683992 399910 684004
rect 468386 683992 468392 684004
rect 399904 683964 468392 683992
rect 399904 683952 399910 683964
rect 468386 683952 468392 683964
rect 468444 683952 468450 684004
rect 401502 683884 401508 683936
rect 401560 683924 401566 683936
rect 476114 683924 476120 683936
rect 401560 683896 476120 683924
rect 401560 683884 401566 683896
rect 476114 683884 476120 683896
rect 476172 683884 476178 683936
rect 409322 683816 409328 683868
rect 409380 683856 409386 683868
rect 497274 683856 497280 683868
rect 409380 683828 497280 683856
rect 409380 683816 409386 683828
rect 497274 683816 497280 683828
rect 497332 683816 497338 683868
rect 393222 683748 393228 683800
rect 393280 683788 393286 683800
rect 499850 683788 499856 683800
rect 393280 683760 499856 683788
rect 393280 683748 393286 683760
rect 499850 683748 499856 683760
rect 499908 683748 499914 683800
rect 524874 683748 524880 683800
rect 524932 683788 524938 683800
rect 582558 683788 582564 683800
rect 524932 683760 582564 683788
rect 524932 683748 524938 683760
rect 582558 683748 582564 683760
rect 582616 683748 582622 683800
rect 405366 683680 405372 683732
rect 405424 683720 405430 683732
rect 437566 683720 437572 683732
rect 405424 683692 437572 683720
rect 405424 683680 405430 683692
rect 437566 683680 437572 683692
rect 437624 683680 437630 683732
rect 468294 683680 468300 683732
rect 468352 683720 468358 683732
rect 579246 683720 579252 683732
rect 468352 683692 579252 683720
rect 468352 683680 468358 683692
rect 579246 683680 579252 683692
rect 579304 683680 579310 683732
rect 377398 683612 377404 683664
rect 377456 683652 377462 683664
rect 422386 683652 422392 683664
rect 377456 683624 422392 683652
rect 377456 683612 377462 683624
rect 422386 683612 422392 683624
rect 422444 683612 422450 683664
rect 441246 683612 441252 683664
rect 441304 683652 441310 683664
rect 554038 683652 554044 683664
rect 441304 683624 554044 683652
rect 441304 683612 441310 683624
rect 554038 683612 554044 683624
rect 554096 683612 554102 683664
rect 438670 683544 438676 683596
rect 438728 683584 438734 683596
rect 567930 683584 567936 683596
rect 438728 683556 567936 683584
rect 438728 683544 438734 683556
rect 567930 683544 567936 683556
rect 567988 683544 567994 683596
rect 406470 683476 406476 683528
rect 406528 683516 406534 683528
rect 552290 683516 552296 683528
rect 406528 683488 552296 683516
rect 406528 683476 406534 683488
rect 552290 683476 552296 683488
rect 552348 683476 552354 683528
rect 407850 683408 407856 683460
rect 407908 683448 407914 683460
rect 553670 683448 553676 683460
rect 407908 683420 553676 683448
rect 407908 683408 407914 683420
rect 553670 683408 553676 683420
rect 553728 683408 553734 683460
rect 406562 683340 406568 683392
rect 406620 683380 406626 683392
rect 553578 683380 553584 683392
rect 406620 683352 553584 683380
rect 406620 683340 406626 683352
rect 553578 683340 553584 683352
rect 553636 683340 553642 683392
rect 403802 683272 403808 683324
rect 403860 683312 403866 683324
rect 555234 683312 555240 683324
rect 403860 683284 555240 683312
rect 403860 683272 403866 683284
rect 555234 683272 555240 683284
rect 555292 683272 555298 683324
rect 416682 683204 416688 683256
rect 416740 683244 416746 683256
rect 571334 683244 571340 683256
rect 416740 683216 571340 683244
rect 416740 683204 416746 683216
rect 571334 683204 571340 683216
rect 571392 683204 571398 683256
rect 404078 683136 404084 683188
rect 404136 683176 404142 683188
rect 580350 683176 580356 683188
rect 404136 683148 580356 683176
rect 404136 683136 404142 683148
rect 580350 683136 580356 683148
rect 580408 683136 580414 683188
rect 529658 682728 529664 682780
rect 529716 682768 529722 682780
rect 551278 682768 551284 682780
rect 529716 682740 551284 682768
rect 529716 682728 529722 682740
rect 551278 682728 551284 682740
rect 551336 682728 551342 682780
rect 408126 682660 408132 682712
rect 408184 682700 408190 682712
rect 553486 682700 553492 682712
rect 408184 682672 553492 682700
rect 408184 682660 408190 682672
rect 553486 682660 553492 682672
rect 553544 682660 553550 682712
rect 364242 682592 364248 682644
rect 364300 682632 364306 682644
rect 546954 682632 546960 682644
rect 364300 682604 546960 682632
rect 364300 682592 364306 682604
rect 546954 682592 546960 682604
rect 547012 682592 547018 682644
rect 3418 682524 3424 682576
rect 3476 682564 3482 682576
rect 550174 682564 550180 682576
rect 3476 682536 550180 682564
rect 3476 682524 3482 682536
rect 550174 682524 550180 682536
rect 550232 682524 550238 682576
rect 402330 682456 402336 682508
rect 402388 682496 402394 682508
rect 441890 682496 441896 682508
rect 402388 682468 441896 682496
rect 402388 682456 402394 682468
rect 441890 682456 441896 682468
rect 441948 682456 441954 682508
rect 507578 682456 507584 682508
rect 507636 682496 507642 682508
rect 553394 682496 553400 682508
rect 507636 682468 553400 682496
rect 507636 682456 507642 682468
rect 553394 682456 553400 682468
rect 553452 682456 553458 682508
rect 402238 682388 402244 682440
rect 402296 682428 402302 682440
rect 458634 682428 458640 682440
rect 402296 682400 458640 682428
rect 402296 682388 402302 682400
rect 458634 682388 458640 682400
rect 458692 682388 458698 682440
rect 477494 682388 477500 682440
rect 477552 682428 477558 682440
rect 566090 682428 566096 682440
rect 477552 682400 566096 682428
rect 477552 682388 477558 682400
rect 566090 682388 566096 682400
rect 566148 682388 566154 682440
rect 403710 682320 403716 682372
rect 403768 682360 403774 682372
rect 463786 682360 463792 682372
rect 403768 682332 463792 682360
rect 403768 682320 403774 682332
rect 463786 682320 463792 682332
rect 463844 682320 463850 682372
rect 502242 682320 502248 682372
rect 502300 682360 502306 682372
rect 560938 682360 560944 682372
rect 502300 682332 560944 682360
rect 502300 682320 502306 682332
rect 560938 682320 560944 682332
rect 560996 682320 561002 682372
rect 373258 682252 373264 682304
rect 373316 682292 373322 682304
rect 439958 682292 439964 682304
rect 373316 682264 439964 682292
rect 373316 682252 373322 682264
rect 439958 682252 439964 682264
rect 440016 682252 440022 682304
rect 447134 682252 447140 682304
rect 447192 682292 447198 682304
rect 509326 682292 509332 682304
rect 447192 682264 509332 682292
rect 447192 682252 447198 682264
rect 509326 682252 509332 682264
rect 509384 682252 509390 682304
rect 517238 682252 517244 682304
rect 517296 682292 517302 682304
rect 574094 682292 574100 682304
rect 517296 682264 574100 682292
rect 517296 682252 517302 682264
rect 574094 682252 574100 682264
rect 574152 682252 574158 682304
rect 385678 682184 385684 682236
rect 385736 682224 385742 682236
rect 480346 682224 480352 682236
rect 385736 682196 480352 682224
rect 385736 682184 385742 682196
rect 480346 682184 480352 682196
rect 480404 682184 480410 682236
rect 512730 682184 512736 682236
rect 512788 682224 512794 682236
rect 575566 682224 575572 682236
rect 512788 682196 575572 682224
rect 512788 682184 512794 682196
rect 575566 682184 575572 682196
rect 575624 682184 575630 682236
rect 360838 682116 360844 682168
rect 360896 682156 360902 682168
rect 429654 682156 429660 682168
rect 360896 682128 429660 682156
rect 360896 682116 360902 682128
rect 429654 682116 429660 682128
rect 429712 682116 429718 682168
rect 442994 682116 443000 682168
rect 443052 682156 443058 682168
rect 458450 682156 458456 682168
rect 443052 682128 458456 682156
rect 443052 682116 443058 682128
rect 458450 682116 458456 682128
rect 458508 682156 458514 682168
rect 554774 682156 554780 682168
rect 458508 682128 554780 682156
rect 458508 682116 458514 682128
rect 554774 682116 554780 682128
rect 554832 682116 554838 682168
rect 398098 682048 398104 682100
rect 398156 682088 398162 682100
rect 524966 682088 524972 682100
rect 398156 682060 524972 682088
rect 398156 682048 398162 682060
rect 524966 682048 524972 682060
rect 525024 682048 525030 682100
rect 549438 682048 549444 682100
rect 549496 682088 549502 682100
rect 577038 682088 577044 682100
rect 549496 682060 577044 682088
rect 549496 682048 549502 682060
rect 577038 682048 577044 682060
rect 577096 682048 577102 682100
rect 549990 681980 549996 682032
rect 550048 682020 550054 682032
rect 570138 682020 570144 682032
rect 550048 681992 570144 682020
rect 550048 681980 550054 681992
rect 570138 681980 570144 681992
rect 570196 681980 570202 682032
rect 387702 681912 387708 681964
rect 387760 681952 387766 681964
rect 534074 681952 534080 681964
rect 387760 681924 534080 681952
rect 387760 681912 387766 681924
rect 534074 681912 534080 681924
rect 534132 681912 534138 681964
rect 535270 681912 535276 681964
rect 535328 681952 535334 681964
rect 568758 681952 568764 681964
rect 535328 681924 568764 681952
rect 535328 681912 535334 681924
rect 568758 681912 568764 681924
rect 568816 681912 568822 681964
rect 403986 681844 403992 681896
rect 404044 681884 404050 681896
rect 580442 681884 580448 681896
rect 404044 681856 580448 681884
rect 404044 681844 404050 681856
rect 580442 681844 580448 681856
rect 580500 681844 580506 681896
rect 537846 681776 537852 681828
rect 537904 681816 537910 681828
rect 571610 681816 571616 681828
rect 537904 681788 571616 681816
rect 537904 681776 537910 681788
rect 571610 681776 571616 681788
rect 571668 681776 571674 681828
rect 499206 681708 499212 681760
rect 499264 681748 499270 681760
rect 517514 681748 517520 681760
rect 499264 681720 517520 681748
rect 499264 681708 499270 681720
rect 517514 681708 517520 681720
rect 517572 681708 517578 681760
rect 541710 681708 541716 681760
rect 541768 681748 541774 681760
rect 571978 681748 571984 681760
rect 541768 681720 571984 681748
rect 541768 681708 541774 681720
rect 571978 681708 571984 681720
rect 572036 681708 572042 681760
rect 400030 681300 400036 681352
rect 400088 681340 400094 681352
rect 580718 681340 580724 681352
rect 400088 681312 580724 681340
rect 400088 681300 400094 681312
rect 580718 681300 580724 681312
rect 580776 681300 580782 681352
rect 517514 681232 517520 681284
rect 517572 681272 517578 681284
rect 580258 681272 580264 681284
rect 517572 681244 580264 681272
rect 517572 681232 517578 681244
rect 580258 681232 580264 681244
rect 580316 681232 580322 681284
rect 174538 681164 174544 681216
rect 174596 681204 174602 681216
rect 461210 681204 461216 681216
rect 174596 681176 461216 681204
rect 174596 681164 174602 681176
rect 461210 681164 461216 681176
rect 461268 681164 461274 681216
rect 501782 681164 501788 681216
rect 501840 681204 501846 681216
rect 576118 681204 576124 681216
rect 501840 681176 576124 681204
rect 501840 681164 501846 681176
rect 576118 681164 576124 681176
rect 576176 681164 576182 681216
rect 407574 681096 407580 681148
rect 407632 681136 407638 681148
rect 442994 681136 443000 681148
rect 407632 681108 443000 681136
rect 407632 681096 407638 681108
rect 442994 681096 443000 681108
rect 443052 681096 443058 681148
rect 496630 681096 496636 681148
rect 496688 681136 496694 681148
rect 575474 681136 575480 681148
rect 496688 681108 575480 681136
rect 496688 681096 496694 681108
rect 575474 681096 575480 681108
rect 575532 681096 575538 681148
rect 408310 681028 408316 681080
rect 408368 681068 408374 681080
rect 447134 681068 447140 681080
rect 408368 681040 447140 681068
rect 408368 681028 408374 681040
rect 447134 681028 447140 681040
rect 447192 681028 447198 681080
rect 484854 681028 484860 681080
rect 484912 681068 484918 681080
rect 570046 681068 570052 681080
rect 484912 681040 570052 681068
rect 484912 681028 484918 681040
rect 570046 681028 570052 681040
rect 570104 681028 570110 681080
rect 342898 680960 342904 681012
rect 342956 681000 342962 681012
rect 432046 681000 432052 681012
rect 342956 680972 432052 681000
rect 342956 680960 342962 680972
rect 432046 680960 432052 680972
rect 432104 680960 432110 681012
rect 434622 680960 434628 681012
rect 434680 681000 434686 681012
rect 550726 681000 550732 681012
rect 434680 680972 550732 681000
rect 434680 680960 434686 680972
rect 550726 680960 550732 680972
rect 550784 680960 550790 681012
rect 409874 680892 409880 680944
rect 409932 680932 409938 680944
rect 552934 680932 552940 680944
rect 409932 680904 552940 680932
rect 409932 680892 409938 680904
rect 552934 680892 552940 680904
rect 552992 680892 552998 680944
rect 408954 680824 408960 680876
rect 409012 680864 409018 680876
rect 552106 680864 552112 680876
rect 409012 680836 552112 680864
rect 409012 680824 409018 680836
rect 552106 680824 552112 680836
rect 552164 680824 552170 680876
rect 406654 680756 406660 680808
rect 406712 680796 406718 680808
rect 551186 680796 551192 680808
rect 406712 680768 551192 680796
rect 406712 680756 406718 680768
rect 551186 680756 551192 680768
rect 551244 680756 551250 680808
rect 406838 680688 406844 680740
rect 406896 680728 406902 680740
rect 552750 680728 552756 680740
rect 406896 680700 552756 680728
rect 406896 680688 406902 680700
rect 552750 680688 552756 680700
rect 552808 680688 552814 680740
rect 406378 680620 406384 680672
rect 406436 680660 406442 680672
rect 555050 680660 555056 680672
rect 406436 680632 555056 680660
rect 406436 680620 406442 680632
rect 555050 680620 555056 680632
rect 555108 680620 555114 680672
rect 399570 680552 399576 680604
rect 399628 680592 399634 680604
rect 550910 680592 550916 680604
rect 399628 680564 550916 680592
rect 399628 680552 399634 680564
rect 550910 680552 550916 680564
rect 550968 680552 550974 680604
rect 400122 680484 400128 680536
rect 400180 680524 400186 680536
rect 552658 680524 552664 680536
rect 400180 680496 552664 680524
rect 400180 680484 400186 680496
rect 552658 680484 552664 680496
rect 552716 680484 552722 680536
rect 409414 680416 409420 680468
rect 409472 680456 409478 680468
rect 424502 680456 424508 680468
rect 409472 680428 424508 680456
rect 409472 680416 409478 680428
rect 424502 680416 424508 680428
rect 424560 680416 424566 680468
rect 399662 680348 399668 680400
rect 399720 680388 399726 680400
rect 427906 680388 427912 680400
rect 399720 680360 427912 680388
rect 399720 680348 399726 680360
rect 427906 680348 427912 680360
rect 427964 680348 427970 680400
rect 439314 680348 439320 680400
rect 439372 680388 439378 680400
rect 551002 680388 551008 680400
rect 439372 680360 551008 680388
rect 439372 680348 439378 680360
rect 551002 680348 551008 680360
rect 551060 680348 551066 680400
rect 437934 680076 437940 680128
rect 437992 680116 437998 680128
rect 446214 680116 446220 680128
rect 437992 680088 446220 680116
rect 437992 680076 437998 680088
rect 446214 680076 446220 680088
rect 446272 680076 446278 680128
rect 441798 680008 441804 680060
rect 441856 680048 441862 680060
rect 445754 680048 445760 680060
rect 441856 680020 445760 680048
rect 441856 680008 441862 680020
rect 445754 680008 445760 680020
rect 445812 680008 445818 680060
rect 435818 679940 435824 679992
rect 435876 679980 435882 679992
rect 446950 679980 446956 679992
rect 435876 679952 446956 679980
rect 435876 679940 435882 679952
rect 446950 679940 446956 679952
rect 447008 679940 447014 679992
rect 441706 679872 441712 679924
rect 441764 679912 441770 679924
rect 445938 679912 445944 679924
rect 441764 679884 445944 679912
rect 441764 679872 441770 679884
rect 445938 679872 445944 679884
rect 445996 679872 446002 679924
rect 465534 679872 465540 679924
rect 465592 679912 465598 679924
rect 467098 679912 467104 679924
rect 465592 679884 467104 679912
rect 465592 679872 465598 679884
rect 467098 679872 467104 679884
rect 467156 679872 467162 679924
rect 411254 679804 411260 679856
rect 411312 679844 411318 679856
rect 421466 679844 421472 679856
rect 411312 679816 421472 679844
rect 411312 679804 411318 679816
rect 421466 679804 421472 679816
rect 421524 679804 421530 679856
rect 434686 679816 446352 679844
rect 413738 679736 413744 679788
rect 413796 679776 413802 679788
rect 415210 679776 415216 679788
rect 413796 679748 415216 679776
rect 413796 679736 413802 679748
rect 415210 679736 415216 679748
rect 415268 679736 415274 679788
rect 415366 679748 425054 679776
rect 409598 679668 409604 679720
rect 409656 679708 409662 679720
rect 415366 679708 415394 679748
rect 409656 679680 415394 679708
rect 409656 679668 409662 679680
rect 415486 679668 415492 679720
rect 415544 679668 415550 679720
rect 425026 679708 425054 679748
rect 434686 679708 434714 679816
rect 442350 679736 442356 679788
rect 442408 679776 442414 679788
rect 442408 679748 445248 679776
rect 442408 679736 442414 679748
rect 425026 679680 434714 679708
rect 443914 679668 443920 679720
rect 443972 679708 443978 679720
rect 443972 679680 445156 679708
rect 443972 679668 443978 679680
rect 415348 679640 415354 679652
rect 408466 679612 415354 679640
rect 406746 679464 406752 679516
rect 406804 679504 406810 679516
rect 408466 679504 408494 679612
rect 415348 679600 415354 679612
rect 415406 679600 415412 679652
rect 415504 679640 415532 679668
rect 415504 679612 425054 679640
rect 414124 679544 414980 679572
rect 406804 679476 408494 679504
rect 406804 679464 406810 679476
rect 411254 679464 411260 679516
rect 411312 679464 411318 679516
rect 413738 679464 413744 679516
rect 413796 679464 413802 679516
rect 405274 679396 405280 679448
rect 405332 679436 405338 679448
rect 411272 679436 411300 679464
rect 405332 679408 411300 679436
rect 405332 679396 405338 679408
rect 396718 679328 396724 679380
rect 396776 679368 396782 679380
rect 413756 679368 413784 679464
rect 396776 679340 413784 679368
rect 396776 679328 396782 679340
rect 399938 679260 399944 679312
rect 399996 679300 400002 679312
rect 414124 679300 414152 679544
rect 414952 679436 414980 679544
rect 415210 679532 415216 679584
rect 415268 679572 415274 679584
rect 415268 679544 421420 679572
rect 415268 679532 415274 679544
rect 414952 679408 415164 679436
rect 399996 679272 414152 679300
rect 399996 679260 400002 679272
rect 358078 679192 358084 679244
rect 358136 679232 358142 679244
rect 415136 679232 415164 679408
rect 421392 679368 421420 679544
rect 421466 679464 421472 679516
rect 421524 679464 421530 679516
rect 425026 679504 425054 679612
rect 437446 679612 445064 679640
rect 432690 679532 432696 679584
rect 432748 679572 432754 679584
rect 437446 679572 437474 679612
rect 432748 679544 437474 679572
rect 432748 679532 432754 679544
rect 432782 679504 432788 679516
rect 425026 679476 432788 679504
rect 432782 679464 432788 679476
rect 432840 679464 432846 679516
rect 432966 679464 432972 679516
rect 433024 679504 433030 679516
rect 435818 679504 435824 679516
rect 433024 679476 435824 679504
rect 433024 679464 433030 679476
rect 435818 679464 435824 679476
rect 435876 679464 435882 679516
rect 437934 679504 437940 679516
rect 437446 679476 437940 679504
rect 421484 679436 421512 679464
rect 437446 679436 437474 679476
rect 437934 679464 437940 679476
rect 437992 679464 437998 679516
rect 441706 679464 441712 679516
rect 441764 679464 441770 679516
rect 441798 679464 441804 679516
rect 441856 679464 441862 679516
rect 442350 679464 442356 679516
rect 442408 679464 442414 679516
rect 443914 679464 443920 679516
rect 443972 679464 443978 679516
rect 421484 679408 437474 679436
rect 441724 679368 441752 679464
rect 421392 679340 441752 679368
rect 441816 679300 441844 679464
rect 420886 679272 441844 679300
rect 420886 679232 420914 679272
rect 442368 679232 442396 679464
rect 358136 679204 413140 679232
rect 415136 679204 420914 679232
rect 425026 679204 442396 679232
rect 358136 679192 358142 679204
rect 395522 679124 395528 679176
rect 395580 679164 395586 679176
rect 395580 679136 411392 679164
rect 395580 679124 395586 679136
rect 9674 679056 9680 679108
rect 9732 679096 9738 679108
rect 408862 679096 408868 679108
rect 9732 679068 408868 679096
rect 9732 679056 9738 679068
rect 408862 679056 408868 679068
rect 408920 679056 408926 679108
rect 3602 678988 3608 679040
rect 3660 679028 3666 679040
rect 411364 679028 411392 679136
rect 413112 679028 413140 679204
rect 425026 679164 425054 679204
rect 3660 679000 411254 679028
rect 411364 679000 412956 679028
rect 3660 678988 3666 679000
rect 411226 678620 411254 679000
rect 412928 678688 412956 679000
rect 413020 679000 413140 679028
rect 416792 679136 425054 679164
rect 429166 679136 435404 679164
rect 413020 678824 413048 679000
rect 416792 678824 416820 679136
rect 429166 679096 429194 679136
rect 413020 678796 416820 678824
rect 416976 679068 429194 679096
rect 416976 678688 417004 679068
rect 420932 679000 433380 679028
rect 420932 678756 420960 679000
rect 412928 678660 417004 678688
rect 420886 678728 420960 678756
rect 420886 678620 420914 678728
rect 411226 678592 420914 678620
rect 433352 678620 433380 679000
rect 435376 678824 435404 679136
rect 443932 678974 443960 679464
rect 445036 679300 445064 679612
rect 444944 679272 445064 679300
rect 444944 679096 444972 679272
rect 445128 679164 445156 679680
rect 445220 679232 445248 679748
rect 446214 679532 446220 679584
rect 446272 679532 446278 679584
rect 446324 679572 446352 679816
rect 466178 679804 466184 679856
rect 466236 679844 466242 679856
rect 466236 679816 471974 679844
rect 466236 679804 466242 679816
rect 462406 679736 462412 679788
rect 462464 679776 462470 679788
rect 467558 679776 467564 679788
rect 462464 679748 467564 679776
rect 462464 679736 462470 679748
rect 467558 679736 467564 679748
rect 467616 679736 467622 679788
rect 462286 679680 467328 679708
rect 462286 679572 462314 679680
rect 467190 679640 467196 679652
rect 446324 679544 462314 679572
rect 465184 679612 467196 679640
rect 445754 679464 445760 679516
rect 445812 679464 445818 679516
rect 445938 679464 445944 679516
rect 445996 679464 446002 679516
rect 445772 679300 445800 679464
rect 445956 679368 445984 679464
rect 446232 679436 446260 679532
rect 447088 679464 447094 679516
rect 447146 679504 447152 679516
rect 462406 679504 462412 679516
rect 447146 679476 462412 679504
rect 447146 679464 447152 679476
rect 462406 679464 462412 679476
rect 462464 679464 462470 679516
rect 465184 679436 465212 679612
rect 467190 679600 467196 679612
rect 467248 679600 467254 679652
rect 467300 679572 467328 679680
rect 471946 679640 471974 679816
rect 473446 679640 473452 679652
rect 471946 679612 473452 679640
rect 473446 679600 473452 679612
rect 473504 679600 473510 679652
rect 552014 679572 552020 679584
rect 465644 679544 466316 679572
rect 467300 679544 552020 679572
rect 465534 679504 465540 679516
rect 446232 679408 465212 679436
rect 465368 679476 465540 679504
rect 465368 679368 465396 679476
rect 465534 679464 465540 679476
rect 465592 679464 465598 679516
rect 465644 679436 465672 679544
rect 466178 679504 466184 679516
rect 445956 679340 465396 679368
rect 465552 679408 465672 679436
rect 466104 679476 466184 679504
rect 465552 679300 465580 679408
rect 445772 679272 465580 679300
rect 466104 679232 466132 679476
rect 466178 679464 466184 679476
rect 466236 679464 466242 679516
rect 466288 679300 466316 679544
rect 552014 679532 552020 679544
rect 552072 679532 552078 679584
rect 467098 679464 467104 679516
rect 467156 679464 467162 679516
rect 467466 679464 467472 679516
rect 467524 679464 467530 679516
rect 467558 679464 467564 679516
rect 467616 679504 467622 679516
rect 552382 679504 552388 679516
rect 467616 679476 552388 679504
rect 467616 679464 467622 679476
rect 552382 679464 552388 679476
rect 552440 679464 552446 679516
rect 467116 679368 467144 679464
rect 467484 679436 467512 679464
rect 557902 679436 557908 679448
rect 467484 679408 557908 679436
rect 557902 679396 557908 679408
rect 557960 679396 557966 679448
rect 553762 679368 553768 679380
rect 467116 679340 553768 679368
rect 553762 679328 553768 679340
rect 553820 679328 553826 679380
rect 580534 679300 580540 679312
rect 466288 679272 580540 679300
rect 580534 679260 580540 679272
rect 580592 679260 580598 679312
rect 445220 679204 466132 679232
rect 580810 679164 580816 679176
rect 445128 679136 580816 679164
rect 580810 679124 580816 679136
rect 580868 679124 580874 679176
rect 579062 679096 579068 679108
rect 444944 679068 579068 679096
rect 579062 679056 579068 679068
rect 579120 679056 579126 679108
rect 550818 679028 550824 679040
rect 444484 679000 550824 679028
rect 444484 678974 444512 679000
rect 550818 678988 550824 679000
rect 550876 678988 550882 679040
rect 552474 678988 552480 679040
rect 552532 679028 552538 679040
rect 582650 679028 582656 679040
rect 552532 679000 582656 679028
rect 552532 678988 552538 679000
rect 582650 678988 582656 679000
rect 582708 678988 582714 679040
rect 443932 678946 444052 678974
rect 435376 678796 438854 678824
rect 438826 678756 438854 678796
rect 444024 678756 444052 678946
rect 438826 678728 444052 678756
rect 444346 678946 444512 678974
rect 444346 678620 444374 678946
rect 552014 678920 552020 678972
rect 552072 678960 552078 678972
rect 552072 678932 552520 678960
rect 552072 678920 552078 678932
rect 552492 678904 552520 678932
rect 552474 678852 552480 678904
rect 552532 678852 552538 678904
rect 433352 678592 444374 678620
rect 407758 678512 407764 678564
rect 407816 678512 407822 678564
rect 407776 678360 407804 678512
rect 407758 678308 407764 678360
rect 407816 678308 407822 678360
rect 165522 678240 165528 678292
rect 165580 678280 165586 678292
rect 169754 678280 169760 678292
rect 165580 678252 169760 678280
rect 165580 678240 165586 678252
rect 169754 678240 169760 678252
rect 169812 678280 169818 678292
rect 337562 678280 337568 678292
rect 169812 678252 337568 678280
rect 169812 678240 169818 678252
rect 337562 678240 337568 678252
rect 337620 678240 337626 678292
rect 407942 678172 407948 678224
rect 408000 678212 408006 678224
rect 408402 678212 408408 678224
rect 408000 678184 408408 678212
rect 408000 678172 408006 678184
rect 408402 678172 408408 678184
rect 408460 678172 408466 678224
rect 325050 677696 325056 677748
rect 325108 677736 325114 677748
rect 343726 677736 343732 677748
rect 325108 677708 343732 677736
rect 325108 677696 325114 677708
rect 343726 677696 343732 677708
rect 343784 677696 343790 677748
rect 153102 677628 153108 677680
rect 153160 677668 153166 677680
rect 171134 677668 171140 677680
rect 153160 677640 171140 677668
rect 153160 677628 153166 677640
rect 171134 677628 171140 677640
rect 171192 677628 171198 677680
rect 325786 677628 325792 677680
rect 325844 677668 325850 677680
rect 353938 677668 353944 677680
rect 325844 677640 353944 677668
rect 325844 677628 325850 677640
rect 353938 677628 353944 677640
rect 353996 677628 354002 677680
rect 552106 677628 552112 677680
rect 552164 677668 552170 677680
rect 572806 677668 572812 677680
rect 552164 677640 572812 677668
rect 552164 677628 552170 677640
rect 572806 677628 572812 677640
rect 572864 677628 572870 677680
rect 7558 677560 7564 677612
rect 7616 677600 7622 677612
rect 407114 677600 407120 677612
rect 7616 677572 407120 677600
rect 7616 677560 7622 677572
rect 407114 677560 407120 677572
rect 407172 677560 407178 677612
rect 552014 677560 552020 677612
rect 552072 677600 552078 677612
rect 579614 677600 579620 677612
rect 552072 677572 579620 677600
rect 552072 677560 552078 677572
rect 579614 677560 579620 677572
rect 579672 677560 579678 677612
rect 337562 676812 337568 676864
rect 337620 676852 337626 676864
rect 400858 676852 400864 676864
rect 337620 676824 400864 676852
rect 337620 676812 337626 676824
rect 400858 676812 400864 676824
rect 400916 676812 400922 676864
rect 552014 674840 552020 674892
rect 552072 674880 552078 674892
rect 574278 674880 574284 674892
rect 552072 674852 574284 674880
rect 552072 674840 552078 674852
rect 574278 674840 574284 674852
rect 574336 674840 574342 674892
rect 552566 674092 552572 674144
rect 552624 674132 552630 674144
rect 552750 674132 552756 674144
rect 552624 674104 552756 674132
rect 552624 674092 552630 674104
rect 552750 674092 552756 674104
rect 552808 674092 552814 674144
rect 552014 672052 552020 672104
rect 552072 672092 552078 672104
rect 571702 672092 571708 672104
rect 552072 672064 571708 672092
rect 552072 672052 552078 672064
rect 571702 672052 571708 672064
rect 571760 672052 571766 672104
rect 552106 671780 552112 671832
rect 552164 671820 552170 671832
rect 552934 671820 552940 671832
rect 552164 671792 552940 671820
rect 552164 671780 552170 671792
rect 552934 671780 552940 671792
rect 552992 671780 552998 671832
rect 342990 670624 342996 670676
rect 343048 670664 343054 670676
rect 407114 670664 407120 670676
rect 343048 670636 407120 670664
rect 343048 670624 343054 670636
rect 407114 670624 407120 670636
rect 407172 670624 407178 670676
rect 552750 669332 552756 669384
rect 552808 669372 552814 669384
rect 563974 669372 563980 669384
rect 552808 669344 563980 669372
rect 552808 669332 552814 669344
rect 563974 669332 563980 669344
rect 564032 669332 564038 669384
rect 367830 667904 367836 667956
rect 367888 667944 367894 667956
rect 407114 667944 407120 667956
rect 367888 667916 407120 667944
rect 367888 667904 367894 667916
rect 407114 667904 407120 667916
rect 407172 667904 407178 667956
rect 551278 667836 551284 667888
rect 551336 667876 551342 667888
rect 552382 667876 552388 667888
rect 551336 667848 552388 667876
rect 551336 667836 551342 667848
rect 552382 667836 552388 667848
rect 552440 667836 552446 667888
rect 404906 666544 404912 666596
rect 404964 666584 404970 666596
rect 407114 666584 407120 666596
rect 404964 666556 407120 666584
rect 404964 666544 404970 666556
rect 407114 666544 407120 666556
rect 407172 666544 407178 666596
rect 364978 665184 364984 665236
rect 365036 665224 365042 665236
rect 407114 665224 407120 665236
rect 365036 665196 407120 665224
rect 365036 665184 365042 665196
rect 407114 665184 407120 665196
rect 407172 665184 407178 665236
rect 397454 663688 397460 663740
rect 397512 663728 397518 663740
rect 407114 663728 407120 663740
rect 397512 663700 407120 663728
rect 397512 663688 397518 663700
rect 407114 663688 407120 663700
rect 407172 663688 407178 663740
rect 388530 661104 388536 661156
rect 388588 661144 388594 661156
rect 407114 661144 407120 661156
rect 388588 661116 407120 661144
rect 388588 661104 388594 661116
rect 407114 661104 407120 661116
rect 407172 661104 407178 661156
rect 381538 661036 381544 661088
rect 381596 661076 381602 661088
rect 407206 661076 407212 661088
rect 381596 661048 407212 661076
rect 381596 661036 381602 661048
rect 407206 661036 407212 661048
rect 407264 661036 407270 661088
rect 553302 656888 553308 656940
rect 553360 656928 553366 656940
rect 563330 656928 563336 656940
rect 553360 656900 563336 656928
rect 553360 656888 553366 656900
rect 563330 656888 563336 656900
rect 563388 656888 563394 656940
rect 399386 655460 399392 655512
rect 399444 655500 399450 655512
rect 407114 655500 407120 655512
rect 399444 655472 407120 655500
rect 399444 655460 399450 655472
rect 407114 655460 407120 655472
rect 407172 655460 407178 655512
rect 383562 654100 383568 654152
rect 383620 654140 383626 654152
rect 407114 654140 407120 654152
rect 383620 654112 407120 654140
rect 383620 654100 383626 654112
rect 407114 654100 407120 654112
rect 407172 654100 407178 654152
rect 380158 652740 380164 652792
rect 380216 652780 380222 652792
rect 407114 652780 407120 652792
rect 380216 652752 407120 652780
rect 380216 652740 380222 652752
rect 407114 652740 407120 652752
rect 407172 652740 407178 652792
rect 553302 652740 553308 652792
rect 553360 652780 553366 652792
rect 560386 652780 560392 652792
rect 553360 652752 560392 652780
rect 553360 652740 553366 652752
rect 560386 652740 560392 652752
rect 560444 652740 560450 652792
rect 394602 651380 394608 651432
rect 394660 651420 394666 651432
rect 407114 651420 407120 651432
rect 394660 651392 407120 651420
rect 394660 651380 394666 651392
rect 407114 651380 407120 651392
rect 407172 651380 407178 651432
rect 400858 651312 400864 651364
rect 400916 651352 400922 651364
rect 407574 651352 407580 651364
rect 400916 651324 407580 651352
rect 400916 651312 400922 651324
rect 407574 651312 407580 651324
rect 407632 651312 407638 651364
rect 402514 648660 402520 648712
rect 402572 648700 402578 648712
rect 407114 648700 407120 648712
rect 402572 648672 407120 648700
rect 402572 648660 402578 648672
rect 407114 648660 407120 648672
rect 407172 648660 407178 648712
rect 347038 648592 347044 648644
rect 347096 648632 347102 648644
rect 407206 648632 407212 648644
rect 347096 648604 407212 648632
rect 347096 648592 347102 648604
rect 407206 648592 407212 648604
rect 407264 648592 407270 648644
rect 553302 648592 553308 648644
rect 553360 648632 553366 648644
rect 561858 648632 561864 648644
rect 553360 648604 561864 648632
rect 553360 648592 553366 648604
rect 561858 648592 561864 648604
rect 561916 648592 561922 648644
rect 552934 646144 552940 646196
rect 552992 646184 552998 646196
rect 556430 646184 556436 646196
rect 552992 646156 556436 646184
rect 552992 646144 552998 646156
rect 556430 646144 556436 646156
rect 556488 646144 556494 646196
rect 552934 644648 552940 644700
rect 552992 644688 552998 644700
rect 556798 644688 556804 644700
rect 552992 644660 556804 644688
rect 552992 644648 552998 644660
rect 556798 644648 556804 644660
rect 556856 644648 556862 644700
rect 403434 644580 403440 644632
rect 403492 644620 403498 644632
rect 407114 644620 407120 644632
rect 403492 644592 407120 644620
rect 403492 644580 403498 644592
rect 407114 644580 407120 644592
rect 407172 644580 407178 644632
rect 384942 644444 384948 644496
rect 385000 644484 385006 644496
rect 407390 644484 407396 644496
rect 385000 644456 407396 644484
rect 385000 644444 385006 644456
rect 407390 644444 407396 644456
rect 407448 644444 407454 644496
rect 553302 644444 553308 644496
rect 553360 644484 553366 644496
rect 565446 644484 565452 644496
rect 553360 644456 565452 644484
rect 553360 644444 553366 644456
rect 565446 644444 565452 644456
rect 565504 644444 565510 644496
rect 393130 643084 393136 643136
rect 393188 643124 393194 643136
rect 407206 643124 407212 643136
rect 393188 643096 407212 643124
rect 393188 643084 393194 643096
rect 407206 643084 407212 643096
rect 407264 643084 407270 643136
rect 552014 642200 552020 642252
rect 552072 642240 552078 642252
rect 555234 642240 555240 642252
rect 552072 642212 555240 642240
rect 552072 642200 552078 642212
rect 555234 642200 555240 642212
rect 555292 642200 555298 642252
rect 390462 641792 390468 641844
rect 390520 641832 390526 641844
rect 407298 641832 407304 641844
rect 390520 641804 407304 641832
rect 390520 641792 390526 641804
rect 407298 641792 407304 641804
rect 407356 641792 407362 641844
rect 344278 641724 344284 641776
rect 344336 641764 344342 641776
rect 407206 641764 407212 641776
rect 344336 641736 407212 641764
rect 344336 641724 344342 641736
rect 407206 641724 407212 641736
rect 407264 641724 407270 641776
rect 358170 640296 358176 640348
rect 358228 640336 358234 640348
rect 407206 640336 407212 640348
rect 358228 640308 407212 640336
rect 358228 640296 358234 640308
rect 407206 640296 407212 640308
rect 407264 640296 407270 640348
rect 552474 637644 552480 637696
rect 552532 637684 552538 637696
rect 563422 637684 563428 637696
rect 552532 637656 563428 637684
rect 552532 637644 552538 637656
rect 563422 637644 563428 637656
rect 563480 637644 563486 637696
rect 405642 637576 405648 637628
rect 405700 637616 405706 637628
rect 407482 637616 407488 637628
rect 405700 637588 407488 637616
rect 405700 637576 405706 637588
rect 407482 637576 407488 637588
rect 407540 637576 407546 637628
rect 552014 637576 552020 637628
rect 552072 637616 552078 637628
rect 564526 637616 564532 637628
rect 552072 637588 564532 637616
rect 552072 637576 552078 637588
rect 564526 637576 564532 637588
rect 564584 637576 564590 637628
rect 391842 636216 391848 636268
rect 391900 636256 391906 636268
rect 407206 636256 407212 636268
rect 391900 636228 407212 636256
rect 391900 636216 391906 636228
rect 407206 636216 407212 636228
rect 407264 636216 407270 636268
rect 387058 633428 387064 633480
rect 387116 633468 387122 633480
rect 407206 633468 407212 633480
rect 387116 633440 407212 633468
rect 387116 633428 387122 633440
rect 407206 633428 407212 633440
rect 407264 633428 407270 633480
rect 369118 632068 369124 632120
rect 369176 632108 369182 632120
rect 407206 632108 407212 632120
rect 369176 632080 407212 632108
rect 369176 632068 369182 632080
rect 407206 632068 407212 632080
rect 407264 632068 407270 632120
rect 556798 632000 556804 632052
rect 556856 632040 556862 632052
rect 580166 632040 580172 632052
rect 556856 632012 580172 632040
rect 556856 632000 556862 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 552014 631728 552020 631780
rect 552072 631768 552078 631780
rect 556522 631768 556528 631780
rect 552072 631740 556528 631768
rect 552072 631728 552078 631740
rect 556522 631728 556528 631740
rect 556580 631728 556586 631780
rect 390370 630640 390376 630692
rect 390428 630680 390434 630692
rect 407206 630680 407212 630692
rect 390428 630652 407212 630680
rect 390428 630640 390434 630652
rect 407206 630640 407212 630652
rect 407264 630640 407270 630692
rect 553302 629280 553308 629332
rect 553360 629320 553366 629332
rect 571426 629320 571432 629332
rect 553360 629292 571432 629320
rect 553360 629280 553366 629292
rect 571426 629280 571432 629292
rect 571484 629280 571490 629332
rect 378962 627920 378968 627972
rect 379020 627960 379026 627972
rect 407206 627960 407212 627972
rect 379020 627932 407212 627960
rect 379020 627920 379026 627932
rect 407206 627920 407212 627932
rect 407264 627920 407270 627972
rect 404722 625336 404728 625388
rect 404780 625376 404786 625388
rect 407390 625376 407396 625388
rect 404780 625348 407396 625376
rect 404780 625336 404786 625348
rect 407390 625336 407396 625348
rect 407448 625336 407454 625388
rect 553302 623772 553308 623824
rect 553360 623812 553366 623824
rect 562502 623812 562508 623824
rect 553360 623784 562508 623812
rect 553360 623772 553366 623784
rect 562502 623772 562508 623784
rect 562560 623772 562566 623824
rect 402606 622412 402612 622464
rect 402664 622452 402670 622464
rect 407206 622452 407212 622464
rect 402664 622424 407212 622452
rect 402664 622412 402670 622424
rect 407206 622412 407212 622424
rect 407264 622412 407270 622464
rect 553302 619624 553308 619676
rect 553360 619664 553366 619676
rect 577498 619664 577504 619676
rect 553360 619636 577504 619664
rect 553360 619624 553366 619636
rect 577498 619624 577504 619636
rect 577556 619624 577562 619676
rect 372062 618264 372068 618316
rect 372120 618304 372126 618316
rect 407206 618304 407212 618316
rect 372120 618276 407212 618304
rect 372120 618264 372126 618276
rect 407206 618264 407212 618276
rect 407264 618264 407270 618316
rect 553302 616836 553308 616888
rect 553360 616876 553366 616888
rect 577590 616876 577596 616888
rect 553360 616848 577596 616876
rect 553360 616836 553366 616848
rect 577590 616836 577596 616848
rect 577648 616836 577654 616888
rect 551278 615884 551284 615936
rect 551336 615924 551342 615936
rect 552658 615924 552664 615936
rect 551336 615896 552664 615924
rect 551336 615884 551342 615896
rect 552658 615884 552664 615896
rect 552716 615884 552722 615936
rect 369302 615476 369308 615528
rect 369360 615516 369366 615528
rect 407298 615516 407304 615528
rect 369360 615488 407304 615516
rect 369360 615476 369366 615488
rect 407298 615476 407304 615488
rect 407356 615476 407362 615528
rect 553302 614116 553308 614168
rect 553360 614156 553366 614168
rect 581178 614156 581184 614168
rect 553360 614128 581184 614156
rect 553360 614116 553366 614128
rect 581178 614116 581184 614128
rect 581236 614116 581242 614168
rect 392854 612756 392860 612808
rect 392912 612796 392918 612808
rect 407206 612796 407212 612808
rect 392912 612768 407212 612796
rect 392912 612756 392918 612768
rect 407206 612756 407212 612768
rect 407264 612756 407270 612808
rect 553302 612756 553308 612808
rect 553360 612796 553366 612808
rect 578878 612796 578884 612808
rect 553360 612768 578884 612796
rect 553360 612756 553366 612768
rect 578878 612756 578884 612768
rect 578936 612756 578942 612808
rect 346302 611328 346308 611380
rect 346360 611368 346366 611380
rect 371326 611368 371332 611380
rect 346360 611340 371332 611368
rect 346360 611328 346366 611340
rect 371326 611328 371332 611340
rect 371384 611328 371390 611380
rect 553302 611328 553308 611380
rect 553360 611368 553366 611380
rect 569954 611368 569960 611380
rect 553360 611340 569960 611368
rect 553360 611328 553366 611340
rect 569954 611328 569960 611340
rect 570012 611328 570018 611380
rect 553302 609968 553308 610020
rect 553360 610008 553366 610020
rect 570690 610008 570696 610020
rect 553360 609980 570696 610008
rect 553360 609968 553366 609980
rect 570690 609968 570696 609980
rect 570748 609968 570754 610020
rect 173802 608608 173808 608660
rect 173860 608648 173866 608660
rect 202138 608648 202144 608660
rect 173860 608620 202144 608648
rect 173860 608608 173866 608620
rect 202138 608608 202144 608620
rect 202196 608608 202202 608660
rect 373350 608608 373356 608660
rect 373408 608648 373414 608660
rect 407206 608648 407212 608660
rect 373408 608620 407212 608648
rect 373408 608608 373414 608620
rect 407206 608608 407212 608620
rect 407264 608608 407270 608660
rect 552474 608608 552480 608660
rect 552532 608648 552538 608660
rect 555694 608648 555700 608660
rect 552532 608620 555700 608648
rect 552532 608608 552538 608620
rect 555694 608608 555700 608620
rect 555752 608608 555758 608660
rect 173802 607180 173808 607232
rect 173860 607220 173866 607232
rect 199378 607220 199384 607232
rect 173860 607192 199384 607220
rect 173860 607180 173866 607192
rect 199378 607180 199384 607192
rect 199436 607180 199442 607232
rect 345106 607180 345112 607232
rect 345164 607220 345170 607232
rect 364334 607220 364340 607232
rect 345164 607192 364340 607220
rect 345164 607180 345170 607192
rect 364334 607180 364340 607192
rect 364392 607180 364398 607232
rect 369210 607180 369216 607232
rect 369268 607220 369274 607232
rect 407206 607220 407212 607232
rect 369268 607192 407212 607220
rect 369268 607180 369274 607192
rect 407206 607180 407212 607192
rect 407264 607180 407270 607232
rect 553302 607180 553308 607232
rect 553360 607220 553366 607232
rect 562042 607220 562048 607232
rect 553360 607192 562048 607220
rect 553360 607180 553366 607192
rect 562042 607180 562048 607192
rect 562100 607180 562106 607232
rect 345566 605820 345572 605872
rect 345624 605860 345630 605872
rect 365806 605860 365812 605872
rect 345624 605832 365812 605860
rect 345624 605820 345630 605832
rect 365806 605820 365812 605832
rect 365864 605820 365870 605872
rect 552014 603916 552020 603968
rect 552072 603956 552078 603968
rect 554774 603956 554780 603968
rect 552072 603928 554780 603956
rect 552072 603916 552078 603928
rect 554774 603916 554780 603928
rect 554832 603916 554838 603968
rect 553302 603100 553308 603152
rect 553360 603140 553366 603152
rect 563146 603140 563152 603152
rect 553360 603112 563152 603140
rect 553360 603100 553366 603112
rect 563146 603100 563152 603112
rect 563204 603100 563210 603152
rect 175918 601672 175924 601724
rect 175976 601712 175982 601724
rect 203058 601712 203064 601724
rect 175976 601684 203064 601712
rect 175976 601672 175982 601684
rect 203058 601672 203064 601684
rect 203116 601672 203122 601724
rect 376018 601672 376024 601724
rect 376076 601712 376082 601724
rect 407298 601712 407304 601724
rect 376076 601684 407304 601712
rect 376076 601672 376082 601684
rect 407298 601672 407304 601684
rect 407356 601672 407362 601724
rect 570598 600924 570604 600976
rect 570656 600964 570662 600976
rect 580902 600964 580908 600976
rect 570656 600936 580908 600964
rect 570656 600924 570662 600936
rect 580902 600924 580908 600936
rect 580960 600924 580966 600976
rect 378870 598952 378876 599004
rect 378928 598992 378934 599004
rect 407298 598992 407304 599004
rect 378928 598964 407304 598992
rect 378928 598952 378934 598964
rect 407298 598952 407304 598964
rect 407356 598952 407362 599004
rect 398650 596164 398656 596216
rect 398708 596204 398714 596216
rect 407298 596204 407304 596216
rect 398708 596176 407304 596204
rect 398708 596164 398714 596176
rect 407298 596164 407304 596176
rect 407356 596164 407362 596216
rect 401410 594804 401416 594856
rect 401468 594844 401474 594856
rect 407298 594844 407304 594856
rect 401468 594816 407304 594844
rect 401468 594804 401474 594816
rect 407298 594804 407304 594816
rect 407356 594804 407362 594856
rect 398558 592016 398564 592068
rect 398616 592056 398622 592068
rect 407298 592056 407304 592068
rect 398616 592028 407304 592056
rect 398616 592016 398622 592028
rect 407298 592016 407304 592028
rect 407356 592016 407362 592068
rect 32674 591948 32680 592000
rect 32732 591988 32738 592000
rect 204898 591988 204904 592000
rect 32732 591960 204904 591988
rect 32732 591948 32738 591960
rect 204898 591948 204904 591960
rect 204956 591948 204962 592000
rect 31570 591336 31576 591388
rect 31628 591376 31634 591388
rect 32398 591376 32404 591388
rect 31628 591348 32404 591376
rect 31628 591336 31634 591348
rect 32398 591336 32404 591348
rect 32456 591336 32462 591388
rect 32858 591336 32864 591388
rect 32916 591376 32922 591388
rect 78858 591376 78864 591388
rect 32916 591348 78864 591376
rect 32916 591336 32922 591348
rect 78858 591336 78864 591348
rect 78916 591336 78922 591388
rect 153654 591336 153660 591388
rect 153712 591376 153718 591388
rect 171318 591376 171324 591388
rect 153712 591348 171324 591376
rect 153712 591336 153718 591348
rect 171318 591336 171324 591348
rect 171376 591336 171382 591388
rect 32766 591268 32772 591320
rect 32824 591308 32830 591320
rect 306282 591308 306288 591320
rect 32824 591280 306288 591308
rect 32824 591268 32830 591280
rect 306282 591268 306288 591280
rect 306340 591268 306346 591320
rect 552014 590792 552020 590844
rect 552072 590832 552078 590844
rect 555786 590832 555792 590844
rect 552072 590804 555792 590832
rect 552072 590792 552078 590804
rect 555786 590792 555792 590804
rect 555844 590792 555850 590844
rect 36998 590656 37004 590708
rect 37056 590696 37062 590708
rect 407298 590696 407304 590708
rect 37056 590668 407304 590696
rect 37056 590656 37062 590668
rect 407298 590656 407304 590668
rect 407356 590656 407362 590708
rect 552474 590656 552480 590708
rect 552532 590696 552538 590708
rect 581086 590696 581092 590708
rect 552532 590668 581092 590696
rect 552532 590656 552538 590668
rect 581086 590656 581092 590668
rect 581144 590656 581150 590708
rect 48958 590248 48964 590300
rect 49016 590288 49022 590300
rect 60366 590288 60372 590300
rect 49016 590260 60372 590288
rect 49016 590248 49022 590260
rect 60366 590248 60372 590260
rect 60424 590248 60430 590300
rect 42610 590180 42616 590232
rect 42668 590220 42674 590232
rect 50062 590220 50068 590232
rect 42668 590192 50068 590220
rect 42668 590180 42674 590192
rect 50062 590180 50068 590192
rect 50120 590180 50126 590232
rect 317414 590180 317420 590232
rect 317472 590220 317478 590232
rect 343726 590220 343732 590232
rect 317472 590192 343732 590220
rect 317472 590180 317478 590192
rect 343726 590180 343732 590192
rect 343784 590180 343790 590232
rect 45278 590112 45284 590164
rect 45336 590152 45342 590164
rect 77294 590152 77300 590164
rect 45336 590124 77300 590152
rect 45336 590112 45342 590124
rect 77294 590112 77300 590124
rect 77352 590112 77358 590164
rect 292758 590112 292764 590164
rect 292816 590152 292822 590164
rect 406470 590152 406476 590164
rect 292816 590124 406476 590152
rect 292816 590112 292822 590124
rect 406470 590112 406476 590124
rect 406528 590112 406534 590164
rect 45094 590044 45100 590096
rect 45152 590084 45158 590096
rect 78674 590084 78680 590096
rect 45152 590056 78680 590084
rect 45152 590044 45158 590056
rect 78674 590044 78680 590056
rect 78732 590044 78738 590096
rect 257338 590044 257344 590096
rect 257396 590084 257402 590096
rect 406562 590084 406568 590096
rect 257396 590056 406568 590084
rect 257396 590044 257402 590056
rect 406562 590044 406568 590056
rect 406620 590044 406626 590096
rect 32858 589976 32864 590028
rect 32916 590016 32922 590028
rect 69014 590016 69020 590028
rect 32916 589988 69020 590016
rect 32916 589976 32922 589988
rect 69014 589976 69020 589988
rect 69072 589976 69078 590028
rect 225138 589976 225144 590028
rect 225196 590016 225202 590028
rect 400122 590016 400128 590028
rect 225196 589988 400128 590016
rect 225196 589976 225202 589988
rect 400122 589976 400128 589988
rect 400180 589976 400186 590028
rect 41230 589908 41236 589960
rect 41288 589948 41294 589960
rect 171134 589948 171140 589960
rect 41288 589920 171140 589948
rect 41288 589908 41294 589920
rect 171134 589908 171140 589920
rect 171192 589908 171198 589960
rect 226426 589908 226432 589960
rect 226484 589948 226490 589960
rect 405090 589948 405096 589960
rect 226484 589920 405096 589948
rect 226484 589908 226490 589920
rect 405090 589908 405096 589920
rect 405148 589908 405154 589960
rect 43714 589840 43720 589892
rect 43772 589880 43778 589892
rect 92474 589880 92480 589892
rect 43772 589852 92480 589880
rect 43772 589840 43778 589852
rect 92474 589840 92480 589852
rect 92532 589840 92538 589892
rect 44634 589772 44640 589824
rect 44692 589812 44698 589824
rect 127342 589812 127348 589824
rect 44692 589784 127348 589812
rect 44692 589772 44698 589784
rect 127342 589772 127348 589784
rect 127400 589772 127406 589824
rect 44726 589704 44732 589756
rect 44784 589744 44790 589756
rect 129734 589744 129740 589756
rect 44784 589716 129740 589744
rect 44784 589704 44790 589716
rect 129734 589704 129740 589716
rect 129792 589704 129798 589756
rect 55858 589636 55864 589688
rect 55916 589676 55922 589688
rect 227070 589676 227076 589688
rect 55916 589648 227076 589676
rect 55916 589636 55922 589648
rect 227070 589636 227076 589648
rect 227128 589636 227134 589688
rect 292114 589636 292120 589688
rect 292172 589676 292178 589688
rect 348510 589676 348516 589688
rect 292172 589648 348516 589676
rect 292172 589636 292178 589648
rect 348510 589636 348516 589648
rect 348568 589636 348574 589688
rect 47578 589568 47584 589620
rect 47636 589608 47642 589620
rect 241514 589608 241520 589620
rect 47636 589580 241520 589608
rect 47636 589568 47642 589580
rect 241514 589568 241520 589580
rect 241572 589568 241578 589620
rect 246666 589568 246672 589620
rect 246724 589608 246730 589620
rect 351178 589608 351184 589620
rect 246724 589580 351184 589608
rect 246724 589568 246730 589580
rect 351178 589568 351184 589580
rect 351236 589568 351242 589620
rect 25774 589500 25780 589552
rect 25832 589540 25838 589552
rect 223022 589540 223028 589552
rect 25832 589512 223028 589540
rect 25832 589500 25838 589512
rect 223022 589500 223028 589512
rect 223080 589500 223086 589552
rect 238386 589500 238392 589552
rect 238444 589540 238450 589552
rect 355042 589540 355048 589552
rect 238444 589512 355048 589540
rect 238444 589500 238450 589512
rect 355042 589500 355048 589512
rect 355100 589500 355106 589552
rect 41138 589432 41144 589484
rect 41196 589472 41202 589484
rect 99926 589472 99932 589484
rect 41196 589444 99932 589472
rect 41196 589432 41202 589444
rect 99926 589432 99932 589444
rect 99984 589432 99990 589484
rect 107562 589432 107568 589484
rect 107620 589472 107626 589484
rect 308398 589472 308404 589484
rect 107620 589444 308404 589472
rect 107620 589432 107626 589444
rect 308398 589432 308404 589444
rect 308456 589432 308462 589484
rect 312078 589432 312084 589484
rect 312136 589472 312142 589484
rect 354766 589472 354772 589484
rect 312136 589444 354772 589472
rect 312136 589432 312142 589444
rect 354766 589432 354772 589444
rect 354824 589432 354830 589484
rect 38378 589364 38384 589416
rect 38436 589404 38442 589416
rect 251174 589404 251180 589416
rect 38436 589376 251180 589404
rect 38436 589364 38442 589376
rect 251174 589364 251180 589376
rect 251232 589364 251238 589416
rect 252370 589364 252376 589416
rect 252428 589404 252434 589416
rect 355134 589404 355140 589416
rect 252428 589376 355140 589404
rect 252428 589364 252434 589376
rect 355134 589364 355140 589376
rect 355192 589364 355198 589416
rect 44910 589296 44916 589348
rect 44968 589336 44974 589348
rect 259454 589336 259460 589348
rect 44968 589308 259460 589336
rect 44968 589296 44974 589308
rect 259454 589296 259460 589308
rect 259512 589296 259518 589348
rect 289538 589296 289544 589348
rect 289596 589336 289602 589348
rect 350810 589336 350816 589348
rect 289596 589308 350816 589336
rect 289596 589296 289602 589308
rect 350810 589296 350816 589308
rect 350868 589296 350874 589348
rect 552014 588956 552020 589008
rect 552072 588996 552078 589008
rect 554866 588996 554872 589008
rect 552072 588968 554872 588996
rect 552072 588956 552078 588968
rect 554866 588956 554872 588968
rect 554924 588956 554930 589008
rect 74810 588616 74816 588668
rect 74868 588656 74874 588668
rect 295978 588656 295984 588668
rect 74868 588628 295984 588656
rect 74868 588616 74874 588628
rect 295978 588616 295984 588628
rect 296036 588616 296042 588668
rect 3510 588548 3516 588600
rect 3568 588588 3574 588600
rect 371970 588588 371976 588600
rect 3568 588560 371976 588588
rect 3568 588548 3574 588560
rect 371970 588548 371976 588560
rect 372028 588548 372034 588600
rect 386322 587868 386328 587920
rect 386380 587908 386386 587920
rect 407298 587908 407304 587920
rect 386380 587880 407304 587908
rect 386380 587868 386386 587880
rect 407298 587868 407304 587880
rect 407356 587868 407362 587920
rect 21818 587800 21824 587852
rect 21876 587840 21882 587852
rect 122558 587840 122564 587852
rect 21876 587812 122564 587840
rect 21876 587800 21882 587812
rect 122558 587800 122564 587812
rect 122616 587800 122622 587852
rect 171686 587800 171692 587852
rect 171744 587840 171750 587852
rect 236086 587840 236092 587852
rect 171744 587812 236092 587840
rect 171744 587800 171750 587812
rect 236086 587800 236092 587812
rect 236144 587800 236150 587852
rect 40954 587732 40960 587784
rect 41012 587772 41018 587784
rect 203610 587772 203616 587784
rect 41012 587744 203616 587772
rect 41012 587732 41018 587744
rect 203610 587732 203616 587744
rect 203668 587732 203674 587784
rect 256050 587732 256056 587784
rect 256108 587772 256114 587784
rect 359274 587772 359280 587784
rect 256108 587744 359280 587772
rect 256108 587732 256114 587744
rect 359274 587732 359280 587744
rect 359332 587732 359338 587784
rect 40862 587664 40868 587716
rect 40920 587704 40926 587716
rect 203518 587704 203524 587716
rect 40920 587676 203524 587704
rect 40920 587664 40926 587676
rect 203518 587664 203524 587676
rect 203576 587664 203582 587716
rect 240594 587664 240600 587716
rect 240652 587704 240658 587716
rect 354674 587704 354680 587716
rect 240652 587676 354680 587704
rect 240652 587664 240658 587676
rect 354674 587664 354680 587676
rect 354732 587664 354738 587716
rect 34882 587596 34888 587648
rect 34940 587636 34946 587648
rect 225322 587636 225328 587648
rect 34940 587608 225328 587636
rect 34940 587596 34946 587608
rect 225322 587596 225328 587608
rect 225380 587596 225386 587648
rect 239306 587596 239312 587648
rect 239364 587636 239370 587648
rect 399846 587636 399852 587648
rect 239364 587608 399852 587636
rect 239364 587596 239370 587608
rect 399846 587596 399852 587608
rect 399904 587596 399910 587648
rect 47026 587528 47032 587580
rect 47084 587568 47090 587580
rect 345014 587568 345020 587580
rect 47084 587540 345020 587568
rect 47084 587528 47090 587540
rect 345014 587528 345020 587540
rect 345072 587528 345078 587580
rect 100846 587460 100852 587512
rect 100904 587500 100910 587512
rect 405274 587500 405280 587512
rect 100904 587472 405280 587500
rect 100904 587460 100910 587472
rect 405274 587460 405280 587472
rect 405332 587460 405338 587512
rect 31570 587392 31576 587444
rect 31628 587432 31634 587444
rect 78674 587432 78680 587444
rect 31628 587404 78680 587432
rect 31628 587392 31634 587404
rect 78674 587392 78680 587404
rect 78732 587392 78738 587444
rect 86034 587392 86040 587444
rect 86092 587432 86098 587444
rect 396718 587432 396724 587444
rect 86092 587404 396724 587432
rect 86092 587392 86098 587404
rect 396718 587392 396724 587404
rect 396776 587392 396782 587444
rect 44082 587324 44088 587376
rect 44140 587364 44146 587376
rect 399754 587364 399760 587376
rect 44140 587336 399760 587364
rect 44140 587324 44146 587336
rect 399754 587324 399760 587336
rect 399812 587324 399818 587376
rect 39942 587256 39948 587308
rect 40000 587296 40006 587308
rect 399938 587296 399944 587308
rect 40000 587268 399944 587296
rect 40000 587256 40006 587268
rect 399938 587256 399944 587268
rect 399996 587256 400002 587308
rect 43990 587188 43996 587240
rect 44048 587228 44054 587240
rect 406930 587228 406936 587240
rect 44048 587200 406936 587228
rect 44048 587188 44054 587200
rect 406930 587188 406936 587200
rect 406988 587188 406994 587240
rect 36722 587120 36728 587172
rect 36780 587160 36786 587172
rect 402514 587160 402520 587172
rect 36780 587132 402520 587160
rect 36780 587120 36786 587132
rect 402514 587120 402520 587132
rect 402572 587120 402578 587172
rect 44818 587052 44824 587104
rect 44876 587092 44882 587104
rect 137278 587092 137284 587104
rect 44876 587064 137284 587092
rect 44876 587052 44882 587064
rect 137278 587052 137284 587064
rect 137336 587052 137342 587104
rect 215478 587052 215484 587104
rect 215536 587092 215542 587104
rect 278958 587092 278964 587104
rect 215536 587064 278964 587092
rect 215536 587052 215542 587064
rect 278958 587052 278964 587064
rect 279016 587052 279022 587104
rect 22738 586984 22744 587036
rect 22796 587024 22802 587036
rect 104894 587024 104900 587036
rect 22796 586996 104900 587024
rect 22796 586984 22802 586996
rect 104894 586984 104900 586996
rect 104952 586984 104958 587036
rect 41966 586508 41972 586560
rect 42024 586548 42030 586560
rect 407298 586548 407304 586560
rect 42024 586520 407304 586548
rect 42024 586508 42030 586520
rect 407298 586508 407304 586520
rect 407356 586508 407362 586560
rect 552014 586508 552020 586560
rect 552072 586548 552078 586560
rect 578970 586548 578976 586560
rect 552072 586520 578976 586548
rect 552072 586508 552078 586520
rect 578970 586508 578976 586520
rect 579028 586508 579034 586560
rect 163314 585896 163320 585948
rect 163372 585936 163378 585948
rect 231854 585936 231860 585948
rect 163372 585908 231860 585936
rect 163372 585896 163378 585908
rect 231854 585896 231860 585908
rect 231912 585896 231918 585948
rect 265066 585896 265072 585948
rect 265124 585936 265130 585948
rect 293954 585936 293960 585948
rect 265124 585908 293960 585936
rect 265124 585896 265130 585908
rect 293954 585896 293960 585908
rect 294012 585896 294018 585948
rect 150434 585828 150440 585880
rect 150492 585868 150498 585880
rect 171226 585868 171232 585880
rect 150492 585840 171232 585868
rect 150492 585828 150498 585840
rect 171226 585828 171232 585840
rect 171284 585828 171290 585880
rect 226610 585828 226616 585880
rect 226668 585868 226674 585880
rect 351454 585868 351460 585880
rect 226668 585840 351460 585868
rect 226668 585828 226674 585840
rect 351454 585828 351460 585840
rect 351512 585828 351518 585880
rect 65426 585760 65432 585812
rect 65484 585800 65490 585812
rect 351086 585800 351092 585812
rect 65484 585772 351092 585800
rect 65484 585760 65490 585772
rect 351086 585760 351092 585772
rect 351144 585760 351150 585812
rect 552014 585148 552020 585200
rect 552072 585188 552078 585200
rect 577222 585188 577228 585200
rect 552072 585160 577228 585188
rect 552072 585148 552078 585160
rect 577222 585148 577228 585160
rect 577280 585148 577286 585200
rect 160094 584468 160100 584520
rect 160152 584508 160158 584520
rect 254118 584508 254124 584520
rect 160152 584480 254124 584508
rect 160152 584468 160158 584480
rect 254118 584468 254124 584480
rect 254176 584468 254182 584520
rect 75730 584400 75736 584452
rect 75788 584440 75794 584452
rect 132494 584440 132500 584452
rect 75788 584412 132500 584440
rect 75788 584400 75794 584412
rect 132494 584400 132500 584412
rect 132552 584400 132558 584452
rect 140774 584400 140780 584452
rect 140832 584440 140838 584452
rect 345106 584440 345112 584452
rect 140832 584412 345112 584440
rect 140832 584400 140838 584412
rect 345106 584400 345112 584412
rect 345164 584400 345170 584452
rect 147214 583040 147220 583092
rect 147272 583080 147278 583092
rect 271874 583080 271880 583092
rect 147272 583052 271880 583080
rect 147272 583040 147278 583052
rect 271874 583040 271880 583052
rect 271932 583040 271938 583092
rect 320450 583040 320456 583092
rect 320508 583080 320514 583092
rect 381538 583080 381544 583092
rect 320508 583052 381544 583080
rect 320508 583040 320514 583052
rect 381538 583040 381544 583052
rect 381596 583040 381602 583092
rect 103422 582972 103428 583024
rect 103480 583012 103486 583024
rect 349614 583012 349620 583024
rect 103480 582984 349620 583012
rect 103480 582972 103486 582984
rect 349614 582972 349620 582984
rect 349672 582972 349678 583024
rect 135622 581748 135628 581800
rect 135680 581788 135686 581800
rect 248506 581788 248512 581800
rect 135680 581760 248512 581788
rect 135680 581748 135686 581760
rect 248506 581748 248512 581760
rect 248564 581748 248570 581800
rect 46658 581680 46664 581732
rect 46716 581720 46722 581732
rect 172606 581720 172612 581732
rect 46716 581692 172612 581720
rect 46716 581680 46722 581692
rect 172606 581680 172612 581692
rect 172664 581680 172670 581732
rect 202874 581680 202880 581732
rect 202932 581720 202938 581732
rect 242894 581720 242900 581732
rect 202932 581692 242900 581720
rect 202932 581680 202938 581692
rect 242894 581680 242900 581692
rect 242952 581680 242958 581732
rect 93762 581612 93768 581664
rect 93820 581652 93826 581664
rect 222194 581652 222200 581664
rect 93820 581624 222200 581652
rect 93820 581612 93826 581624
rect 222194 581612 222200 581624
rect 222252 581612 222258 581664
rect 277302 581612 277308 581664
rect 277360 581652 277366 581664
rect 350718 581652 350724 581664
rect 277360 581624 350724 581652
rect 277360 581612 277366 581624
rect 350718 581612 350724 581624
rect 350776 581612 350782 581664
rect 43898 580456 43904 580508
rect 43956 580496 43962 580508
rect 117314 580496 117320 580508
rect 43956 580468 117320 580496
rect 43956 580456 43962 580468
rect 117314 580456 117320 580468
rect 117372 580456 117378 580508
rect 204898 580456 204904 580508
rect 204956 580496 204962 580508
rect 250438 580496 250444 580508
rect 204956 580468 250444 580496
rect 204956 580456 204962 580468
rect 250438 580456 250444 580468
rect 250496 580456 250502 580508
rect 205542 580388 205548 580440
rect 205600 580428 205606 580440
rect 278590 580428 278596 580440
rect 205600 580400 278596 580428
rect 205600 580388 205606 580400
rect 278590 580388 278596 580400
rect 278648 580388 278654 580440
rect 297910 580388 297916 580440
rect 297968 580428 297974 580440
rect 347038 580428 347044 580440
rect 297968 580400 347044 580428
rect 297968 580388 297974 580400
rect 347038 580388 347044 580400
rect 347096 580388 347102 580440
rect 117314 580320 117320 580372
rect 117372 580360 117378 580372
rect 233234 580360 233240 580372
rect 117372 580332 233240 580360
rect 117372 580320 117378 580332
rect 233234 580320 233240 580332
rect 233292 580320 233298 580372
rect 239950 580320 239956 580372
rect 240008 580360 240014 580372
rect 350350 580360 350356 580372
rect 240008 580332 350356 580360
rect 240008 580320 240014 580332
rect 350350 580320 350356 580332
rect 350408 580320 350414 580372
rect 202138 580252 202144 580304
rect 202196 580292 202202 580304
rect 349890 580292 349896 580304
rect 202196 580264 349896 580292
rect 202196 580252 202202 580264
rect 349890 580252 349896 580264
rect 349948 580252 349954 580304
rect 383286 579640 383292 579692
rect 383344 579680 383350 579692
rect 407298 579680 407304 579692
rect 383344 579652 407304 579680
rect 383344 579640 383350 579652
rect 407298 579640 407304 579652
rect 407356 579640 407362 579692
rect 158622 578960 158628 579012
rect 158680 579000 158686 579012
rect 270218 579000 270224 579012
rect 158680 578972 270224 579000
rect 158680 578960 158686 578972
rect 270218 578960 270224 578972
rect 270276 578960 270282 579012
rect 282822 578960 282828 579012
rect 282880 579000 282886 579012
rect 350626 579000 350632 579012
rect 282880 578972 350632 579000
rect 282880 578960 282886 578972
rect 350626 578960 350632 578972
rect 350684 578960 350690 579012
rect 46382 578892 46388 578944
rect 46440 578932 46446 578944
rect 299474 578932 299480 578944
rect 46440 578904 299480 578932
rect 46440 578892 46446 578904
rect 299474 578892 299480 578904
rect 299532 578892 299538 578944
rect 552014 578212 552020 578264
rect 552072 578252 552078 578264
rect 563606 578252 563612 578264
rect 552072 578224 563612 578252
rect 552072 578212 552078 578224
rect 563606 578212 563612 578224
rect 563664 578212 563670 578264
rect 140682 577668 140688 577720
rect 140740 577708 140746 577720
rect 163958 577708 163964 577720
rect 140740 577680 163964 577708
rect 140740 577668 140746 577680
rect 163958 577668 163964 577680
rect 164016 577668 164022 577720
rect 230290 577668 230296 577720
rect 230348 577708 230354 577720
rect 306374 577708 306380 577720
rect 230348 577680 306380 577708
rect 230348 577668 230354 577680
rect 306374 577668 306380 577680
rect 306432 577668 306438 577720
rect 82630 577600 82636 577652
rect 82688 577640 82694 577652
rect 147858 577640 147864 577652
rect 82688 577612 147864 577640
rect 82688 577600 82694 577612
rect 147858 577600 147864 577612
rect 147916 577600 147922 577652
rect 154574 577600 154580 577652
rect 154632 577640 154638 577652
rect 251266 577640 251272 577652
rect 154632 577612 251272 577640
rect 154632 577600 154638 577612
rect 251266 577600 251272 577612
rect 251324 577600 251330 577652
rect 46842 577532 46848 577584
rect 46900 577572 46906 577584
rect 235994 577572 236000 577584
rect 46900 577544 236000 577572
rect 46900 577532 46906 577544
rect 235994 577532 236000 577544
rect 236052 577532 236058 577584
rect 240042 577532 240048 577584
rect 240100 577572 240106 577584
rect 349246 577572 349252 577584
rect 240100 577544 349252 577572
rect 240100 577532 240106 577544
rect 349246 577532 349252 577544
rect 349304 577532 349310 577584
rect 31386 577464 31392 577516
rect 31444 577504 31450 577516
rect 348050 577504 348056 577516
rect 31444 577476 348056 577504
rect 31444 577464 31450 577476
rect 348050 577464 348056 577476
rect 348108 577464 348114 577516
rect 552014 577464 552020 577516
rect 552072 577504 552078 577516
rect 556154 577504 556160 577516
rect 552072 577476 556160 577504
rect 552072 577464 552078 577476
rect 556154 577464 556160 577476
rect 556212 577464 556218 577516
rect 360930 576852 360936 576904
rect 360988 576892 360994 576904
rect 407298 576892 407304 576904
rect 360988 576864 407304 576892
rect 360988 576852 360994 576864
rect 407298 576852 407304 576864
rect 407356 576852 407362 576904
rect 308398 576240 308404 576292
rect 308456 576280 308462 576292
rect 330202 576280 330208 576292
rect 308456 576252 330208 576280
rect 308456 576240 308462 576252
rect 330202 576240 330208 576252
rect 330260 576240 330266 576292
rect 49050 576172 49056 576224
rect 49108 576212 49114 576224
rect 220814 576212 220820 576224
rect 49108 576184 220820 576212
rect 49108 576172 49114 576184
rect 220814 576172 220820 576184
rect 220872 576172 220878 576224
rect 270402 576172 270408 576224
rect 270460 576212 270466 576224
rect 307018 576212 307024 576224
rect 270460 576184 307024 576212
rect 270460 576172 270466 576184
rect 307018 576172 307024 576184
rect 307076 576172 307082 576224
rect 307754 576172 307760 576224
rect 307812 576212 307818 576224
rect 343634 576212 343640 576224
rect 307812 576184 343640 576212
rect 307812 576172 307818 576184
rect 343634 576172 343640 576184
rect 343692 576172 343698 576224
rect 81342 576104 81348 576156
rect 81400 576144 81406 576156
rect 347774 576144 347780 576156
rect 81400 576116 347780 576144
rect 81400 576104 81406 576116
rect 347774 576104 347780 576116
rect 347832 576104 347838 576156
rect 552014 575492 552020 575544
rect 552072 575532 552078 575544
rect 560570 575532 560576 575544
rect 552072 575504 560576 575532
rect 552072 575492 552078 575504
rect 560570 575492 560576 575504
rect 560628 575492 560634 575544
rect 264790 574948 264796 575000
rect 264848 574988 264854 575000
rect 354950 574988 354956 575000
rect 264848 574960 354956 574988
rect 264848 574948 264854 574960
rect 354950 574948 354956 574960
rect 355008 574948 355014 575000
rect 113082 574880 113088 574932
rect 113140 574920 113146 574932
rect 211706 574920 211712 574932
rect 113140 574892 211712 574920
rect 113140 574880 113146 574892
rect 211706 574880 211712 574892
rect 211764 574880 211770 574932
rect 237282 574880 237288 574932
rect 237340 574920 237346 574932
rect 347958 574920 347964 574932
rect 237340 574892 347964 574920
rect 237340 574880 237346 574892
rect 347958 574880 347964 574892
rect 348016 574880 348022 574932
rect 88242 574812 88248 574864
rect 88300 574852 88306 574864
rect 349430 574852 349436 574864
rect 88300 574824 349436 574852
rect 88300 574812 88306 574824
rect 349430 574812 349436 574824
rect 349488 574812 349494 574864
rect 3602 574744 3608 574796
rect 3660 574784 3666 574796
rect 384666 574784 384672 574796
rect 3660 574756 384672 574784
rect 3660 574744 3666 574756
rect 384666 574744 384672 574756
rect 384724 574744 384730 574796
rect 552014 574064 552020 574116
rect 552072 574104 552078 574116
rect 563514 574104 563520 574116
rect 552072 574076 563520 574104
rect 552072 574064 552078 574076
rect 563514 574064 563520 574076
rect 563572 574064 563578 574116
rect 45370 573588 45376 573640
rect 45428 573628 45434 573640
rect 223574 573628 223580 573640
rect 45428 573600 223580 573628
rect 45428 573588 45434 573600
rect 223574 573588 223580 573600
rect 223632 573588 223638 573640
rect 157242 573520 157248 573572
rect 157300 573560 157306 573572
rect 347866 573560 347872 573572
rect 157300 573532 347872 573560
rect 157300 573520 157306 573532
rect 347866 573520 347872 573532
rect 347924 573520 347930 573572
rect 95142 573452 95148 573504
rect 95200 573492 95206 573504
rect 331490 573492 331496 573504
rect 95200 573464 331496 573492
rect 95200 573452 95206 573464
rect 331490 573452 331496 573464
rect 331548 573452 331554 573504
rect 82722 573384 82728 573436
rect 82780 573424 82786 573436
rect 349798 573424 349804 573436
rect 82780 573396 349804 573424
rect 82780 573384 82786 573396
rect 349798 573384 349804 573396
rect 349856 573384 349862 573436
rect 52730 573316 52736 573368
rect 52788 573356 52794 573368
rect 404998 573356 405004 573368
rect 52788 573328 405004 573356
rect 52788 573316 52794 573328
rect 404998 573316 405004 573328
rect 405056 573316 405062 573368
rect 405366 572704 405372 572756
rect 405424 572744 405430 572756
rect 407666 572744 407672 572756
rect 405424 572716 407672 572744
rect 405424 572704 405430 572716
rect 407666 572704 407672 572716
rect 407724 572704 407730 572756
rect 552014 572704 552020 572756
rect 552072 572744 552078 572756
rect 582926 572744 582932 572756
rect 552072 572716 582932 572744
rect 552072 572704 552078 572716
rect 582926 572704 582932 572716
rect 582984 572704 582990 572756
rect 245838 572092 245844 572144
rect 245896 572132 245902 572144
rect 344278 572132 344284 572144
rect 245896 572104 344284 572132
rect 245896 572092 245902 572104
rect 344278 572092 344284 572104
rect 344336 572092 344342 572144
rect 245562 572024 245568 572076
rect 245620 572064 245626 572076
rect 353294 572064 353300 572076
rect 245620 572036 353300 572064
rect 245620 572024 245626 572036
rect 353294 572024 353300 572036
rect 353352 572024 353358 572076
rect 31478 571956 31484 572008
rect 31536 571996 31542 572008
rect 349154 571996 349160 572008
rect 31536 571968 349160 571996
rect 31536 571956 31542 571968
rect 349154 571956 349160 571968
rect 349212 571956 349218 572008
rect 236178 571344 236184 571396
rect 236236 571384 236242 571396
rect 363598 571384 363604 571396
rect 236236 571356 363604 571384
rect 236236 571344 236242 571356
rect 363598 571344 363604 571356
rect 363656 571344 363662 571396
rect 363690 571344 363696 571396
rect 363748 571384 363754 571396
rect 407298 571384 407304 571396
rect 363748 571356 407304 571384
rect 363748 571344 363754 571356
rect 407298 571344 407304 571356
rect 407356 571344 407362 571396
rect 264882 571208 264888 571260
rect 264940 571248 264946 571260
rect 350902 571248 350908 571260
rect 264940 571220 350908 571248
rect 264940 571208 264946 571220
rect 350902 571208 350908 571220
rect 350960 571208 350966 571260
rect 257890 571140 257896 571192
rect 257948 571180 257954 571192
rect 349338 571180 349344 571192
rect 257948 571152 349344 571180
rect 257948 571140 257954 571152
rect 349338 571140 349344 571152
rect 349396 571140 349402 571192
rect 230198 571072 230204 571124
rect 230256 571112 230262 571124
rect 361666 571112 361672 571124
rect 230256 571084 361672 571112
rect 230256 571072 230262 571084
rect 361666 571072 361672 571084
rect 361724 571072 361730 571124
rect 203886 571004 203892 571056
rect 203944 571044 203950 571056
rect 352558 571044 352564 571056
rect 203944 571016 352564 571044
rect 203944 571004 203950 571016
rect 352558 571004 352564 571016
rect 352616 571004 352622 571056
rect 84102 570936 84108 570988
rect 84160 570976 84166 570988
rect 237374 570976 237380 570988
rect 84160 570948 237380 570976
rect 84160 570936 84166 570948
rect 237374 570936 237380 570948
rect 237432 570936 237438 570988
rect 248322 570936 248328 570988
rect 248380 570976 248386 570988
rect 349706 570976 349712 570988
rect 248380 570948 349712 570976
rect 248380 570936 248386 570948
rect 349706 570936 349712 570948
rect 349764 570936 349770 570988
rect 46566 570868 46572 570920
rect 46624 570908 46630 570920
rect 260834 570908 260840 570920
rect 46624 570880 260840 570908
rect 46624 570868 46630 570880
rect 260834 570868 260840 570880
rect 260892 570868 260898 570920
rect 263502 570868 263508 570920
rect 263560 570908 263566 570920
rect 360194 570908 360200 570920
rect 263560 570880 360200 570908
rect 263560 570868 263566 570880
rect 360194 570868 360200 570880
rect 360252 570868 360258 570920
rect 46198 570800 46204 570852
rect 46256 570840 46262 570852
rect 296714 570840 296720 570852
rect 46256 570812 296720 570840
rect 46256 570800 46262 570812
rect 296714 570800 296720 570812
rect 296772 570800 296778 570852
rect 91002 570732 91008 570784
rect 91060 570772 91066 570784
rect 348142 570772 348148 570784
rect 91060 570744 348148 570772
rect 91060 570732 91066 570744
rect 348142 570732 348148 570744
rect 348200 570732 348206 570784
rect 60642 570664 60648 570716
rect 60700 570704 60706 570716
rect 352190 570704 352196 570716
rect 60700 570676 352196 570704
rect 60700 570664 60706 570676
rect 352190 570664 352196 570676
rect 352248 570664 352254 570716
rect 67542 570596 67548 570648
rect 67600 570636 67606 570648
rect 378134 570636 378140 570648
rect 67600 570608 378140 570636
rect 67600 570596 67606 570608
rect 378134 570596 378140 570608
rect 378192 570596 378198 570648
rect 290918 569916 290924 569968
rect 290976 569956 290982 569968
rect 368474 569956 368480 569968
rect 290976 569928 368480 569956
rect 290976 569916 290982 569928
rect 368474 569916 368480 569928
rect 368532 569916 368538 569968
rect 234522 569508 234528 569560
rect 234580 569548 234586 569560
rect 348234 569548 348240 569560
rect 234580 569520 348240 569548
rect 234580 569508 234586 569520
rect 348234 569508 348240 569520
rect 348292 569508 348298 569560
rect 230382 569440 230388 569492
rect 230440 569480 230446 569492
rect 352006 569480 352012 569492
rect 230440 569452 352012 569480
rect 230440 569440 230446 569452
rect 352006 569440 352012 569452
rect 352064 569440 352070 569492
rect 47670 569372 47676 569424
rect 47728 569412 47734 569424
rect 133874 569412 133880 569424
rect 47728 569384 133880 569412
rect 47728 569372 47734 569384
rect 133874 569372 133880 569384
rect 133932 569372 133938 569424
rect 229002 569372 229008 569424
rect 229060 569412 229066 569424
rect 356146 569412 356152 569424
rect 229060 569384 356152 569412
rect 229060 569372 229066 569384
rect 356146 569372 356152 569384
rect 356204 569372 356210 569424
rect 46474 569304 46480 569356
rect 46532 569344 46538 569356
rect 249794 569344 249800 569356
rect 46532 569316 249800 569344
rect 46532 569304 46538 569316
rect 249794 569304 249800 569316
rect 249852 569304 249858 569356
rect 257982 569304 257988 569356
rect 258040 569344 258046 569356
rect 353386 569344 353392 569356
rect 258040 569316 353392 569344
rect 258040 569304 258046 569316
rect 353386 569304 353392 569316
rect 353444 569304 353450 569356
rect 119982 569236 119988 569288
rect 120040 569276 120046 569288
rect 352650 569276 352656 569288
rect 120040 569248 352656 569276
rect 120040 569236 120046 569248
rect 352650 569236 352656 569248
rect 352708 569236 352714 569288
rect 115842 569168 115848 569220
rect 115900 569208 115906 569220
rect 353846 569208 353852 569220
rect 115900 569180 353852 569208
rect 115900 569168 115906 569180
rect 353846 569168 353852 569180
rect 353904 569168 353910 569220
rect 303982 568896 303988 568948
rect 304040 568936 304046 568948
rect 366358 568936 366364 568948
rect 304040 568908 366364 568936
rect 304040 568896 304046 568908
rect 366358 568896 366364 568908
rect 366416 568896 366422 568948
rect 265158 568828 265164 568880
rect 265216 568868 265222 568880
rect 357434 568868 357440 568880
rect 265216 568840 357440 568868
rect 265216 568828 265222 568840
rect 357434 568828 357440 568840
rect 357492 568828 357498 568880
rect 222010 568760 222016 568812
rect 222068 568800 222074 568812
rect 371234 568800 371240 568812
rect 222068 568772 371240 568800
rect 222068 568760 222074 568772
rect 371234 568760 371240 568772
rect 371292 568760 371298 568812
rect 198182 568692 198188 568744
rect 198240 568732 198246 568744
rect 357526 568732 357532 568744
rect 198240 568704 357532 568732
rect 198240 568692 198246 568704
rect 357526 568692 357532 568704
rect 357584 568692 357590 568744
rect 188522 568624 188528 568676
rect 188580 568664 188586 568676
rect 377490 568664 377496 568676
rect 188580 568636 377496 568664
rect 188580 568624 188586 568636
rect 377490 568624 377496 568636
rect 377548 568624 377554 568676
rect 36538 568556 36544 568608
rect 36596 568596 36602 568608
rect 407298 568596 407304 568608
rect 36596 568568 407304 568596
rect 36596 568556 36602 568568
rect 407298 568556 407304 568568
rect 407356 568556 407362 568608
rect 329650 568148 329656 568200
rect 329708 568188 329714 568200
rect 363046 568188 363052 568200
rect 329708 568160 363052 568188
rect 329708 568148 329714 568160
rect 363046 568148 363052 568160
rect 363104 568148 363110 568200
rect 259270 568080 259276 568132
rect 259328 568120 259334 568132
rect 348602 568120 348608 568132
rect 259328 568092 348608 568120
rect 259328 568080 259334 568092
rect 348602 568080 348608 568092
rect 348660 568080 348666 568132
rect 204162 568012 204168 568064
rect 204220 568052 204226 568064
rect 350994 568052 351000 568064
rect 204220 568024 351000 568052
rect 204220 568012 204226 568024
rect 350994 568012 351000 568024
rect 351052 568012 351058 568064
rect 203794 567944 203800 567996
rect 203852 567984 203858 567996
rect 356422 567984 356428 567996
rect 203852 567956 356428 567984
rect 203852 567944 203858 567956
rect 356422 567944 356428 567956
rect 356480 567944 356486 567996
rect 203978 567876 203984 567928
rect 204036 567916 204042 567928
rect 358998 567916 359004 567928
rect 204036 567888 359004 567916
rect 204036 567876 204042 567888
rect 358998 567876 359004 567888
rect 359056 567876 359062 567928
rect 46290 567808 46296 567860
rect 46348 567848 46354 567860
rect 234614 567848 234620 567860
rect 46348 567820 234620 567848
rect 46348 567808 46354 567820
rect 234614 567808 234620 567820
rect 234672 567808 234678 567860
rect 244182 567808 244188 567860
rect 244240 567848 244246 567860
rect 352282 567848 352288 567860
rect 244240 567820 352288 567848
rect 244240 567808 244246 567820
rect 352282 567808 352288 567820
rect 352340 567808 352346 567860
rect 289170 567604 289176 567656
rect 289228 567644 289234 567656
rect 373994 567644 374000 567656
rect 289228 567616 374000 567644
rect 289228 567604 289234 567616
rect 373994 567604 374000 567616
rect 374052 567604 374058 567656
rect 263226 567536 263232 567588
rect 263284 567576 263290 567588
rect 351914 567576 351920 567588
rect 263284 567548 351920 567576
rect 263284 567536 263290 567548
rect 351914 567536 351920 567548
rect 351972 567536 351978 567588
rect 241330 567468 241336 567520
rect 241388 567508 241394 567520
rect 358538 567508 358544 567520
rect 241388 567480 358544 567508
rect 241388 567468 241394 567480
rect 358538 567468 358544 567480
rect 358596 567468 358602 567520
rect 238662 567400 238668 567452
rect 238720 567440 238726 567452
rect 356054 567440 356060 567452
rect 238720 567412 356060 567440
rect 238720 567400 238726 567412
rect 356054 567400 356060 567412
rect 356112 567400 356118 567452
rect 131206 567332 131212 567384
rect 131264 567372 131270 567384
rect 354030 567372 354036 567384
rect 131264 567344 354036 567372
rect 131264 567332 131270 567344
rect 354030 567332 354036 567344
rect 354088 567332 354094 567384
rect 109954 567264 109960 567316
rect 110012 567304 110018 567316
rect 368198 567304 368204 567316
rect 110012 567276 368204 567304
rect 110012 567264 110018 567276
rect 368198 567264 368204 567276
rect 368256 567264 368262 567316
rect 553118 567264 553124 567316
rect 553176 567304 553182 567316
rect 559282 567304 559288 567316
rect 553176 567276 559288 567304
rect 553176 567264 553182 567276
rect 559282 567264 559288 567276
rect 559340 567264 559346 567316
rect 26050 567196 26056 567248
rect 26108 567236 26114 567248
rect 352098 567236 352104 567248
rect 26108 567208 352104 567236
rect 26108 567196 26114 567208
rect 352098 567196 352104 567208
rect 352156 567196 352162 567248
rect 374914 567196 374920 567248
rect 374972 567236 374978 567248
rect 407390 567236 407396 567248
rect 374972 567208 407396 567236
rect 374972 567196 374978 567208
rect 407390 567196 407396 567208
rect 407448 567196 407454 567248
rect 553302 567196 553308 567248
rect 553360 567236 553366 567248
rect 560478 567236 560484 567248
rect 553360 567208 560484 567236
rect 553360 567196 553366 567208
rect 560478 567196 560484 567208
rect 560536 567196 560542 567248
rect 329742 566720 329748 566772
rect 329800 566760 329806 566772
rect 353754 566760 353760 566772
rect 329800 566732 353760 566760
rect 329800 566720 329806 566732
rect 353754 566720 353760 566732
rect 353812 566720 353818 566772
rect 75638 566652 75644 566704
rect 75696 566692 75702 566704
rect 225414 566692 225420 566704
rect 75696 566664 225420 566692
rect 75696 566652 75702 566664
rect 225414 566652 225420 566664
rect 225472 566652 225478 566704
rect 253842 566652 253848 566704
rect 253900 566692 253906 566704
rect 349522 566692 349528 566704
rect 253900 566664 349528 566692
rect 253900 566652 253906 566664
rect 349522 566652 349528 566664
rect 349580 566652 349586 566704
rect 46750 566584 46756 566636
rect 46808 566624 46814 566636
rect 175918 566624 175924 566636
rect 46808 566596 175924 566624
rect 46808 566584 46814 566596
rect 175918 566584 175924 566596
rect 175976 566584 175982 566636
rect 204070 566584 204076 566636
rect 204128 566624 204134 566636
rect 353570 566624 353576 566636
rect 204128 566596 353576 566624
rect 204128 566584 204134 566596
rect 353570 566584 353576 566596
rect 353628 566584 353634 566636
rect 89622 566516 89628 566568
rect 89680 566556 89686 566568
rect 253934 566556 253940 566568
rect 89680 566528 253940 566556
rect 89680 566516 89686 566528
rect 253934 566516 253940 566528
rect 253992 566516 253998 566568
rect 262122 566516 262128 566568
rect 262180 566556 262186 566568
rect 348326 566556 348332 566568
rect 262180 566528 348332 566556
rect 262180 566516 262186 566528
rect 348326 566516 348332 566528
rect 348384 566516 348390 566568
rect 39574 566448 39580 566500
rect 39632 566488 39638 566500
rect 62206 566488 62212 566500
rect 39632 566460 62212 566488
rect 39632 566448 39638 566460
rect 62206 566448 62212 566460
rect 62264 566448 62270 566500
rect 125502 566448 125508 566500
rect 125560 566488 125566 566500
rect 353478 566488 353484 566500
rect 125560 566460 353484 566488
rect 125560 566448 125566 566460
rect 353478 566448 353484 566460
rect 353536 566448 353542 566500
rect 336274 566176 336280 566228
rect 336332 566216 336338 566228
rect 382918 566216 382924 566228
rect 336332 566188 382924 566216
rect 336332 566176 336338 566188
rect 382918 566176 382924 566188
rect 382976 566176 382982 566228
rect 233786 566108 233792 566160
rect 233844 566148 233850 566160
rect 347590 566148 347596 566160
rect 233844 566120 347596 566148
rect 233844 566108 233850 566120
rect 347590 566108 347596 566120
rect 347648 566108 347654 566160
rect 273162 566040 273168 566092
rect 273220 566080 273226 566092
rect 387794 566080 387800 566092
rect 273220 566052 387800 566080
rect 273220 566040 273226 566052
rect 387794 566040 387800 566052
rect 387852 566040 387858 566092
rect 40770 565972 40776 566024
rect 40828 566012 40834 566024
rect 372246 566012 372252 566024
rect 40828 565984 372252 566012
rect 40828 565972 40834 565984
rect 372246 565972 372252 565984
rect 372304 565972 372310 566024
rect 35618 565904 35624 565956
rect 35676 565944 35682 565956
rect 370682 565944 370688 565956
rect 35676 565916 370688 565944
rect 35676 565904 35682 565916
rect 370682 565904 370688 565916
rect 370740 565904 370746 565956
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 17218 565876 17224 565888
rect 3292 565848 17224 565876
rect 3292 565836 3298 565848
rect 17218 565836 17224 565848
rect 17276 565836 17282 565888
rect 34422 565836 34428 565888
rect 34480 565876 34486 565888
rect 380710 565876 380716 565888
rect 34480 565848 380716 565876
rect 34480 565836 34486 565848
rect 380710 565836 380716 565848
rect 380768 565836 380774 565888
rect 551462 565836 551468 565888
rect 551520 565876 551526 565888
rect 552474 565876 552480 565888
rect 551520 565848 552480 565876
rect 551520 565836 551526 565848
rect 552474 565836 552480 565848
rect 552532 565836 552538 565888
rect 31202 565360 31208 565412
rect 31260 565400 31266 565412
rect 404998 565400 405004 565412
rect 31260 565372 405004 565400
rect 31260 565360 31266 565372
rect 404998 565360 405004 565372
rect 405056 565360 405062 565412
rect 110322 565292 110328 565344
rect 110380 565332 110386 565344
rect 219710 565332 219716 565344
rect 110380 565304 219716 565332
rect 110380 565292 110386 565304
rect 219710 565292 219716 565304
rect 219768 565292 219774 565344
rect 242802 565292 242808 565344
rect 242860 565332 242866 565344
rect 281534 565332 281540 565344
rect 242860 565304 281540 565332
rect 242860 565292 242866 565304
rect 281534 565292 281540 565304
rect 281592 565292 281598 565344
rect 42150 565224 42156 565276
rect 42208 565264 42214 565276
rect 172514 565264 172520 565276
rect 42208 565236 172520 565264
rect 42208 565224 42214 565236
rect 172514 565224 172520 565236
rect 172572 565224 172578 565276
rect 199378 565224 199384 565276
rect 199436 565264 199442 565276
rect 243630 565264 243636 565276
rect 199436 565236 243636 565264
rect 199436 565224 199442 565236
rect 243630 565224 243636 565236
rect 243688 565224 243694 565276
rect 315942 565224 315948 565276
rect 316000 565264 316006 565276
rect 376110 565264 376116 565276
rect 316000 565236 376116 565264
rect 316000 565224 316006 565236
rect 376110 565224 376116 565236
rect 376168 565224 376174 565276
rect 87690 565156 87696 565208
rect 87748 565196 87754 565208
rect 244274 565196 244280 565208
rect 87748 565168 244280 565196
rect 87748 565156 87754 565168
rect 244274 565156 244280 565168
rect 244332 565156 244338 565208
rect 269850 565156 269856 565208
rect 269908 565196 269914 565208
rect 387242 565196 387248 565208
rect 269908 565168 387248 565196
rect 269908 565156 269914 565168
rect 387242 565156 387248 565168
rect 387300 565156 387306 565208
rect 42426 565088 42432 565140
rect 42484 565128 42490 565140
rect 51074 565128 51080 565140
rect 42484 565100 51080 565128
rect 42484 565088 42490 565100
rect 51074 565088 51080 565100
rect 51132 565088 51138 565140
rect 64782 565088 64788 565140
rect 64840 565128 64846 565140
rect 247034 565128 247040 565140
rect 64840 565100 247040 565128
rect 64840 565088 64846 565100
rect 247034 565088 247040 565100
rect 247092 565088 247098 565140
rect 251818 565088 251824 565140
rect 251876 565128 251882 565140
rect 369486 565128 369492 565140
rect 251876 565100 369492 565128
rect 251876 565088 251882 565100
rect 369486 565088 369492 565100
rect 369544 565088 369550 565140
rect 36906 565020 36912 565072
rect 36964 565060 36970 565072
rect 111886 565060 111892 565072
rect 36964 565032 111892 565060
rect 36964 565020 36970 565032
rect 111886 565020 111892 565032
rect 111944 565020 111950 565072
rect 235074 565020 235080 565072
rect 235132 565060 235138 565072
rect 355410 565060 355416 565072
rect 235132 565032 355416 565060
rect 235132 565020 235138 565032
rect 355410 565020 355416 565032
rect 355468 565020 355474 565072
rect 40678 564952 40684 565004
rect 40736 564992 40742 565004
rect 162302 564992 162308 565004
rect 40736 564964 162308 564992
rect 40736 564952 40742 564964
rect 162302 564952 162308 564964
rect 162360 564952 162366 565004
rect 255130 564952 255136 565004
rect 255188 564992 255194 565004
rect 388438 564992 388444 565004
rect 255188 564964 388444 564992
rect 255188 564952 255194 564964
rect 388438 564952 388444 564964
rect 388496 564952 388502 565004
rect 35342 564884 35348 564936
rect 35400 564924 35406 564936
rect 168558 564924 168564 564936
rect 35400 564896 168564 564924
rect 35400 564884 35406 564896
rect 168558 564884 168564 564896
rect 168616 564884 168622 564936
rect 232498 564884 232504 564936
rect 232556 564924 232562 564936
rect 369946 564924 369952 564936
rect 232556 564896 369952 564924
rect 232556 564884 232562 564896
rect 369946 564884 369952 564896
rect 370004 564884 370010 564936
rect 33962 564816 33968 564868
rect 34020 564856 34026 564868
rect 244918 564856 244924 564868
rect 34020 564828 244924 564856
rect 34020 564816 34026 564828
rect 244918 564816 244924 564828
rect 244976 564816 244982 564868
rect 248322 564816 248328 564868
rect 248380 564856 248386 564868
rect 391382 564856 391388 564868
rect 248380 564828 391388 564856
rect 248380 564816 248386 564828
rect 391382 564816 391388 564828
rect 391440 564816 391446 564868
rect 34974 564748 34980 564800
rect 35032 564788 35038 564800
rect 124950 564788 124956 564800
rect 35032 564760 124956 564788
rect 35032 564748 35038 564760
rect 124950 564748 124956 564760
rect 125008 564748 125014 564800
rect 146202 564748 146208 564800
rect 146260 564788 146266 564800
rect 358814 564788 358820 564800
rect 146260 564760 358820 564788
rect 146260 564748 146266 564760
rect 358814 564748 358820 564760
rect 358872 564748 358878 564800
rect 19242 564680 19248 564732
rect 19300 564720 19306 564732
rect 301406 564720 301412 564732
rect 19300 564692 301412 564720
rect 19300 564680 19306 564692
rect 301406 564680 301412 564692
rect 301464 564680 301470 564732
rect 314930 564680 314936 564732
rect 314988 564720 314994 564732
rect 377582 564720 377588 564732
rect 314988 564692 377588 564720
rect 314988 564680 314994 564692
rect 377582 564680 377588 564692
rect 377640 564680 377646 564732
rect 47854 564612 47860 564664
rect 47912 564652 47918 564664
rect 58986 564652 58992 564664
rect 47912 564624 58992 564652
rect 47912 564612 47918 564624
rect 58986 564612 58992 564624
rect 59044 564612 59050 564664
rect 62482 564612 62488 564664
rect 62540 564652 62546 564664
rect 400858 564652 400864 564664
rect 62540 564624 400864 564652
rect 62540 564612 62546 564624
rect 400858 564612 400864 564624
rect 400916 564612 400922 564664
rect 39850 564544 39856 564596
rect 39908 564584 39914 564596
rect 381722 564584 381728 564596
rect 39908 564556 381728 564584
rect 39908 564544 39914 564556
rect 381722 564544 381728 564556
rect 381780 564544 381786 564596
rect 36630 564476 36636 564528
rect 36688 564516 36694 564528
rect 405182 564516 405188 564528
rect 36688 564488 405188 564516
rect 36688 564476 36694 564488
rect 405182 564476 405188 564488
rect 405240 564476 405246 564528
rect 322106 564408 322112 564460
rect 322164 564448 322170 564460
rect 356330 564448 356336 564460
rect 322164 564420 356336 564448
rect 322164 564408 322170 564420
rect 356330 564408 356336 564420
rect 356388 564408 356394 564460
rect 404630 564408 404636 564460
rect 404688 564448 404694 564460
rect 407390 564448 407396 564460
rect 404688 564420 407396 564448
rect 404688 564408 404694 564420
rect 407390 564408 407396 564420
rect 407448 564408 407454 564460
rect 553302 564408 553308 564460
rect 553360 564448 553366 564460
rect 563698 564448 563704 564460
rect 553360 564420 563704 564448
rect 553360 564408 553366 564420
rect 563698 564408 563704 564420
rect 563756 564408 563762 564460
rect 43438 564068 43444 564120
rect 43496 564108 43502 564120
rect 407850 564108 407856 564120
rect 43496 564080 407856 564108
rect 43496 564068 43502 564080
rect 407850 564068 407856 564080
rect 407908 564068 407914 564120
rect 45186 564000 45192 564052
rect 45244 564040 45250 564052
rect 89714 564040 89720 564052
rect 45244 564012 89720 564040
rect 45244 564000 45250 564012
rect 89714 564000 89720 564012
rect 89772 564000 89778 564052
rect 42058 563932 42064 563984
rect 42116 563972 42122 563984
rect 86954 563972 86960 563984
rect 42116 563944 86960 563972
rect 42116 563932 42122 563944
rect 86954 563932 86960 563944
rect 87012 563932 87018 563984
rect 39666 563864 39672 563916
rect 39724 563904 39730 563916
rect 85574 563904 85580 563916
rect 39724 563876 85580 563904
rect 39724 563864 39730 563876
rect 85574 563864 85580 563876
rect 85632 563864 85638 563916
rect 324682 563864 324688 563916
rect 324740 563904 324746 563916
rect 354858 563904 354864 563916
rect 324740 563876 354864 563904
rect 324740 563864 324746 563876
rect 354858 563864 354864 563876
rect 354916 563864 354922 563916
rect 37090 563796 37096 563848
rect 37148 563836 37154 563848
rect 84194 563836 84200 563848
rect 37148 563808 84200 563836
rect 37148 563796 37154 563808
rect 84194 563796 84200 563808
rect 84252 563796 84258 563848
rect 179690 563796 179696 563848
rect 179748 563836 179754 563848
rect 258074 563836 258080 563848
rect 179748 563808 258080 563836
rect 179748 563796 179754 563808
rect 258074 563796 258080 563808
rect 258132 563796 258138 563848
rect 266262 563796 266268 563848
rect 266320 563836 266326 563848
rect 346486 563836 346492 563848
rect 266320 563808 346492 563836
rect 266320 563796 266326 563808
rect 346486 563796 346492 563808
rect 346544 563796 346550 563848
rect 34146 563728 34152 563780
rect 34204 563768 34210 563780
rect 81434 563768 81440 563780
rect 34204 563740 81440 563768
rect 34204 563728 34210 563740
rect 81434 563728 81440 563740
rect 81492 563728 81498 563780
rect 108298 563728 108304 563780
rect 108356 563768 108362 563780
rect 230474 563768 230480 563780
rect 108356 563740 230480 563768
rect 108356 563728 108362 563740
rect 230474 563728 230480 563740
rect 230532 563728 230538 563780
rect 260742 563728 260748 563780
rect 260800 563768 260806 563780
rect 343726 563768 343732 563780
rect 260800 563740 343732 563768
rect 260800 563728 260806 563740
rect 343726 563728 343732 563740
rect 343784 563728 343790 563780
rect 43622 563660 43628 563712
rect 43680 563700 43686 563712
rect 91094 563700 91100 563712
rect 43680 563672 91100 563700
rect 43680 563660 43686 563672
rect 91094 563660 91100 563672
rect 91152 563660 91158 563712
rect 208026 563660 208032 563712
rect 208084 563700 208090 563712
rect 354122 563700 354128 563712
rect 208084 563672 354128 563700
rect 208084 563660 208090 563672
rect 354122 563660 354128 563672
rect 354180 563660 354186 563712
rect 217778 563592 217784 563644
rect 217836 563632 217842 563644
rect 370958 563632 370964 563644
rect 217836 563604 370964 563632
rect 217836 563592 217842 563604
rect 370958 563592 370964 563604
rect 371016 563592 371022 563644
rect 39298 563524 39304 563576
rect 39356 563564 39362 563576
rect 86310 563564 86316 563576
rect 39356 563536 86316 563564
rect 39356 563524 39362 563536
rect 86310 563524 86316 563536
rect 86368 563524 86374 563576
rect 224218 563524 224224 563576
rect 224276 563564 224282 563576
rect 390002 563564 390008 563576
rect 224276 563536 390008 563564
rect 224276 563524 224282 563536
rect 390002 563524 390008 563536
rect 390060 563524 390066 563576
rect 38102 563456 38108 563508
rect 38160 563496 38166 563508
rect 191374 563496 191380 563508
rect 38160 563468 191380 563496
rect 38160 563456 38166 563468
rect 191374 563456 191380 563468
rect 191432 563456 191438 563508
rect 224770 563456 224776 563508
rect 224828 563496 224834 563508
rect 395430 563496 395436 563508
rect 224828 563468 395436 563496
rect 224828 563456 224834 563468
rect 395430 563456 395436 563468
rect 395488 563456 395494 563508
rect 179138 563388 179144 563440
rect 179196 563428 179202 563440
rect 381538 563428 381544 563440
rect 179196 563400 381544 563428
rect 179196 563388 179202 563400
rect 381538 563388 381544 563400
rect 381596 563388 381602 563440
rect 24762 563320 24768 563372
rect 24820 563360 24826 563372
rect 255498 563360 255504 563372
rect 24820 563332 255504 563360
rect 24820 563320 24826 563332
rect 255498 563320 255504 563332
rect 255556 563320 255562 563372
rect 307754 563320 307760 563372
rect 307812 563360 307818 563372
rect 308490 563360 308496 563372
rect 307812 563332 308496 563360
rect 307812 563320 307818 563332
rect 308490 563320 308496 563332
rect 308548 563320 308554 563372
rect 313090 563320 313096 563372
rect 313148 563360 313154 563372
rect 361574 563360 361580 563372
rect 313148 563332 361580 563360
rect 313148 563320 313154 563332
rect 361574 563320 361580 563332
rect 361632 563320 361638 563372
rect 24486 563252 24492 563304
rect 24544 563292 24550 563304
rect 255682 563292 255688 563304
rect 24544 563264 255688 563292
rect 24544 563252 24550 563264
rect 255682 563252 255688 563264
rect 255740 563252 255746 563304
rect 260742 563252 260748 563304
rect 260800 563292 260806 563304
rect 372614 563292 372620 563304
rect 260800 563264 372620 563292
rect 260800 563252 260806 563264
rect 372614 563252 372620 563264
rect 372672 563252 372678 563304
rect 24302 563184 24308 563236
rect 24360 563224 24366 563236
rect 325970 563224 325976 563236
rect 24360 563196 325976 563224
rect 24360 563184 24366 563196
rect 325970 563184 325976 563196
rect 326028 563184 326034 563236
rect 334986 563184 334992 563236
rect 335044 563224 335050 563236
rect 367094 563224 367100 563236
rect 335044 563196 367100 563224
rect 335044 563184 335050 563196
rect 367094 563184 367100 563196
rect 367152 563184 367158 563236
rect 32490 563116 32496 563168
rect 32548 563156 32554 563168
rect 395614 563156 395620 563168
rect 32548 563128 395620 563156
rect 32548 563116 32554 563128
rect 395614 563116 395620 563128
rect 395672 563116 395678 563168
rect 45002 563048 45008 563100
rect 45060 563088 45066 563100
rect 181070 563088 181076 563100
rect 45060 563060 181076 563088
rect 45060 563048 45066 563060
rect 181070 563048 181076 563060
rect 181128 563048 181134 563100
rect 340138 563048 340144 563100
rect 340196 563088 340202 563100
rect 354214 563088 354220 563100
rect 340196 563060 354220 563088
rect 340196 563048 340202 563060
rect 354214 563048 354220 563060
rect 354272 563048 354278 563100
rect 338022 562980 338028 563032
rect 338080 563020 338086 563032
rect 342898 563020 342904 563032
rect 338080 562992 342904 563020
rect 338080 562980 338086 562992
rect 342898 562980 342904 562992
rect 342956 562980 342962 563032
rect 70302 562640 70308 562692
rect 70360 562680 70366 562692
rect 91278 562680 91284 562692
rect 70360 562652 91284 562680
rect 70360 562640 70366 562652
rect 91278 562640 91284 562652
rect 91336 562640 91342 562692
rect 201402 562640 201408 562692
rect 201460 562680 201466 562692
rect 379054 562680 379060 562692
rect 201460 562652 379060 562680
rect 201460 562640 201466 562652
rect 379054 562640 379060 562652
rect 379112 562640 379118 562692
rect 22922 562572 22928 562624
rect 22980 562612 22986 562624
rect 65702 562612 65708 562624
rect 22980 562584 65708 562612
rect 22980 562572 22986 562584
rect 65702 562572 65708 562584
rect 65760 562572 65766 562624
rect 90818 562572 90824 562624
rect 90876 562612 90882 562624
rect 171778 562612 171784 562624
rect 90876 562584 171784 562612
rect 90876 562572 90882 562584
rect 171778 562572 171784 562584
rect 171836 562572 171842 562624
rect 317966 562572 317972 562624
rect 318024 562612 318030 562624
rect 365254 562612 365260 562624
rect 318024 562584 365260 562612
rect 318024 562572 318030 562584
rect 365254 562572 365260 562584
rect 365312 562572 365318 562624
rect 47210 562504 47216 562556
rect 47268 562544 47274 562556
rect 74534 562544 74540 562556
rect 47268 562516 74540 562544
rect 47268 562504 47274 562516
rect 74534 562504 74540 562516
rect 74592 562504 74598 562556
rect 76650 562504 76656 562556
rect 76708 562544 76714 562556
rect 174538 562544 174544 562556
rect 76708 562516 174544 562544
rect 76708 562504 76714 562516
rect 174538 562504 174544 562516
rect 174596 562504 174602 562556
rect 304074 562504 304080 562556
rect 304132 562544 304138 562556
rect 363782 562544 363788 562556
rect 304132 562516 363788 562544
rect 304132 562504 304138 562516
rect 363782 562504 363788 562516
rect 363840 562504 363846 562556
rect 41874 562436 41880 562488
rect 41932 562476 41938 562488
rect 50338 562476 50344 562488
rect 41932 562448 50344 562476
rect 41932 562436 41938 562448
rect 50338 562436 50344 562448
rect 50396 562436 50402 562488
rect 58986 562436 58992 562488
rect 59044 562476 59050 562488
rect 164326 562476 164332 562488
rect 59044 562448 164332 562476
rect 59044 562436 59050 562448
rect 164326 562436 164332 562448
rect 164384 562436 164390 562488
rect 203150 562436 203156 562488
rect 203208 562476 203214 562488
rect 340138 562476 340144 562488
rect 203208 562448 340144 562476
rect 203208 562436 203214 562448
rect 340138 562436 340144 562448
rect 340196 562436 340202 562488
rect 47302 562368 47308 562420
rect 47360 562408 47366 562420
rect 75914 562408 75920 562420
rect 47360 562380 75920 562408
rect 47360 562368 47366 562380
rect 75914 562368 75920 562380
rect 75972 562368 75978 562420
rect 157794 562368 157800 562420
rect 157852 562408 157858 562420
rect 303982 562408 303988 562420
rect 157852 562380 303988 562408
rect 157852 562368 157858 562380
rect 303982 562368 303988 562380
rect 304040 562368 304046 562420
rect 305914 562368 305920 562420
rect 305972 562408 305978 562420
rect 365070 562408 365076 562420
rect 305972 562380 365076 562408
rect 305972 562368 305978 562380
rect 365070 562368 365076 562380
rect 365128 562368 365134 562420
rect 39758 562300 39764 562352
rect 39816 562340 39822 562352
rect 81618 562340 81624 562352
rect 39816 562312 81624 562340
rect 39816 562300 39822 562312
rect 81618 562300 81624 562312
rect 81676 562300 81682 562352
rect 148778 562300 148784 562352
rect 148836 562340 148842 562352
rect 336182 562340 336188 562352
rect 148836 562312 336188 562340
rect 148836 562300 148842 562312
rect 336182 562300 336188 562312
rect 336240 562300 336246 562352
rect 35802 562232 35808 562284
rect 35860 562272 35866 562284
rect 83734 562272 83740 562284
rect 35860 562244 83740 562272
rect 35860 562232 35866 562244
rect 83734 562232 83740 562244
rect 83792 562232 83798 562284
rect 278314 562232 278320 562284
rect 278372 562272 278378 562284
rect 347222 562272 347228 562284
rect 278372 562244 347228 562272
rect 278372 562232 278378 562244
rect 347222 562232 347228 562244
rect 347280 562232 347286 562284
rect 36262 562164 36268 562216
rect 36320 562204 36326 562216
rect 94774 562204 94780 562216
rect 36320 562176 94780 562204
rect 36320 562164 36326 562176
rect 94774 562164 94780 562176
rect 94832 562164 94838 562216
rect 243538 562164 243544 562216
rect 243596 562204 243602 562216
rect 363874 562204 363880 562216
rect 243596 562176 363880 562204
rect 243596 562164 243602 562176
rect 363874 562164 363880 562176
rect 363932 562164 363938 562216
rect 43346 562096 43352 562148
rect 43404 562136 43410 562148
rect 50246 562136 50252 562148
rect 43404 562108 50252 562136
rect 43404 562096 43410 562108
rect 50246 562096 50252 562108
rect 50304 562096 50310 562148
rect 50338 562096 50344 562148
rect 50396 562136 50402 562148
rect 99374 562136 99380 562148
rect 50396 562108 99380 562136
rect 50396 562096 50402 562108
rect 99374 562096 99380 562108
rect 99432 562096 99438 562148
rect 260282 562096 260288 562148
rect 260340 562136 260346 562148
rect 387334 562136 387340 562148
rect 260340 562108 387340 562136
rect 260340 562096 260346 562108
rect 387334 562096 387340 562108
rect 387392 562096 387398 562148
rect 38286 562028 38292 562080
rect 38344 562068 38350 562080
rect 45830 562068 45836 562080
rect 38344 562040 45836 562068
rect 38344 562028 38350 562040
rect 45830 562028 45836 562040
rect 45888 562028 45894 562080
rect 46014 562028 46020 562080
rect 46072 562068 46078 562080
rect 105078 562068 105084 562080
rect 46072 562040 105084 562068
rect 46072 562028 46078 562040
rect 105078 562028 105084 562040
rect 105136 562028 105142 562080
rect 214466 562028 214472 562080
rect 214524 562068 214530 562080
rect 347314 562068 347320 562080
rect 214524 562040 347320 562068
rect 214524 562028 214530 562040
rect 347314 562028 347320 562040
rect 347372 562028 347378 562080
rect 347682 562028 347688 562080
rect 347740 562068 347746 562080
rect 391198 562068 391204 562080
rect 347740 562040 391204 562068
rect 347740 562028 347746 562040
rect 391198 562028 391204 562040
rect 391256 562028 391262 562080
rect 20622 561960 20628 562012
rect 20680 562000 20686 562012
rect 43346 562000 43352 562012
rect 20680 561972 43352 562000
rect 20680 561960 20686 561972
rect 43346 561960 43352 561972
rect 43404 561960 43410 562012
rect 48222 561960 48228 562012
rect 48280 562000 48286 562012
rect 49050 562000 49056 562012
rect 48280 561972 49056 562000
rect 48280 561960 48286 561972
rect 49050 561960 49056 561972
rect 49108 561960 49114 562012
rect 52822 561960 52828 562012
rect 52880 562000 52886 562012
rect 138014 562000 138020 562012
rect 52880 561972 138020 562000
rect 52880 561960 52886 561972
rect 138014 561960 138020 561972
rect 138072 561960 138078 562012
rect 250438 561960 250444 562012
rect 250496 562000 250502 562012
rect 403618 562000 403624 562012
rect 250496 561972 403624 562000
rect 250496 561960 250502 561972
rect 403618 561960 403624 561972
rect 403676 561960 403682 562012
rect 22830 561892 22836 561944
rect 22888 561932 22894 561944
rect 113450 561932 113456 561944
rect 22888 561904 113456 561932
rect 22888 561892 22894 561904
rect 113450 561892 113456 561904
rect 113508 561892 113514 561944
rect 186866 561892 186872 561944
rect 186924 561932 186930 561944
rect 340138 561932 340144 561944
rect 186924 561904 340144 561932
rect 186924 561892 186930 561904
rect 340138 561892 340144 561904
rect 340196 561892 340202 561944
rect 24394 561824 24400 561876
rect 24452 561864 24458 561876
rect 51534 561864 51540 561876
rect 24452 561836 51540 561864
rect 24452 561824 24458 561836
rect 51534 561824 51540 561836
rect 51592 561824 51598 561876
rect 51994 561824 52000 561876
rect 52052 561864 52058 561876
rect 181622 561864 181628 561876
rect 52052 561836 181628 561864
rect 52052 561824 52058 561836
rect 181622 561824 181628 561836
rect 181680 561824 181686 561876
rect 192570 561824 192576 561876
rect 192628 561864 192634 561876
rect 365714 561864 365720 561876
rect 192628 561836 365720 561864
rect 192628 561824 192634 561836
rect 365714 561824 365720 561836
rect 365772 561824 365778 561876
rect 41322 561756 41328 561808
rect 41380 561796 41386 561808
rect 193858 561796 193864 561808
rect 41380 561768 193864 561796
rect 41380 561756 41386 561768
rect 193858 561756 193864 561768
rect 193916 561756 193922 561808
rect 340046 561756 340052 561808
rect 340104 561796 340110 561808
rect 358354 561796 358360 561808
rect 340104 561768 358360 561796
rect 340104 561756 340110 561768
rect 358354 561756 358360 561768
rect 358412 561756 358418 561808
rect 31478 561688 31484 561740
rect 31536 561728 31542 561740
rect 138566 561728 138572 561740
rect 31536 561700 138572 561728
rect 31536 561688 31542 561700
rect 138566 561688 138572 561700
rect 138624 561688 138630 561740
rect 140498 561688 140504 561740
rect 140556 561728 140562 561740
rect 319162 561728 319168 561740
rect 140556 561700 319168 561728
rect 140556 561688 140562 561700
rect 319162 561688 319168 561700
rect 319220 561688 319226 561740
rect 325602 561688 325608 561740
rect 325660 561728 325666 561740
rect 355226 561728 355232 561740
rect 325660 561700 355232 561728
rect 325660 561688 325666 561700
rect 355226 561688 355232 561700
rect 355284 561688 355290 561740
rect 47118 561552 47124 561604
rect 47176 561592 47182 561604
rect 66254 561592 66260 561604
rect 47176 561564 66260 561592
rect 47176 561552 47182 561564
rect 66254 561552 66260 561564
rect 66312 561552 66318 561604
rect 29914 561484 29920 561536
rect 29972 561524 29978 561536
rect 51166 561524 51172 561536
rect 29972 561496 51172 561524
rect 29972 561484 29978 561496
rect 51166 561484 51172 561496
rect 51224 561484 51230 561536
rect 47486 561416 47492 561468
rect 47544 561456 47550 561468
rect 73154 561456 73160 561468
rect 47544 561428 73160 561456
rect 47544 561416 47550 561428
rect 73154 561416 73160 561428
rect 73212 561416 73218 561468
rect 21726 561348 21732 561400
rect 21784 561388 21790 561400
rect 53834 561388 53840 561400
rect 21784 561360 53840 561388
rect 21784 561348 21790 561360
rect 53834 561348 53840 561360
rect 53892 561348 53898 561400
rect 35526 561280 35532 561332
rect 35584 561320 35590 561332
rect 67726 561320 67732 561332
rect 35584 561292 67732 561320
rect 35584 561280 35590 561292
rect 67726 561280 67732 561292
rect 67784 561280 67790 561332
rect 25590 561212 25596 561264
rect 25648 561252 25654 561264
rect 58066 561252 58072 561264
rect 25648 561224 58072 561252
rect 25648 561212 25654 561224
rect 58066 561212 58072 561224
rect 58124 561212 58130 561264
rect 28718 561144 28724 561196
rect 28776 561184 28782 561196
rect 62114 561184 62120 561196
rect 28776 561156 62120 561184
rect 28776 561144 28782 561156
rect 62114 561144 62120 561156
rect 62172 561144 62178 561196
rect 307662 561144 307668 561196
rect 307720 561184 307726 561196
rect 355318 561184 355324 561196
rect 307720 561156 355324 561184
rect 307720 561144 307726 561156
rect 355318 561144 355324 561156
rect 355376 561144 355382 561196
rect 27246 561076 27252 561128
rect 27304 561116 27310 561128
rect 60826 561116 60832 561128
rect 27304 561088 60832 561116
rect 27304 561076 27310 561088
rect 60826 561076 60832 561088
rect 60884 561076 60890 561128
rect 337562 561076 337568 561128
rect 337620 561116 337626 561128
rect 405274 561116 405280 561128
rect 337620 561088 405280 561116
rect 337620 561076 337626 561088
rect 405274 561076 405280 561088
rect 405332 561076 405338 561128
rect 38194 561008 38200 561060
rect 38252 561048 38258 561060
rect 71774 561048 71780 561060
rect 38252 561020 71780 561048
rect 38252 561008 38258 561020
rect 71774 561008 71780 561020
rect 71832 561008 71838 561060
rect 315666 561008 315672 561060
rect 315724 561048 315730 561060
rect 395338 561048 395344 561060
rect 315724 561020 395344 561048
rect 315724 561008 315730 561020
rect 395338 561008 395344 561020
rect 395396 561008 395402 561060
rect 34054 560940 34060 560992
rect 34112 560980 34118 560992
rect 67634 560980 67640 560992
rect 34112 560952 67640 560980
rect 34112 560940 34118 560952
rect 67634 560940 67640 560952
rect 67692 560940 67698 560992
rect 299382 560940 299388 560992
rect 299440 560980 299446 560992
rect 380250 560980 380256 560992
rect 299440 560952 380256 560980
rect 299440 560940 299446 560952
rect 380250 560940 380256 560952
rect 380308 560940 380314 560992
rect 287882 560872 287888 560924
rect 287940 560912 287946 560924
rect 374638 560912 374644 560924
rect 287940 560884 374644 560912
rect 287940 560872 287946 560884
rect 374638 560872 374644 560884
rect 374696 560872 374702 560924
rect 244826 560804 244832 560856
rect 244884 560844 244890 560856
rect 376846 560844 376852 560856
rect 244884 560816 376852 560844
rect 244884 560804 244890 560816
rect 376846 560804 376852 560816
rect 376904 560804 376910 560856
rect 240962 560736 240968 560788
rect 241020 560776 241026 560788
rect 376754 560776 376760 560788
rect 241020 560748 376760 560776
rect 241020 560736 241026 560748
rect 376754 560736 376760 560748
rect 376812 560736 376818 560788
rect 235810 560668 235816 560720
rect 235868 560708 235874 560720
rect 396718 560708 396724 560720
rect 235868 560680 396724 560708
rect 235868 560668 235874 560680
rect 396718 560668 396724 560680
rect 396776 560668 396782 560720
rect 183002 560600 183008 560652
rect 183060 560640 183066 560652
rect 394050 560640 394056 560652
rect 183060 560612 394056 560640
rect 183060 560600 183066 560612
rect 394050 560600 394056 560612
rect 394108 560600 394114 560652
rect 116578 560532 116584 560584
rect 116636 560572 116642 560584
rect 358630 560572 358636 560584
rect 116636 560544 358636 560572
rect 116636 560532 116642 560544
rect 358630 560532 358636 560544
rect 358688 560532 358694 560584
rect 32766 560464 32772 560516
rect 32824 560504 32830 560516
rect 381814 560504 381820 560516
rect 32824 560476 381820 560504
rect 32824 560464 32830 560476
rect 381814 560464 381820 560476
rect 381872 560464 381878 560516
rect 39482 560396 39488 560448
rect 39540 560436 39546 560448
rect 395890 560436 395896 560448
rect 39540 560408 395896 560436
rect 39540 560396 39546 560408
rect 395890 560396 395896 560408
rect 395948 560396 395954 560448
rect 43530 560328 43536 560380
rect 43588 560368 43594 560380
rect 405090 560368 405096 560380
rect 43588 560340 405096 560368
rect 43588 560328 43594 560340
rect 405090 560328 405096 560340
rect 405148 560328 405154 560380
rect 553302 560328 553308 560380
rect 553360 560368 553366 560380
rect 566734 560368 566740 560380
rect 553360 560340 566740 560368
rect 553360 560328 553366 560340
rect 566734 560328 566740 560340
rect 566792 560328 566798 560380
rect 37826 560260 37832 560312
rect 37884 560300 37890 560312
rect 407390 560300 407396 560312
rect 37884 560272 407396 560300
rect 37884 560260 37890 560272
rect 407390 560260 407396 560272
rect 407448 560260 407454 560312
rect 553118 560260 553124 560312
rect 553176 560300 553182 560312
rect 568022 560300 568028 560312
rect 553176 560272 568028 560300
rect 553176 560260 553182 560272
rect 568022 560260 568028 560272
rect 568080 560260 568086 560312
rect 347590 560192 347596 560244
rect 347648 560232 347654 560244
rect 351270 560232 351276 560244
rect 347648 560204 351276 560232
rect 347648 560192 347654 560204
rect 351270 560192 351276 560204
rect 351328 560192 351334 560244
rect 52822 560028 52828 560040
rect 41386 560000 52828 560028
rect 39390 559580 39396 559632
rect 39448 559620 39454 559632
rect 41386 559620 41414 560000
rect 52822 559988 52828 560000
rect 52880 559988 52886 560040
rect 319162 559988 319168 560040
rect 319220 560028 319226 560040
rect 319220 560000 345014 560028
rect 319220 559988 319226 560000
rect 45738 559920 45744 559972
rect 45796 559960 45802 559972
rect 48866 559960 48872 559972
rect 45796 559932 48872 559960
rect 45796 559920 45802 559932
rect 48866 559920 48872 559932
rect 48924 559920 48930 559972
rect 51994 559920 52000 559972
rect 52052 559920 52058 559972
rect 148962 559960 148968 559972
rect 142126 559932 148968 559960
rect 39448 559592 41414 559620
rect 39448 559580 39454 559592
rect 36814 559512 36820 559564
rect 36872 559552 36878 559564
rect 52012 559552 52040 559920
rect 36872 559524 52040 559552
rect 36872 559512 36878 559524
rect 41046 558900 41052 558952
rect 41104 558940 41110 558952
rect 142126 558940 142154 559932
rect 148962 559920 148968 559932
rect 149020 559920 149026 559972
rect 327718 559920 327724 559972
rect 327776 559920 327782 559972
rect 336642 559920 336648 559972
rect 336700 559920 336706 559972
rect 340690 559920 340696 559972
rect 340748 559920 340754 559972
rect 327736 559008 327764 559920
rect 336660 559076 336688 559920
rect 340708 559484 340736 559920
rect 344986 559552 345014 560000
rect 347222 559920 347228 559972
rect 347280 559920 347286 559972
rect 347314 559920 347320 559972
rect 347372 559960 347378 559972
rect 347372 559932 354674 559960
rect 347372 559920 347378 559932
rect 347240 559892 347268 559920
rect 347240 559864 349844 559892
rect 349816 559620 349844 559864
rect 354646 559688 354674 559932
rect 389174 559688 389180 559700
rect 354646 559660 389180 559688
rect 389174 559648 389180 559660
rect 389232 559648 389238 559700
rect 407942 559620 407948 559632
rect 349816 559592 407948 559620
rect 407942 559580 407948 559592
rect 408000 559580 408006 559632
rect 407666 559552 407672 559564
rect 344986 559524 407672 559552
rect 407666 559512 407672 559524
rect 407724 559512 407730 559564
rect 349982 559484 349988 559496
rect 340708 559456 349988 559484
rect 349982 559444 349988 559456
rect 350040 559444 350046 559496
rect 364426 559076 364432 559088
rect 336660 559048 364432 559076
rect 364426 559036 364432 559048
rect 364484 559036 364490 559088
rect 356238 559008 356244 559020
rect 327736 558980 356244 559008
rect 356238 558968 356244 558980
rect 356296 558968 356302 559020
rect 41104 558912 142154 558940
rect 41104 558900 41110 558912
rect 349982 558900 349988 558952
rect 350040 558940 350046 558952
rect 380526 558940 380532 558952
rect 350040 558912 380532 558940
rect 350040 558900 350046 558912
rect 380526 558900 380532 558912
rect 380584 558900 380590 558952
rect 552934 557948 552940 558000
rect 552992 557988 552998 558000
rect 556614 557988 556620 558000
rect 552992 557960 556620 557988
rect 552992 557948 552998 557960
rect 556614 557948 556620 557960
rect 556672 557948 556678 558000
rect 553302 557540 553308 557592
rect 553360 557580 553366 557592
rect 568666 557580 568672 557592
rect 553360 557552 568672 557580
rect 553360 557540 553366 557552
rect 568666 557540 568672 557552
rect 568724 557540 568730 557592
rect 405274 557200 405280 557252
rect 405332 557240 405338 557252
rect 407666 557240 407672 557252
rect 405332 557212 407672 557240
rect 405332 557200 405338 557212
rect 407666 557200 407672 557212
rect 407724 557200 407730 557252
rect 553302 556520 553308 556572
rect 553360 556560 553366 556572
rect 559742 556560 559748 556572
rect 553360 556532 559748 556560
rect 553360 556520 553366 556532
rect 559742 556520 559748 556532
rect 559800 556520 559806 556572
rect 44542 556180 44548 556232
rect 44600 556220 44606 556232
rect 46106 556220 46112 556232
rect 44600 556192 46112 556220
rect 44600 556180 44606 556192
rect 46106 556180 46112 556192
rect 46164 556180 46170 556232
rect 394510 556180 394516 556232
rect 394568 556220 394574 556232
rect 407390 556220 407396 556232
rect 394568 556192 407396 556220
rect 394568 556180 394574 556192
rect 407390 556180 407396 556192
rect 407448 556180 407454 556232
rect 553302 556180 553308 556232
rect 553360 556220 553366 556232
rect 573542 556220 573548 556232
rect 553360 556192 573548 556220
rect 553360 556180 553366 556192
rect 573542 556180 573548 556192
rect 573600 556180 573606 556232
rect 350442 554684 350448 554736
rect 350500 554724 350506 554736
rect 353294 554724 353300 554736
rect 350500 554696 353300 554724
rect 350500 554684 350506 554696
rect 353294 554684 353300 554696
rect 353352 554684 353358 554736
rect 552014 553664 552020 553716
rect 552072 553704 552078 553716
rect 555142 553704 555148 553716
rect 552072 553676 555148 553704
rect 552072 553664 552078 553676
rect 555142 553664 555148 553676
rect 555200 553664 555206 553716
rect 407850 552644 407856 552696
rect 407908 552684 407914 552696
rect 408310 552684 408316 552696
rect 407908 552656 408316 552684
rect 407908 552644 407914 552656
rect 408310 552644 408316 552656
rect 408368 552644 408374 552696
rect 387610 552032 387616 552084
rect 387668 552072 387674 552084
rect 407482 552072 407488 552084
rect 387668 552044 407488 552072
rect 387668 552032 387674 552044
rect 407482 552032 407488 552044
rect 407540 552032 407546 552084
rect 351362 551964 351368 552016
rect 351420 552004 351426 552016
rect 407390 552004 407396 552016
rect 351420 551976 407396 552004
rect 351420 551964 351426 551976
rect 407390 551964 407396 551976
rect 407448 551964 407454 552016
rect 41782 551148 41788 551200
rect 41840 551188 41846 551200
rect 46106 551188 46112 551200
rect 41840 551160 46112 551188
rect 41840 551148 41846 551160
rect 46106 551148 46112 551160
rect 46164 551148 46170 551200
rect 350442 551080 350448 551132
rect 350500 551120 350506 551132
rect 356790 551120 356796 551132
rect 350500 551092 356796 551120
rect 350500 551080 350506 551092
rect 356790 551080 356796 551092
rect 356848 551080 356854 551132
rect 42334 550808 42340 550860
rect 42392 550848 42398 550860
rect 46106 550848 46112 550860
rect 42392 550820 46112 550848
rect 42392 550808 42398 550820
rect 46106 550808 46112 550820
rect 46164 550808 46170 550860
rect 552014 550808 552020 550860
rect 552072 550848 552078 550860
rect 555234 550848 555240 550860
rect 552072 550820 555240 550848
rect 552072 550808 552078 550820
rect 555234 550808 555240 550820
rect 555292 550808 555298 550860
rect 404170 550604 404176 550656
rect 404228 550644 404234 550656
rect 407390 550644 407396 550656
rect 404228 550616 407396 550644
rect 404228 550604 404234 550616
rect 407390 550604 407396 550616
rect 407448 550604 407454 550656
rect 553302 550604 553308 550656
rect 553360 550644 553366 550656
rect 562594 550644 562600 550656
rect 553360 550616 562600 550644
rect 553360 550604 553366 550616
rect 562594 550604 562600 550616
rect 562652 550604 562658 550656
rect 30190 549244 30196 549296
rect 30248 549284 30254 549296
rect 46106 549284 46112 549296
rect 30248 549256 46112 549284
rect 30248 549244 30254 549256
rect 46106 549244 46112 549256
rect 46164 549244 46170 549296
rect 358446 549244 358452 549296
rect 358504 549284 358510 549296
rect 407390 549284 407396 549296
rect 358504 549256 407396 549284
rect 358504 549244 358510 549256
rect 407390 549244 407396 549256
rect 407448 549244 407454 549296
rect 553302 549244 553308 549296
rect 553360 549284 553366 549296
rect 574186 549284 574192 549296
rect 553360 549256 574192 549284
rect 553360 549244 553366 549256
rect 574186 549244 574192 549256
rect 574244 549244 574250 549296
rect 350166 549176 350172 549228
rect 350224 549216 350230 549228
rect 352098 549216 352104 549228
rect 350224 549188 352104 549216
rect 350224 549176 350230 549188
rect 352098 549176 352104 549188
rect 352156 549176 352162 549228
rect 405182 549176 405188 549228
rect 405240 549216 405246 549228
rect 407482 549216 407488 549228
rect 405240 549188 407488 549216
rect 405240 549176 405246 549188
rect 407482 549176 407488 549188
rect 407540 549176 407546 549228
rect 30282 547884 30288 547936
rect 30340 547924 30346 547936
rect 46106 547924 46112 547936
rect 30340 547896 46112 547924
rect 30340 547884 30346 547896
rect 46106 547884 46112 547896
rect 46164 547884 46170 547936
rect 350442 546592 350448 546644
rect 350500 546632 350506 546644
rect 384298 546632 384304 546644
rect 350500 546604 384304 546632
rect 350500 546592 350506 546604
rect 384298 546592 384304 546604
rect 384356 546592 384362 546644
rect 371878 546524 371884 546576
rect 371936 546564 371942 546576
rect 407390 546564 407396 546576
rect 371936 546536 407396 546564
rect 371936 546524 371942 546536
rect 407390 546524 407396 546536
rect 407448 546524 407454 546576
rect 350258 546456 350264 546508
rect 350316 546496 350322 546508
rect 385954 546496 385960 546508
rect 350316 546468 385960 546496
rect 350316 546456 350322 546468
rect 385954 546456 385960 546468
rect 386012 546456 386018 546508
rect 551370 546456 551376 546508
rect 551428 546496 551434 546508
rect 552014 546496 552020 546508
rect 551428 546468 552020 546496
rect 551428 546456 551434 546468
rect 552014 546456 552020 546468
rect 552072 546456 552078 546508
rect 46106 545980 46112 546032
rect 46164 546020 46170 546032
rect 46750 546020 46756 546032
rect 46164 545992 46756 546020
rect 46164 545980 46170 545992
rect 46750 545980 46756 545992
rect 46808 545980 46814 546032
rect 34330 545096 34336 545148
rect 34388 545136 34394 545148
rect 46750 545136 46756 545148
rect 34388 545108 46756 545136
rect 34388 545096 34394 545108
rect 46750 545096 46756 545108
rect 46808 545096 46814 545148
rect 405182 543804 405188 543856
rect 405240 543844 405246 543856
rect 407482 543844 407488 543856
rect 405240 543816 407488 543844
rect 405240 543804 405246 543816
rect 407482 543804 407488 543816
rect 407540 543804 407546 543856
rect 552566 543804 552572 543856
rect 552624 543844 552630 543856
rect 555142 543844 555148 543856
rect 552624 543816 555148 543844
rect 552624 543804 552630 543816
rect 555142 543804 555148 543816
rect 555200 543804 555206 543856
rect 43070 543736 43076 543788
rect 43128 543776 43134 543788
rect 46750 543776 46756 543788
rect 43128 543748 46756 543776
rect 43128 543736 43134 543748
rect 46750 543736 46756 543748
rect 46808 543736 46814 543788
rect 389818 543736 389824 543788
rect 389876 543776 389882 543788
rect 407390 543776 407396 543788
rect 389876 543748 407396 543776
rect 389876 543736 389882 543748
rect 407390 543736 407396 543748
rect 407448 543736 407454 543788
rect 350442 542376 350448 542428
rect 350500 542416 350506 542428
rect 398374 542416 398380 542428
rect 350500 542388 398380 542416
rect 350500 542376 350506 542388
rect 398374 542376 398380 542388
rect 398432 542376 398438 542428
rect 354030 542308 354036 542360
rect 354088 542348 354094 542360
rect 407390 542348 407396 542360
rect 354088 542320 407396 542348
rect 354088 542308 354094 542320
rect 407390 542308 407396 542320
rect 407448 542308 407454 542360
rect 22002 540948 22008 541000
rect 22060 540988 22066 541000
rect 46750 540988 46756 541000
rect 22060 540960 46756 540988
rect 22060 540948 22066 540960
rect 46750 540948 46756 540960
rect 46808 540948 46814 541000
rect 553302 539656 553308 539708
rect 553360 539696 553366 539708
rect 562226 539696 562232 539708
rect 553360 539668 562232 539696
rect 553360 539656 553366 539668
rect 562226 539656 562232 539668
rect 562284 539656 562290 539708
rect 553118 539588 553124 539640
rect 553176 539628 553182 539640
rect 567286 539628 567292 539640
rect 553176 539600 567292 539628
rect 553176 539588 553182 539600
rect 567286 539588 567292 539600
rect 567344 539588 567350 539640
rect 350442 538228 350448 538280
rect 350500 538268 350506 538280
rect 365162 538268 365168 538280
rect 350500 538240 365168 538268
rect 350500 538228 350506 538240
rect 365162 538228 365168 538240
rect 365220 538228 365226 538280
rect 43438 538160 43444 538212
rect 43496 538200 43502 538212
rect 46750 538200 46756 538212
rect 43496 538172 46756 538200
rect 43496 538160 43502 538172
rect 46750 538160 46756 538172
rect 46808 538160 46814 538212
rect 350442 536800 350448 536852
rect 350500 536840 350506 536852
rect 386414 536840 386420 536852
rect 350500 536812 386420 536840
rect 350500 536800 350506 536812
rect 386414 536800 386420 536812
rect 386472 536800 386478 536852
rect 553302 535440 553308 535492
rect 553360 535480 553366 535492
rect 560754 535480 560760 535492
rect 553360 535452 560760 535480
rect 553360 535440 553366 535452
rect 560754 535440 560760 535452
rect 560812 535440 560818 535492
rect 350442 534080 350448 534132
rect 350500 534120 350506 534132
rect 362218 534120 362224 534132
rect 350500 534092 362224 534120
rect 350500 534080 350506 534092
rect 362218 534080 362224 534092
rect 362276 534080 362282 534132
rect 391290 534080 391296 534132
rect 391348 534120 391354 534132
rect 407298 534120 407304 534132
rect 391348 534092 407304 534120
rect 391348 534080 391354 534092
rect 407298 534080 407304 534092
rect 407356 534080 407362 534132
rect 553302 534080 553308 534132
rect 553360 534120 553366 534132
rect 581454 534120 581460 534132
rect 553360 534092 581460 534120
rect 553360 534080 553366 534092
rect 581454 534080 581460 534092
rect 581512 534080 581518 534132
rect 350258 532788 350264 532840
rect 350316 532828 350322 532840
rect 358906 532828 358912 532840
rect 350316 532800 358912 532828
rect 350316 532788 350322 532800
rect 358906 532788 358912 532800
rect 358964 532788 358970 532840
rect 27430 532720 27436 532772
rect 27488 532760 27494 532772
rect 46750 532760 46756 532772
rect 27488 532732 46756 532760
rect 27488 532720 27494 532732
rect 46750 532720 46756 532732
rect 46808 532720 46814 532772
rect 350442 532720 350448 532772
rect 350500 532760 350506 532772
rect 386138 532760 386144 532772
rect 350500 532732 386144 532760
rect 350500 532720 350506 532732
rect 386138 532720 386144 532732
rect 386196 532720 386202 532772
rect 395706 532720 395712 532772
rect 395764 532760 395770 532772
rect 407298 532760 407304 532772
rect 395764 532732 407304 532760
rect 395764 532720 395770 532732
rect 407298 532720 407304 532732
rect 407356 532720 407362 532772
rect 552382 532516 552388 532568
rect 552440 532556 552446 532568
rect 553670 532556 553676 532568
rect 552440 532528 553676 532556
rect 552440 532516 552446 532528
rect 553670 532516 553676 532528
rect 553728 532516 553734 532568
rect 25866 531292 25872 531344
rect 25924 531332 25930 531344
rect 46750 531332 46756 531344
rect 25924 531304 46756 531332
rect 25924 531292 25930 531304
rect 46750 531292 46756 531304
rect 46808 531292 46814 531344
rect 350442 531292 350448 531344
rect 350500 531332 350506 531344
rect 353662 531332 353668 531344
rect 350500 531304 353668 531332
rect 350500 531292 350506 531304
rect 353662 531292 353668 531304
rect 353720 531292 353726 531344
rect 401318 531292 401324 531344
rect 401376 531332 401382 531344
rect 407298 531332 407304 531344
rect 401376 531304 407304 531332
rect 401376 531292 401382 531304
rect 407298 531292 407304 531304
rect 407356 531292 407362 531344
rect 552382 530476 552388 530528
rect 552440 530516 552446 530528
rect 553762 530516 553768 530528
rect 552440 530488 553768 530516
rect 552440 530476 552446 530488
rect 553762 530476 553768 530488
rect 553820 530476 553826 530528
rect 553302 530272 553308 530324
rect 553360 530312 553366 530324
rect 557994 530312 558000 530324
rect 553360 530284 558000 530312
rect 553360 530272 553366 530284
rect 557994 530272 558000 530284
rect 558052 530272 558058 530324
rect 18966 529932 18972 529984
rect 19024 529972 19030 529984
rect 46750 529972 46756 529984
rect 19024 529944 46756 529972
rect 19024 529932 19030 529944
rect 46750 529932 46756 529944
rect 46808 529932 46814 529984
rect 350442 529932 350448 529984
rect 350500 529972 350506 529984
rect 380434 529972 380440 529984
rect 350500 529944 380440 529972
rect 350500 529932 350506 529944
rect 380434 529932 380440 529944
rect 380492 529932 380498 529984
rect 40402 528572 40408 528624
rect 40460 528612 40466 528624
rect 46106 528612 46112 528624
rect 40460 528584 46112 528612
rect 40460 528572 40466 528584
rect 46106 528572 46112 528584
rect 46164 528572 46170 528624
rect 350442 527144 350448 527196
rect 350500 527184 350506 527196
rect 366450 527184 366456 527196
rect 350500 527156 366456 527184
rect 350500 527144 350506 527156
rect 366450 527144 366456 527156
rect 366508 527144 366514 527196
rect 553302 527144 553308 527196
rect 553360 527184 553366 527196
rect 566274 527184 566280 527196
rect 553360 527156 566280 527184
rect 553360 527144 553366 527156
rect 566274 527144 566280 527156
rect 566332 527144 566338 527196
rect 407114 526464 407120 526516
rect 407172 526504 407178 526516
rect 407298 526504 407304 526516
rect 407172 526476 407304 526504
rect 407172 526464 407178 526476
rect 407298 526464 407304 526476
rect 407356 526464 407362 526516
rect 552382 526260 552388 526312
rect 552440 526300 552446 526312
rect 553762 526300 553768 526312
rect 552440 526272 553768 526300
rect 552440 526260 552446 526272
rect 553762 526260 553768 526272
rect 553820 526260 553826 526312
rect 350442 525920 350448 525972
rect 350500 525960 350506 525972
rect 356882 525960 356888 525972
rect 350500 525932 356888 525960
rect 350500 525920 350506 525932
rect 356882 525920 356888 525932
rect 356940 525920 356946 525972
rect 400122 525784 400128 525836
rect 400180 525824 400186 525836
rect 407298 525824 407304 525836
rect 400180 525796 407304 525824
rect 400180 525784 400186 525796
rect 407298 525784 407304 525796
rect 407356 525784 407362 525836
rect 44082 525716 44088 525768
rect 44140 525756 44146 525768
rect 46750 525756 46756 525768
rect 44140 525728 46756 525756
rect 44140 525716 44146 525728
rect 46750 525716 46756 525728
rect 46808 525716 46814 525768
rect 570690 525716 570696 525768
rect 570748 525756 570754 525768
rect 580166 525756 580172 525768
rect 570748 525728 580172 525756
rect 570748 525716 570754 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 46014 524424 46020 524476
rect 46072 524464 46078 524476
rect 47578 524464 47584 524476
rect 46072 524436 47584 524464
rect 46072 524424 46078 524436
rect 47578 524424 47584 524436
rect 47636 524424 47642 524476
rect 395982 524424 395988 524476
rect 396040 524464 396046 524476
rect 407114 524464 407120 524476
rect 396040 524436 407120 524464
rect 396040 524424 396046 524436
rect 407114 524424 407120 524436
rect 407172 524424 407178 524476
rect 350258 524356 350264 524408
rect 350316 524396 350322 524408
rect 353754 524396 353760 524408
rect 350316 524368 353760 524396
rect 350316 524356 350322 524368
rect 353754 524356 353760 524368
rect 353812 524356 353818 524408
rect 350442 522996 350448 523048
rect 350500 523036 350506 523048
rect 369394 523036 369400 523048
rect 350500 523008 369400 523036
rect 350500 522996 350506 523008
rect 369394 522996 369400 523008
rect 369452 522996 369458 523048
rect 385862 522996 385868 523048
rect 385920 523036 385926 523048
rect 407298 523036 407304 523048
rect 385920 523008 407304 523036
rect 385920 522996 385926 523008
rect 407298 522996 407304 523008
rect 407356 522996 407362 523048
rect 383010 522928 383016 522980
rect 383068 522968 383074 522980
rect 407114 522968 407120 522980
rect 383068 522940 407120 522968
rect 383068 522928 383074 522940
rect 407114 522928 407120 522940
rect 407172 522928 407178 522980
rect 407482 522928 407488 522980
rect 407540 522968 407546 522980
rect 409138 522968 409144 522980
rect 407540 522940 409144 522968
rect 407540 522928 407546 522940
rect 409138 522928 409144 522940
rect 409196 522928 409202 522980
rect 402698 521636 402704 521688
rect 402756 521676 402762 521688
rect 407390 521676 407396 521688
rect 402756 521648 407396 521676
rect 402756 521636 402762 521648
rect 407390 521636 407396 521648
rect 407448 521636 407454 521688
rect 40954 521500 40960 521552
rect 41012 521540 41018 521552
rect 46290 521540 46296 521552
rect 41012 521512 46296 521540
rect 41012 521500 41018 521512
rect 46290 521500 46296 521512
rect 46348 521500 46354 521552
rect 23290 520344 23296 520396
rect 23348 520384 23354 520396
rect 45554 520384 45560 520396
rect 23348 520356 45560 520384
rect 23348 520344 23354 520356
rect 45554 520344 45560 520356
rect 45612 520344 45618 520396
rect 17862 520276 17868 520328
rect 17920 520316 17926 520328
rect 45646 520316 45652 520328
rect 17920 520288 45652 520316
rect 17920 520276 17926 520288
rect 45646 520276 45652 520288
rect 45704 520276 45710 520328
rect 350166 520276 350172 520328
rect 350224 520316 350230 520328
rect 352098 520316 352104 520328
rect 350224 520288 352104 520316
rect 350224 520276 350230 520288
rect 352098 520276 352104 520288
rect 352156 520276 352162 520328
rect 552014 520276 552020 520328
rect 552072 520316 552078 520328
rect 571518 520316 571524 520328
rect 552072 520288 571524 520316
rect 552072 520276 552078 520288
rect 571518 520276 571524 520288
rect 571576 520276 571582 520328
rect 45830 519528 45836 519580
rect 45888 519568 45894 519580
rect 46014 519568 46020 519580
rect 45888 519540 46020 519568
rect 45888 519528 45894 519540
rect 46014 519528 46020 519540
rect 46072 519528 46078 519580
rect 552014 519256 552020 519308
rect 552072 519296 552078 519308
rect 553670 519296 553676 519308
rect 552072 519268 553676 519296
rect 552072 519256 552078 519268
rect 553670 519256 553676 519268
rect 553728 519256 553734 519308
rect 552014 518984 552020 519036
rect 552072 519024 552078 519036
rect 564710 519024 564716 519036
rect 552072 518996 564716 519024
rect 552072 518984 552078 518996
rect 564710 518984 564716 518996
rect 564768 518984 564774 519036
rect 350442 517556 350448 517608
rect 350500 517596 350506 517608
rect 381630 517596 381636 517608
rect 350500 517568 381636 517596
rect 350500 517556 350506 517568
rect 381630 517556 381636 517568
rect 381688 517556 381694 517608
rect 388254 517556 388260 517608
rect 388312 517596 388318 517608
rect 407114 517596 407120 517608
rect 388312 517568 407120 517596
rect 388312 517556 388318 517568
rect 407114 517556 407120 517568
rect 407172 517556 407178 517608
rect 373442 517488 373448 517540
rect 373500 517528 373506 517540
rect 407298 517528 407304 517540
rect 373500 517500 407304 517528
rect 373500 517488 373506 517500
rect 407298 517488 407304 517500
rect 407356 517488 407362 517540
rect 350258 516196 350264 516248
rect 350316 516236 350322 516248
rect 387150 516236 387156 516248
rect 350316 516208 387156 516236
rect 350316 516196 350322 516208
rect 387150 516196 387156 516208
rect 387208 516196 387214 516248
rect 397362 516196 397368 516248
rect 397420 516236 397426 516248
rect 407114 516236 407120 516248
rect 397420 516208 407120 516236
rect 397420 516196 397426 516208
rect 407114 516196 407120 516208
rect 407172 516196 407178 516248
rect 34238 516128 34244 516180
rect 34296 516168 34302 516180
rect 45554 516168 45560 516180
rect 34296 516140 45560 516168
rect 34296 516128 34302 516140
rect 45554 516128 45560 516140
rect 45612 516128 45618 516180
rect 350442 516128 350448 516180
rect 350500 516168 350506 516180
rect 361850 516168 361856 516180
rect 350500 516140 361856 516168
rect 350500 516128 350506 516140
rect 361850 516128 361856 516140
rect 361908 516128 361914 516180
rect 370498 516128 370504 516180
rect 370556 516168 370562 516180
rect 407298 516168 407304 516180
rect 370556 516140 407304 516168
rect 370556 516128 370562 516140
rect 407298 516128 407304 516140
rect 407356 516128 407362 516180
rect 552014 516128 552020 516180
rect 552072 516168 552078 516180
rect 570782 516168 570788 516180
rect 552072 516140 570788 516168
rect 552072 516128 552078 516140
rect 570782 516128 570788 516140
rect 570840 516128 570846 516180
rect 405090 516060 405096 516112
rect 405148 516100 405154 516112
rect 407574 516100 407580 516112
rect 405148 516072 407580 516100
rect 405148 516060 405154 516072
rect 407574 516060 407580 516072
rect 407632 516060 407638 516112
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 26970 514808 26976 514820
rect 3476 514780 26976 514808
rect 3476 514768 3482 514780
rect 26970 514768 26976 514780
rect 27028 514768 27034 514820
rect 38562 514768 38568 514820
rect 38620 514808 38626 514820
rect 45554 514808 45560 514820
rect 38620 514780 45560 514808
rect 38620 514768 38626 514780
rect 45554 514768 45560 514780
rect 45612 514768 45618 514820
rect 552014 514768 552020 514820
rect 552072 514808 552078 514820
rect 564802 514808 564808 514820
rect 552072 514780 564808 514808
rect 552072 514768 552078 514780
rect 564802 514768 564808 514780
rect 564860 514768 564866 514820
rect 45830 514020 45836 514072
rect 45888 514060 45894 514072
rect 46106 514060 46112 514072
rect 45888 514032 46112 514060
rect 45888 514020 45894 514032
rect 46106 514020 46112 514032
rect 46164 514020 46170 514072
rect 350258 513408 350264 513460
rect 350316 513448 350322 513460
rect 353754 513448 353760 513460
rect 350316 513420 353760 513448
rect 350316 513408 350322 513420
rect 353754 513408 353760 513420
rect 353812 513408 353818 513460
rect 38010 513340 38016 513392
rect 38068 513380 38074 513392
rect 46198 513380 46204 513392
rect 38068 513352 46204 513380
rect 38068 513340 38074 513352
rect 46198 513340 46204 513352
rect 46256 513340 46262 513392
rect 350442 513340 350448 513392
rect 350500 513380 350506 513392
rect 394142 513380 394148 513392
rect 350500 513352 394148 513380
rect 350500 513340 350506 513352
rect 394142 513340 394148 513352
rect 394200 513340 394206 513392
rect 389910 513272 389916 513324
rect 389968 513312 389974 513324
rect 407114 513312 407120 513324
rect 389968 513284 407120 513312
rect 389968 513272 389974 513284
rect 407114 513272 407120 513284
rect 407172 513272 407178 513324
rect 377674 511980 377680 512032
rect 377732 512020 377738 512032
rect 407114 512020 407120 512032
rect 377732 511992 407120 512020
rect 377732 511980 377738 511992
rect 407114 511980 407120 511992
rect 407172 511980 407178 512032
rect 39850 510552 39856 510604
rect 39908 510592 39914 510604
rect 46750 510592 46756 510604
rect 39908 510564 46756 510592
rect 39908 510552 39914 510564
rect 46750 510552 46756 510564
rect 46808 510552 46814 510604
rect 553302 509600 553308 509652
rect 553360 509640 553366 509652
rect 559834 509640 559840 509652
rect 553360 509612 559840 509640
rect 553360 509600 553366 509612
rect 559834 509600 559840 509612
rect 559892 509600 559898 509652
rect 44910 509260 44916 509312
rect 44968 509300 44974 509312
rect 46198 509300 46204 509312
rect 44968 509272 46204 509300
rect 44968 509260 44974 509272
rect 46198 509260 46204 509272
rect 46256 509260 46262 509312
rect 389910 509260 389916 509312
rect 389968 509300 389974 509312
rect 407114 509300 407120 509312
rect 389968 509272 407120 509300
rect 389968 509260 389974 509272
rect 407114 509260 407120 509272
rect 407172 509260 407178 509312
rect 350442 509192 350448 509244
rect 350500 509232 350506 509244
rect 406378 509232 406384 509244
rect 350500 509204 406384 509232
rect 350500 509192 350506 509204
rect 406378 509192 406384 509204
rect 406436 509192 406442 509244
rect 40678 508308 40684 508360
rect 40736 508348 40742 508360
rect 44910 508348 44916 508360
rect 40736 508320 44916 508348
rect 40736 508308 40742 508320
rect 44910 508308 44916 508320
rect 44968 508308 44974 508360
rect 350442 506472 350448 506524
rect 350500 506512 350506 506524
rect 375374 506512 375380 506524
rect 350500 506484 375380 506512
rect 350500 506472 350506 506484
rect 375374 506472 375380 506484
rect 375432 506472 375438 506524
rect 350258 506404 350264 506456
rect 350316 506444 350322 506456
rect 399570 506444 399576 506456
rect 350316 506416 399576 506444
rect 350316 506404 350322 506416
rect 399570 506404 399576 506416
rect 399628 506404 399634 506456
rect 553302 506404 553308 506456
rect 553360 506444 553366 506456
rect 570598 506444 570604 506456
rect 553360 506416 570604 506444
rect 553360 506404 553366 506416
rect 570598 506404 570604 506416
rect 570656 506404 570662 506456
rect 19150 505112 19156 505164
rect 19208 505152 19214 505164
rect 46750 505152 46756 505164
rect 19208 505124 46756 505152
rect 19208 505112 19214 505124
rect 46750 505112 46756 505124
rect 46808 505112 46814 505164
rect 350442 505112 350448 505164
rect 350500 505152 350506 505164
rect 383102 505152 383108 505164
rect 350500 505124 383108 505152
rect 350500 505112 350506 505124
rect 383102 505112 383108 505124
rect 383160 505112 383166 505164
rect 350442 503684 350448 503736
rect 350500 503724 350506 503736
rect 360286 503724 360292 503736
rect 350500 503696 360292 503724
rect 350500 503684 350506 503696
rect 360286 503684 360292 503696
rect 360344 503684 360350 503736
rect 553302 503684 553308 503736
rect 553360 503724 553366 503736
rect 574554 503724 574560 503736
rect 553360 503696 574560 503724
rect 553360 503684 553366 503696
rect 574554 503684 574560 503696
rect 574612 503684 574618 503736
rect 553302 502392 553308 502444
rect 553360 502432 553366 502444
rect 557718 502432 557724 502444
rect 553360 502404 557724 502432
rect 553360 502392 553366 502404
rect 557718 502392 557724 502404
rect 557776 502392 557782 502444
rect 39942 502052 39948 502104
rect 40000 502092 40006 502104
rect 45830 502092 45836 502104
rect 40000 502064 45836 502092
rect 40000 502052 40006 502064
rect 45830 502052 45836 502064
rect 45888 502052 45894 502104
rect 553302 501304 553308 501356
rect 553360 501344 553366 501356
rect 559190 501344 559196 501356
rect 553360 501316 559196 501344
rect 553360 501304 553366 501316
rect 559190 501304 559196 501316
rect 559248 501304 559254 501356
rect 553302 500964 553308 501016
rect 553360 501004 553366 501016
rect 574922 501004 574928 501016
rect 553360 500976 574928 501004
rect 553360 500964 553366 500976
rect 574922 500964 574928 500976
rect 574980 500964 574986 501016
rect 40862 500896 40868 500948
rect 40920 500936 40926 500948
rect 46750 500936 46756 500948
rect 40920 500908 46756 500936
rect 40920 500896 40926 500908
rect 46750 500896 46756 500908
rect 46808 500896 46814 500948
rect 402422 500896 402428 500948
rect 402480 500936 402486 500948
rect 407114 500936 407120 500948
rect 402480 500908 407120 500936
rect 402480 500896 402486 500908
rect 407114 500896 407120 500908
rect 407172 500896 407178 500948
rect 553302 499808 553308 499860
rect 553360 499848 553366 499860
rect 557626 499848 557632 499860
rect 553360 499820 557632 499848
rect 553360 499808 553366 499820
rect 557626 499808 557632 499820
rect 557684 499808 557690 499860
rect 350442 499536 350448 499588
rect 350500 499576 350506 499588
rect 384758 499576 384764 499588
rect 350500 499548 384764 499576
rect 350500 499536 350506 499548
rect 384758 499536 384764 499548
rect 384816 499536 384822 499588
rect 553302 498448 553308 498500
rect 553360 498488 553366 498500
rect 557534 498488 557540 498500
rect 553360 498460 557540 498488
rect 553360 498448 553366 498460
rect 557534 498448 557540 498460
rect 557592 498448 557598 498500
rect 350442 498176 350448 498228
rect 350500 498216 350506 498228
rect 354030 498216 354036 498228
rect 350500 498188 354036 498216
rect 350500 498176 350506 498188
rect 354030 498176 354036 498188
rect 354088 498176 354094 498228
rect 42518 498108 42524 498160
rect 42576 498148 42582 498160
rect 45830 498148 45836 498160
rect 42576 498120 45836 498148
rect 42576 498108 42582 498120
rect 45830 498108 45836 498120
rect 45888 498108 45894 498160
rect 46014 497020 46020 497072
rect 46072 497060 46078 497072
rect 46382 497060 46388 497072
rect 46072 497032 46388 497060
rect 46072 497020 46078 497032
rect 46382 497020 46388 497032
rect 46440 497020 46446 497072
rect 384482 496816 384488 496868
rect 384540 496856 384546 496868
rect 407114 496856 407120 496868
rect 384540 496828 407120 496856
rect 384540 496816 384546 496828
rect 407114 496816 407120 496828
rect 407172 496816 407178 496868
rect 40770 496748 40776 496800
rect 40828 496788 40834 496800
rect 46750 496788 46756 496800
rect 40828 496760 46756 496788
rect 40828 496748 40834 496760
rect 46750 496748 46756 496760
rect 46808 496748 46814 496800
rect 39114 495456 39120 495508
rect 39172 495496 39178 495508
rect 46382 495496 46388 495508
rect 39172 495468 46388 495496
rect 39172 495456 39178 495468
rect 46382 495456 46388 495468
rect 46440 495456 46446 495508
rect 350442 495456 350448 495508
rect 350500 495496 350506 495508
rect 386046 495496 386052 495508
rect 350500 495468 386052 495496
rect 350500 495456 350506 495468
rect 386046 495456 386052 495468
rect 386104 495456 386110 495508
rect 401134 495456 401140 495508
rect 401192 495496 401198 495508
rect 407114 495496 407120 495508
rect 401192 495468 407120 495496
rect 401192 495456 401198 495468
rect 407114 495456 407120 495468
rect 407172 495456 407178 495508
rect 41966 495388 41972 495440
rect 42024 495428 42030 495440
rect 46750 495428 46756 495440
rect 42024 495400 46756 495428
rect 42024 495388 42030 495400
rect 46750 495388 46756 495400
rect 46808 495388 46814 495440
rect 350442 493416 350448 493468
rect 350500 493456 350506 493468
rect 351270 493456 351276 493468
rect 350500 493428 351276 493456
rect 350500 493416 350506 493428
rect 351270 493416 351276 493428
rect 351328 493416 351334 493468
rect 23198 492668 23204 492720
rect 23256 492708 23262 492720
rect 46750 492708 46756 492720
rect 23256 492680 46756 492708
rect 23256 492668 23262 492680
rect 46750 492668 46756 492680
rect 46808 492668 46814 492720
rect 384390 492668 384396 492720
rect 384448 492708 384454 492720
rect 407114 492708 407120 492720
rect 384448 492680 407120 492708
rect 384448 492668 384454 492680
rect 407114 492668 407120 492680
rect 407172 492668 407178 492720
rect 552658 492668 552664 492720
rect 552716 492708 552722 492720
rect 563790 492708 563796 492720
rect 552716 492680 563796 492708
rect 552716 492668 552722 492680
rect 563790 492668 563796 492680
rect 563848 492668 563854 492720
rect 350258 491376 350264 491428
rect 350316 491416 350322 491428
rect 359090 491416 359096 491428
rect 350316 491388 359096 491416
rect 350316 491376 350322 491388
rect 359090 491376 359096 491388
rect 359148 491376 359154 491428
rect 350442 491308 350448 491360
rect 350500 491348 350506 491360
rect 367922 491348 367928 491360
rect 350500 491320 367928 491348
rect 350500 491308 350506 491320
rect 367922 491308 367928 491320
rect 367980 491308 367986 491360
rect 40862 489948 40868 490000
rect 40920 489988 40926 490000
rect 46750 489988 46756 490000
rect 40920 489960 46756 489988
rect 40920 489948 40926 489960
rect 46750 489948 46756 489960
rect 46808 489948 46814 490000
rect 350442 489948 350448 490000
rect 350500 489988 350506 490000
rect 379514 489988 379520 490000
rect 350500 489960 379520 489988
rect 350500 489948 350506 489960
rect 379514 489948 379520 489960
rect 379572 489948 379578 490000
rect 381906 489948 381912 490000
rect 381964 489988 381970 490000
rect 407114 489988 407120 490000
rect 381964 489960 407120 489988
rect 381964 489948 381970 489960
rect 407114 489948 407120 489960
rect 407172 489948 407178 490000
rect 28626 489880 28632 489932
rect 28684 489920 28690 489932
rect 46382 489920 46388 489932
rect 28684 489892 46388 489920
rect 28684 489880 28690 489892
rect 46382 489880 46388 489892
rect 46440 489880 46446 489932
rect 350258 489880 350264 489932
rect 350316 489920 350322 489932
rect 392762 489920 392768 489932
rect 350316 489892 392768 489920
rect 350316 489880 350322 489892
rect 392762 489880 392768 489892
rect 392820 489880 392826 489932
rect 42610 489812 42616 489864
rect 42668 489852 42674 489864
rect 46750 489852 46756 489864
rect 42668 489824 46756 489852
rect 42668 489812 42674 489824
rect 46750 489812 46756 489824
rect 46808 489812 46814 489864
rect 350166 489812 350172 489864
rect 350224 489852 350230 489864
rect 352282 489852 352288 489864
rect 350224 489824 352288 489852
rect 350224 489812 350230 489824
rect 352282 489812 352288 489824
rect 352340 489812 352346 489864
rect 553302 488860 553308 488912
rect 553360 488900 553366 488912
rect 559098 488900 559104 488912
rect 553360 488872 559104 488900
rect 553360 488860 553366 488872
rect 559098 488860 559104 488872
rect 559156 488860 559162 488912
rect 393038 488588 393044 488640
rect 393096 488628 393102 488640
rect 407298 488628 407304 488640
rect 393096 488600 407304 488628
rect 393096 488588 393102 488600
rect 407298 488588 407304 488600
rect 407356 488588 407362 488640
rect 384574 488520 384580 488572
rect 384632 488560 384638 488572
rect 407114 488560 407120 488572
rect 384632 488532 407120 488560
rect 384632 488520 384638 488532
rect 407114 488520 407120 488532
rect 407172 488520 407178 488572
rect 350258 488452 350264 488504
rect 350316 488492 350322 488504
rect 372062 488492 372068 488504
rect 350316 488464 372068 488492
rect 350316 488452 350322 488464
rect 372062 488452 372068 488464
rect 372120 488452 372126 488504
rect 44634 488180 44640 488232
rect 44692 488220 44698 488232
rect 46382 488220 46388 488232
rect 44692 488192 46388 488220
rect 44692 488180 44698 488192
rect 46382 488180 46388 488192
rect 46440 488180 46446 488232
rect 401226 487160 401232 487212
rect 401284 487200 401290 487212
rect 407114 487200 407120 487212
rect 401284 487172 407120 487200
rect 401284 487160 401290 487172
rect 407114 487160 407120 487172
rect 407172 487160 407178 487212
rect 553302 487160 553308 487212
rect 553360 487200 553366 487212
rect 572898 487200 572904 487212
rect 553360 487172 572904 487200
rect 553360 487160 553366 487172
rect 572898 487160 572904 487172
rect 572956 487160 572962 487212
rect 39850 485800 39856 485852
rect 39908 485840 39914 485852
rect 46750 485840 46756 485852
rect 39908 485812 46756 485840
rect 39908 485800 39914 485812
rect 46750 485800 46756 485812
rect 46808 485800 46814 485852
rect 394326 485800 394332 485852
rect 394384 485840 394390 485852
rect 407114 485840 407120 485852
rect 394384 485812 407120 485840
rect 394384 485800 394390 485812
rect 407114 485800 407120 485812
rect 407172 485800 407178 485852
rect 21634 484372 21640 484424
rect 21692 484412 21698 484424
rect 46750 484412 46756 484424
rect 21692 484384 46756 484412
rect 21692 484372 21698 484384
rect 46750 484372 46756 484384
rect 46808 484372 46814 484424
rect 349982 484372 349988 484424
rect 350040 484412 350046 484424
rect 352282 484412 352288 484424
rect 350040 484384 352288 484412
rect 350040 484372 350046 484384
rect 352282 484372 352288 484384
rect 352340 484372 352346 484424
rect 373534 484372 373540 484424
rect 373592 484412 373598 484424
rect 407114 484412 407120 484424
rect 373592 484384 407120 484412
rect 373592 484372 373598 484384
rect 407114 484372 407120 484384
rect 407172 484372 407178 484424
rect 387426 483080 387432 483132
rect 387484 483120 387490 483132
rect 407114 483120 407120 483132
rect 387484 483092 407120 483120
rect 387484 483080 387490 483092
rect 407114 483080 407120 483092
rect 407172 483080 407178 483132
rect 19058 483012 19064 483064
rect 19116 483052 19122 483064
rect 46750 483052 46756 483064
rect 19116 483024 46756 483052
rect 19116 483012 19122 483024
rect 46750 483012 46756 483024
rect 46808 483012 46814 483064
rect 350258 483012 350264 483064
rect 350316 483052 350322 483064
rect 377766 483052 377772 483064
rect 350316 483024 377772 483052
rect 350316 483012 350322 483024
rect 377766 483012 377772 483024
rect 377824 483012 377830 483064
rect 552658 483012 552664 483064
rect 552716 483052 552722 483064
rect 574370 483052 574376 483064
rect 552716 483024 574376 483052
rect 552716 483012 552722 483024
rect 574370 483012 574376 483024
rect 574428 483012 574434 483064
rect 350442 481652 350448 481704
rect 350500 481692 350506 481704
rect 370038 481692 370044 481704
rect 350500 481664 370044 481692
rect 350500 481652 350506 481664
rect 370038 481652 370044 481664
rect 370096 481652 370102 481704
rect 402790 481652 402796 481704
rect 402848 481692 402854 481704
rect 407114 481692 407120 481704
rect 402848 481664 407120 481692
rect 402848 481652 402854 481664
rect 407114 481652 407120 481664
rect 407172 481652 407178 481704
rect 41874 480428 41880 480480
rect 41932 480468 41938 480480
rect 45830 480468 45836 480480
rect 41932 480440 45836 480468
rect 41932 480428 41938 480440
rect 45830 480428 45836 480440
rect 45888 480428 45894 480480
rect 350258 480292 350264 480344
rect 350316 480332 350322 480344
rect 366082 480332 366088 480344
rect 350316 480304 366088 480332
rect 350316 480292 350322 480304
rect 366082 480292 366088 480304
rect 366140 480292 366146 480344
rect 350442 480224 350448 480276
rect 350500 480264 350506 480276
rect 370130 480264 370136 480276
rect 350500 480236 370136 480264
rect 350500 480224 350506 480236
rect 370130 480224 370136 480236
rect 370188 480224 370194 480276
rect 383010 478864 383016 478916
rect 383068 478904 383074 478916
rect 407114 478904 407120 478916
rect 383068 478876 407120 478904
rect 383068 478864 383074 478876
rect 407114 478864 407120 478876
rect 407172 478864 407178 478916
rect 44726 478660 44732 478712
rect 44784 478700 44790 478712
rect 46658 478700 46664 478712
rect 44784 478672 46664 478700
rect 44784 478660 44790 478672
rect 46658 478660 46664 478672
rect 46716 478660 46722 478712
rect 553302 477504 553308 477556
rect 553360 477544 553366 477556
rect 562410 477544 562416 477556
rect 553360 477516 562416 477544
rect 553360 477504 553366 477516
rect 562410 477504 562416 477516
rect 562468 477504 562474 477556
rect 348510 476212 348516 476264
rect 348568 476252 348574 476264
rect 349798 476252 349804 476264
rect 348568 476224 349804 476252
rect 348568 476212 348574 476224
rect 349798 476212 349804 476224
rect 349856 476212 349862 476264
rect 350166 476144 350172 476196
rect 350224 476184 350230 476196
rect 361942 476184 361948 476196
rect 350224 476156 361948 476184
rect 350224 476144 350230 476156
rect 361942 476144 361948 476156
rect 362000 476144 362006 476196
rect 23106 476076 23112 476128
rect 23164 476116 23170 476128
rect 46750 476116 46756 476128
rect 23164 476088 46756 476116
rect 23164 476076 23170 476088
rect 46750 476076 46756 476088
rect 46808 476076 46814 476128
rect 350258 476076 350264 476128
rect 350316 476116 350322 476128
rect 370590 476116 370596 476128
rect 350316 476088 370596 476116
rect 350316 476076 350322 476088
rect 370590 476076 370596 476088
rect 370648 476076 370654 476128
rect 403342 474784 403348 474836
rect 403400 474824 403406 474836
rect 407298 474824 407304 474836
rect 403400 474796 407304 474824
rect 403400 474784 403406 474796
rect 407298 474784 407304 474796
rect 407356 474784 407362 474836
rect 552566 474784 552572 474836
rect 552624 474824 552630 474836
rect 561122 474824 561128 474836
rect 552624 474796 561128 474824
rect 552624 474784 552630 474796
rect 561122 474784 561128 474796
rect 561180 474784 561186 474836
rect 399570 474716 399576 474768
rect 399628 474756 399634 474768
rect 407114 474756 407120 474768
rect 399628 474728 407120 474756
rect 399628 474716 399634 474728
rect 407114 474716 407120 474728
rect 407172 474716 407178 474768
rect 553302 474716 553308 474768
rect 553360 474756 553366 474768
rect 561950 474756 561956 474768
rect 553360 474728 561956 474756
rect 553360 474716 553366 474728
rect 561950 474716 561956 474728
rect 562008 474716 562014 474768
rect 45094 474648 45100 474700
rect 45152 474688 45158 474700
rect 46474 474688 46480 474700
rect 45152 474660 46480 474688
rect 45152 474648 45158 474660
rect 46474 474648 46480 474660
rect 46532 474648 46538 474700
rect 43530 474580 43536 474632
rect 43588 474620 43594 474632
rect 46566 474620 46572 474632
rect 43588 474592 46572 474620
rect 43588 474580 43594 474592
rect 46566 474580 46572 474592
rect 46624 474580 46630 474632
rect 394418 473424 394424 473476
rect 394476 473464 394482 473476
rect 407114 473464 407120 473476
rect 394476 473436 407120 473464
rect 394476 473424 394482 473436
rect 407114 473424 407120 473436
rect 407172 473424 407178 473476
rect 350258 473356 350264 473408
rect 350316 473396 350322 473408
rect 352374 473396 352380 473408
rect 350316 473368 352380 473396
rect 350316 473356 350322 473368
rect 352374 473356 352380 473368
rect 352432 473356 352438 473408
rect 372062 473356 372068 473408
rect 372120 473396 372126 473408
rect 407298 473396 407304 473408
rect 372120 473368 407304 473396
rect 372120 473356 372126 473368
rect 407298 473356 407304 473368
rect 407356 473356 407362 473408
rect 350442 471996 350448 472048
rect 350500 472036 350506 472048
rect 353938 472036 353944 472048
rect 350500 472008 353944 472036
rect 350500 471996 350506 472008
rect 353938 471996 353944 472008
rect 353996 471996 354002 472048
rect 553302 470568 553308 470620
rect 553360 470608 553366 470620
rect 567838 470608 567844 470620
rect 553360 470580 567844 470608
rect 553360 470568 553366 470580
rect 567838 470568 567844 470580
rect 567896 470568 567902 470620
rect 570690 470568 570696 470620
rect 570748 470608 570754 470620
rect 580166 470608 580172 470620
rect 570748 470580 580172 470608
rect 570748 470568 570754 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 33594 469208 33600 469260
rect 33652 469248 33658 469260
rect 46750 469248 46756 469260
rect 33652 469220 46756 469248
rect 33652 469208 33658 469220
rect 46750 469208 46756 469220
rect 46808 469208 46814 469260
rect 361022 469208 361028 469260
rect 361080 469248 361086 469260
rect 407114 469248 407120 469260
rect 361080 469220 407120 469248
rect 361080 469208 361086 469220
rect 407114 469208 407120 469220
rect 407172 469208 407178 469260
rect 553302 469208 553308 469260
rect 553360 469248 553366 469260
rect 577314 469248 577320 469260
rect 553360 469220 577320 469248
rect 553360 469208 553366 469220
rect 577314 469208 577320 469220
rect 577372 469208 577378 469260
rect 404078 469140 404084 469192
rect 404136 469180 404142 469192
rect 407298 469180 407304 469192
rect 404136 469152 407304 469180
rect 404136 469140 404142 469152
rect 407298 469140 407304 469152
rect 407356 469140 407362 469192
rect 40770 467916 40776 467968
rect 40828 467956 40834 467968
rect 46750 467956 46756 467968
rect 40828 467928 46756 467956
rect 40828 467916 40834 467928
rect 46750 467916 46756 467928
rect 46808 467916 46814 467968
rect 23014 467848 23020 467900
rect 23072 467888 23078 467900
rect 46566 467888 46572 467900
rect 23072 467860 46572 467888
rect 23072 467848 23078 467860
rect 46566 467848 46572 467860
rect 46624 467848 46630 467900
rect 388898 467848 388904 467900
rect 388956 467888 388962 467900
rect 407114 467888 407120 467900
rect 388956 467860 407120 467888
rect 388956 467848 388962 467860
rect 407114 467848 407120 467860
rect 407172 467848 407178 467900
rect 350442 466420 350448 466472
rect 350500 466460 350506 466472
rect 392578 466460 392584 466472
rect 350500 466432 392584 466460
rect 350500 466420 350506 466432
rect 392578 466420 392584 466432
rect 392636 466420 392642 466472
rect 553302 466420 553308 466472
rect 553360 466460 553366 466472
rect 567470 466460 567476 466472
rect 553360 466432 567476 466460
rect 553360 466420 553366 466432
rect 567470 466420 567476 466432
rect 567528 466420 567534 466472
rect 350258 466352 350264 466404
rect 350316 466392 350322 466404
rect 403802 466392 403808 466404
rect 350316 466364 403808 466392
rect 350316 466352 350322 466364
rect 403802 466352 403808 466364
rect 403860 466352 403866 466404
rect 397270 465060 397276 465112
rect 397328 465100 397334 465112
rect 407114 465100 407120 465112
rect 397328 465072 407120 465100
rect 397328 465060 397334 465072
rect 407114 465060 407120 465072
rect 407172 465060 407178 465112
rect 552014 465060 552020 465112
rect 552072 465100 552078 465112
rect 575934 465100 575940 465112
rect 552072 465072 575940 465100
rect 552072 465060 552078 465072
rect 575934 465060 575940 465072
rect 575992 465060 575998 465112
rect 40586 464108 40592 464160
rect 40644 464148 40650 464160
rect 46750 464148 46756 464160
rect 40644 464120 46756 464148
rect 40644 464108 40650 464120
rect 46750 464108 46756 464120
rect 46808 464108 46814 464160
rect 552014 463904 552020 463956
rect 552072 463944 552078 463956
rect 556246 463944 556252 463956
rect 552072 463916 556252 463944
rect 552072 463904 552078 463916
rect 556246 463904 556252 463916
rect 556304 463904 556310 463956
rect 18874 463700 18880 463752
rect 18932 463740 18938 463752
rect 45646 463740 45652 463752
rect 18932 463712 45652 463740
rect 18932 463700 18938 463712
rect 45646 463700 45652 463712
rect 45704 463700 45710 463752
rect 383194 463700 383200 463752
rect 383252 463740 383258 463752
rect 407114 463740 407120 463752
rect 383252 463712 407120 463740
rect 383252 463700 383258 463712
rect 407114 463700 407120 463712
rect 407172 463700 407178 463752
rect 35618 463632 35624 463684
rect 35676 463672 35682 463684
rect 46750 463672 46756 463684
rect 35676 463644 46756 463672
rect 35676 463632 35682 463644
rect 46750 463632 46756 463644
rect 46808 463632 46814 463684
rect 350442 462476 350448 462528
rect 350500 462516 350506 462528
rect 395798 462516 395804 462528
rect 350500 462488 395804 462516
rect 350500 462476 350506 462488
rect 395798 462476 395804 462488
rect 395856 462476 395862 462528
rect 350258 462408 350264 462460
rect 350316 462448 350322 462460
rect 376294 462448 376300 462460
rect 350316 462420 376300 462448
rect 350316 462408 350322 462420
rect 376294 462408 376300 462420
rect 376352 462408 376358 462460
rect 392670 462408 392676 462460
rect 392728 462448 392734 462460
rect 407114 462448 407120 462460
rect 392728 462420 407120 462448
rect 392728 462408 392734 462420
rect 407114 462408 407120 462420
rect 407172 462408 407178 462460
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 19978 462380 19984 462392
rect 3568 462352 19984 462380
rect 3568 462340 3574 462352
rect 19978 462340 19984 462352
rect 20036 462340 20042 462392
rect 394234 462340 394240 462392
rect 394292 462380 394298 462392
rect 407298 462380 407304 462392
rect 394292 462352 407304 462380
rect 394292 462340 394298 462352
rect 407298 462340 407304 462352
rect 407356 462340 407362 462392
rect 552014 462340 552020 462392
rect 552072 462380 552078 462392
rect 573082 462380 573088 462392
rect 552072 462352 573088 462380
rect 552072 462340 552078 462352
rect 573082 462340 573088 462352
rect 573140 462340 573146 462392
rect 350442 461048 350448 461100
rect 350500 461088 350506 461100
rect 362954 461088 362960 461100
rect 350500 461060 362960 461088
rect 350500 461048 350506 461060
rect 362954 461048 362960 461060
rect 363012 461048 363018 461100
rect 350258 460980 350264 461032
rect 350316 461020 350322 461032
rect 364518 461020 364524 461032
rect 350316 460992 364524 461020
rect 350316 460980 350322 460992
rect 364518 460980 364524 460992
rect 364576 460980 364582 461032
rect 21910 460912 21916 460964
rect 21968 460952 21974 460964
rect 46750 460952 46756 460964
rect 21968 460924 46756 460952
rect 21968 460912 21974 460924
rect 46750 460912 46756 460924
rect 46808 460912 46814 460964
rect 362310 460912 362316 460964
rect 362368 460952 362374 460964
rect 407114 460952 407120 460964
rect 362368 460924 407120 460952
rect 362368 460912 362374 460924
rect 407114 460912 407120 460924
rect 407172 460912 407178 460964
rect 39482 460844 39488 460896
rect 39540 460884 39546 460896
rect 46566 460884 46572 460896
rect 39540 460856 46572 460884
rect 39540 460844 39546 460856
rect 46566 460844 46572 460856
rect 46624 460844 46630 460896
rect 350442 459552 350448 459604
rect 350500 459592 350506 459604
rect 396902 459592 396908 459604
rect 350500 459564 396908 459592
rect 350500 459552 350506 459564
rect 396902 459552 396908 459564
rect 396960 459552 396966 459604
rect 552014 459552 552020 459604
rect 552072 459592 552078 459604
rect 560846 459592 560852 459604
rect 552072 459564 560852 459592
rect 552072 459552 552078 459564
rect 560846 459552 560852 459564
rect 560904 459552 560910 459604
rect 552014 459008 552020 459060
rect 552072 459048 552078 459060
rect 553854 459048 553860 459060
rect 552072 459020 553860 459048
rect 552072 459008 552078 459020
rect 553854 459008 553860 459020
rect 553912 459008 553918 459060
rect 31386 458192 31392 458244
rect 31444 458232 31450 458244
rect 46750 458232 46756 458244
rect 31444 458204 46756 458232
rect 31444 458192 31450 458204
rect 46750 458192 46756 458204
rect 46808 458192 46814 458244
rect 403894 458192 403900 458244
rect 403952 458232 403958 458244
rect 407114 458232 407120 458244
rect 403952 458204 407120 458232
rect 403952 458192 403958 458204
rect 407114 458192 407120 458204
rect 407172 458192 407178 458244
rect 350442 456832 350448 456884
rect 350500 456872 350506 456884
rect 367186 456872 367192 456884
rect 350500 456844 367192 456872
rect 350500 456832 350506 456844
rect 367186 456832 367192 456844
rect 367244 456832 367250 456884
rect 350258 456764 350264 456816
rect 350316 456804 350322 456816
rect 375466 456804 375472 456816
rect 350316 456776 375472 456804
rect 350316 456764 350322 456776
rect 375466 456764 375472 456776
rect 375524 456764 375530 456816
rect 391474 456764 391480 456816
rect 391532 456804 391538 456816
rect 407114 456804 407120 456816
rect 391532 456776 407120 456804
rect 391532 456764 391538 456776
rect 407114 456764 407120 456776
rect 407172 456764 407178 456816
rect 552014 456764 552020 456816
rect 552072 456804 552078 456816
rect 576210 456804 576216 456816
rect 552072 456776 576216 456804
rect 552072 456764 552078 456776
rect 576210 456764 576216 456776
rect 576268 456764 576274 456816
rect 43990 456696 43996 456748
rect 44048 456736 44054 456748
rect 46750 456736 46756 456748
rect 44048 456708 46756 456736
rect 44048 456696 44054 456708
rect 46750 456696 46756 456708
rect 46808 456696 46814 456748
rect 386046 456696 386052 456748
rect 386104 456736 386110 456748
rect 407298 456736 407304 456748
rect 386104 456708 407304 456736
rect 386104 456696 386110 456708
rect 407298 456696 407304 456708
rect 407356 456696 407362 456748
rect 552014 456016 552020 456068
rect 552072 456056 552078 456068
rect 553946 456056 553952 456068
rect 552072 456028 553952 456056
rect 552072 456016 552078 456028
rect 553946 456016 553952 456028
rect 554004 456016 554010 456068
rect 348970 455336 348976 455388
rect 349028 455376 349034 455388
rect 350534 455376 350540 455388
rect 349028 455348 350540 455376
rect 349028 455336 349034 455348
rect 350534 455336 350540 455348
rect 350592 455336 350598 455388
rect 369486 455336 369492 455388
rect 369544 455376 369550 455388
rect 407114 455376 407120 455388
rect 369544 455348 407120 455376
rect 369544 455336 369550 455348
rect 407114 455336 407120 455348
rect 407172 455336 407178 455388
rect 350442 454044 350448 454096
rect 350500 454084 350506 454096
rect 380618 454084 380624 454096
rect 350500 454056 380624 454084
rect 350500 454044 350506 454056
rect 380618 454044 380624 454056
rect 380676 454044 380682 454096
rect 405274 454044 405280 454096
rect 405332 454084 405338 454096
rect 407666 454084 407672 454096
rect 405332 454056 407672 454084
rect 405332 454044 405338 454056
rect 407666 454044 407672 454056
rect 407724 454044 407730 454096
rect 553302 454044 553308 454096
rect 553360 454084 553366 454096
rect 565906 454084 565912 454096
rect 553360 454056 565912 454084
rect 553360 454044 553366 454056
rect 565906 454044 565912 454056
rect 565964 454044 565970 454096
rect 552842 452752 552848 452804
rect 552900 452792 552906 452804
rect 556338 452792 556344 452804
rect 552900 452764 556344 452792
rect 552900 452752 552906 452764
rect 556338 452752 556344 452764
rect 556396 452752 556402 452804
rect 366542 452616 366548 452668
rect 366600 452656 366606 452668
rect 407114 452656 407120 452668
rect 366600 452628 407120 452656
rect 366600 452616 366606 452628
rect 407114 452616 407120 452628
rect 407172 452616 407178 452668
rect 350442 451256 350448 451308
rect 350500 451296 350506 451308
rect 386046 451296 386052 451308
rect 350500 451268 386052 451296
rect 350500 451256 350506 451268
rect 386046 451256 386052 451268
rect 386104 451256 386110 451308
rect 400950 451256 400956 451308
rect 401008 451296 401014 451308
rect 407114 451296 407120 451308
rect 401008 451268 407120 451296
rect 401008 451256 401014 451268
rect 407114 451256 407120 451268
rect 407172 451256 407178 451308
rect 34422 451188 34428 451240
rect 34480 451228 34486 451240
rect 46750 451228 46756 451240
rect 34480 451200 46756 451228
rect 34480 451188 34486 451200
rect 46750 451188 46756 451200
rect 46808 451188 46814 451240
rect 350442 449896 350448 449948
rect 350500 449936 350506 449948
rect 362494 449936 362500 449948
rect 350500 449908 362500 449936
rect 350500 449896 350506 449908
rect 362494 449896 362500 449908
rect 362552 449896 362558 449948
rect 553302 449896 553308 449948
rect 553360 449936 553366 449948
rect 578326 449936 578332 449948
rect 553360 449908 578332 449936
rect 553360 449896 553366 449908
rect 578326 449896 578332 449908
rect 578384 449896 578390 449948
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 17310 448576 17316 448588
rect 3200 448548 17316 448576
rect 3200 448536 3206 448548
rect 17310 448536 17316 448548
rect 17368 448536 17374 448588
rect 383470 448536 383476 448588
rect 383528 448576 383534 448588
rect 407114 448576 407120 448588
rect 383528 448548 407120 448576
rect 383528 448536 383534 448548
rect 407114 448536 407120 448548
rect 407172 448536 407178 448588
rect 552566 448536 552572 448588
rect 552624 448576 552630 448588
rect 575658 448576 575664 448588
rect 552624 448548 575664 448576
rect 552624 448536 552630 448548
rect 575658 448536 575664 448548
rect 575716 448536 575722 448588
rect 348878 447108 348884 447160
rect 348936 447148 348942 447160
rect 349154 447148 349160 447160
rect 348936 447120 349160 447148
rect 348936 447108 348942 447120
rect 349154 447108 349160 447120
rect 349212 447108 349218 447160
rect 350442 447108 350448 447160
rect 350500 447148 350506 447160
rect 367278 447148 367284 447160
rect 350500 447120 367284 447148
rect 350500 447108 350506 447120
rect 367278 447108 367284 447120
rect 367336 447108 367342 447160
rect 403526 447108 403532 447160
rect 403584 447148 403590 447160
rect 407298 447148 407304 447160
rect 403584 447120 407304 447148
rect 403584 447108 403590 447120
rect 407298 447108 407304 447120
rect 407356 447108 407362 447160
rect 395614 447040 395620 447092
rect 395672 447080 395678 447092
rect 407114 447080 407120 447092
rect 395672 447052 407120 447080
rect 395672 447040 395678 447052
rect 407114 447040 407120 447052
rect 407172 447040 407178 447092
rect 29638 445748 29644 445800
rect 29696 445788 29702 445800
rect 46750 445788 46756 445800
rect 29696 445760 46756 445788
rect 29696 445748 29702 445760
rect 46750 445748 46756 445760
rect 46808 445748 46814 445800
rect 350258 445748 350264 445800
rect 350316 445788 350322 445800
rect 370774 445788 370780 445800
rect 350316 445760 370780 445788
rect 350316 445748 350322 445760
rect 370774 445748 370780 445760
rect 370832 445748 370838 445800
rect 552566 445748 552572 445800
rect 552624 445788 552630 445800
rect 566366 445788 566372 445800
rect 552624 445760 566372 445788
rect 552624 445748 552630 445760
rect 566366 445748 566372 445760
rect 566424 445748 566430 445800
rect 350442 445680 350448 445732
rect 350500 445720 350506 445732
rect 399662 445720 399668 445732
rect 350500 445692 399668 445720
rect 350500 445680 350506 445692
rect 399662 445680 399668 445692
rect 399720 445680 399726 445732
rect 373626 445612 373632 445664
rect 373684 445652 373690 445664
rect 407114 445652 407120 445664
rect 373684 445624 407120 445652
rect 373684 445612 373690 445624
rect 407114 445612 407120 445624
rect 407172 445612 407178 445664
rect 27062 444388 27068 444440
rect 27120 444428 27126 444440
rect 46750 444428 46756 444440
rect 27120 444400 46756 444428
rect 27120 444388 27126 444400
rect 46750 444388 46756 444400
rect 46808 444388 46814 444440
rect 552566 444388 552572 444440
rect 552624 444428 552630 444440
rect 581270 444428 581276 444440
rect 552624 444400 581276 444428
rect 552624 444388 552630 444400
rect 581270 444388 581276 444400
rect 581328 444388 581334 444440
rect 38470 442960 38476 443012
rect 38528 443000 38534 443012
rect 46750 443000 46756 443012
rect 38528 442972 46756 443000
rect 38528 442960 38534 442972
rect 46750 442960 46756 442972
rect 46808 442960 46814 443012
rect 553302 442960 553308 443012
rect 553360 443000 553366 443012
rect 569126 443000 569132 443012
rect 553360 442972 569132 443000
rect 553360 442960 553366 442972
rect 569126 442960 569132 442972
rect 569184 442960 569190 443012
rect 362402 441600 362408 441652
rect 362460 441640 362466 441652
rect 407114 441640 407120 441652
rect 362460 441612 407120 441640
rect 362460 441600 362466 441612
rect 407114 441600 407120 441612
rect 407172 441600 407178 441652
rect 395890 441532 395896 441584
rect 395948 441572 395954 441584
rect 407298 441572 407304 441584
rect 395948 441544 407304 441572
rect 395948 441532 395954 441544
rect 407298 441532 407304 441544
rect 407356 441532 407362 441584
rect 350442 440240 350448 440292
rect 350500 440280 350506 440292
rect 395614 440280 395620 440292
rect 350500 440252 395620 440280
rect 350500 440240 350506 440252
rect 395614 440240 395620 440252
rect 395672 440240 395678 440292
rect 40678 438948 40684 439000
rect 40736 438988 40742 439000
rect 46750 438988 46756 439000
rect 40736 438960 46756 438988
rect 40736 438948 40742 438960
rect 46750 438948 46756 438960
rect 46808 438948 46814 439000
rect 41690 438880 41696 438932
rect 41748 438920 41754 438932
rect 46014 438920 46020 438932
rect 41748 438892 46020 438920
rect 41748 438880 41754 438892
rect 46014 438880 46020 438892
rect 46072 438880 46078 438932
rect 386230 438880 386236 438932
rect 386288 438920 386294 438932
rect 407114 438920 407120 438932
rect 386288 438892 407120 438920
rect 386288 438880 386294 438892
rect 407114 438880 407120 438892
rect 407172 438880 407178 438932
rect 404998 438812 405004 438864
rect 405056 438852 405062 438864
rect 407482 438852 407488 438864
rect 405056 438824 407488 438852
rect 405056 438812 405062 438824
rect 407482 438812 407488 438824
rect 407540 438812 407546 438864
rect 562410 437588 562416 437640
rect 562468 437628 562474 437640
rect 563238 437628 563244 437640
rect 562468 437600 563244 437628
rect 562468 437588 562474 437600
rect 563238 437588 563244 437600
rect 563296 437588 563302 437640
rect 350258 437452 350264 437504
rect 350316 437492 350322 437504
rect 398466 437492 398472 437504
rect 350316 437464 398472 437492
rect 350316 437452 350322 437464
rect 398466 437452 398472 437464
rect 398524 437452 398530 437504
rect 553302 437452 553308 437504
rect 553360 437492 553366 437504
rect 562318 437492 562324 437504
rect 553360 437464 562324 437492
rect 553360 437452 553366 437464
rect 562318 437452 562324 437464
rect 562376 437452 562382 437504
rect 350442 437384 350448 437436
rect 350500 437424 350506 437436
rect 403710 437424 403716 437436
rect 350500 437396 403716 437424
rect 350500 437384 350506 437396
rect 403710 437384 403716 437396
rect 403768 437384 403774 437436
rect 553026 437384 553032 437436
rect 553084 437424 553090 437436
rect 556890 437424 556896 437436
rect 553084 437396 556896 437424
rect 553084 437384 553090 437396
rect 556890 437384 556896 437396
rect 556948 437384 556954 437436
rect 348878 436296 348884 436348
rect 348936 436336 348942 436348
rect 349154 436336 349160 436348
rect 348936 436308 349160 436336
rect 348936 436296 348942 436308
rect 349154 436296 349160 436308
rect 349212 436296 349218 436348
rect 43530 436092 43536 436144
rect 43588 436132 43594 436144
rect 46750 436132 46756 436144
rect 43588 436104 46756 436132
rect 43588 436092 43594 436104
rect 46750 436092 46756 436104
rect 46808 436092 46814 436144
rect 397178 436092 397184 436144
rect 397236 436132 397242 436144
rect 407114 436132 407120 436144
rect 397236 436104 407120 436132
rect 397236 436092 397242 436104
rect 407114 436092 407120 436104
rect 407172 436092 407178 436144
rect 553302 436092 553308 436144
rect 553360 436132 553366 436144
rect 577682 436132 577688 436144
rect 553360 436104 577688 436132
rect 553360 436092 553366 436104
rect 577682 436092 577688 436104
rect 577740 436092 577746 436144
rect 553026 435956 553032 436008
rect 553084 435996 553090 436008
rect 553302 435996 553308 436008
rect 553084 435968 553308 435996
rect 553084 435956 553090 435968
rect 553302 435956 553308 435968
rect 553360 435956 553366 436008
rect 350442 434800 350448 434852
rect 350500 434840 350506 434852
rect 370222 434840 370228 434852
rect 350500 434812 370228 434840
rect 350500 434800 350506 434812
rect 370222 434800 370228 434812
rect 370280 434800 370286 434852
rect 43990 434732 43996 434784
rect 44048 434772 44054 434784
rect 46750 434772 46756 434784
rect 44048 434744 46756 434772
rect 44048 434732 44054 434744
rect 46750 434732 46756 434744
rect 46808 434732 46814 434784
rect 363966 434732 363972 434784
rect 364024 434772 364030 434784
rect 407114 434772 407120 434784
rect 364024 434744 407120 434772
rect 364024 434732 364030 434744
rect 407114 434732 407120 434744
rect 407172 434732 407178 434784
rect 33870 433304 33876 433356
rect 33928 433344 33934 433356
rect 46750 433344 46756 433356
rect 33928 433316 46756 433344
rect 33928 433304 33934 433316
rect 46750 433304 46756 433316
rect 46808 433304 46814 433356
rect 42518 431944 42524 431996
rect 42576 431984 42582 431996
rect 46750 431984 46756 431996
rect 42576 431956 46756 431984
rect 42576 431944 42582 431956
rect 46750 431944 46756 431956
rect 46808 431944 46814 431996
rect 577590 431740 577596 431792
rect 577648 431780 577654 431792
rect 579890 431780 579896 431792
rect 577648 431752 579896 431780
rect 577648 431740 577654 431752
rect 579890 431740 579896 431752
rect 579948 431740 579954 431792
rect 350442 430652 350448 430704
rect 350500 430692 350506 430704
rect 373810 430692 373816 430704
rect 350500 430664 373816 430692
rect 350500 430652 350506 430664
rect 373810 430652 373816 430664
rect 373868 430652 373874 430704
rect 350258 430584 350264 430636
rect 350316 430624 350322 430636
rect 396994 430624 397000 430636
rect 350316 430596 397000 430624
rect 350316 430584 350322 430596
rect 396994 430584 397000 430596
rect 397052 430584 397058 430636
rect 552198 430176 552204 430228
rect 552256 430216 552262 430228
rect 555050 430216 555056 430228
rect 552256 430188 555056 430216
rect 552256 430176 552262 430188
rect 555050 430176 555056 430188
rect 555108 430176 555114 430228
rect 402606 429224 402612 429276
rect 402664 429264 402670 429276
rect 407114 429264 407120 429276
rect 402664 429236 407120 429264
rect 402664 429224 402670 429236
rect 407114 429224 407120 429236
rect 407172 429224 407178 429276
rect 40494 427864 40500 427916
rect 40552 427904 40558 427916
rect 46658 427904 46664 427916
rect 40552 427876 46664 427904
rect 40552 427864 40558 427876
rect 46658 427864 46664 427876
rect 46716 427864 46722 427916
rect 396626 427864 396632 427916
rect 396684 427904 396690 427916
rect 407114 427904 407120 427916
rect 396684 427876 407120 427904
rect 396684 427864 396690 427876
rect 407114 427864 407120 427876
rect 407172 427864 407178 427916
rect 33778 427796 33784 427848
rect 33836 427836 33842 427848
rect 46750 427836 46756 427848
rect 33836 427808 46756 427836
rect 33836 427796 33842 427808
rect 46750 427796 46756 427808
rect 46808 427796 46814 427848
rect 350442 427796 350448 427848
rect 350500 427836 350506 427848
rect 375006 427836 375012 427848
rect 350500 427808 375012 427836
rect 350500 427796 350506 427808
rect 375006 427796 375012 427808
rect 375064 427796 375070 427848
rect 553026 427796 553032 427848
rect 553084 427836 553090 427848
rect 563882 427836 563888 427848
rect 553084 427808 563888 427836
rect 553084 427796 553090 427808
rect 563882 427796 563888 427808
rect 563940 427796 563946 427848
rect 369486 426572 369492 426624
rect 369544 426612 369550 426624
rect 407206 426612 407212 426624
rect 369544 426584 407212 426612
rect 369544 426572 369550 426584
rect 407206 426572 407212 426584
rect 407264 426572 407270 426624
rect 361114 426504 361120 426556
rect 361172 426544 361178 426556
rect 407114 426544 407120 426556
rect 361172 426516 407120 426544
rect 361172 426504 361178 426516
rect 407114 426504 407120 426516
rect 407172 426504 407178 426556
rect 350442 426436 350448 426488
rect 350500 426476 350506 426488
rect 399662 426476 399668 426488
rect 350500 426448 399668 426476
rect 350500 426436 350506 426448
rect 399662 426436 399668 426448
rect 399720 426436 399726 426488
rect 553026 426436 553032 426488
rect 553084 426476 553090 426488
rect 577130 426476 577136 426488
rect 553084 426448 577136 426476
rect 553084 426436 553090 426448
rect 577130 426436 577136 426448
rect 577188 426436 577194 426488
rect 43438 425076 43444 425128
rect 43496 425116 43502 425128
rect 45646 425116 45652 425128
rect 43496 425088 45652 425116
rect 43496 425076 43502 425088
rect 45646 425076 45652 425088
rect 45704 425076 45710 425128
rect 350442 425076 350448 425128
rect 350500 425116 350506 425128
rect 359182 425116 359188 425128
rect 350500 425088 359188 425116
rect 350500 425076 350506 425088
rect 359182 425076 359188 425088
rect 359240 425076 359246 425128
rect 553026 425076 553032 425128
rect 553084 425116 553090 425128
rect 569494 425116 569500 425128
rect 553084 425088 569500 425116
rect 553084 425076 553090 425088
rect 569494 425076 569500 425088
rect 569552 425076 569558 425128
rect 553026 423716 553032 423768
rect 553084 423756 553090 423768
rect 570598 423756 570604 423768
rect 553084 423728 570604 423756
rect 553084 423716 553090 423728
rect 570598 423716 570604 423728
rect 570656 423716 570662 423768
rect 24118 423648 24124 423700
rect 24176 423688 24182 423700
rect 46750 423688 46756 423700
rect 24176 423660 46756 423688
rect 24176 423648 24182 423660
rect 46750 423648 46756 423660
rect 46808 423648 46814 423700
rect 374822 423648 374828 423700
rect 374880 423688 374886 423700
rect 407114 423688 407120 423700
rect 374880 423660 407120 423688
rect 374880 423648 374886 423660
rect 407114 423648 407120 423660
rect 407172 423648 407178 423700
rect 552934 423648 552940 423700
rect 552992 423688 552998 423700
rect 574830 423688 574836 423700
rect 552992 423660 574836 423688
rect 552992 423648 552998 423660
rect 574830 423648 574836 423660
rect 574888 423648 574894 423700
rect 350442 422288 350448 422340
rect 350500 422328 350506 422340
rect 376570 422328 376576 422340
rect 350500 422300 376576 422328
rect 350500 422288 350506 422300
rect 376570 422288 376576 422300
rect 376628 422288 376634 422340
rect 393866 422288 393872 422340
rect 393924 422328 393930 422340
rect 407114 422328 407120 422340
rect 393924 422300 407120 422328
rect 393924 422288 393930 422300
rect 407114 422288 407120 422300
rect 407172 422288 407178 422340
rect 349982 420996 349988 421048
rect 350040 421036 350046 421048
rect 352466 421036 352472 421048
rect 350040 421008 352472 421036
rect 350040 420996 350046 421008
rect 352466 420996 352472 421008
rect 352524 420996 352530 421048
rect 552198 420996 552204 421048
rect 552256 421036 552262 421048
rect 554958 421036 554964 421048
rect 552256 421008 554964 421036
rect 552256 420996 552262 421008
rect 554958 420996 554964 421008
rect 555016 420996 555022 421048
rect 35158 420928 35164 420980
rect 35216 420968 35222 420980
rect 45646 420968 45652 420980
rect 35216 420940 45652 420968
rect 35216 420928 35222 420940
rect 45646 420928 45652 420940
rect 45704 420928 45710 420980
rect 350442 420928 350448 420980
rect 350500 420968 350506 420980
rect 383378 420968 383384 420980
rect 350500 420940 383384 420968
rect 350500 420928 350506 420940
rect 383378 420928 383384 420940
rect 383436 420928 383442 420980
rect 570782 420180 570788 420232
rect 570840 420220 570846 420232
rect 580442 420220 580448 420232
rect 570840 420192 580448 420220
rect 570840 420180 570846 420192
rect 580442 420180 580448 420192
rect 580500 420180 580506 420232
rect 553026 420112 553032 420164
rect 553084 420152 553090 420164
rect 559558 420152 559564 420164
rect 553084 420124 559564 420152
rect 553084 420112 553090 420124
rect 559558 420112 559564 420124
rect 559616 420112 559622 420164
rect 28350 419568 28356 419620
rect 28408 419608 28414 419620
rect 45646 419608 45652 419620
rect 28408 419580 45652 419608
rect 28408 419568 28414 419580
rect 45646 419568 45652 419580
rect 45704 419568 45710 419620
rect 350442 419568 350448 419620
rect 350500 419608 350506 419620
rect 368566 419608 368572 419620
rect 350500 419580 368572 419608
rect 350500 419568 350506 419580
rect 368566 419568 368572 419580
rect 368624 419568 368630 419620
rect 369578 419568 369584 419620
rect 369636 419608 369642 419620
rect 407206 419608 407212 419620
rect 369636 419580 407212 419608
rect 369636 419568 369642 419580
rect 407206 419568 407212 419580
rect 407264 419568 407270 419620
rect 26786 419500 26792 419552
rect 26844 419540 26850 419552
rect 45922 419540 45928 419552
rect 26844 419512 45928 419540
rect 26844 419500 26850 419512
rect 45922 419500 45928 419512
rect 45980 419500 45986 419552
rect 356974 419500 356980 419552
rect 357032 419540 357038 419552
rect 407114 419540 407120 419552
rect 357032 419512 407120 419540
rect 357032 419500 357038 419512
rect 407114 419500 407120 419512
rect 407172 419500 407178 419552
rect 350442 418208 350448 418260
rect 350500 418248 350506 418260
rect 381998 418248 382004 418260
rect 350500 418220 382004 418248
rect 350500 418208 350506 418220
rect 381998 418208 382004 418220
rect 382056 418208 382062 418260
rect 39482 418140 39488 418192
rect 39540 418180 39546 418192
rect 45922 418180 45928 418192
rect 39540 418152 45928 418180
rect 39540 418140 39546 418152
rect 45922 418140 45928 418152
rect 45980 418140 45986 418192
rect 372338 418140 372344 418192
rect 372396 418180 372402 418192
rect 407114 418180 407120 418192
rect 372396 418152 407120 418180
rect 372396 418140 372402 418152
rect 407114 418140 407120 418152
rect 407172 418140 407178 418192
rect 350442 416780 350448 416832
rect 350500 416820 350506 416832
rect 379146 416820 379152 416832
rect 350500 416792 379152 416820
rect 350500 416780 350506 416792
rect 379146 416780 379152 416792
rect 379204 416780 379210 416832
rect 380710 416712 380716 416764
rect 380768 416752 380774 416764
rect 407114 416752 407120 416764
rect 380768 416724 407120 416752
rect 380768 416712 380774 416724
rect 407114 416712 407120 416724
rect 407172 416712 407178 416764
rect 553026 416032 553032 416084
rect 553084 416072 553090 416084
rect 559466 416072 559472 416084
rect 553084 416044 559472 416072
rect 553084 416032 553090 416044
rect 559466 416032 559472 416044
rect 559524 416032 559530 416084
rect 28810 415488 28816 415540
rect 28868 415528 28874 415540
rect 45646 415528 45652 415540
rect 28868 415500 45652 415528
rect 28868 415488 28874 415500
rect 45646 415488 45652 415500
rect 45704 415488 45710 415540
rect 24210 415420 24216 415472
rect 24268 415460 24274 415472
rect 45922 415460 45928 415472
rect 24268 415432 45928 415460
rect 24268 415420 24274 415432
rect 45922 415420 45928 415432
rect 45980 415420 45986 415472
rect 553026 415420 553032 415472
rect 553084 415460 553090 415472
rect 579706 415460 579712 415472
rect 553084 415432 579712 415460
rect 553084 415420 553090 415432
rect 579706 415420 579712 415432
rect 579764 415420 579770 415472
rect 350442 414060 350448 414112
rect 350500 414100 350506 414112
rect 374730 414100 374736 414112
rect 350500 414072 374736 414100
rect 350500 414060 350506 414072
rect 374730 414060 374736 414072
rect 374788 414060 374794 414112
rect 20162 413992 20168 414044
rect 20220 414032 20226 414044
rect 46750 414032 46756 414044
rect 20220 414004 46756 414032
rect 20220 413992 20226 414004
rect 46750 413992 46756 414004
rect 46808 413992 46814 414044
rect 350258 413992 350264 414044
rect 350316 414032 350322 414044
rect 376478 414032 376484 414044
rect 350316 414004 376484 414032
rect 350316 413992 350322 414004
rect 376478 413992 376484 414004
rect 376536 413992 376542 414044
rect 388990 413992 388996 414044
rect 389048 414032 389054 414044
rect 407114 414032 407120 414044
rect 389048 414004 407120 414032
rect 389048 413992 389054 414004
rect 407114 413992 407120 414004
rect 407172 413992 407178 414044
rect 552382 412768 552388 412820
rect 552440 412808 552446 412820
rect 555326 412808 555332 412820
rect 552440 412780 555332 412808
rect 552440 412768 552446 412780
rect 555326 412768 555332 412780
rect 555384 412768 555390 412820
rect 553026 412632 553032 412684
rect 553084 412672 553090 412684
rect 580074 412672 580080 412684
rect 553084 412644 580080 412672
rect 553084 412632 553090 412644
rect 580074 412632 580080 412644
rect 580132 412632 580138 412684
rect 35618 411272 35624 411324
rect 35676 411312 35682 411324
rect 46750 411312 46756 411324
rect 35676 411284 46756 411312
rect 35676 411272 35682 411284
rect 46750 411272 46756 411284
rect 46808 411272 46814 411324
rect 350442 411272 350448 411324
rect 350500 411312 350506 411324
rect 375098 411312 375104 411324
rect 350500 411284 375104 411312
rect 350500 411272 350506 411284
rect 375098 411272 375104 411284
rect 375156 411272 375162 411324
rect 395890 411272 395896 411324
rect 395948 411312 395954 411324
rect 407114 411312 407120 411324
rect 395948 411284 407120 411312
rect 395948 411272 395954 411284
rect 407114 411272 407120 411284
rect 407172 411272 407178 411324
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 32490 411244 32496 411256
rect 3016 411216 32496 411244
rect 3016 411204 3022 411216
rect 32490 411204 32496 411216
rect 32548 411204 32554 411256
rect 359550 409844 359556 409896
rect 359608 409884 359614 409896
rect 407114 409884 407120 409896
rect 359608 409856 407120 409884
rect 359608 409844 359614 409856
rect 407114 409844 407120 409856
rect 407172 409844 407178 409896
rect 553026 409844 553032 409896
rect 553084 409884 553090 409896
rect 570230 409884 570236 409896
rect 553084 409856 570236 409884
rect 553084 409844 553090 409856
rect 570230 409844 570236 409856
rect 570288 409844 570294 409896
rect 399938 408484 399944 408536
rect 399996 408524 400002 408536
rect 407114 408524 407120 408536
rect 399996 408496 407120 408524
rect 399996 408484 400002 408496
rect 407114 408484 407120 408496
rect 407172 408484 407178 408536
rect 348970 407736 348976 407788
rect 349028 407776 349034 407788
rect 350166 407776 350172 407788
rect 349028 407748 350172 407776
rect 349028 407736 349034 407748
rect 350166 407736 350172 407748
rect 350224 407736 350230 407788
rect 21450 407124 21456 407176
rect 21508 407164 21514 407176
rect 46750 407164 46756 407176
rect 21508 407136 46756 407164
rect 21508 407124 21514 407136
rect 46750 407124 46756 407136
rect 46808 407124 46814 407176
rect 368014 405696 368020 405748
rect 368072 405736 368078 405748
rect 407114 405736 407120 405748
rect 368072 405708 407120 405736
rect 368072 405696 368078 405708
rect 407114 405696 407120 405708
rect 407172 405696 407178 405748
rect 400030 405628 400036 405680
rect 400088 405668 400094 405680
rect 407206 405668 407212 405680
rect 400088 405640 407212 405668
rect 400088 405628 400094 405640
rect 407206 405628 407212 405640
rect 407264 405628 407270 405680
rect 553026 405628 553032 405680
rect 553084 405668 553090 405680
rect 579154 405668 579160 405680
rect 553084 405640 579160 405668
rect 553084 405628 553090 405640
rect 579154 405628 579160 405640
rect 579212 405628 579218 405680
rect 350258 404404 350264 404456
rect 350316 404444 350322 404456
rect 364610 404444 364616 404456
rect 350316 404416 364616 404444
rect 350316 404404 350322 404416
rect 364610 404404 364616 404416
rect 364668 404404 364674 404456
rect 350442 404336 350448 404388
rect 350500 404376 350506 404388
rect 368290 404376 368296 404388
rect 350500 404348 368296 404376
rect 350500 404336 350506 404348
rect 368290 404336 368296 404348
rect 368348 404336 368354 404388
rect 553026 403656 553032 403708
rect 553084 403696 553090 403708
rect 557810 403696 557816 403708
rect 553084 403668 557816 403696
rect 553084 403656 553090 403668
rect 557810 403656 557816 403668
rect 557868 403656 557874 403708
rect 41966 402976 41972 403028
rect 42024 403016 42030 403028
rect 46750 403016 46756 403028
rect 42024 402988 46756 403016
rect 42024 402976 42030 402988
rect 46750 402976 46756 402988
rect 46808 402976 46814 403028
rect 553026 402976 553032 403028
rect 553084 403016 553090 403028
rect 579890 403016 579896 403028
rect 553084 402988 579896 403016
rect 553084 402976 553090 402988
rect 579890 402976 579896 402988
rect 579948 402976 579954 403028
rect 42150 402092 42156 402144
rect 42208 402132 42214 402144
rect 44174 402132 44180 402144
rect 42208 402104 44180 402132
rect 42208 402092 42214 402104
rect 44174 402092 44180 402104
rect 44232 402092 44238 402144
rect 42150 400188 42156 400240
rect 42208 400228 42214 400240
rect 46750 400228 46756 400240
rect 42208 400200 46756 400228
rect 42208 400188 42214 400200
rect 46750 400188 46756 400200
rect 46808 400188 46814 400240
rect 350442 400188 350448 400240
rect 350500 400228 350506 400240
rect 372154 400228 372160 400240
rect 350500 400200 372160 400228
rect 350500 400188 350506 400200
rect 372154 400188 372160 400200
rect 372212 400188 372218 400240
rect 404998 400188 405004 400240
rect 405056 400228 405062 400240
rect 407482 400228 407488 400240
rect 405056 400200 407488 400228
rect 405056 400188 405062 400200
rect 407482 400188 407488 400200
rect 407540 400188 407546 400240
rect 553026 400188 553032 400240
rect 553084 400228 553090 400240
rect 582742 400228 582748 400240
rect 553084 400200 582748 400228
rect 553084 400188 553090 400200
rect 582742 400188 582748 400200
rect 582800 400188 582806 400240
rect 403986 400120 403992 400172
rect 404044 400160 404050 400172
rect 407114 400160 407120 400172
rect 404044 400132 407120 400160
rect 404044 400120 404050 400132
rect 407114 400120 407120 400132
rect 407172 400120 407178 400172
rect 20438 398828 20444 398880
rect 20496 398868 20502 398880
rect 46750 398868 46756 398880
rect 20496 398840 46756 398868
rect 20496 398828 20502 398840
rect 46750 398828 46756 398840
rect 46808 398828 46814 398880
rect 350442 398828 350448 398880
rect 350500 398868 350506 398880
rect 360470 398868 360476 398880
rect 350500 398840 360476 398868
rect 350500 398828 350506 398840
rect 360470 398828 360476 398840
rect 360528 398828 360534 398880
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 17402 397508 17408 397520
rect 3568 397480 17408 397508
rect 3568 397468 3574 397480
rect 17402 397468 17408 397480
rect 17460 397468 17466 397520
rect 350442 397468 350448 397520
rect 350500 397508 350506 397520
rect 388714 397508 388720 397520
rect 350500 397480 388720 397508
rect 350500 397468 350506 397480
rect 388714 397468 388720 397480
rect 388772 397468 388778 397520
rect 392946 397468 392952 397520
rect 393004 397508 393010 397520
rect 407114 397508 407120 397520
rect 393004 397480 407120 397508
rect 393004 397468 393010 397480
rect 407114 397468 407120 397480
rect 407172 397468 407178 397520
rect 349798 396788 349804 396840
rect 349856 396828 349862 396840
rect 352650 396828 352656 396840
rect 349856 396800 352656 396828
rect 349856 396788 349862 396800
rect 352650 396788 352656 396800
rect 352708 396788 352714 396840
rect 350442 396040 350448 396092
rect 350500 396080 350506 396092
rect 382734 396080 382740 396092
rect 350500 396052 382740 396080
rect 350500 396040 350506 396052
rect 382734 396040 382740 396052
rect 382792 396040 382798 396092
rect 349890 395972 349896 396024
rect 349948 396012 349954 396024
rect 351178 396012 351184 396024
rect 349948 395984 351184 396012
rect 349948 395972 349954 395984
rect 351178 395972 351184 395984
rect 351236 395972 351242 396024
rect 400030 394748 400036 394800
rect 400088 394788 400094 394800
rect 407206 394788 407212 394800
rect 400088 394760 407212 394788
rect 400088 394748 400094 394760
rect 407206 394748 407212 394760
rect 407264 394748 407270 394800
rect 20530 394680 20536 394732
rect 20588 394720 20594 394732
rect 46750 394720 46756 394732
rect 20588 394692 46756 394720
rect 20588 394680 20594 394692
rect 46750 394680 46756 394692
rect 46808 394680 46814 394732
rect 350258 394680 350264 394732
rect 350316 394720 350322 394732
rect 352834 394720 352840 394732
rect 350316 394692 352840 394720
rect 350316 394680 350322 394692
rect 352834 394680 352840 394692
rect 352892 394680 352898 394732
rect 382182 394680 382188 394732
rect 382240 394720 382246 394732
rect 407114 394720 407120 394732
rect 382240 394692 407120 394720
rect 382240 394680 382246 394692
rect 407114 394680 407120 394692
rect 407172 394680 407178 394732
rect 553026 394680 553032 394732
rect 553084 394720 553090 394732
rect 581730 394720 581736 394732
rect 553084 394692 581736 394720
rect 553084 394680 553090 394692
rect 581730 394680 581736 394692
rect 581788 394680 581794 394732
rect 350442 394612 350448 394664
rect 350500 394652 350506 394664
rect 392854 394652 392860 394664
rect 350500 394624 392860 394652
rect 350500 394612 350506 394624
rect 392854 394612 392860 394624
rect 392912 394612 392918 394664
rect 552198 393728 552204 393780
rect 552256 393768 552262 393780
rect 554958 393768 554964 393780
rect 552256 393740 554964 393768
rect 552256 393728 552262 393740
rect 554958 393728 554964 393740
rect 555016 393728 555022 393780
rect 390094 393320 390100 393372
rect 390152 393360 390158 393372
rect 407114 393360 407120 393372
rect 390152 393332 407120 393360
rect 390152 393320 390158 393332
rect 407114 393320 407120 393332
rect 407172 393320 407178 393372
rect 37918 392028 37924 392080
rect 37976 392068 37982 392080
rect 46014 392068 46020 392080
rect 37976 392040 46020 392068
rect 37976 392028 37982 392040
rect 46014 392028 46020 392040
rect 46072 392028 46078 392080
rect 25682 391960 25688 392012
rect 25740 392000 25746 392012
rect 46106 392000 46112 392012
rect 25740 391972 46112 392000
rect 25740 391960 25746 391972
rect 46106 391960 46112 391972
rect 46164 391960 46170 392012
rect 348878 391960 348884 392012
rect 348936 392000 348942 392012
rect 349338 392000 349344 392012
rect 348936 391972 349344 392000
rect 348936 391960 348942 391972
rect 349338 391960 349344 391972
rect 349396 391960 349402 392012
rect 350442 391960 350448 392012
rect 350500 392000 350506 392012
rect 402422 392000 402428 392012
rect 350500 391972 402428 392000
rect 350500 391960 350506 391972
rect 402422 391960 402428 391972
rect 402480 391960 402486 392012
rect 377858 390600 377864 390652
rect 377916 390640 377922 390652
rect 407206 390640 407212 390652
rect 377916 390612 407212 390640
rect 377916 390600 377922 390612
rect 407206 390600 407212 390612
rect 407264 390600 407270 390652
rect 553026 390600 553032 390652
rect 553084 390640 553090 390652
rect 581638 390640 581644 390652
rect 553084 390612 581644 390640
rect 553084 390600 553090 390612
rect 581638 390600 581644 390612
rect 581696 390600 581702 390652
rect 349614 390532 349620 390584
rect 349672 390572 349678 390584
rect 351270 390572 351276 390584
rect 349672 390544 351276 390572
rect 349672 390532 349678 390544
rect 351270 390532 351276 390544
rect 351328 390532 351334 390584
rect 368106 390532 368112 390584
rect 368164 390572 368170 390584
rect 407114 390572 407120 390584
rect 368164 390544 407120 390572
rect 368164 390532 368170 390544
rect 407114 390532 407120 390544
rect 407172 390532 407178 390584
rect 350442 390464 350448 390516
rect 350500 390504 350506 390516
rect 395522 390504 395528 390516
rect 350500 390476 395528 390504
rect 350500 390464 350506 390476
rect 395522 390464 395528 390476
rect 395580 390464 395586 390516
rect 17770 389172 17776 389224
rect 17828 389212 17834 389224
rect 46474 389212 46480 389224
rect 17828 389184 46480 389212
rect 17828 389172 17834 389184
rect 46474 389172 46480 389184
rect 46532 389172 46538 389224
rect 350258 389172 350264 389224
rect 350316 389212 350322 389224
rect 373718 389212 373724 389224
rect 350316 389184 373724 389212
rect 350316 389172 350322 389184
rect 373718 389172 373724 389184
rect 373776 389172 373782 389224
rect 391750 389172 391756 389224
rect 391808 389212 391814 389224
rect 407114 389212 407120 389224
rect 391808 389184 407120 389212
rect 391808 389172 391814 389184
rect 407114 389172 407120 389184
rect 407172 389172 407178 389224
rect 553026 389172 553032 389224
rect 553084 389212 553090 389224
rect 570414 389212 570420 389224
rect 553084 389184 570420 389212
rect 553084 389172 553090 389184
rect 570414 389172 570420 389184
rect 570472 389172 570478 389224
rect 350442 387812 350448 387864
rect 350500 387852 350506 387864
rect 377950 387852 377956 387864
rect 350500 387824 377956 387852
rect 350500 387812 350506 387824
rect 377950 387812 377956 387824
rect 378008 387812 378014 387864
rect 553026 387812 553032 387864
rect 553084 387852 553090 387864
rect 579798 387852 579804 387864
rect 553084 387824 579804 387852
rect 553084 387812 553090 387824
rect 579798 387812 579804 387824
rect 579856 387812 579862 387864
rect 350258 387744 350264 387796
rect 350316 387784 350322 387796
rect 400950 387784 400956 387796
rect 350316 387756 400956 387784
rect 350316 387744 350322 387756
rect 400950 387744 400956 387756
rect 401008 387744 401014 387796
rect 29822 386384 29828 386436
rect 29880 386424 29886 386436
rect 46474 386424 46480 386436
rect 29880 386396 46480 386424
rect 29880 386384 29886 386396
rect 46474 386384 46480 386396
rect 46532 386384 46538 386436
rect 553026 386384 553032 386436
rect 553084 386424 553090 386436
rect 561030 386424 561036 386436
rect 553084 386396 561036 386424
rect 553084 386384 553090 386396
rect 561030 386384 561036 386396
rect 561088 386384 561094 386436
rect 32398 386316 32404 386368
rect 32456 386356 32462 386368
rect 46106 386356 46112 386368
rect 32456 386328 46112 386356
rect 32456 386316 32462 386328
rect 46106 386316 46112 386328
rect 46164 386316 46170 386368
rect 350442 386316 350448 386368
rect 350500 386356 350506 386368
rect 352190 386356 352196 386368
rect 350500 386328 352196 386356
rect 350500 386316 350506 386328
rect 352190 386316 352196 386328
rect 352248 386316 352254 386368
rect 368198 386316 368204 386368
rect 368256 386356 368262 386368
rect 407114 386356 407120 386368
rect 368256 386328 407120 386356
rect 368256 386316 368262 386328
rect 407114 386316 407120 386328
rect 407172 386316 407178 386368
rect 36170 385024 36176 385076
rect 36228 385064 36234 385076
rect 46474 385064 46480 385076
rect 36228 385036 46480 385064
rect 36228 385024 36234 385036
rect 46474 385024 46480 385036
rect 46532 385024 46538 385076
rect 553026 385024 553032 385076
rect 553084 385064 553090 385076
rect 562134 385064 562140 385076
rect 553084 385036 562140 385064
rect 553084 385024 553090 385036
rect 562134 385024 562140 385036
rect 562192 385024 562198 385076
rect 349062 384956 349068 385008
rect 349120 384996 349126 385008
rect 352650 384996 352656 385008
rect 349120 384968 352656 384996
rect 349120 384956 349126 384968
rect 352650 384956 352656 384968
rect 352708 384956 352714 385008
rect 350442 384276 350448 384328
rect 350500 384316 350506 384328
rect 359274 384316 359280 384328
rect 350500 384288 359280 384316
rect 350500 384276 350506 384288
rect 359274 384276 359280 384288
rect 359332 384276 359338 384328
rect 403158 383936 403164 383988
rect 403216 383976 403222 383988
rect 407114 383976 407120 383988
rect 403216 383948 407120 383976
rect 403216 383936 403222 383948
rect 407114 383936 407120 383948
rect 407172 383936 407178 383988
rect 36722 383596 36728 383648
rect 36780 383636 36786 383648
rect 46474 383636 46480 383648
rect 36780 383608 46480 383636
rect 36780 383596 36786 383608
rect 46474 383596 46480 383608
rect 46532 383596 46538 383648
rect 350258 382236 350264 382288
rect 350316 382276 350322 382288
rect 400950 382276 400956 382288
rect 350316 382248 400956 382276
rect 350316 382236 350322 382248
rect 400950 382236 400956 382248
rect 401008 382236 401014 382288
rect 402514 382236 402520 382288
rect 402572 382276 402578 382288
rect 407114 382276 407120 382288
rect 402572 382248 407120 382276
rect 402572 382236 402578 382248
rect 407114 382236 407120 382248
rect 407172 382236 407178 382288
rect 553026 381488 553032 381540
rect 553084 381528 553090 381540
rect 558086 381528 558092 381540
rect 553084 381500 558092 381528
rect 553084 381488 553090 381500
rect 558086 381488 558092 381500
rect 558144 381488 558150 381540
rect 46474 381080 46480 381132
rect 46532 381120 46538 381132
rect 46842 381120 46848 381132
rect 46532 381092 46848 381120
rect 46532 381080 46538 381092
rect 46842 381080 46848 381092
rect 46900 381080 46906 381132
rect 36446 380944 36452 380996
rect 36504 380984 36510 380996
rect 45002 380984 45008 380996
rect 36504 380956 45008 380984
rect 36504 380944 36510 380956
rect 45002 380944 45008 380956
rect 45060 380944 45066 380996
rect 350074 380944 350080 380996
rect 350132 380984 350138 380996
rect 380894 380984 380900 380996
rect 350132 380956 380900 380984
rect 350132 380944 350138 380956
rect 380894 380944 380900 380956
rect 380952 380944 380958 380996
rect 28442 380876 28448 380928
rect 28500 380916 28506 380928
rect 46842 380916 46848 380928
rect 28500 380888 46848 380916
rect 28500 380876 28506 380888
rect 46842 380876 46848 380888
rect 46900 380876 46906 380928
rect 350258 380876 350264 380928
rect 350316 380916 350322 380928
rect 385586 380916 385592 380928
rect 350316 380888 385592 380916
rect 350316 380876 350322 380888
rect 385586 380876 385592 380888
rect 385644 380876 385650 380928
rect 395522 380876 395528 380928
rect 395580 380916 395586 380928
rect 407114 380916 407120 380928
rect 395580 380888 407120 380916
rect 395580 380876 395586 380888
rect 407114 380876 407120 380888
rect 407172 380876 407178 380928
rect 31294 379516 31300 379568
rect 31352 379556 31358 379568
rect 46842 379556 46848 379568
rect 31352 379528 46848 379556
rect 31352 379516 31358 379528
rect 46842 379516 46848 379528
rect 46900 379516 46906 379568
rect 408126 378768 408132 378820
rect 408184 378808 408190 378820
rect 409322 378808 409328 378820
rect 408184 378780 409328 378808
rect 408184 378768 408190 378780
rect 409322 378768 409328 378780
rect 409380 378768 409386 378820
rect 553026 378292 553032 378344
rect 553084 378332 553090 378344
rect 557902 378332 557908 378344
rect 553084 378304 557908 378332
rect 553084 378292 553090 378304
rect 557902 378292 557908 378304
rect 557960 378292 557966 378344
rect 392854 378156 392860 378208
rect 392912 378196 392918 378208
rect 407114 378196 407120 378208
rect 392912 378168 407120 378196
rect 392912 378156 392918 378168
rect 407114 378156 407120 378168
rect 407172 378156 407178 378208
rect 572070 378156 572076 378208
rect 572128 378196 572134 378208
rect 580166 378196 580172 378208
rect 572128 378168 580172 378196
rect 572128 378156 572134 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 350074 378088 350080 378140
rect 350132 378128 350138 378140
rect 352558 378128 352564 378140
rect 350132 378100 352564 378128
rect 350132 378088 350138 378100
rect 352558 378088 352564 378100
rect 352616 378088 352622 378140
rect 350258 376728 350264 376780
rect 350316 376768 350322 376780
rect 408494 376768 408500 376780
rect 350316 376740 408500 376768
rect 350316 376728 350322 376740
rect 408494 376728 408500 376740
rect 408552 376728 408558 376780
rect 553026 376728 553032 376780
rect 553084 376768 553090 376780
rect 582834 376768 582840 376780
rect 553084 376740 582840 376768
rect 553084 376728 553090 376740
rect 582834 376728 582840 376740
rect 582892 376728 582898 376780
rect 350074 375368 350080 375420
rect 350132 375408 350138 375420
rect 403710 375408 403716 375420
rect 350132 375380 403716 375408
rect 350132 375368 350138 375380
rect 403710 375368 403716 375380
rect 403768 375368 403774 375420
rect 350258 375300 350264 375352
rect 350316 375340 350322 375352
rect 374914 375340 374920 375352
rect 350316 375312 374920 375340
rect 350316 375300 350322 375312
rect 374914 375300 374920 375312
rect 374972 375300 374978 375352
rect 552198 372648 552204 372700
rect 552256 372688 552262 372700
rect 555050 372688 555056 372700
rect 552256 372660 555056 372688
rect 552256 372648 552262 372660
rect 555050 372648 555056 372660
rect 555108 372648 555114 372700
rect 28258 372580 28264 372632
rect 28316 372620 28322 372632
rect 46842 372620 46848 372632
rect 28316 372592 46848 372620
rect 28316 372580 28322 372592
rect 46842 372580 46848 372592
rect 46900 372580 46906 372632
rect 350258 372580 350264 372632
rect 350316 372620 350322 372632
rect 374914 372620 374920 372632
rect 350316 372592 374920 372620
rect 350316 372580 350322 372592
rect 374914 372580 374920 372592
rect 374972 372580 374978 372632
rect 397086 372580 397092 372632
rect 397144 372620 397150 372632
rect 407114 372620 407120 372632
rect 397144 372592 407120 372620
rect 397144 372580 397150 372592
rect 407114 372580 407120 372592
rect 407172 372580 407178 372632
rect 29730 371220 29736 371272
rect 29788 371260 29794 371272
rect 46842 371260 46848 371272
rect 29788 371232 46848 371260
rect 29788 371220 29794 371232
rect 46842 371220 46848 371232
rect 46900 371220 46906 371272
rect 350258 371220 350264 371272
rect 350316 371260 350322 371272
rect 380710 371260 380716 371272
rect 350316 371232 380716 371260
rect 350316 371220 350322 371232
rect 380710 371220 380716 371232
rect 380768 371220 380774 371272
rect 43806 371152 43812 371204
rect 43864 371192 43870 371204
rect 45646 371192 45652 371204
rect 43864 371164 45652 371192
rect 43864 371152 43870 371164
rect 45646 371152 45652 371164
rect 45704 371152 45710 371204
rect 350074 371152 350080 371204
rect 350132 371192 350138 371204
rect 356422 371192 356428 371204
rect 350132 371164 356428 371192
rect 350132 371152 350138 371164
rect 356422 371152 356428 371164
rect 356480 371152 356486 371204
rect 362494 371152 362500 371204
rect 362552 371192 362558 371204
rect 407114 371192 407120 371204
rect 362552 371164 407120 371192
rect 362552 371152 362558 371164
rect 407114 371152 407120 371164
rect 407172 371152 407178 371204
rect 553026 369860 553032 369912
rect 553084 369900 553090 369912
rect 560662 369900 560668 369912
rect 553084 369872 560668 369900
rect 553084 369860 553090 369872
rect 560662 369860 560668 369872
rect 560720 369860 560726 369912
rect 407666 369112 407672 369164
rect 407724 369152 407730 369164
rect 408126 369152 408132 369164
rect 407724 369124 408132 369152
rect 407724 369112 407730 369124
rect 408126 369112 408132 369124
rect 408184 369112 408190 369164
rect 552198 368568 552204 368620
rect 552256 368608 552262 368620
rect 555418 368608 555424 368620
rect 552256 368580 555424 368608
rect 552256 368568 552262 368580
rect 555418 368568 555424 368580
rect 555476 368568 555482 368620
rect 43806 368500 43812 368552
rect 43864 368540 43870 368552
rect 46842 368540 46848 368552
rect 43864 368512 46848 368540
rect 43864 368500 43870 368512
rect 46842 368500 46848 368512
rect 46900 368500 46906 368552
rect 553026 368500 553032 368552
rect 553084 368540 553090 368552
rect 572990 368540 572996 368552
rect 553084 368512 572996 368540
rect 553084 368500 553090 368512
rect 572990 368500 572996 368512
rect 573048 368500 573054 368552
rect 349062 368432 349068 368484
rect 349120 368472 349126 368484
rect 349338 368472 349344 368484
rect 349120 368444 349344 368472
rect 349120 368432 349126 368444
rect 349338 368432 349344 368444
rect 349396 368432 349402 368484
rect 552014 367956 552020 368008
rect 552072 367996 552078 368008
rect 553762 367996 553768 368008
rect 552072 367968 553768 367996
rect 552072 367956 552078 367968
rect 553762 367956 553768 367968
rect 553820 367956 553826 368008
rect 32122 367072 32128 367124
rect 32180 367112 32186 367124
rect 46842 367112 46848 367124
rect 32180 367084 46848 367112
rect 32180 367072 32186 367084
rect 46842 367072 46848 367084
rect 46900 367072 46906 367124
rect 32766 367004 32772 367056
rect 32824 367044 32830 367056
rect 46014 367044 46020 367056
rect 32824 367016 46020 367044
rect 32824 367004 32830 367016
rect 46014 367004 46020 367016
rect 46072 367004 46078 367056
rect 553026 365780 553032 365832
rect 553084 365820 553090 365832
rect 567562 365820 567568 365832
rect 553084 365792 567568 365820
rect 553084 365780 553090 365792
rect 567562 365780 567568 365792
rect 567620 365780 567626 365832
rect 552934 365712 552940 365764
rect 552992 365752 552998 365764
rect 578418 365752 578424 365764
rect 552992 365724 578424 365752
rect 552992 365712 552998 365724
rect 578418 365712 578424 365724
rect 578476 365712 578482 365764
rect 552014 365168 552020 365220
rect 552072 365208 552078 365220
rect 554130 365208 554136 365220
rect 552072 365180 554136 365208
rect 552072 365168 552078 365180
rect 554130 365168 554136 365180
rect 554188 365168 554194 365220
rect 27154 362924 27160 362976
rect 27212 362964 27218 362976
rect 46842 362964 46848 362976
rect 27212 362936 46848 362964
rect 27212 362924 27218 362936
rect 46842 362924 46848 362936
rect 46900 362924 46906 362976
rect 350074 362924 350080 362976
rect 350132 362964 350138 362976
rect 352558 362964 352564 362976
rect 350132 362936 352564 362964
rect 350132 362924 350138 362936
rect 352558 362924 352564 362936
rect 352616 362924 352622 362976
rect 45278 361496 45284 361548
rect 45336 361536 45342 361548
rect 46474 361536 46480 361548
rect 45336 361508 46480 361536
rect 45336 361496 45342 361508
rect 46474 361496 46480 361508
rect 46532 361496 46538 361548
rect 370774 361496 370780 361548
rect 370832 361536 370838 361548
rect 407114 361536 407120 361548
rect 370832 361508 407120 361536
rect 370832 361496 370838 361508
rect 407114 361496 407120 361508
rect 407172 361496 407178 361548
rect 553026 360408 553032 360460
rect 553084 360448 553090 360460
rect 557902 360448 557908 360460
rect 553084 360420 557908 360448
rect 553084 360408 553090 360420
rect 557902 360408 557908 360420
rect 557960 360408 557966 360460
rect 366634 360204 366640 360256
rect 366692 360244 366698 360256
rect 407114 360244 407120 360256
rect 366692 360216 407120 360244
rect 366692 360204 366698 360216
rect 407114 360204 407120 360216
rect 407172 360204 407178 360256
rect 552934 360204 552940 360256
rect 552992 360244 552998 360256
rect 574738 360244 574744 360256
rect 552992 360216 574744 360244
rect 552992 360204 552998 360216
rect 574738 360204 574744 360216
rect 574796 360204 574802 360256
rect 350258 358776 350264 358828
rect 350316 358816 350322 358828
rect 363138 358816 363144 358828
rect 350316 358788 363144 358816
rect 350316 358776 350322 358788
rect 363138 358776 363144 358788
rect 363196 358776 363202 358828
rect 37826 358708 37832 358760
rect 37884 358748 37890 358760
rect 46842 358748 46848 358760
rect 37884 358720 46848 358748
rect 37884 358708 37890 358720
rect 46842 358708 46848 358720
rect 46900 358708 46906 358760
rect 553026 358708 553032 358760
rect 553084 358748 553090 358760
rect 572070 358748 572076 358760
rect 553084 358720 572076 358748
rect 553084 358708 553090 358720
rect 572070 358708 572076 358720
rect 572128 358708 572134 358760
rect 350258 357960 350264 358012
rect 350316 358000 350322 358012
rect 355502 358000 355508 358012
rect 350316 357972 355508 358000
rect 350316 357960 350322 357972
rect 355502 357960 355508 357972
rect 355560 357960 355566 358012
rect 46474 357756 46480 357808
rect 46532 357796 46538 357808
rect 46842 357796 46848 357808
rect 46532 357768 46848 357796
rect 46532 357756 46538 357768
rect 46842 357756 46848 357768
rect 46900 357756 46906 357808
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 28074 357456 28080 357468
rect 3200 357428 28080 357456
rect 3200 357416 3206 357428
rect 28074 357416 28080 357428
rect 28132 357416 28138 357468
rect 552934 357416 552940 357468
rect 552992 357456 552998 357468
rect 573266 357456 573272 357468
rect 552992 357428 573272 357456
rect 552992 357416 552998 357428
rect 573266 357416 573272 357428
rect 573324 357416 573330 357468
rect 369670 356192 369676 356244
rect 369728 356232 369734 356244
rect 407114 356232 407120 356244
rect 369728 356204 407120 356232
rect 369728 356192 369734 356204
rect 407114 356192 407120 356204
rect 407172 356192 407178 356244
rect 350258 356124 350264 356176
rect 350316 356164 350322 356176
rect 378226 356164 378232 356176
rect 350316 356136 378232 356164
rect 350316 356124 350322 356136
rect 378226 356124 378232 356136
rect 378284 356124 378290 356176
rect 350258 355988 350264 356040
rect 350316 356028 350322 356040
rect 396810 356028 396816 356040
rect 350316 356000 396816 356028
rect 350316 355988 350322 356000
rect 396810 355988 396816 356000
rect 396868 355988 396874 356040
rect 37826 354696 37832 354748
rect 37884 354736 37890 354748
rect 46474 354736 46480 354748
rect 37884 354708 46480 354736
rect 37884 354696 37890 354708
rect 46474 354696 46480 354708
rect 46532 354696 46538 354748
rect 350258 354696 350264 354748
rect 350316 354736 350322 354748
rect 359642 354736 359648 354748
rect 350316 354708 359648 354736
rect 350316 354696 350322 354708
rect 359642 354696 359648 354708
rect 359700 354696 359706 354748
rect 553026 354696 553032 354748
rect 553084 354736 553090 354748
rect 568114 354736 568120 354748
rect 553084 354708 568120 354736
rect 553084 354696 553090 354708
rect 568114 354696 568120 354708
rect 568172 354696 568178 354748
rect 376386 353268 376392 353320
rect 376444 353308 376450 353320
rect 407114 353308 407120 353320
rect 376444 353280 407120 353308
rect 376444 353268 376450 353280
rect 407114 353268 407120 353280
rect 407172 353268 407178 353320
rect 553026 353268 553032 353320
rect 553084 353308 553090 353320
rect 575842 353308 575848 353320
rect 553084 353280 575848 353308
rect 553084 353268 553090 353280
rect 575842 353268 575848 353280
rect 575900 353268 575906 353320
rect 36538 353200 36544 353252
rect 36596 353240 36602 353252
rect 46474 353240 46480 353252
rect 36596 353212 46480 353240
rect 36596 353200 36602 353212
rect 46474 353200 46480 353212
rect 46532 353200 46538 353252
rect 398834 351976 398840 352028
rect 398892 352016 398898 352028
rect 407114 352016 407120 352028
rect 398892 351988 407120 352016
rect 398892 351976 398898 351988
rect 407114 351976 407120 351988
rect 407172 351976 407178 352028
rect 388806 351908 388812 351960
rect 388864 351948 388870 351960
rect 407206 351948 407212 351960
rect 388864 351920 407212 351948
rect 388864 351908 388870 351920
rect 407206 351908 407212 351920
rect 407264 351908 407270 351960
rect 553118 350888 553124 350940
rect 553176 350928 553182 350940
rect 558178 350928 558184 350940
rect 553176 350900 558184 350928
rect 553176 350888 553182 350900
rect 558178 350888 558184 350900
rect 558236 350888 558242 350940
rect 350258 350548 350264 350600
rect 350316 350588 350322 350600
rect 362034 350588 362040 350600
rect 350316 350560 362040 350588
rect 350316 350548 350322 350560
rect 362034 350548 362040 350560
rect 362092 350548 362098 350600
rect 384850 350548 384856 350600
rect 384908 350588 384914 350600
rect 407114 350588 407120 350600
rect 384908 350560 407120 350588
rect 384908 350548 384914 350560
rect 407114 350548 407120 350560
rect 407172 350548 407178 350600
rect 552842 350548 552848 350600
rect 552900 350588 552906 350600
rect 583018 350588 583024 350600
rect 552900 350560 583024 350588
rect 552900 350548 552906 350560
rect 583018 350548 583024 350560
rect 583076 350548 583082 350600
rect 350074 349188 350080 349240
rect 350132 349228 350138 349240
rect 364058 349228 364064 349240
rect 350132 349200 364064 349228
rect 350132 349188 350138 349200
rect 364058 349188 364064 349200
rect 364116 349188 364122 349240
rect 21542 349120 21548 349172
rect 21600 349160 21606 349172
rect 46474 349160 46480 349172
rect 21600 349132 46480 349160
rect 21600 349120 21606 349132
rect 46474 349120 46480 349132
rect 46532 349120 46538 349172
rect 350258 349120 350264 349172
rect 350316 349160 350322 349172
rect 365438 349160 365444 349172
rect 350316 349132 365444 349160
rect 350316 349120 350322 349132
rect 365438 349120 365444 349132
rect 365496 349120 365502 349172
rect 372430 349120 372436 349172
rect 372488 349160 372494 349172
rect 407114 349160 407120 349172
rect 372488 349132 407120 349160
rect 372488 349120 372494 349132
rect 407114 349120 407120 349132
rect 407172 349120 407178 349172
rect 553118 349120 553124 349172
rect 553176 349160 553182 349172
rect 583478 349160 583484 349172
rect 553176 349132 583484 349160
rect 553176 349120 553182 349132
rect 583478 349120 583484 349132
rect 583536 349120 583542 349172
rect 553118 346468 553124 346520
rect 553176 346508 553182 346520
rect 575750 346508 575756 346520
rect 553176 346480 575756 346508
rect 553176 346468 553182 346480
rect 575750 346468 575756 346480
rect 575808 346468 575814 346520
rect 29546 346400 29552 346452
rect 29604 346440 29610 346452
rect 46474 346440 46480 346452
rect 29604 346412 46480 346440
rect 29604 346400 29610 346412
rect 46474 346400 46480 346412
rect 46532 346400 46538 346452
rect 392394 346400 392400 346452
rect 392452 346440 392458 346452
rect 407114 346440 407120 346452
rect 392452 346412 407120 346440
rect 392452 346400 392458 346412
rect 407114 346400 407120 346412
rect 407172 346400 407178 346452
rect 553026 346400 553032 346452
rect 553084 346440 553090 346452
rect 578694 346440 578700 346452
rect 553084 346412 578700 346440
rect 553084 346400 553090 346412
rect 578694 346400 578700 346412
rect 578752 346400 578758 346452
rect 3510 345108 3516 345160
rect 3568 345148 3574 345160
rect 29454 345148 29460 345160
rect 3568 345120 29460 345148
rect 3568 345108 3574 345120
rect 29454 345108 29460 345120
rect 29512 345108 29518 345160
rect 20346 345040 20352 345092
rect 20404 345080 20410 345092
rect 46474 345080 46480 345092
rect 20404 345052 46480 345080
rect 20404 345040 20410 345052
rect 46474 345040 46480 345052
rect 46532 345040 46538 345092
rect 350258 345040 350264 345092
rect 350316 345080 350322 345092
rect 379606 345080 379612 345092
rect 350316 345052 379612 345080
rect 350316 345040 350322 345052
rect 379606 345040 379612 345052
rect 379664 345040 379670 345092
rect 376570 344972 376576 345024
rect 376628 345012 376634 345024
rect 407114 345012 407120 345024
rect 376628 344984 407120 345012
rect 376628 344972 376634 344984
rect 407114 344972 407120 344984
rect 407172 344972 407178 345024
rect 350258 343680 350264 343732
rect 350316 343720 350322 343732
rect 361298 343720 361304 343732
rect 350316 343692 361304 343720
rect 350316 343680 350322 343692
rect 361298 343680 361304 343692
rect 361356 343680 361362 343732
rect 350074 343612 350080 343664
rect 350132 343652 350138 343664
rect 382826 343652 382832 343664
rect 350132 343624 382832 343652
rect 350132 343612 350138 343624
rect 382826 343612 382832 343624
rect 382884 343612 382890 343664
rect 553026 343000 553032 343052
rect 553084 343040 553090 343052
rect 556706 343040 556712 343052
rect 553084 343012 556712 343040
rect 553084 343000 553090 343012
rect 556706 343000 556712 343012
rect 556764 343000 556770 343052
rect 552014 342796 552020 342848
rect 552072 342836 552078 342848
rect 553670 342836 553676 342848
rect 552072 342808 553676 342836
rect 552072 342796 552078 342808
rect 553670 342796 553676 342808
rect 553728 342796 553734 342848
rect 398006 342252 398012 342304
rect 398064 342292 398070 342304
rect 407114 342292 407120 342304
rect 398064 342264 407120 342292
rect 398064 342252 398070 342264
rect 407114 342252 407120 342264
rect 407172 342252 407178 342304
rect 370774 339464 370780 339516
rect 370832 339504 370838 339516
rect 407114 339504 407120 339516
rect 370832 339476 407120 339504
rect 370832 339464 370838 339476
rect 407114 339464 407120 339476
rect 407172 339464 407178 339516
rect 391658 338104 391664 338156
rect 391716 338144 391722 338156
rect 407114 338144 407120 338156
rect 391716 338116 407120 338144
rect 391716 338104 391722 338116
rect 407114 338104 407120 338116
rect 407172 338104 407178 338156
rect 553118 338104 553124 338156
rect 553176 338144 553182 338156
rect 569218 338144 569224 338156
rect 553176 338116 569224 338144
rect 553176 338104 553182 338116
rect 569218 338104 569224 338116
rect 569276 338104 569282 338156
rect 25406 336744 25412 336796
rect 25464 336784 25470 336796
rect 46474 336784 46480 336796
rect 25464 336756 46480 336784
rect 25464 336744 25470 336756
rect 46474 336744 46480 336756
rect 46532 336744 46538 336796
rect 372246 336676 372252 336728
rect 372304 336716 372310 336728
rect 407114 336716 407120 336728
rect 372304 336688 407120 336716
rect 372304 336676 372310 336688
rect 407114 336676 407120 336688
rect 407172 336676 407178 336728
rect 553026 335316 553032 335368
rect 553084 335356 553090 335368
rect 566458 335356 566464 335368
rect 553084 335328 566464 335356
rect 553084 335316 553090 335328
rect 566458 335316 566464 335328
rect 566516 335316 566522 335368
rect 553118 335248 553124 335300
rect 553176 335288 553182 335300
rect 566182 335288 566188 335300
rect 553176 335260 566188 335288
rect 553176 335248 553182 335260
rect 566182 335248 566188 335260
rect 566240 335248 566246 335300
rect 350350 334024 350356 334076
rect 350408 334064 350414 334076
rect 357066 334064 357072 334076
rect 350408 334036 357072 334064
rect 350408 334024 350414 334036
rect 357066 334024 357072 334036
rect 357124 334024 357130 334076
rect 350350 332596 350356 332648
rect 350408 332636 350414 332648
rect 359274 332636 359280 332648
rect 350408 332608 359280 332636
rect 350408 332596 350414 332608
rect 359274 332596 359280 332608
rect 359332 332596 359338 332648
rect 32674 331168 32680 331220
rect 32732 331208 32738 331220
rect 46474 331208 46480 331220
rect 32732 331180 46480 331208
rect 32732 331168 32738 331180
rect 46474 331168 46480 331180
rect 46532 331168 46538 331220
rect 350350 329808 350356 329860
rect 350408 329848 350414 329860
rect 374086 329848 374092 329860
rect 350408 329820 374092 329848
rect 350408 329808 350414 329820
rect 374086 329808 374092 329820
rect 374144 329808 374150 329860
rect 400766 329808 400772 329860
rect 400824 329848 400830 329860
rect 407114 329848 407120 329860
rect 400824 329820 407120 329848
rect 400824 329808 400830 329820
rect 407114 329808 407120 329820
rect 407172 329808 407178 329860
rect 31018 328448 31024 328500
rect 31076 328488 31082 328500
rect 46474 328488 46480 328500
rect 31076 328460 46480 328488
rect 31076 328448 31082 328460
rect 46474 328448 46480 328460
rect 46532 328448 46538 328500
rect 350350 328448 350356 328500
rect 350408 328488 350414 328500
rect 370866 328488 370872 328500
rect 350408 328460 370872 328488
rect 350408 328448 350414 328460
rect 370866 328448 370872 328460
rect 370924 328448 370930 328500
rect 379238 328448 379244 328500
rect 379296 328488 379302 328500
rect 407114 328488 407120 328500
rect 379296 328460 407120 328488
rect 379296 328448 379302 328460
rect 407114 328448 407120 328460
rect 407172 328448 407178 328500
rect 553026 327156 553032 327208
rect 553084 327196 553090 327208
rect 570506 327196 570512 327208
rect 553084 327168 570512 327196
rect 553084 327156 553090 327168
rect 570506 327156 570512 327168
rect 570564 327156 570570 327208
rect 362494 327088 362500 327140
rect 362552 327128 362558 327140
rect 407114 327128 407120 327140
rect 362552 327100 407120 327128
rect 362552 327088 362558 327100
rect 407114 327088 407120 327100
rect 407172 327088 407178 327140
rect 553118 327088 553124 327140
rect 553176 327128 553182 327140
rect 578786 327128 578792 327140
rect 553176 327100 578792 327128
rect 553176 327088 553182 327100
rect 578786 327088 578792 327100
rect 578844 327088 578850 327140
rect 46290 327020 46296 327072
rect 46348 327060 46354 327072
rect 46934 327060 46940 327072
rect 46348 327032 46940 327060
rect 46348 327020 46354 327032
rect 46934 327020 46940 327032
rect 46992 327020 46998 327072
rect 553026 325728 553032 325780
rect 553084 325768 553090 325780
rect 581362 325768 581368 325780
rect 553084 325740 581368 325768
rect 553084 325728 553090 325740
rect 581362 325728 581368 325740
rect 581420 325728 581426 325780
rect 350350 325660 350356 325712
rect 350408 325700 350414 325712
rect 364702 325700 364708 325712
rect 350408 325672 364708 325700
rect 350408 325660 350414 325672
rect 364702 325660 364708 325672
rect 364760 325660 364766 325712
rect 376570 325660 376576 325712
rect 376628 325700 376634 325712
rect 407114 325700 407120 325712
rect 376628 325672 407120 325700
rect 376628 325660 376634 325672
rect 407114 325660 407120 325672
rect 407172 325660 407178 325712
rect 553118 325660 553124 325712
rect 553176 325700 553182 325712
rect 583570 325700 583576 325712
rect 553176 325672 583576 325700
rect 553176 325660 553182 325672
rect 583570 325660 583576 325672
rect 583628 325660 583634 325712
rect 31202 325592 31208 325644
rect 31260 325632 31266 325644
rect 46474 325632 46480 325644
rect 31260 325604 46480 325632
rect 31260 325592 31266 325604
rect 46474 325592 46480 325604
rect 46532 325592 46538 325644
rect 370682 325592 370688 325644
rect 370740 325632 370746 325644
rect 407206 325632 407212 325644
rect 370740 325604 407212 325632
rect 370740 325592 370746 325604
rect 407206 325592 407212 325604
rect 407264 325592 407270 325644
rect 574922 325592 574928 325644
rect 574980 325632 574986 325644
rect 580166 325632 580172 325644
rect 574980 325604 580172 325632
rect 574980 325592 574986 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 43346 323484 43352 323536
rect 43404 323524 43410 323536
rect 44634 323524 44640 323536
rect 43404 323496 44640 323524
rect 43404 323484 43410 323496
rect 44634 323484 44640 323496
rect 44692 323484 44698 323536
rect 46290 323144 46296 323196
rect 46348 323184 46354 323196
rect 46842 323184 46848 323196
rect 46348 323156 46848 323184
rect 46348 323144 46354 323156
rect 46842 323144 46848 323156
rect 46900 323144 46906 323196
rect 399846 323008 399852 323060
rect 399904 323048 399910 323060
rect 407206 323048 407212 323060
rect 399904 323020 407212 323048
rect 399904 323008 399910 323020
rect 407206 323008 407212 323020
rect 407264 323008 407270 323060
rect 36538 322940 36544 322992
rect 36596 322980 36602 322992
rect 46842 322980 46848 322992
rect 36596 322952 46848 322980
rect 36596 322940 36602 322952
rect 46842 322940 46848 322952
rect 46900 322940 46906 322992
rect 373902 322940 373908 322992
rect 373960 322980 373966 322992
rect 407114 322980 407120 322992
rect 373960 322952 407120 322980
rect 373960 322940 373966 322952
rect 407114 322940 407120 322952
rect 407172 322940 407178 322992
rect 44910 322872 44916 322924
rect 44968 322912 44974 322924
rect 45738 322912 45744 322924
rect 44968 322884 45744 322912
rect 44968 322872 44974 322884
rect 45738 322872 45744 322884
rect 45796 322872 45802 322924
rect 358630 322872 358636 322924
rect 358688 322912 358694 322924
rect 407206 322912 407212 322924
rect 358688 322884 407212 322912
rect 358688 322872 358694 322884
rect 407206 322872 407212 322884
rect 407264 322872 407270 322924
rect 364702 322804 364708 322856
rect 364760 322844 364766 322856
rect 407114 322844 407120 322856
rect 364760 322816 407120 322844
rect 364760 322804 364766 322816
rect 407114 322804 407120 322816
rect 407172 322804 407178 322856
rect 552014 322328 552020 322380
rect 552072 322368 552078 322380
rect 553670 322368 553676 322380
rect 552072 322340 553676 322368
rect 552072 322328 552078 322340
rect 553670 322328 553676 322340
rect 553728 322328 553734 322380
rect 43346 321580 43352 321632
rect 43404 321620 43410 321632
rect 46842 321620 46848 321632
rect 43404 321592 46848 321620
rect 43404 321580 43410 321592
rect 46842 321580 46848 321592
rect 46900 321580 46906 321632
rect 350350 321580 350356 321632
rect 350408 321620 350414 321632
rect 373166 321620 373172 321632
rect 350408 321592 373172 321620
rect 350408 321580 350414 321592
rect 373166 321580 373172 321592
rect 373224 321580 373230 321632
rect 42242 321512 42248 321564
rect 42300 321552 42306 321564
rect 46474 321552 46480 321564
rect 42300 321524 46480 321552
rect 42300 321512 42306 321524
rect 46474 321512 46480 321524
rect 46532 321512 46538 321564
rect 32398 320152 32404 320204
rect 32456 320192 32462 320204
rect 46842 320192 46848 320204
rect 32456 320164 46848 320192
rect 32456 320152 32462 320164
rect 46842 320152 46848 320164
rect 46900 320152 46906 320204
rect 350350 320152 350356 320204
rect 350408 320192 350414 320204
rect 379330 320192 379336 320204
rect 350408 320164 379336 320192
rect 350408 320152 350414 320164
rect 379330 320152 379336 320164
rect 379388 320152 379394 320204
rect 405090 320152 405096 320204
rect 405148 320192 405154 320204
rect 407298 320192 407304 320204
rect 405148 320164 407304 320192
rect 405148 320152 405154 320164
rect 407298 320152 407304 320164
rect 407356 320152 407362 320204
rect 350258 320084 350264 320136
rect 350316 320124 350322 320136
rect 383286 320124 383292 320136
rect 350316 320096 383292 320124
rect 350316 320084 350322 320096
rect 383286 320084 383292 320096
rect 383344 320084 383350 320136
rect 42242 318928 42248 318980
rect 42300 318968 42306 318980
rect 46842 318968 46848 318980
rect 42300 318940 46848 318968
rect 42300 318928 42306 318940
rect 46842 318928 46848 318940
rect 46900 318928 46906 318980
rect 350350 318792 350356 318844
rect 350408 318832 350414 318844
rect 382642 318832 382648 318844
rect 350408 318804 382648 318832
rect 350408 318792 350414 318804
rect 382642 318792 382648 318804
rect 382700 318792 382706 318844
rect 552750 317568 552756 317620
rect 552808 317608 552814 317620
rect 559374 317608 559380 317620
rect 552808 317580 559380 317608
rect 552808 317568 552814 317580
rect 559374 317568 559380 317580
rect 559432 317568 559438 317620
rect 553118 317500 553124 317552
rect 553176 317540 553182 317552
rect 566182 317540 566188 317552
rect 553176 317512 566188 317540
rect 553176 317500 553182 317512
rect 566182 317500 566188 317512
rect 566240 317500 566246 317552
rect 350350 317432 350356 317484
rect 350408 317472 350414 317484
rect 370682 317472 370688 317484
rect 350408 317444 370688 317472
rect 350408 317432 350414 317444
rect 370682 317432 370688 317444
rect 370740 317432 370746 317484
rect 553026 317432 553032 317484
rect 553084 317472 553090 317484
rect 579982 317472 579988 317484
rect 553084 317444 579988 317472
rect 553084 317432 553090 317444
rect 579982 317432 579988 317444
rect 580040 317432 580046 317484
rect 553118 316004 553124 316056
rect 553176 316044 553182 316056
rect 576302 316044 576308 316056
rect 553176 316016 576308 316044
rect 553176 316004 553182 316016
rect 576302 316004 576308 316016
rect 576360 316004 576366 316056
rect 350350 315936 350356 315988
rect 350408 315976 350414 315988
rect 390094 315976 390100 315988
rect 350408 315948 390100 315976
rect 350408 315936 350414 315948
rect 390094 315936 390100 315948
rect 390152 315936 390158 315988
rect 25498 314644 25504 314696
rect 25556 314684 25562 314696
rect 46290 314684 46296 314696
rect 25556 314656 46296 314684
rect 25556 314644 25562 314656
rect 46290 314644 46296 314656
rect 46348 314644 46354 314696
rect 406194 314644 406200 314696
rect 406252 314684 406258 314696
rect 407114 314684 407120 314696
rect 406252 314656 407120 314684
rect 406252 314644 406258 314656
rect 407114 314644 407120 314656
rect 407172 314644 407178 314696
rect 553118 314644 553124 314696
rect 553176 314684 553182 314696
rect 571794 314684 571800 314696
rect 553176 314656 571800 314684
rect 553176 314644 553182 314656
rect 571794 314644 571800 314656
rect 571852 314644 571858 314696
rect 553026 313284 553032 313336
rect 553084 313324 553090 313336
rect 583110 313324 583116 313336
rect 553084 313296 583116 313324
rect 553084 313284 553090 313296
rect 583110 313284 583116 313296
rect 583168 313284 583174 313336
rect 553118 313216 553124 313268
rect 553176 313256 553182 313268
rect 566090 313256 566096 313268
rect 553176 313228 566096 313256
rect 553176 313216 553182 313228
rect 566090 313216 566096 313228
rect 566148 313216 566154 313268
rect 350350 311856 350356 311908
rect 350408 311896 350414 311908
rect 390278 311896 390284 311908
rect 350408 311868 390284 311896
rect 350408 311856 350414 311868
rect 390278 311856 390284 311868
rect 390336 311856 390342 311908
rect 403802 310564 403808 310616
rect 403860 310604 403866 310616
rect 407114 310604 407120 310616
rect 403860 310576 407120 310604
rect 403860 310564 403866 310576
rect 407114 310564 407120 310576
rect 407172 310564 407178 310616
rect 553118 310564 553124 310616
rect 553176 310604 553182 310616
rect 572070 310604 572076 310616
rect 553176 310576 572076 310604
rect 553176 310564 553182 310576
rect 572070 310564 572076 310576
rect 572128 310564 572134 310616
rect 28534 310496 28540 310548
rect 28592 310536 28598 310548
rect 46106 310536 46112 310548
rect 28592 310508 46112 310536
rect 28592 310496 28598 310508
rect 46106 310496 46112 310508
rect 46164 310496 46170 310548
rect 392486 310496 392492 310548
rect 392544 310536 392550 310548
rect 407206 310536 407212 310548
rect 392544 310508 407212 310536
rect 392544 310496 392550 310508
rect 407206 310496 407212 310508
rect 407264 310496 407270 310548
rect 553026 310496 553032 310548
rect 553084 310536 553090 310548
rect 573450 310536 573456 310548
rect 553084 310508 573456 310536
rect 553084 310496 553090 310508
rect 573450 310496 573456 310508
rect 573508 310496 573514 310548
rect 36630 310428 36636 310480
rect 36688 310468 36694 310480
rect 46290 310468 46296 310480
rect 36688 310440 46296 310468
rect 36688 310428 36694 310440
rect 46290 310428 46296 310440
rect 46348 310428 46354 310480
rect 350166 310428 350172 310480
rect 350224 310468 350230 310480
rect 350534 310468 350540 310480
rect 350224 310440 350540 310468
rect 350224 310428 350230 310440
rect 350534 310428 350540 310440
rect 350592 310428 350598 310480
rect 394142 310428 394148 310480
rect 394200 310468 394206 310480
rect 407114 310468 407120 310480
rect 394200 310440 407120 310468
rect 394200 310428 394206 310440
rect 407114 310428 407120 310440
rect 407172 310428 407178 310480
rect 33686 309136 33692 309188
rect 33744 309176 33750 309188
rect 46106 309176 46112 309188
rect 33744 309148 46112 309176
rect 33744 309136 33750 309148
rect 46106 309136 46112 309148
rect 46164 309136 46170 309188
rect 553118 309136 553124 309188
rect 553176 309176 553182 309188
rect 577406 309176 577412 309188
rect 553176 309148 577412 309176
rect 553176 309136 553182 309148
rect 577406 309136 577412 309148
rect 577464 309136 577470 309188
rect 375190 307844 375196 307896
rect 375248 307884 375254 307896
rect 407114 307884 407120 307896
rect 375248 307856 407120 307884
rect 375248 307844 375254 307856
rect 407114 307844 407120 307856
rect 407172 307844 407178 307896
rect 350350 307776 350356 307828
rect 350408 307816 350414 307828
rect 390094 307816 390100 307828
rect 350408 307788 390100 307816
rect 350408 307776 350414 307788
rect 390094 307776 390100 307788
rect 390152 307776 390158 307828
rect 553118 307776 553124 307828
rect 553176 307816 553182 307828
rect 575014 307816 575020 307828
rect 553176 307788 575020 307816
rect 553176 307776 553182 307788
rect 575014 307776 575020 307788
rect 575072 307776 575078 307828
rect 364058 307708 364064 307760
rect 364116 307748 364122 307760
rect 407114 307748 407120 307760
rect 364116 307720 407120 307748
rect 364116 307708 364122 307720
rect 407114 307708 407120 307720
rect 407172 307708 407178 307760
rect 407574 307436 407580 307488
rect 407632 307476 407638 307488
rect 407942 307476 407948 307488
rect 407632 307448 407948 307476
rect 407632 307436 407638 307448
rect 407942 307436 407948 307448
rect 408000 307436 408006 307488
rect 552014 307436 552020 307488
rect 552072 307476 552078 307488
rect 553946 307476 553952 307488
rect 552072 307448 553952 307476
rect 552072 307436 552078 307448
rect 553946 307436 553952 307448
rect 554004 307436 554010 307488
rect 396534 307028 396540 307080
rect 396592 307068 396598 307080
rect 409230 307068 409236 307080
rect 396592 307040 409236 307068
rect 396592 307028 396598 307040
rect 409230 307028 409236 307040
rect 409288 307028 409294 307080
rect 552198 305464 552204 305516
rect 552256 305504 552262 305516
rect 555510 305504 555516 305516
rect 552256 305476 555516 305504
rect 552256 305464 552262 305476
rect 555510 305464 555516 305476
rect 555568 305464 555574 305516
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 26694 305028 26700 305040
rect 3568 305000 26700 305028
rect 3568 304988 3574 305000
rect 26694 304988 26700 305000
rect 26752 304988 26758 305040
rect 396810 304988 396816 305040
rect 396868 305028 396874 305040
rect 407114 305028 407120 305040
rect 396868 305000 407120 305028
rect 396868 304988 396874 305000
rect 407114 304988 407120 305000
rect 407172 304988 407178 305040
rect 553118 304988 553124 305040
rect 553176 305028 553182 305040
rect 583202 305028 583208 305040
rect 553176 305000 583208 305028
rect 553176 304988 553182 305000
rect 583202 304988 583208 305000
rect 583260 304988 583266 305040
rect 391566 304240 391572 304292
rect 391624 304280 391630 304292
rect 407574 304280 407580 304292
rect 391624 304252 407580 304280
rect 391624 304240 391630 304252
rect 407574 304240 407580 304252
rect 407632 304240 407638 304292
rect 350442 303696 350448 303748
rect 350500 303736 350506 303748
rect 369762 303736 369768 303748
rect 350500 303708 369768 303736
rect 350500 303696 350506 303708
rect 369762 303696 369768 303708
rect 369820 303696 369826 303748
rect 365346 303628 365352 303680
rect 365404 303668 365410 303680
rect 407114 303668 407120 303680
rect 365404 303640 407120 303668
rect 365404 303628 365410 303640
rect 407114 303628 407120 303640
rect 407172 303628 407178 303680
rect 350166 302268 350172 302320
rect 350224 302308 350230 302320
rect 350902 302308 350908 302320
rect 350224 302280 350908 302308
rect 350224 302268 350230 302280
rect 350902 302268 350908 302280
rect 350960 302268 350966 302320
rect 22554 302200 22560 302252
rect 22612 302240 22618 302252
rect 46382 302240 46388 302252
rect 22612 302212 46388 302240
rect 22612 302200 22618 302212
rect 46382 302200 46388 302212
rect 46440 302200 46446 302252
rect 350442 302200 350448 302252
rect 350500 302240 350506 302252
rect 382090 302240 382096 302252
rect 350500 302212 382096 302240
rect 350500 302200 350506 302212
rect 382090 302200 382096 302212
rect 382148 302200 382154 302252
rect 43714 302132 43720 302184
rect 43772 302172 43778 302184
rect 46290 302172 46296 302184
rect 43772 302144 46296 302172
rect 43772 302132 43778 302144
rect 46290 302132 46296 302144
rect 46348 302132 46354 302184
rect 350442 300908 350448 300960
rect 350500 300948 350506 300960
rect 372246 300948 372252 300960
rect 350500 300920 372252 300948
rect 350500 300908 350506 300920
rect 372246 300908 372252 300920
rect 372304 300908 372310 300960
rect 388346 300908 388352 300960
rect 388404 300948 388410 300960
rect 407114 300948 407120 300960
rect 388404 300920 407120 300948
rect 388404 300908 388410 300920
rect 407114 300908 407120 300920
rect 407172 300908 407178 300960
rect 553026 300908 553032 300960
rect 553084 300948 553090 300960
rect 566550 300948 566556 300960
rect 553084 300920 566556 300948
rect 553084 300908 553090 300920
rect 566550 300908 566556 300920
rect 566608 300908 566614 300960
rect 21266 300840 21272 300892
rect 21324 300880 21330 300892
rect 46382 300880 46388 300892
rect 21324 300852 46388 300880
rect 21324 300840 21330 300852
rect 46382 300840 46388 300852
rect 46440 300840 46446 300892
rect 366726 300840 366732 300892
rect 366784 300880 366790 300892
rect 407206 300880 407212 300892
rect 366784 300852 407212 300880
rect 366784 300840 366790 300852
rect 407206 300840 407212 300852
rect 407264 300840 407270 300892
rect 553118 300840 553124 300892
rect 553176 300880 553182 300892
rect 574462 300880 574468 300892
rect 553176 300852 574468 300880
rect 553176 300840 553182 300852
rect 574462 300840 574468 300852
rect 574520 300840 574526 300892
rect 350442 299548 350448 299600
rect 350500 299588 350506 299600
rect 379422 299588 379428 299600
rect 350500 299560 379428 299588
rect 350500 299548 350506 299560
rect 379422 299548 379428 299560
rect 379480 299548 379486 299600
rect 361206 299480 361212 299532
rect 361264 299520 361270 299532
rect 407114 299520 407120 299532
rect 361264 299492 407120 299520
rect 361264 299480 361270 299492
rect 407114 299480 407120 299492
rect 407172 299480 407178 299532
rect 553118 299480 553124 299532
rect 553176 299520 553182 299532
rect 574922 299520 574928 299532
rect 553176 299492 574928 299520
rect 553176 299480 553182 299492
rect 574922 299480 574928 299492
rect 574980 299480 574986 299532
rect 36630 298528 36636 298580
rect 36688 298568 36694 298580
rect 39390 298568 39396 298580
rect 36688 298540 39396 298568
rect 36688 298528 36694 298540
rect 39390 298528 39396 298540
rect 39448 298528 39454 298580
rect 20254 298120 20260 298172
rect 20312 298160 20318 298172
rect 46382 298160 46388 298172
rect 20312 298132 46388 298160
rect 20312 298120 20318 298132
rect 46382 298120 46388 298132
rect 46440 298120 46446 298172
rect 350442 298120 350448 298172
rect 350500 298160 350506 298172
rect 384114 298160 384120 298172
rect 350500 298132 384120 298160
rect 350500 298120 350506 298132
rect 384114 298120 384120 298132
rect 384172 298120 384178 298172
rect 365254 297372 365260 297424
rect 365312 297412 365318 297424
rect 375282 297412 375288 297424
rect 365312 297384 375288 297412
rect 365312 297372 365318 297384
rect 375282 297372 375288 297384
rect 375340 297372 375346 297424
rect 39390 296692 39396 296744
rect 39448 296732 39454 296744
rect 46382 296732 46388 296744
rect 39448 296704 46388 296732
rect 39448 296692 39454 296704
rect 46382 296692 46388 296704
rect 46440 296692 46446 296744
rect 553118 296692 553124 296744
rect 553176 296732 553182 296744
rect 573358 296732 573364 296744
rect 553176 296704 573364 296732
rect 553176 296692 553182 296704
rect 573358 296692 573364 296704
rect 573416 296692 573422 296744
rect 350442 296624 350448 296676
rect 350500 296664 350506 296676
rect 363046 296664 363052 296676
rect 350500 296636 363052 296664
rect 350500 296624 350506 296636
rect 363046 296624 363052 296636
rect 363104 296624 363110 296676
rect 349246 295740 349252 295792
rect 349304 295780 349310 295792
rect 350810 295780 350816 295792
rect 349304 295752 350816 295780
rect 349304 295740 349310 295752
rect 350810 295740 350816 295752
rect 350868 295740 350874 295792
rect 406102 295400 406108 295452
rect 406160 295440 406166 295452
rect 407850 295440 407856 295452
rect 406160 295412 407856 295440
rect 406160 295400 406166 295412
rect 407850 295400 407856 295412
rect 407908 295400 407914 295452
rect 350442 295332 350448 295384
rect 350500 295372 350506 295384
rect 365254 295372 365260 295384
rect 350500 295344 365260 295372
rect 350500 295332 350506 295344
rect 365254 295332 365260 295344
rect 365312 295332 365318 295384
rect 399754 295332 399760 295384
rect 399812 295372 399818 295384
rect 407114 295372 407120 295384
rect 399812 295344 407120 295372
rect 399812 295332 399818 295344
rect 407114 295332 407120 295344
rect 407172 295332 407178 295384
rect 350350 294040 350356 294092
rect 350408 294080 350414 294092
rect 350810 294080 350816 294092
rect 350408 294052 350816 294080
rect 350408 294040 350414 294052
rect 350810 294040 350816 294052
rect 350868 294040 350874 294092
rect 43254 293972 43260 294024
rect 43312 294012 43318 294024
rect 44174 294012 44180 294024
rect 43312 293984 44180 294012
rect 43312 293972 43318 293984
rect 44174 293972 44180 293984
rect 44232 293972 44238 294024
rect 350442 293972 350448 294024
rect 350500 294012 350506 294024
rect 363046 294012 363052 294024
rect 350500 293984 363052 294012
rect 350500 293972 350506 293984
rect 363046 293972 363052 293984
rect 363104 293972 363110 294024
rect 35250 293904 35256 293956
rect 35308 293944 35314 293956
rect 46106 293944 46112 293956
rect 35308 293916 46112 293944
rect 35308 293904 35314 293916
rect 46106 293904 46112 293916
rect 46164 293904 46170 293956
rect 552014 293088 552020 293140
rect 552072 293128 552078 293140
rect 553762 293128 553768 293140
rect 552072 293100 553768 293128
rect 552072 293088 552078 293100
rect 553762 293088 553768 293100
rect 553820 293088 553826 293140
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 17494 292584 17500 292596
rect 3568 292556 17500 292584
rect 3568 292544 3574 292556
rect 17494 292544 17500 292556
rect 17552 292544 17558 292596
rect 32490 292544 32496 292596
rect 32548 292584 32554 292596
rect 46382 292584 46388 292596
rect 32548 292556 46388 292584
rect 32548 292544 32554 292556
rect 46382 292544 46388 292556
rect 46440 292544 46446 292596
rect 364058 292544 364064 292596
rect 364116 292584 364122 292596
rect 407206 292584 407212 292596
rect 364116 292556 407212 292584
rect 364116 292544 364122 292556
rect 407206 292544 407212 292556
rect 407264 292544 407270 292596
rect 371970 292476 371976 292528
rect 372028 292516 372034 292528
rect 407114 292516 407120 292528
rect 372028 292488 407120 292516
rect 372028 292476 372034 292488
rect 407114 292476 407120 292488
rect 407172 292476 407178 292528
rect 402698 292408 402704 292460
rect 402756 292448 402762 292460
rect 407206 292448 407212 292460
rect 402756 292420 407212 292448
rect 402756 292408 402762 292420
rect 407206 292408 407212 292420
rect 407264 292408 407270 292460
rect 552014 291728 552020 291780
rect 552072 291768 552078 291780
rect 554038 291768 554044 291780
rect 552072 291740 554044 291768
rect 552072 291728 552078 291740
rect 554038 291728 554044 291740
rect 554096 291728 554102 291780
rect 43714 291184 43720 291236
rect 43772 291224 43778 291236
rect 46382 291224 46388 291236
rect 43772 291196 46388 291224
rect 43772 291184 43778 291196
rect 46382 291184 46388 291196
rect 46440 291184 46446 291236
rect 553118 291184 553124 291236
rect 553176 291224 553182 291236
rect 583294 291224 583300 291236
rect 553176 291196 583300 291224
rect 553176 291184 553182 291196
rect 583294 291184 583300 291196
rect 583352 291184 583358 291236
rect 373626 290436 373632 290488
rect 373684 290476 373690 290488
rect 403526 290476 403532 290488
rect 373684 290448 403532 290476
rect 373684 290436 373690 290448
rect 403526 290436 403532 290448
rect 403584 290436 403590 290488
rect 553118 289824 553124 289876
rect 553176 289864 553182 289876
rect 566090 289864 566096 289876
rect 553176 289836 566096 289864
rect 553176 289824 553182 289836
rect 566090 289824 566096 289836
rect 566148 289824 566154 289876
rect 402146 288464 402152 288516
rect 402204 288504 402210 288516
rect 407114 288504 407120 288516
rect 402204 288476 407120 288504
rect 402204 288464 402210 288476
rect 407114 288464 407120 288476
rect 407172 288464 407178 288516
rect 553026 288464 553032 288516
rect 553084 288504 553090 288516
rect 564986 288504 564992 288516
rect 553084 288476 564992 288504
rect 553084 288464 553090 288476
rect 564986 288464 564992 288476
rect 565044 288464 565050 288516
rect 350442 288396 350448 288448
rect 350500 288436 350506 288448
rect 403526 288436 403532 288448
rect 350500 288408 403532 288436
rect 350500 288396 350506 288408
rect 403526 288396 403532 288408
rect 403584 288396 403590 288448
rect 404906 288396 404912 288448
rect 404964 288436 404970 288448
rect 407298 288436 407304 288448
rect 404964 288408 407304 288436
rect 404964 288396 404970 288408
rect 407298 288396 407304 288408
rect 407356 288396 407362 288448
rect 553118 288396 553124 288448
rect 553176 288436 553182 288448
rect 578510 288436 578516 288448
rect 553176 288408 578516 288436
rect 553176 288396 553182 288408
rect 578510 288396 578516 288408
rect 578568 288396 578574 288448
rect 401134 288328 401140 288380
rect 401192 288368 401198 288380
rect 402698 288368 402704 288380
rect 401192 288340 402704 288368
rect 401192 288328 401198 288340
rect 402698 288328 402704 288340
rect 402756 288328 402762 288380
rect 350442 287104 350448 287156
rect 350500 287144 350506 287156
rect 357158 287144 357164 287156
rect 350500 287116 357164 287144
rect 350500 287104 350506 287116
rect 357158 287104 357164 287116
rect 357216 287104 357222 287156
rect 401134 287104 401140 287156
rect 401192 287144 401198 287156
rect 407114 287144 407120 287156
rect 401192 287116 407120 287144
rect 401192 287104 401198 287116
rect 407114 287104 407120 287116
rect 407172 287104 407178 287156
rect 380802 287036 380808 287088
rect 380860 287076 380866 287088
rect 407206 287076 407212 287088
rect 380860 287048 407212 287076
rect 380860 287036 380866 287048
rect 407206 287036 407212 287048
rect 407264 287036 407270 287088
rect 553118 287036 553124 287088
rect 553176 287076 553182 287088
rect 570322 287076 570328 287088
rect 553176 287048 570328 287076
rect 553176 287036 553182 287048
rect 570322 287036 570328 287048
rect 570380 287036 570386 287088
rect 390186 285744 390192 285796
rect 390244 285784 390250 285796
rect 407114 285784 407120 285796
rect 390244 285756 407120 285784
rect 390244 285744 390250 285756
rect 407114 285744 407120 285756
rect 407172 285744 407178 285796
rect 28166 285676 28172 285728
rect 28224 285716 28230 285728
rect 46382 285716 46388 285728
rect 28224 285688 46388 285716
rect 28224 285676 28230 285688
rect 46382 285676 46388 285688
rect 46440 285676 46446 285728
rect 350442 285676 350448 285728
rect 350500 285716 350506 285728
rect 401042 285716 401048 285728
rect 350500 285688 401048 285716
rect 350500 285676 350506 285688
rect 401042 285676 401048 285688
rect 401100 285676 401106 285728
rect 350350 285608 350356 285660
rect 350408 285648 350414 285660
rect 400766 285648 400772 285660
rect 350408 285620 400772 285648
rect 350408 285608 350414 285620
rect 400766 285608 400772 285620
rect 400824 285608 400830 285660
rect 393038 284928 393044 284980
rect 393096 284968 393102 284980
rect 394142 284968 394148 284980
rect 393096 284940 394148 284968
rect 393096 284928 393102 284940
rect 394142 284928 394148 284940
rect 394200 284928 394206 284980
rect 43622 284656 43628 284708
rect 43680 284696 43686 284708
rect 45646 284696 45652 284708
rect 43680 284668 45652 284696
rect 43680 284656 43686 284668
rect 45646 284656 45652 284668
rect 45704 284656 45710 284708
rect 384206 284316 384212 284368
rect 384264 284356 384270 284368
rect 407114 284356 407120 284368
rect 384264 284328 407120 284356
rect 384264 284316 384270 284328
rect 407114 284316 407120 284328
rect 407172 284316 407178 284368
rect 365438 284248 365444 284300
rect 365496 284288 365502 284300
rect 407206 284288 407212 284300
rect 365496 284260 407212 284288
rect 365496 284248 365502 284260
rect 407206 284248 407212 284260
rect 407264 284248 407270 284300
rect 553118 283568 553124 283620
rect 553176 283608 553182 283620
rect 566182 283608 566188 283620
rect 553176 283580 566188 283608
rect 553176 283568 553182 283580
rect 566182 283568 566188 283580
rect 566240 283568 566246 283620
rect 393038 282888 393044 282940
rect 393096 282928 393102 282940
rect 407114 282928 407120 282940
rect 393096 282900 407120 282928
rect 393096 282888 393102 282900
rect 407114 282888 407120 282900
rect 407172 282888 407178 282940
rect 566182 282888 566188 282940
rect 566240 282928 566246 282940
rect 566642 282928 566648 282940
rect 566240 282900 566648 282928
rect 566240 282888 566246 282900
rect 566642 282888 566648 282900
rect 566700 282888 566706 282940
rect 553118 282820 553124 282872
rect 553176 282860 553182 282872
rect 565998 282860 566004 282872
rect 553176 282832 566004 282860
rect 553176 282820 553182 282832
rect 565998 282820 566004 282832
rect 566056 282820 566062 282872
rect 348510 281936 348516 281988
rect 348568 281976 348574 281988
rect 350166 281976 350172 281988
rect 348568 281948 350172 281976
rect 348568 281936 348574 281948
rect 350166 281936 350172 281948
rect 350224 281936 350230 281988
rect 39206 281664 39212 281716
rect 39264 281704 39270 281716
rect 44818 281704 44824 281716
rect 39264 281676 44824 281704
rect 39264 281664 39270 281676
rect 44818 281664 44824 281676
rect 44876 281664 44882 281716
rect 32582 281596 32588 281648
rect 32640 281636 32646 281648
rect 46842 281636 46848 281648
rect 32640 281608 46848 281636
rect 32640 281596 32646 281608
rect 46842 281596 46848 281608
rect 46900 281596 46906 281648
rect 24026 281528 24032 281580
rect 24084 281568 24090 281580
rect 45646 281568 45652 281580
rect 24084 281540 45652 281568
rect 24084 281528 24090 281540
rect 45646 281528 45652 281540
rect 45704 281528 45710 281580
rect 387518 281460 387524 281512
rect 387576 281500 387582 281512
rect 387794 281500 387800 281512
rect 387576 281472 387800 281500
rect 387576 281460 387582 281472
rect 387794 281460 387800 281472
rect 387852 281460 387858 281512
rect 553118 280236 553124 280288
rect 553176 280276 553182 280288
rect 566826 280276 566832 280288
rect 553176 280248 566832 280276
rect 553176 280236 553182 280248
rect 566826 280236 566832 280248
rect 566884 280236 566890 280288
rect 553026 280168 553032 280220
rect 553084 280208 553090 280220
rect 571886 280208 571892 280220
rect 553084 280180 571892 280208
rect 553084 280168 553090 280180
rect 571886 280168 571892 280180
rect 571944 280168 571950 280220
rect 553118 280100 553124 280152
rect 553176 280140 553182 280152
rect 566274 280140 566280 280152
rect 553176 280112 566280 280140
rect 553176 280100 553182 280112
rect 566274 280100 566280 280112
rect 566332 280100 566338 280152
rect 349062 279012 349068 279064
rect 349120 279052 349126 279064
rect 350810 279052 350816 279064
rect 349120 279024 350816 279052
rect 349120 279012 349126 279024
rect 350810 279012 350816 279024
rect 350868 279012 350874 279064
rect 400766 278808 400772 278860
rect 400824 278848 400830 278860
rect 407114 278848 407120 278860
rect 400824 278820 407120 278848
rect 400824 278808 400830 278820
rect 407114 278808 407120 278820
rect 407172 278808 407178 278860
rect 553118 278808 553124 278860
rect 553176 278848 553182 278860
rect 557074 278848 557080 278860
rect 553176 278820 557080 278848
rect 553176 278808 553182 278820
rect 557074 278808 557080 278820
rect 557132 278808 557138 278860
rect 388162 278740 388168 278792
rect 388220 278780 388226 278792
rect 407206 278780 407212 278792
rect 388220 278752 407212 278780
rect 388220 278740 388226 278752
rect 407206 278740 407212 278752
rect 407264 278740 407270 278792
rect 25314 277380 25320 277432
rect 25372 277420 25378 277432
rect 46842 277420 46848 277432
rect 25372 277392 46848 277420
rect 25372 277380 25378 277392
rect 46842 277380 46848 277392
rect 46900 277380 46906 277432
rect 350442 277380 350448 277432
rect 350500 277420 350506 277432
rect 381446 277420 381452 277432
rect 350500 277392 381452 277420
rect 350500 277380 350506 277392
rect 381446 277380 381452 277392
rect 381504 277380 381510 277432
rect 553118 277380 553124 277432
rect 553176 277420 553182 277432
rect 567378 277420 567384 277432
rect 553176 277392 567384 277420
rect 553176 277380 553182 277392
rect 567378 277380 567384 277392
rect 567436 277380 567442 277432
rect 380526 277312 380532 277364
rect 380584 277352 380590 277364
rect 407114 277352 407120 277364
rect 380584 277324 407120 277352
rect 380584 277312 380590 277324
rect 407114 277312 407120 277324
rect 407172 277312 407178 277364
rect 408402 276768 408408 276820
rect 408460 276808 408466 276820
rect 409138 276808 409144 276820
rect 408460 276780 409144 276808
rect 408460 276768 408466 276780
rect 409138 276768 409144 276780
rect 409196 276768 409202 276820
rect 553026 276088 553032 276140
rect 553084 276128 553090 276140
rect 556798 276128 556804 276140
rect 553084 276100 556804 276128
rect 553084 276088 553090 276100
rect 556798 276088 556804 276100
rect 556856 276088 556862 276140
rect 46474 276020 46480 276072
rect 46532 276060 46538 276072
rect 47578 276060 47584 276072
rect 46532 276032 47584 276060
rect 46532 276020 46538 276032
rect 47578 276020 47584 276032
rect 47636 276020 47642 276072
rect 350442 275952 350448 276004
rect 350500 275992 350506 276004
rect 388530 275992 388536 276004
rect 350500 275964 388536 275992
rect 350500 275952 350506 275964
rect 388530 275952 388536 275964
rect 388588 275952 388594 276004
rect 384666 275884 384672 275936
rect 384724 275924 384730 275936
rect 407114 275924 407120 275936
rect 384724 275896 407120 275924
rect 384724 275884 384730 275896
rect 407114 275884 407120 275896
rect 407172 275884 407178 275936
rect 46474 274660 46480 274712
rect 46532 274700 46538 274712
rect 47302 274700 47308 274712
rect 46532 274672 47308 274700
rect 46532 274660 46538 274672
rect 47302 274660 47308 274672
rect 47360 274660 47366 274712
rect 351362 274660 351368 274712
rect 351420 274700 351426 274712
rect 354122 274700 354128 274712
rect 351420 274672 354128 274700
rect 351420 274660 351426 274672
rect 354122 274660 354128 274672
rect 354180 274660 354186 274712
rect 376662 274660 376668 274712
rect 376720 274700 376726 274712
rect 379514 274700 379520 274712
rect 376720 274672 379520 274700
rect 376720 274660 376726 274672
rect 379514 274660 379520 274672
rect 379572 274660 379578 274712
rect 553118 274660 553124 274712
rect 553176 274700 553182 274712
rect 565078 274700 565084 274712
rect 553176 274672 565084 274700
rect 553176 274660 553182 274672
rect 565078 274660 565084 274672
rect 565136 274660 565142 274712
rect 350442 273300 350448 273352
rect 350500 273340 350506 273352
rect 364702 273340 364708 273352
rect 350500 273312 364708 273340
rect 350500 273300 350506 273312
rect 364702 273300 364708 273312
rect 364760 273300 364766 273352
rect 32674 273232 32680 273284
rect 32732 273272 32738 273284
rect 46842 273272 46848 273284
rect 32732 273244 46848 273272
rect 32732 273232 32738 273244
rect 46842 273232 46848 273244
rect 46900 273232 46906 273284
rect 350350 273232 350356 273284
rect 350408 273272 350414 273284
rect 393774 273272 393780 273284
rect 350408 273244 393780 273272
rect 350408 273232 350414 273244
rect 393774 273232 393780 273244
rect 393832 273232 393838 273284
rect 553118 273232 553124 273284
rect 553176 273272 553182 273284
rect 576026 273272 576032 273284
rect 553176 273244 576032 273272
rect 553176 273232 553182 273244
rect 576026 273232 576032 273244
rect 576084 273232 576090 273284
rect 575014 273164 575020 273216
rect 575072 273204 575078 273216
rect 580166 273204 580172 273216
rect 575072 273176 580172 273204
rect 575072 273164 575078 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 46474 272552 46480 272604
rect 46532 272592 46538 272604
rect 46842 272592 46848 272604
rect 46532 272564 46848 272592
rect 46532 272552 46538 272564
rect 46842 272552 46848 272564
rect 46900 272552 46906 272604
rect 407482 272552 407488 272604
rect 407540 272592 407546 272604
rect 407758 272592 407764 272604
rect 407540 272564 407764 272592
rect 407540 272552 407546 272564
rect 407758 272552 407764 272564
rect 407816 272552 407822 272604
rect 405366 271804 405372 271856
rect 405424 271844 405430 271856
rect 407114 271844 407120 271856
rect 405424 271816 407120 271844
rect 405424 271804 405430 271816
rect 407114 271804 407120 271816
rect 407172 271804 407178 271856
rect 553118 270512 553124 270564
rect 553176 270552 553182 270564
rect 578602 270552 578608 270564
rect 553176 270524 578608 270552
rect 553176 270512 553182 270524
rect 578602 270512 578608 270524
rect 578660 270512 578666 270564
rect 350442 270444 350448 270496
rect 350500 270484 350506 270496
rect 378962 270484 378968 270496
rect 350500 270456 378968 270484
rect 350500 270444 350506 270456
rect 378962 270444 378968 270456
rect 379020 270444 379026 270496
rect 36814 269764 36820 269816
rect 36872 269804 36878 269816
rect 45554 269804 45560 269816
rect 36872 269776 45560 269804
rect 36872 269764 36878 269776
rect 45554 269764 45560 269776
rect 45612 269764 45618 269816
rect 358630 269084 358636 269136
rect 358688 269124 358694 269136
rect 407114 269124 407120 269136
rect 358688 269096 407120 269124
rect 358688 269084 358694 269096
rect 407114 269084 407120 269096
rect 407172 269084 407178 269136
rect 350442 269016 350448 269068
rect 350500 269056 350506 269068
rect 378134 269056 378140 269068
rect 350500 269028 378140 269056
rect 350500 269016 350506 269028
rect 378134 269016 378140 269028
rect 378192 269016 378198 269068
rect 33962 268336 33968 268388
rect 34020 268376 34026 268388
rect 47118 268376 47124 268388
rect 34020 268348 47124 268376
rect 34020 268336 34026 268348
rect 47118 268336 47124 268348
rect 47176 268336 47182 268388
rect 36814 267792 36820 267844
rect 36872 267832 36878 267844
rect 46382 267832 46388 267844
rect 36872 267804 46388 267832
rect 36872 267792 36878 267804
rect 46382 267792 46388 267804
rect 46440 267792 46446 267844
rect 30926 267724 30932 267776
rect 30984 267764 30990 267776
rect 46474 267764 46480 267776
rect 30984 267736 46480 267764
rect 30984 267724 30990 267736
rect 46474 267724 46480 267736
rect 46532 267724 46538 267776
rect 401962 267724 401968 267776
rect 402020 267764 402026 267776
rect 407114 267764 407120 267776
rect 402020 267736 407120 267764
rect 402020 267724 402026 267736
rect 407114 267724 407120 267736
rect 407172 267724 407178 267776
rect 45462 266364 45468 266416
rect 45520 266404 45526 266416
rect 46934 266404 46940 266416
rect 45520 266376 46940 266404
rect 45520 266364 45526 266376
rect 46934 266364 46940 266376
rect 46992 266364 46998 266416
rect 350442 266364 350448 266416
rect 350500 266404 350506 266416
rect 378962 266404 378968 266416
rect 350500 266376 378968 266404
rect 350500 266364 350506 266376
rect 378962 266364 378968 266376
rect 379020 266364 379026 266416
rect 405366 266364 405372 266416
rect 405424 266404 405430 266416
rect 407758 266404 407764 266416
rect 405424 266376 407764 266404
rect 405424 266364 405430 266376
rect 407758 266364 407764 266376
rect 407816 266364 407822 266416
rect 553118 266364 553124 266416
rect 553176 266404 553182 266416
rect 574646 266404 574652 266416
rect 553176 266376 574652 266404
rect 553176 266364 553182 266376
rect 574646 266364 574652 266376
rect 574704 266364 574710 266416
rect 552014 265208 552020 265260
rect 552072 265248 552078 265260
rect 554222 265248 554228 265260
rect 552072 265220 554228 265248
rect 552072 265208 552078 265220
rect 554222 265208 554228 265220
rect 554280 265208 554286 265260
rect 350442 263644 350448 263696
rect 350500 263684 350506 263696
rect 371418 263684 371424 263696
rect 350500 263656 371424 263684
rect 350500 263644 350506 263656
rect 371418 263644 371424 263656
rect 371476 263644 371482 263696
rect 360378 263576 360384 263628
rect 360436 263616 360442 263628
rect 407114 263616 407120 263628
rect 360436 263588 407120 263616
rect 360436 263576 360442 263588
rect 407114 263576 407120 263588
rect 407172 263576 407178 263628
rect 553118 263576 553124 263628
rect 553176 263616 553182 263628
rect 564434 263616 564440 263628
rect 553176 263588 564440 263616
rect 553176 263576 553182 263588
rect 564434 263576 564440 263588
rect 564492 263576 564498 263628
rect 552014 263168 552020 263220
rect 552072 263208 552078 263220
rect 554774 263208 554780 263220
rect 552072 263180 554780 263208
rect 552072 263168 552078 263180
rect 554774 263168 554780 263180
rect 554832 263168 554838 263220
rect 394142 262896 394148 262948
rect 394200 262936 394206 262948
rect 395154 262936 395160 262948
rect 394200 262908 395160 262936
rect 394200 262896 394206 262908
rect 395154 262896 395160 262908
rect 395212 262896 395218 262948
rect 389082 262624 389088 262676
rect 389140 262664 389146 262676
rect 392394 262664 392400 262676
rect 389140 262636 392400 262664
rect 389140 262624 389146 262636
rect 392394 262624 392400 262636
rect 392452 262624 392458 262676
rect 364150 262216 364156 262268
rect 364208 262256 364214 262268
rect 407114 262256 407120 262268
rect 364208 262228 407120 262256
rect 364208 262216 364214 262228
rect 407114 262216 407120 262228
rect 407172 262216 407178 262268
rect 349062 262148 349068 262200
rect 349120 262188 349126 262200
rect 349982 262188 349988 262200
rect 349120 262160 349988 262188
rect 349120 262148 349126 262160
rect 349982 262148 349988 262160
rect 350040 262148 350046 262200
rect 350442 262148 350448 262200
rect 350500 262188 350506 262200
rect 360378 262188 360384 262200
rect 350500 262160 360384 262188
rect 350500 262148 350506 262160
rect 360378 262148 360384 262160
rect 360436 262148 360442 262200
rect 394142 261536 394148 261588
rect 394200 261576 394206 261588
rect 395706 261576 395712 261588
rect 394200 261548 395712 261576
rect 394200 261536 394206 261548
rect 395706 261536 395712 261548
rect 395764 261536 395770 261588
rect 351822 261400 351828 261452
rect 351880 261440 351886 261452
rect 355134 261440 355140 261452
rect 351880 261412 355140 261440
rect 351880 261400 351886 261412
rect 355134 261400 355140 261412
rect 355192 261400 355198 261452
rect 404814 261128 404820 261180
rect 404872 261168 404878 261180
rect 407482 261168 407488 261180
rect 404872 261140 407488 261168
rect 404872 261128 404878 261140
rect 407482 261128 407488 261140
rect 407540 261128 407546 261180
rect 407574 261128 407580 261180
rect 407632 261128 407638 261180
rect 407592 260976 407620 261128
rect 407574 260924 407580 260976
rect 407632 260924 407638 260976
rect 380526 260856 380532 260908
rect 380584 260896 380590 260908
rect 407114 260896 407120 260908
rect 380584 260868 407120 260896
rect 380584 260856 380590 260868
rect 407114 260856 407120 260868
rect 407172 260856 407178 260908
rect 552014 260856 552020 260908
rect 552072 260896 552078 260908
rect 568574 260896 568580 260908
rect 552072 260868 568580 260896
rect 552072 260856 552078 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 552842 260380 552848 260432
rect 552900 260420 552906 260432
rect 553026 260420 553032 260432
rect 552900 260392 553032 260420
rect 552900 260380 552906 260392
rect 553026 260380 553032 260392
rect 553084 260380 553090 260432
rect 552106 259496 552112 259548
rect 552164 259536 552170 259548
rect 569034 259536 569040 259548
rect 552164 259508 569040 259536
rect 552164 259496 552170 259508
rect 569034 259496 569040 259508
rect 569092 259496 569098 259548
rect 395706 259428 395712 259480
rect 395764 259468 395770 259480
rect 407114 259468 407120 259480
rect 395764 259440 407120 259468
rect 395764 259428 395770 259440
rect 407114 259428 407120 259440
rect 407172 259428 407178 259480
rect 552014 259428 552020 259480
rect 552072 259468 552078 259480
rect 583386 259468 583392 259480
rect 552072 259440 583392 259468
rect 552072 259428 552078 259440
rect 583386 259428 583392 259440
rect 583444 259428 583450 259480
rect 552106 258136 552112 258188
rect 552164 258176 552170 258188
rect 560294 258176 560300 258188
rect 552164 258148 560300 258176
rect 552164 258136 552170 258148
rect 560294 258136 560300 258148
rect 560352 258136 560358 258188
rect 44450 258068 44456 258120
rect 44508 258108 44514 258120
rect 46014 258108 46020 258120
rect 44508 258080 46020 258108
rect 44508 258068 44514 258080
rect 46014 258068 46020 258080
rect 46072 258068 46078 258120
rect 350442 258068 350448 258120
rect 350500 258108 350506 258120
rect 386966 258108 386972 258120
rect 350500 258080 386972 258108
rect 350500 258068 350506 258080
rect 386966 258068 386972 258080
rect 387024 258068 387030 258120
rect 552014 258068 552020 258120
rect 552072 258108 552078 258120
rect 568942 258108 568948 258120
rect 552072 258080 568948 258108
rect 552072 258068 552078 258080
rect 568942 258068 568948 258080
rect 569000 258068 569006 258120
rect 37182 257320 37188 257372
rect 37240 257360 37246 257372
rect 45646 257360 45652 257372
rect 37240 257332 45652 257360
rect 37240 257320 37246 257332
rect 45646 257320 45652 257332
rect 45704 257320 45710 257372
rect 402514 257320 402520 257372
rect 402572 257360 402578 257372
rect 406562 257360 406568 257372
rect 402572 257332 406568 257360
rect 402572 257320 402578 257332
rect 406562 257320 406568 257332
rect 406620 257320 406626 257372
rect 46842 257184 46848 257236
rect 46900 257224 46906 257236
rect 47394 257224 47400 257236
rect 46900 257196 47400 257224
rect 46900 257184 46906 257196
rect 47394 257184 47400 257196
rect 47452 257184 47458 257236
rect 399386 256776 399392 256828
rect 399444 256816 399450 256828
rect 407114 256816 407120 256828
rect 399444 256788 407120 256816
rect 399444 256776 399450 256788
rect 407114 256776 407120 256788
rect 407172 256776 407178 256828
rect 45462 256708 45468 256760
rect 45520 256748 45526 256760
rect 46014 256748 46020 256760
rect 45520 256720 46020 256748
rect 45520 256708 45526 256720
rect 46014 256708 46020 256720
rect 46072 256708 46078 256760
rect 371970 256708 371976 256760
rect 372028 256748 372034 256760
rect 407206 256748 407212 256760
rect 372028 256720 407212 256748
rect 372028 256708 372034 256720
rect 407206 256708 407212 256720
rect 407264 256708 407270 256760
rect 552014 256708 552020 256760
rect 552072 256748 552078 256760
rect 565814 256748 565820 256760
rect 552072 256720 565820 256748
rect 552072 256708 552078 256720
rect 565814 256708 565820 256720
rect 565872 256708 565878 256760
rect 35066 255960 35072 256012
rect 35124 256000 35130 256012
rect 36630 256000 36636 256012
rect 35124 255972 36636 256000
rect 35124 255960 35130 255972
rect 36630 255960 36636 255972
rect 36688 255960 36694 256012
rect 375006 255960 375012 256012
rect 375064 256000 375070 256012
rect 384666 256000 384672 256012
rect 375064 255972 384672 256000
rect 375064 255960 375070 255972
rect 384666 255960 384672 255972
rect 384724 255960 384730 256012
rect 387334 255960 387340 256012
rect 387392 256000 387398 256012
rect 391106 256000 391112 256012
rect 387392 255972 391112 256000
rect 387392 255960 387398 255972
rect 391106 255960 391112 255972
rect 391164 255960 391170 256012
rect 402054 255960 402060 256012
rect 402112 256000 402118 256012
rect 407482 256000 407488 256012
rect 402112 255972 407488 256000
rect 402112 255960 402118 255972
rect 407482 255960 407488 255972
rect 407540 255960 407546 256012
rect 349890 255416 349896 255468
rect 349948 255456 349954 255468
rect 350534 255456 350540 255468
rect 349948 255428 350540 255456
rect 349948 255416 349954 255428
rect 350534 255416 350540 255428
rect 350592 255416 350598 255468
rect 350350 255348 350356 255400
rect 350408 255388 350414 255400
rect 391014 255388 391020 255400
rect 350408 255360 391020 255388
rect 350408 255348 350414 255360
rect 391014 255348 391020 255360
rect 391072 255348 391078 255400
rect 350442 255280 350448 255332
rect 350500 255320 350506 255332
rect 397914 255320 397920 255332
rect 350500 255292 397920 255320
rect 350500 255280 350506 255292
rect 397914 255280 397920 255292
rect 397972 255280 397978 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 26878 255252 26884 255264
rect 3200 255224 26884 255252
rect 3200 255212 3206 255224
rect 26878 255212 26884 255224
rect 26936 255212 26942 255264
rect 405182 255212 405188 255264
rect 405240 255252 405246 255264
rect 407482 255252 407488 255264
rect 405240 255224 407488 255252
rect 405240 255212 405246 255224
rect 407482 255212 407488 255224
rect 407540 255212 407546 255264
rect 406746 253988 406752 254040
rect 406804 254028 406810 254040
rect 407298 254028 407304 254040
rect 406804 254000 407304 254028
rect 406804 253988 406810 254000
rect 407298 253988 407304 254000
rect 407356 253988 407362 254040
rect 552106 253988 552112 254040
rect 552164 254028 552170 254040
rect 566182 254028 566188 254040
rect 552164 254000 566188 254028
rect 552164 253988 552170 254000
rect 566182 253988 566188 254000
rect 566240 253988 566246 254040
rect 36630 253920 36636 253972
rect 36688 253960 36694 253972
rect 46842 253960 46848 253972
rect 36688 253932 46848 253960
rect 36688 253920 36694 253932
rect 46842 253920 46848 253932
rect 46900 253920 46906 253972
rect 350442 253920 350448 253972
rect 350500 253960 350506 253972
rect 355686 253960 355692 253972
rect 350500 253932 355692 253960
rect 350500 253920 350506 253932
rect 355686 253920 355692 253932
rect 355744 253920 355750 253972
rect 387334 253920 387340 253972
rect 387392 253960 387398 253972
rect 407114 253960 407120 253972
rect 387392 253932 407120 253960
rect 387392 253920 387398 253932
rect 407114 253920 407120 253932
rect 407172 253920 407178 253972
rect 552014 253920 552020 253972
rect 552072 253960 552078 253972
rect 573174 253960 573180 253972
rect 552072 253932 573180 253960
rect 552072 253920 552078 253932
rect 573174 253920 573180 253932
rect 573232 253920 573238 253972
rect 36446 253648 36452 253700
rect 36504 253688 36510 253700
rect 43162 253688 43168 253700
rect 36504 253660 43168 253688
rect 36504 253648 36510 253660
rect 43162 253648 43168 253660
rect 43220 253648 43226 253700
rect 43622 253648 43628 253700
rect 43680 253688 43686 253700
rect 44818 253688 44824 253700
rect 43680 253660 44824 253688
rect 43680 253648 43686 253660
rect 44818 253648 44824 253660
rect 44876 253648 44882 253700
rect 354122 253444 354128 253496
rect 354180 253484 354186 253496
rect 355042 253484 355048 253496
rect 354180 253456 355048 253484
rect 354180 253444 354186 253456
rect 355042 253444 355048 253456
rect 355100 253444 355106 253496
rect 402146 253172 402152 253224
rect 402204 253212 402210 253224
rect 409230 253212 409236 253224
rect 402204 253184 409236 253212
rect 402204 253172 402210 253184
rect 409230 253172 409236 253184
rect 409288 253172 409294 253224
rect 553118 252560 553124 252612
rect 553176 252600 553182 252612
rect 570782 252600 570788 252612
rect 553176 252572 570788 252600
rect 553176 252560 553182 252572
rect 570782 252560 570788 252572
rect 570840 252560 570846 252612
rect 552658 252492 552664 252544
rect 552716 252532 552722 252544
rect 553946 252532 553952 252544
rect 552716 252504 553952 252532
rect 552716 252492 552722 252504
rect 553946 252492 553952 252504
rect 554004 252492 554010 252544
rect 361298 251812 361304 251864
rect 361356 251852 361362 251864
rect 378686 251852 378692 251864
rect 361356 251824 378692 251852
rect 361356 251812 361362 251824
rect 378686 251812 378692 251824
rect 378744 251812 378750 251864
rect 402514 251200 402520 251252
rect 402572 251240 402578 251252
rect 407114 251240 407120 251252
rect 402572 251212 407120 251240
rect 402572 251200 402578 251212
rect 407114 251200 407120 251212
rect 407172 251200 407178 251252
rect 553118 251200 553124 251252
rect 553176 251240 553182 251252
rect 561674 251240 561680 251252
rect 553176 251212 561680 251240
rect 553176 251200 553182 251212
rect 561674 251200 561680 251212
rect 561732 251200 561738 251252
rect 402882 251132 402888 251184
rect 402940 251172 402946 251184
rect 407206 251172 407212 251184
rect 402940 251144 407212 251172
rect 402940 251132 402946 251144
rect 407206 251132 407212 251144
rect 407264 251132 407270 251184
rect 361298 249840 361304 249892
rect 361356 249880 361362 249892
rect 407114 249880 407120 249892
rect 361356 249852 407120 249880
rect 361356 249840 361362 249852
rect 407114 249840 407120 249852
rect 407172 249840 407178 249892
rect 552658 249840 552664 249892
rect 552716 249880 552722 249892
rect 553394 249880 553400 249892
rect 552716 249852 553400 249880
rect 552716 249840 552722 249852
rect 553394 249840 553400 249852
rect 553452 249840 553458 249892
rect 350442 249772 350448 249824
rect 350500 249812 350506 249824
rect 400674 249812 400680 249824
rect 350500 249784 400680 249812
rect 350500 249772 350506 249784
rect 400674 249772 400680 249784
rect 400732 249772 400738 249824
rect 552014 249772 552020 249824
rect 552072 249812 552078 249824
rect 552072 249784 553440 249812
rect 552072 249772 552078 249784
rect 553412 249756 553440 249784
rect 553394 249704 553400 249756
rect 553452 249704 553458 249756
rect 405550 248752 405556 248804
rect 405608 248792 405614 248804
rect 407758 248792 407764 248804
rect 405608 248764 407764 248792
rect 405608 248752 405614 248764
rect 407758 248752 407764 248764
rect 407816 248752 407822 248804
rect 350442 248412 350448 248464
rect 350500 248452 350506 248464
rect 402146 248452 402152 248464
rect 350500 248424 402152 248452
rect 350500 248412 350506 248424
rect 402146 248412 402152 248424
rect 402204 248412 402210 248464
rect 349522 248140 349528 248192
rect 349580 248180 349586 248192
rect 351454 248180 351460 248192
rect 349580 248152 351460 248180
rect 349580 248140 349586 248152
rect 351454 248140 351460 248152
rect 351512 248140 351518 248192
rect 37182 247664 37188 247716
rect 37240 247704 37246 247716
rect 45554 247704 45560 247716
rect 37240 247676 45560 247704
rect 37240 247664 37246 247676
rect 45554 247664 45560 247676
rect 45612 247664 45618 247716
rect 552934 247664 552940 247716
rect 552992 247704 552998 247716
rect 567194 247704 567200 247716
rect 552992 247676 567200 247704
rect 552992 247664 552998 247676
rect 567194 247664 567200 247676
rect 567252 247664 567258 247716
rect 36446 247052 36452 247104
rect 36504 247092 36510 247104
rect 46842 247092 46848 247104
rect 36504 247064 46848 247092
rect 36504 247052 36510 247064
rect 46842 247052 46848 247064
rect 46900 247052 46906 247104
rect 351454 247052 351460 247104
rect 351512 247092 351518 247104
rect 353846 247092 353852 247104
rect 351512 247064 353852 247092
rect 351512 247052 351518 247064
rect 353846 247052 353852 247064
rect 353904 247052 353910 247104
rect 404262 247052 404268 247104
rect 404320 247092 404326 247104
rect 404814 247092 404820 247104
rect 404320 247064 404820 247092
rect 404320 247052 404326 247064
rect 404814 247052 404820 247064
rect 404872 247052 404878 247104
rect 404998 247052 405004 247104
rect 405056 247092 405062 247104
rect 406286 247092 406292 247104
rect 405056 247064 406292 247092
rect 405056 247052 405062 247064
rect 406286 247052 406292 247064
rect 406344 247052 406350 247104
rect 553118 247052 553124 247104
rect 553176 247092 553182 247104
rect 561674 247092 561680 247104
rect 553176 247064 561680 247092
rect 553176 247052 553182 247064
rect 561674 247052 561680 247064
rect 561732 247052 561738 247104
rect 404998 245828 405004 245880
rect 405056 245868 405062 245880
rect 406378 245868 406384 245880
rect 405056 245840 406384 245868
rect 405056 245828 405062 245840
rect 406378 245828 406384 245840
rect 406436 245828 406442 245880
rect 405182 245760 405188 245812
rect 405240 245800 405246 245812
rect 406470 245800 406476 245812
rect 405240 245772 406476 245800
rect 405240 245760 405246 245772
rect 406470 245760 406476 245772
rect 406528 245760 406534 245812
rect 406746 245760 406752 245812
rect 406804 245800 406810 245812
rect 407574 245800 407580 245812
rect 406804 245772 407580 245800
rect 406804 245760 406810 245772
rect 407574 245760 407580 245772
rect 407632 245760 407638 245812
rect 395246 245692 395252 245744
rect 395304 245732 395310 245744
rect 407114 245732 407120 245744
rect 395304 245704 407120 245732
rect 395304 245692 395310 245704
rect 407114 245692 407120 245704
rect 407172 245692 407178 245744
rect 552198 245692 552204 245744
rect 552256 245732 552262 245744
rect 564894 245732 564900 245744
rect 552256 245704 564900 245732
rect 552256 245692 552262 245704
rect 564894 245692 564900 245704
rect 564952 245692 564958 245744
rect 350442 245624 350448 245676
rect 350500 245664 350506 245676
rect 359366 245664 359372 245676
rect 350500 245636 359372 245664
rect 350500 245624 350506 245636
rect 359366 245624 359372 245636
rect 359424 245624 359430 245676
rect 375006 245624 375012 245676
rect 375064 245664 375070 245676
rect 407206 245664 407212 245676
rect 375064 245636 407212 245664
rect 375064 245624 375070 245636
rect 407206 245624 407212 245636
rect 407264 245624 407270 245676
rect 553118 245624 553124 245676
rect 553176 245664 553182 245676
rect 572254 245664 572260 245676
rect 553176 245636 572260 245664
rect 553176 245624 553182 245636
rect 572254 245624 572260 245636
rect 572312 245624 572318 245676
rect 45462 245556 45468 245608
rect 45520 245596 45526 245608
rect 46014 245596 46020 245608
rect 45520 245568 46020 245596
rect 45520 245556 45526 245568
rect 46014 245556 46020 245568
rect 46072 245556 46078 245608
rect 382918 245556 382924 245608
rect 382976 245596 382982 245608
rect 385494 245596 385500 245608
rect 382976 245568 385500 245596
rect 382976 245556 382982 245568
rect 385494 245556 385500 245568
rect 385552 245556 385558 245608
rect 400122 245556 400128 245608
rect 400180 245596 400186 245608
rect 408954 245596 408960 245608
rect 400180 245568 408960 245596
rect 400180 245556 400186 245568
rect 408954 245556 408960 245568
rect 409012 245556 409018 245608
rect 44818 245488 44824 245540
rect 44876 245528 44882 245540
rect 45922 245528 45928 245540
rect 44876 245500 45928 245528
rect 44876 245488 44882 245500
rect 45922 245488 45928 245500
rect 45980 245488 45986 245540
rect 44634 245420 44640 245472
rect 44692 245460 44698 245472
rect 45646 245460 45652 245472
rect 44692 245432 45652 245460
rect 44692 245420 44698 245432
rect 45646 245420 45652 245432
rect 45704 245420 45710 245472
rect 44634 245284 44640 245336
rect 44692 245324 44698 245336
rect 45738 245324 45744 245336
rect 44692 245296 45744 245324
rect 44692 245284 44698 245296
rect 45738 245284 45744 245296
rect 45796 245284 45802 245336
rect 45646 245216 45652 245268
rect 45704 245216 45710 245268
rect 45664 245064 45692 245216
rect 45646 245012 45652 245064
rect 45704 245012 45710 245064
rect 349982 244876 349988 244928
rect 350040 244916 350046 244928
rect 358722 244916 358728 244928
rect 350040 244888 358728 244916
rect 350040 244876 350046 244888
rect 358722 244876 358728 244888
rect 358780 244876 358786 244928
rect 404906 244672 404912 244724
rect 404964 244712 404970 244724
rect 406378 244712 406384 244724
rect 404964 244684 406384 244712
rect 404964 244672 404970 244684
rect 406378 244672 406384 244684
rect 406436 244672 406442 244724
rect 389726 244332 389732 244384
rect 389784 244372 389790 244384
rect 407114 244372 407120 244384
rect 389784 244344 407120 244372
rect 389784 244332 389790 244344
rect 407114 244332 407120 244344
rect 407172 244332 407178 244384
rect 350442 244264 350448 244316
rect 350500 244304 350506 244316
rect 392394 244304 392400 244316
rect 350500 244276 392400 244304
rect 350500 244264 350506 244276
rect 392394 244264 392400 244276
rect 392452 244264 392458 244316
rect 405458 244264 405464 244316
rect 405516 244304 405522 244316
rect 407298 244304 407304 244316
rect 405516 244276 407304 244304
rect 405516 244264 405522 244276
rect 407298 244264 407304 244276
rect 407356 244264 407362 244316
rect 407758 244264 407764 244316
rect 407816 244304 407822 244316
rect 408494 244304 408500 244316
rect 407816 244276 408500 244304
rect 407816 244264 407822 244276
rect 408494 244264 408500 244276
rect 408552 244264 408558 244316
rect 409046 244264 409052 244316
rect 409104 244304 409110 244316
rect 409414 244304 409420 244316
rect 409104 244276 409420 244304
rect 409104 244264 409110 244276
rect 409414 244264 409420 244276
rect 409472 244264 409478 244316
rect 553118 244264 553124 244316
rect 553176 244304 553182 244316
rect 577590 244304 577596 244316
rect 553176 244276 577596 244304
rect 553176 244264 553182 244276
rect 577590 244264 577596 244276
rect 577648 244264 577654 244316
rect 351822 244196 351828 244248
rect 351880 244236 351886 244248
rect 355134 244236 355140 244248
rect 351880 244208 355140 244236
rect 351880 244196 351886 244208
rect 355134 244196 355140 244208
rect 355192 244196 355198 244248
rect 395890 243516 395896 243568
rect 395948 243556 395954 243568
rect 408862 243556 408868 243568
rect 395948 243528 408868 243556
rect 395948 243516 395954 243528
rect 408862 243516 408868 243528
rect 408920 243516 408926 243568
rect 350442 242904 350448 242956
rect 350500 242944 350506 242956
rect 382918 242944 382924 242956
rect 350500 242916 382924 242944
rect 350500 242904 350506 242916
rect 382918 242904 382924 242916
rect 382976 242904 382982 242956
rect 375098 242836 375104 242888
rect 375156 242876 375162 242888
rect 407114 242876 407120 242888
rect 375156 242848 407120 242876
rect 375156 242836 375162 242848
rect 407114 242836 407120 242848
rect 407172 242836 407178 242888
rect 550358 241476 550364 241528
rect 550416 241516 550422 241528
rect 552106 241516 552112 241528
rect 550416 241488 552112 241516
rect 550416 241476 550422 241488
rect 552106 241476 552112 241488
rect 552164 241476 552170 241528
rect 378686 241272 378692 241324
rect 378744 241312 378750 241324
rect 581454 241312 581460 241324
rect 378744 241284 581460 241312
rect 378744 241272 378750 241284
rect 581454 241272 581460 241284
rect 581512 241272 581518 241324
rect 381722 241204 381728 241256
rect 381780 241244 381786 241256
rect 576302 241244 576308 241256
rect 381780 241216 576308 241244
rect 381780 241204 381786 241216
rect 576302 241204 576308 241216
rect 576360 241204 576366 241256
rect 405366 241136 405372 241188
rect 405424 241176 405430 241188
rect 569126 241176 569132 241188
rect 405424 241148 569132 241176
rect 405424 241136 405430 241148
rect 569126 241136 569132 241148
rect 569184 241136 569190 241188
rect 409506 241068 409512 241120
rect 409564 241108 409570 241120
rect 571702 241108 571708 241120
rect 409564 241080 571708 241108
rect 409564 241068 409570 241080
rect 571702 241068 571708 241080
rect 571760 241068 571766 241120
rect 401962 240728 401968 240780
rect 402020 240768 402026 240780
rect 560294 240768 560300 240780
rect 402020 240740 528554 240768
rect 402020 240728 402026 240740
rect 409506 240592 409512 240644
rect 409564 240632 409570 240644
rect 410150 240632 410156 240644
rect 409564 240604 410156 240632
rect 409564 240592 409570 240604
rect 410150 240592 410156 240604
rect 410208 240592 410214 240644
rect 528526 240632 528554 240740
rect 557506 240740 560300 240768
rect 537662 240632 537668 240644
rect 528526 240604 537668 240632
rect 537662 240592 537668 240604
rect 537720 240592 537726 240644
rect 550542 240524 550548 240576
rect 550600 240564 550606 240576
rect 557506 240564 557534 240740
rect 560294 240728 560300 240740
rect 560352 240728 560358 240780
rect 550600 240536 557534 240564
rect 550600 240524 550606 240536
rect 549990 240252 549996 240304
rect 550048 240292 550054 240304
rect 550450 240292 550456 240304
rect 550048 240264 550456 240292
rect 550048 240252 550054 240264
rect 550450 240252 550456 240264
rect 550508 240252 550514 240304
rect 549254 240184 549260 240236
rect 549312 240224 549318 240236
rect 552474 240224 552480 240236
rect 549312 240196 552480 240224
rect 549312 240184 549318 240196
rect 552474 240184 552480 240196
rect 552532 240184 552538 240236
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 32214 240156 32220 240168
rect 3108 240128 32220 240156
rect 3108 240116 3114 240128
rect 32214 240116 32220 240128
rect 32272 240116 32278 240168
rect 549530 240116 549536 240168
rect 549588 240156 549594 240168
rect 550266 240156 550272 240168
rect 549588 240128 550272 240156
rect 549588 240116 549594 240128
rect 550266 240116 550272 240128
rect 550324 240116 550330 240168
rect 550450 240116 550456 240168
rect 550508 240156 550514 240168
rect 554130 240156 554136 240168
rect 550508 240128 554136 240156
rect 550508 240116 550514 240128
rect 554130 240116 554136 240128
rect 554188 240116 554194 240168
rect 391566 240048 391572 240100
rect 391624 240088 391630 240100
rect 566366 240088 566372 240100
rect 391624 240060 566372 240088
rect 391624 240048 391630 240060
rect 566366 240048 566372 240060
rect 566424 240048 566430 240100
rect 395522 239980 395528 240032
rect 395580 240020 395586 240032
rect 396074 240020 396080 240032
rect 395580 239992 396080 240020
rect 395580 239980 395586 239992
rect 396074 239980 396080 239992
rect 396132 239980 396138 240032
rect 400950 239980 400956 240032
rect 401008 240020 401014 240032
rect 573450 240020 573456 240032
rect 401008 239992 573456 240020
rect 401008 239980 401014 239992
rect 573450 239980 573456 239992
rect 573508 239980 573514 240032
rect 397362 239912 397368 239964
rect 397420 239952 397426 239964
rect 568574 239952 568580 239964
rect 397420 239924 568580 239952
rect 397420 239912 397426 239924
rect 568574 239912 568580 239924
rect 568632 239912 568638 239964
rect 396902 239844 396908 239896
rect 396960 239884 396966 239896
rect 564434 239884 564440 239896
rect 396960 239856 564440 239884
rect 396960 239844 396966 239856
rect 564434 239844 564440 239856
rect 564492 239844 564498 239896
rect 402146 239776 402152 239828
rect 402204 239816 402210 239828
rect 567470 239816 567476 239828
rect 402204 239788 567476 239816
rect 402204 239776 402210 239788
rect 567470 239776 567476 239788
rect 567528 239776 567534 239828
rect 349062 239708 349068 239760
rect 349120 239748 349126 239760
rect 349890 239748 349896 239760
rect 349120 239720 349896 239748
rect 349120 239708 349126 239720
rect 349890 239708 349896 239720
rect 349948 239708 349954 239760
rect 408954 239708 408960 239760
rect 409012 239748 409018 239760
rect 566642 239748 566648 239760
rect 409012 239720 566648 239748
rect 409012 239708 409018 239720
rect 566642 239708 566648 239720
rect 566700 239708 566706 239760
rect 409046 239640 409052 239692
rect 409104 239680 409110 239692
rect 552014 239680 552020 239692
rect 409104 239652 552020 239680
rect 409104 239640 409110 239652
rect 552014 239640 552020 239652
rect 552072 239640 552078 239692
rect 409414 239572 409420 239624
rect 409472 239612 409478 239624
rect 550450 239612 550456 239624
rect 409472 239584 550456 239612
rect 409472 239572 409478 239584
rect 550450 239572 550456 239584
rect 550508 239572 550514 239624
rect 552750 239572 552756 239624
rect 552808 239612 552814 239624
rect 561674 239612 561680 239624
rect 552808 239584 561680 239612
rect 552808 239572 552814 239584
rect 561674 239572 561680 239584
rect 561732 239572 561738 239624
rect 549070 239504 549076 239556
rect 549128 239544 549134 239556
rect 568758 239544 568764 239556
rect 549128 239516 568764 239544
rect 549128 239504 549134 239516
rect 568758 239504 568764 239516
rect 568816 239504 568822 239556
rect 382734 239436 382740 239488
rect 382792 239476 382798 239488
rect 547782 239476 547788 239488
rect 382792 239448 547788 239476
rect 382792 239436 382798 239448
rect 547782 239436 547788 239448
rect 547840 239436 547846 239488
rect 552842 239436 552848 239488
rect 552900 239476 552906 239488
rect 577682 239476 577688 239488
rect 552900 239448 577688 239476
rect 552900 239436 552906 239448
rect 577682 239436 577688 239448
rect 577740 239436 577746 239488
rect 350258 239368 350264 239420
rect 350316 239408 350322 239420
rect 547230 239408 547236 239420
rect 350316 239380 547236 239408
rect 350316 239368 350322 239380
rect 547230 239368 547236 239380
rect 547288 239368 547294 239420
rect 547414 239368 547420 239420
rect 547472 239408 547478 239420
rect 547472 239380 567194 239408
rect 547472 239368 547478 239380
rect 567166 239340 567194 239380
rect 569310 239368 569316 239420
rect 569368 239408 569374 239420
rect 571794 239408 571800 239420
rect 569368 239380 571800 239408
rect 569368 239368 569374 239380
rect 571794 239368 571800 239380
rect 571852 239368 571858 239420
rect 574922 239340 574928 239352
rect 567166 239312 574928 239340
rect 574922 239300 574928 239312
rect 574980 239300 574986 239352
rect 350442 238960 350448 239012
rect 350500 239000 350506 239012
rect 457438 239000 457444 239012
rect 350500 238972 457444 239000
rect 350500 238960 350506 238972
rect 457438 238960 457444 238972
rect 457496 238960 457502 239012
rect 535270 238960 535276 239012
rect 535328 239000 535334 239012
rect 551370 239000 551376 239012
rect 535328 238972 551376 239000
rect 535328 238960 535334 238972
rect 551370 238960 551376 238972
rect 551428 238960 551434 239012
rect 381446 238892 381452 238944
rect 381504 238932 381510 238944
rect 463142 238932 463148 238944
rect 381504 238904 463148 238932
rect 381504 238892 381510 238904
rect 463142 238892 463148 238904
rect 463200 238892 463206 238944
rect 506658 238892 506664 238944
rect 506716 238932 506722 238944
rect 555326 238932 555332 238944
rect 506716 238904 555332 238932
rect 506716 238892 506722 238904
rect 555326 238892 555332 238904
rect 555384 238892 555390 238944
rect 350350 238824 350356 238876
rect 350408 238864 350414 238876
rect 355226 238864 355232 238876
rect 350408 238836 355232 238864
rect 350408 238824 350414 238836
rect 355226 238824 355232 238836
rect 355284 238824 355290 238876
rect 405550 238824 405556 238876
rect 405608 238864 405614 238876
rect 504358 238864 504364 238876
rect 405608 238836 504364 238864
rect 405608 238824 405614 238836
rect 504358 238824 504364 238836
rect 504416 238824 504422 238876
rect 505646 238824 505652 238876
rect 505704 238864 505710 238876
rect 570690 238864 570696 238876
rect 505704 238836 570696 238864
rect 505704 238824 505710 238836
rect 570690 238824 570696 238836
rect 570748 238824 570754 238876
rect 350442 238756 350448 238808
rect 350500 238796 350506 238808
rect 386874 238796 386880 238808
rect 350500 238768 386880 238796
rect 350500 238756 350506 238768
rect 386874 238756 386880 238768
rect 386932 238756 386938 238808
rect 398190 238756 398196 238808
rect 398248 238796 398254 238808
rect 427814 238796 427820 238808
rect 398248 238768 427820 238796
rect 398248 238756 398254 238768
rect 427814 238756 427820 238768
rect 427872 238756 427878 238808
rect 436738 238756 436744 238808
rect 436796 238796 436802 238808
rect 551094 238796 551100 238808
rect 436796 238768 551100 238796
rect 436796 238756 436802 238768
rect 551094 238756 551100 238768
rect 551152 238756 551158 238808
rect 36998 238688 37004 238740
rect 37056 238728 37062 238740
rect 46658 238728 46664 238740
rect 37056 238700 46664 238728
rect 37056 238688 37062 238700
rect 46658 238688 46664 238700
rect 46716 238688 46722 238740
rect 403526 238688 403532 238740
rect 403584 238728 403590 238740
rect 545574 238728 545580 238740
rect 403584 238700 545580 238728
rect 403584 238688 403590 238700
rect 545574 238688 545580 238700
rect 545632 238688 545638 238740
rect 547782 238688 547788 238740
rect 547840 238728 547846 238740
rect 564802 238728 564808 238740
rect 547840 238700 564808 238728
rect 547840 238688 547846 238700
rect 564802 238688 564808 238700
rect 564860 238688 564866 238740
rect 390002 238620 390008 238672
rect 390060 238660 390066 238672
rect 528830 238660 528836 238672
rect 390060 238632 528836 238660
rect 390060 238620 390066 238632
rect 528830 238620 528836 238632
rect 528888 238620 528894 238672
rect 532050 238620 532056 238672
rect 532108 238660 532114 238672
rect 558178 238660 558184 238672
rect 532108 238632 558184 238660
rect 532108 238620 532114 238632
rect 558178 238620 558184 238632
rect 558236 238620 558242 238672
rect 399662 238552 399668 238604
rect 399720 238592 399726 238604
rect 440234 238592 440240 238604
rect 399720 238564 440240 238592
rect 399720 238552 399726 238564
rect 440234 238552 440240 238564
rect 440292 238552 440298 238604
rect 447042 238552 447048 238604
rect 447100 238592 447106 238604
rect 570506 238592 570512 238604
rect 447100 238564 570512 238592
rect 447100 238552 447106 238564
rect 570506 238552 570512 238564
rect 570564 238552 570570 238604
rect 395430 238484 395436 238536
rect 395488 238524 395494 238536
rect 416682 238524 416688 238536
rect 395488 238496 416688 238524
rect 395488 238484 395494 238496
rect 416682 238484 416688 238496
rect 416740 238484 416746 238536
rect 497918 238484 497924 238536
rect 497976 238524 497982 238536
rect 556890 238524 556896 238536
rect 497976 238496 556896 238524
rect 497976 238484 497982 238496
rect 556890 238484 556896 238496
rect 556948 238484 556954 238536
rect 398742 238416 398748 238468
rect 398800 238456 398806 238468
rect 432230 238456 432236 238468
rect 398800 238428 432236 238456
rect 398800 238416 398806 238428
rect 432230 238416 432236 238428
rect 432288 238416 432294 238468
rect 445110 238416 445116 238468
rect 445168 238456 445174 238468
rect 554222 238456 554228 238468
rect 445168 238428 554228 238456
rect 445168 238416 445174 238428
rect 554222 238416 554228 238428
rect 554280 238416 554286 238468
rect 392762 238348 392768 238400
rect 392820 238388 392826 238400
rect 454126 238388 454132 238400
rect 392820 238360 454132 238388
rect 392820 238348 392826 238360
rect 454126 238348 454132 238360
rect 454184 238348 454190 238400
rect 457346 238348 457352 238400
rect 457404 238388 457410 238400
rect 551278 238388 551284 238400
rect 457404 238360 551284 238388
rect 457404 238348 457410 238360
rect 551278 238348 551284 238360
rect 551336 238348 551342 238400
rect 409322 238280 409328 238332
rect 409380 238320 409386 238332
rect 442534 238320 442540 238332
rect 409380 238292 442540 238320
rect 409380 238280 409386 238292
rect 442534 238280 442540 238292
rect 442592 238280 442598 238332
rect 470594 238280 470600 238332
rect 470652 238320 470658 238332
rect 556430 238320 556436 238332
rect 470652 238292 556436 238320
rect 470652 238280 470658 238292
rect 556430 238280 556436 238292
rect 556488 238280 556494 238332
rect 401042 238212 401048 238264
rect 401100 238252 401106 238264
rect 428366 238252 428372 238264
rect 401100 238224 428372 238252
rect 401100 238212 401106 238224
rect 428366 238212 428372 238224
rect 428424 238212 428430 238264
rect 472618 238212 472624 238264
rect 472676 238252 472682 238264
rect 550818 238252 550824 238264
rect 472676 238224 550824 238252
rect 472676 238212 472682 238224
rect 550818 238212 550824 238224
rect 550876 238212 550882 238264
rect 403618 238144 403624 238196
rect 403676 238184 403682 238196
rect 422570 238184 422576 238196
rect 403676 238156 422576 238184
rect 403676 238144 403682 238156
rect 422570 238144 422576 238156
rect 422628 238184 422634 238196
rect 423582 238184 423588 238196
rect 422628 238156 423588 238184
rect 422628 238144 422634 238156
rect 423582 238144 423588 238156
rect 423640 238144 423646 238196
rect 476390 238144 476396 238196
rect 476448 238184 476454 238196
rect 554774 238184 554780 238196
rect 476448 238156 554780 238184
rect 476448 238144 476454 238156
rect 554774 238144 554780 238156
rect 554832 238144 554838 238196
rect 421282 238076 421288 238128
rect 421340 238116 421346 238128
rect 543918 238116 543924 238128
rect 421340 238088 543924 238116
rect 421340 238076 421346 238088
rect 543918 238076 543924 238088
rect 543976 238076 543982 238128
rect 36998 238008 37004 238060
rect 37056 238048 37062 238060
rect 45738 238048 45744 238060
rect 37056 238020 45744 238048
rect 37056 238008 37062 238020
rect 45738 238008 45744 238020
rect 45796 238008 45802 238060
rect 414842 238008 414848 238060
rect 414900 238048 414906 238060
rect 541158 238048 541164 238060
rect 414900 238020 541164 238048
rect 414900 238008 414906 238020
rect 541158 238008 541164 238020
rect 541216 238008 541222 238060
rect 549162 238008 549168 238060
rect 549220 238048 549226 238060
rect 583662 238048 583668 238060
rect 549220 238020 583668 238048
rect 549220 238008 549226 238020
rect 583662 238008 583668 238020
rect 583720 238008 583726 238060
rect 416682 237940 416688 237992
rect 416740 237980 416746 237992
rect 490558 237980 490564 237992
rect 416740 237952 490564 237980
rect 416740 237940 416746 237952
rect 490558 237940 490564 237952
rect 490616 237980 490622 237992
rect 491110 237980 491116 237992
rect 490616 237952 491116 237980
rect 490616 237940 490622 237952
rect 491110 237940 491116 237952
rect 491168 237940 491174 237992
rect 501782 237940 501788 237992
rect 501840 237980 501846 237992
rect 547598 237980 547604 237992
rect 501840 237952 547604 237980
rect 501840 237940 501846 237952
rect 547598 237940 547604 237952
rect 547656 237940 547662 237992
rect 423582 237872 423588 237924
rect 423640 237912 423646 237924
rect 482922 237912 482928 237924
rect 423640 237884 482928 237912
rect 423640 237872 423646 237884
rect 482922 237872 482928 237884
rect 482980 237872 482986 237924
rect 528186 237872 528192 237924
rect 528244 237912 528250 237924
rect 560386 237912 560392 237924
rect 528244 237884 560392 237912
rect 528244 237872 528250 237884
rect 560386 237872 560392 237884
rect 560444 237872 560450 237924
rect 391382 237804 391388 237856
rect 391440 237844 391446 237856
rect 515306 237844 515312 237856
rect 391440 237816 515312 237844
rect 391440 237804 391446 237816
rect 515306 237804 515312 237816
rect 515364 237804 515370 237856
rect 544194 237736 544200 237788
rect 544252 237776 544258 237788
rect 560294 237776 560300 237788
rect 544252 237748 560300 237776
rect 544252 237736 544258 237748
rect 560294 237736 560300 237748
rect 560352 237736 560358 237788
rect 529842 237600 529848 237652
rect 529900 237640 529906 237652
rect 547690 237640 547696 237652
rect 529900 237612 547696 237640
rect 529900 237600 529906 237612
rect 547690 237600 547696 237612
rect 547748 237600 547754 237652
rect 541894 237464 541900 237516
rect 541952 237504 541958 237516
rect 549622 237504 549628 237516
rect 541952 237476 549628 237504
rect 541952 237464 541958 237476
rect 549622 237464 549628 237476
rect 549680 237464 549686 237516
rect 413554 237396 413560 237448
rect 413612 237436 413618 237448
rect 414014 237436 414020 237448
rect 413612 237408 414020 237436
rect 413612 237396 413618 237408
rect 414014 237396 414020 237408
rect 414072 237396 414078 237448
rect 482922 237396 482928 237448
rect 482980 237436 482986 237448
rect 483750 237436 483756 237448
rect 482980 237408 483756 237436
rect 482980 237396 482986 237408
rect 483750 237396 483756 237408
rect 483808 237396 483814 237448
rect 547138 237396 547144 237448
rect 547196 237436 547202 237448
rect 547874 237436 547880 237448
rect 547196 237408 547880 237436
rect 547196 237396 547202 237408
rect 547874 237396 547880 237408
rect 547932 237396 547938 237448
rect 560938 237396 560944 237448
rect 560996 237436 561002 237448
rect 561766 237436 561772 237448
rect 560996 237408 561772 237436
rect 560996 237396 561002 237408
rect 561766 237396 561772 237408
rect 561824 237396 561830 237448
rect 350442 237328 350448 237380
rect 350500 237368 350506 237380
rect 370774 237368 370780 237380
rect 350500 237340 370780 237368
rect 350500 237328 350506 237340
rect 370774 237328 370780 237340
rect 370832 237328 370838 237380
rect 391106 237328 391112 237380
rect 391164 237368 391170 237380
rect 583478 237368 583484 237380
rect 391164 237340 583484 237368
rect 391164 237328 391170 237340
rect 583478 237328 583484 237340
rect 583536 237328 583542 237380
rect 385586 237260 385592 237312
rect 385644 237300 385650 237312
rect 573082 237300 573088 237312
rect 385644 237272 573088 237300
rect 385644 237260 385650 237272
rect 573082 237260 573088 237272
rect 573140 237260 573146 237312
rect 394510 237192 394516 237244
rect 394568 237232 394574 237244
rect 580442 237232 580448 237244
rect 394568 237204 580448 237232
rect 394568 237192 394574 237204
rect 580442 237192 580448 237204
rect 580500 237192 580506 237244
rect 395154 237124 395160 237176
rect 395212 237164 395218 237176
rect 578694 237164 578700 237176
rect 395212 237136 578700 237164
rect 395212 237124 395218 237136
rect 578694 237124 578700 237136
rect 578752 237124 578758 237176
rect 384666 237056 384672 237108
rect 384724 237096 384730 237108
rect 567194 237096 567200 237108
rect 384724 237068 567200 237096
rect 384724 237056 384730 237068
rect 567194 237056 567200 237068
rect 567252 237056 567258 237108
rect 389082 236988 389088 237040
rect 389140 237028 389146 237040
rect 569218 237028 569224 237040
rect 389140 237000 569224 237028
rect 389140 236988 389146 237000
rect 569218 236988 569224 237000
rect 569276 236988 569282 237040
rect 405458 236920 405464 236972
rect 405516 236960 405522 236972
rect 582926 236960 582932 236972
rect 405516 236932 582932 236960
rect 405516 236920 405522 236932
rect 582926 236920 582932 236932
rect 582984 236920 582990 236972
rect 402054 236852 402060 236904
rect 402112 236892 402118 236904
rect 574554 236892 574560 236904
rect 402112 236864 574560 236892
rect 402112 236852 402118 236864
rect 574554 236852 574560 236864
rect 574612 236852 574618 236904
rect 398374 236784 398380 236836
rect 398432 236824 398438 236836
rect 552198 236824 552204 236836
rect 398432 236796 552204 236824
rect 398432 236784 398438 236796
rect 552198 236784 552204 236796
rect 552256 236784 552262 236836
rect 560294 236784 560300 236836
rect 560352 236824 560358 236836
rect 560938 236824 560944 236836
rect 560352 236796 560944 236824
rect 560352 236784 560358 236796
rect 560938 236784 560944 236796
rect 560996 236784 561002 236836
rect 395798 236716 395804 236768
rect 395856 236756 395862 236768
rect 532694 236756 532700 236768
rect 395856 236728 532700 236756
rect 395856 236716 395862 236728
rect 532694 236716 532700 236728
rect 532752 236716 532758 236768
rect 547506 236716 547512 236768
rect 547564 236756 547570 236768
rect 567286 236756 567292 236768
rect 547564 236728 567292 236756
rect 547564 236716 547570 236728
rect 567286 236716 567292 236728
rect 567344 236716 567350 236768
rect 417418 236648 417424 236700
rect 417476 236688 417482 236700
rect 550634 236688 550640 236700
rect 417476 236660 550640 236688
rect 417476 236648 417482 236660
rect 550634 236648 550640 236660
rect 550692 236648 550698 236700
rect 404630 236580 404636 236632
rect 404688 236620 404694 236632
rect 514754 236620 514760 236632
rect 404688 236592 514760 236620
rect 404688 236580 404694 236592
rect 514754 236580 514760 236592
rect 514812 236580 514818 236632
rect 478598 236512 478604 236564
rect 478656 236552 478662 236564
rect 550910 236552 550916 236564
rect 478656 236524 550916 236552
rect 478656 236512 478662 236524
rect 550910 236512 550916 236524
rect 550968 236512 550974 236564
rect 499206 236444 499212 236496
rect 499264 236484 499270 236496
rect 555418 236484 555424 236496
rect 499264 236456 555424 236484
rect 499264 236444 499270 236456
rect 555418 236444 555424 236456
rect 555476 236444 555482 236496
rect 42702 235968 42708 236020
rect 42760 236008 42766 236020
rect 43254 236008 43260 236020
rect 42760 235980 43260 236008
rect 42760 235968 42766 235980
rect 43254 235968 43260 235980
rect 43312 235968 43318 236020
rect 396534 235900 396540 235952
rect 396592 235940 396598 235952
rect 580350 235940 580356 235952
rect 396592 235912 580356 235940
rect 396592 235900 396598 235912
rect 580350 235900 580356 235912
rect 580408 235900 580414 235952
rect 404262 235832 404268 235884
rect 404320 235872 404326 235884
rect 549990 235872 549996 235884
rect 404320 235844 549996 235872
rect 404320 235832 404326 235844
rect 549990 235832 549996 235844
rect 550048 235832 550054 235884
rect 474642 235764 474648 235816
rect 474700 235804 474706 235816
rect 541618 235804 541624 235816
rect 474700 235776 541624 235804
rect 474700 235764 474706 235776
rect 541618 235764 541624 235776
rect 541676 235764 541682 235816
rect 481542 235696 481548 235748
rect 481600 235736 481606 235748
rect 570506 235736 570512 235748
rect 481600 235708 570512 235736
rect 481600 235696 481606 235708
rect 570506 235696 570512 235708
rect 570564 235696 570570 235748
rect 393774 235628 393780 235680
rect 393832 235668 393838 235680
rect 527542 235668 527548 235680
rect 393832 235640 527548 235668
rect 393832 235628 393838 235640
rect 527542 235628 527548 235640
rect 527600 235628 527606 235680
rect 528738 235628 528744 235680
rect 528796 235668 528802 235680
rect 568758 235668 568764 235680
rect 528796 235640 568764 235668
rect 528796 235628 528802 235640
rect 568758 235628 568764 235640
rect 568816 235628 568822 235680
rect 370682 235560 370688 235612
rect 370740 235600 370746 235612
rect 511442 235600 511448 235612
rect 370740 235572 511448 235600
rect 370740 235560 370746 235572
rect 511442 235560 511448 235572
rect 511500 235560 511506 235612
rect 524322 235560 524328 235612
rect 524380 235600 524386 235612
rect 564986 235600 564992 235612
rect 524380 235572 564992 235600
rect 524380 235560 524386 235572
rect 564986 235560 564992 235572
rect 565044 235560 565050 235612
rect 430298 235492 430304 235544
rect 430356 235532 430362 235544
rect 573266 235532 573272 235544
rect 430356 235504 573272 235532
rect 430356 235492 430362 235504
rect 573266 235492 573272 235504
rect 573324 235492 573330 235544
rect 395982 235424 395988 235476
rect 396040 235464 396046 235476
rect 565170 235464 565176 235476
rect 396040 235436 565176 235464
rect 396040 235424 396046 235436
rect 565170 235424 565176 235436
rect 565228 235424 565234 235476
rect 385034 235356 385040 235408
rect 385092 235396 385098 235408
rect 556522 235396 556528 235408
rect 385092 235368 556528 235396
rect 385092 235356 385098 235368
rect 556522 235356 556528 235368
rect 556580 235356 556586 235408
rect 376938 235288 376944 235340
rect 376996 235328 377002 235340
rect 555234 235328 555240 235340
rect 376996 235300 555240 235328
rect 376996 235288 377002 235300
rect 555234 235288 555240 235300
rect 555292 235288 555298 235340
rect 378134 235220 378140 235272
rect 378192 235260 378198 235272
rect 559558 235260 559564 235272
rect 378192 235232 559564 235260
rect 378192 235220 378198 235232
rect 559558 235220 559564 235232
rect 559616 235220 559622 235272
rect 493410 235152 493416 235204
rect 493468 235192 493474 235204
rect 557994 235192 558000 235204
rect 493468 235164 558000 235192
rect 493468 235152 493474 235164
rect 557994 235152 558000 235164
rect 558052 235152 558058 235204
rect 488626 235084 488632 235136
rect 488684 235124 488690 235136
rect 551278 235124 551284 235136
rect 488684 235096 551284 235124
rect 488684 235084 488690 235096
rect 551278 235084 551284 235096
rect 551336 235084 551342 235136
rect 491202 235016 491208 235068
rect 491260 235056 491266 235068
rect 552106 235056 552112 235068
rect 491260 235028 552112 235056
rect 491260 235016 491266 235028
rect 552106 235016 552112 235028
rect 552164 235016 552170 235068
rect 44082 234812 44088 234864
rect 44140 234852 44146 234864
rect 45922 234852 45928 234864
rect 44140 234824 45928 234852
rect 44140 234812 44146 234824
rect 45922 234812 45928 234824
rect 45980 234812 45986 234864
rect 30834 234608 30840 234660
rect 30892 234648 30898 234660
rect 46658 234648 46664 234660
rect 30892 234620 46664 234648
rect 30892 234608 30898 234620
rect 46658 234608 46664 234620
rect 46716 234608 46722 234660
rect 350442 234608 350448 234660
rect 350500 234648 350506 234660
rect 360378 234648 360384 234660
rect 350500 234620 360384 234648
rect 350500 234608 350506 234620
rect 360378 234608 360384 234620
rect 360436 234608 360442 234660
rect 453482 234540 453488 234592
rect 453540 234580 453546 234592
rect 571610 234580 571616 234592
rect 453540 234552 571616 234580
rect 453540 234540 453546 234552
rect 571610 234540 571616 234552
rect 571668 234540 571674 234592
rect 436738 234472 436744 234524
rect 436796 234512 436802 234524
rect 559282 234512 559288 234524
rect 436796 234484 559288 234512
rect 436796 234472 436802 234484
rect 559282 234472 559288 234484
rect 559340 234472 559346 234524
rect 456702 234404 456708 234456
rect 456760 234444 456766 234456
rect 580442 234444 580448 234456
rect 456760 234416 580448 234444
rect 456760 234404 456766 234416
rect 580442 234404 580448 234416
rect 580500 234404 580506 234456
rect 401134 234336 401140 234388
rect 401192 234376 401198 234388
rect 541710 234376 541716 234388
rect 401192 234348 541716 234376
rect 401192 234336 401198 234348
rect 541710 234336 541716 234348
rect 541768 234336 541774 234388
rect 400766 234268 400772 234320
rect 400824 234308 400830 234320
rect 545206 234308 545212 234320
rect 400824 234280 545212 234308
rect 400824 234268 400830 234280
rect 545206 234268 545212 234280
rect 545264 234268 545270 234320
rect 393866 234200 393872 234252
rect 393924 234240 393930 234252
rect 544838 234240 544844 234252
rect 393924 234212 544844 234240
rect 393924 234200 393930 234212
rect 544838 234200 544844 234212
rect 544896 234200 544902 234252
rect 394234 234132 394240 234184
rect 394292 234172 394298 234184
rect 544378 234172 544384 234184
rect 394292 234144 544384 234172
rect 394292 234132 394298 234144
rect 544378 234132 544384 234144
rect 544436 234132 544442 234184
rect 388162 234064 388168 234116
rect 388220 234104 388226 234116
rect 552474 234104 552480 234116
rect 388220 234076 552480 234104
rect 388220 234064 388226 234076
rect 552474 234064 552480 234076
rect 552532 234064 552538 234116
rect 43898 233996 43904 234048
rect 43956 234036 43962 234048
rect 45922 234036 45928 234048
rect 43956 234008 45928 234036
rect 43956 233996 43962 234008
rect 45922 233996 45928 234008
rect 45980 233996 45986 234048
rect 398006 233996 398012 234048
rect 398064 234036 398070 234048
rect 578694 234036 578700 234048
rect 398064 234008 578700 234036
rect 398064 233996 398070 234008
rect 578694 233996 578700 234008
rect 578752 233996 578758 234048
rect 349982 233928 349988 233980
rect 350040 233968 350046 233980
rect 541434 233968 541440 233980
rect 350040 233940 541440 233968
rect 350040 233928 350046 233940
rect 541434 233928 541440 233940
rect 541492 233928 541498 233980
rect 543826 233928 543832 233980
rect 543884 233968 543890 233980
rect 544286 233968 544292 233980
rect 543884 233940 544292 233968
rect 543884 233928 543890 233940
rect 544286 233928 544292 233940
rect 544344 233928 544350 233980
rect 355594 233860 355600 233912
rect 355652 233900 355658 233912
rect 554038 233900 554044 233912
rect 355652 233872 554044 233900
rect 355652 233860 355658 233872
rect 554038 233860 554044 233872
rect 554096 233860 554102 233912
rect 409966 233792 409972 233844
rect 410024 233832 410030 233844
rect 410334 233832 410340 233844
rect 410024 233804 410340 233832
rect 410024 233792 410030 233804
rect 410334 233792 410340 233804
rect 410392 233792 410398 233844
rect 418798 233792 418804 233844
rect 418856 233832 418862 233844
rect 419994 233832 420000 233844
rect 418856 233804 420000 233832
rect 418856 233792 418862 233804
rect 419994 233792 420000 233804
rect 420052 233792 420058 233844
rect 461210 233792 461216 233844
rect 461268 233832 461274 233844
rect 562226 233832 562232 233844
rect 461268 233804 562232 233832
rect 461268 233792 461274 233804
rect 562226 233792 562232 233804
rect 562284 233792 562290 233844
rect 409690 233724 409696 233776
rect 409748 233764 409754 233776
rect 491294 233764 491300 233776
rect 409748 233736 491300 233764
rect 409748 233724 409754 233736
rect 491294 233724 491300 233736
rect 491352 233724 491358 233776
rect 406194 233656 406200 233708
rect 406252 233696 406258 233708
rect 472802 233696 472808 233708
rect 406252 233668 472808 233696
rect 406252 233656 406258 233668
rect 472802 233656 472808 233668
rect 472860 233656 472866 233708
rect 45462 233384 45468 233436
rect 45520 233424 45526 233436
rect 45738 233424 45744 233436
rect 45520 233396 45744 233424
rect 45520 233384 45526 233396
rect 45738 233384 45744 233396
rect 45796 233384 45802 233436
rect 349062 233180 349068 233232
rect 349120 233220 349126 233232
rect 349706 233220 349712 233232
rect 349120 233192 349712 233220
rect 349120 233180 349126 233192
rect 349706 233180 349712 233192
rect 349764 233180 349770 233232
rect 390370 233180 390376 233232
rect 390428 233220 390434 233232
rect 580166 233220 580172 233232
rect 390428 233192 580172 233220
rect 390428 233180 390434 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 401502 233112 401508 233164
rect 401560 233152 401566 233164
rect 540422 233152 540428 233164
rect 401560 233124 540428 233152
rect 401560 233112 401566 233124
rect 540422 233112 540428 233124
rect 540480 233112 540486 233164
rect 407574 233044 407580 233096
rect 407632 233084 407638 233096
rect 548518 233084 548524 233096
rect 407632 233056 548524 233084
rect 407632 233044 407638 233056
rect 548518 233044 548524 233056
rect 548576 233044 548582 233096
rect 400030 232976 400036 233028
rect 400088 233016 400094 233028
rect 542538 233016 542544 233028
rect 400088 232988 542544 233016
rect 400088 232976 400094 232988
rect 542538 232976 542544 232988
rect 542596 232976 542602 233028
rect 387610 232908 387616 232960
rect 387668 232948 387674 232960
rect 538858 232948 538864 232960
rect 387668 232920 538864 232948
rect 387668 232908 387674 232920
rect 538858 232908 538864 232920
rect 538916 232908 538922 232960
rect 399846 232840 399852 232892
rect 399904 232880 399910 232892
rect 555602 232880 555608 232892
rect 399904 232852 555608 232880
rect 399904 232840 399910 232852
rect 555602 232840 555608 232852
rect 555660 232840 555666 232892
rect 394602 232772 394608 232824
rect 394660 232812 394666 232824
rect 556982 232812 556988 232824
rect 394660 232784 556988 232812
rect 394660 232772 394666 232784
rect 556982 232772 556988 232784
rect 557040 232772 557046 232824
rect 394326 232704 394332 232756
rect 394384 232744 394390 232756
rect 558178 232744 558184 232756
rect 394384 232716 558184 232744
rect 394384 232704 394390 232716
rect 558178 232704 558184 232716
rect 558236 232704 558242 232756
rect 383562 232636 383568 232688
rect 383620 232676 383626 232688
rect 549898 232676 549904 232688
rect 383620 232648 549904 232676
rect 383620 232636 383626 232648
rect 549898 232636 549904 232648
rect 549956 232636 549962 232688
rect 396810 232568 396816 232620
rect 396868 232608 396874 232620
rect 566642 232608 566648 232620
rect 396868 232580 566648 232608
rect 396868 232568 396874 232580
rect 566642 232568 566648 232580
rect 566700 232568 566706 232620
rect 383470 232500 383476 232552
rect 383528 232540 383534 232552
rect 580350 232540 580356 232552
rect 383528 232512 580356 232540
rect 383528 232500 383534 232512
rect 580350 232500 580356 232512
rect 580408 232500 580414 232552
rect 403434 232432 403440 232484
rect 403492 232472 403498 232484
rect 416774 232472 416780 232484
rect 403492 232444 416780 232472
rect 403492 232432 403498 232444
rect 416774 232432 416780 232444
rect 416832 232432 416838 232484
rect 452562 232432 452568 232484
rect 452620 232472 452626 232484
rect 569126 232472 569132 232484
rect 452620 232444 569132 232472
rect 452620 232432 452626 232444
rect 569126 232432 569132 232444
rect 569184 232432 569190 232484
rect 460934 232364 460940 232416
rect 460992 232404 460998 232416
rect 564802 232404 564808 232416
rect 460992 232376 564808 232404
rect 460992 232364 460998 232376
rect 564802 232364 564808 232376
rect 564860 232364 564866 232416
rect 491110 232296 491116 232348
rect 491168 232336 491174 232348
rect 566274 232336 566280 232348
rect 491168 232308 566280 232336
rect 491168 232296 491174 232308
rect 566274 232296 566280 232308
rect 566332 232296 566338 232348
rect 580166 232228 580172 232280
rect 580224 232268 580230 232280
rect 580442 232268 580448 232280
rect 580224 232240 580448 232268
rect 580224 232228 580230 232240
rect 580442 232228 580448 232240
rect 580500 232228 580506 232280
rect 33962 231820 33968 231872
rect 34020 231860 34026 231872
rect 45554 231860 45560 231872
rect 34020 231832 45560 231860
rect 34020 231820 34026 231832
rect 45554 231820 45560 231832
rect 45612 231820 45618 231872
rect 350442 231820 350448 231872
rect 350500 231860 350506 231872
rect 353846 231860 353852 231872
rect 350500 231832 353852 231860
rect 350500 231820 350506 231832
rect 353846 231820 353852 231832
rect 353904 231820 353910 231872
rect 358538 231752 358544 231804
rect 358596 231792 358602 231804
rect 358998 231792 359004 231804
rect 358596 231764 359004 231792
rect 358596 231752 358602 231764
rect 358998 231752 359004 231764
rect 359056 231752 359062 231804
rect 405642 231208 405648 231260
rect 405700 231248 405706 231260
rect 444466 231248 444472 231260
rect 405700 231220 444472 231248
rect 405700 231208 405706 231220
rect 444466 231208 444472 231220
rect 444524 231208 444530 231260
rect 373810 231140 373816 231192
rect 373868 231180 373874 231192
rect 429194 231180 429200 231192
rect 373868 231152 429200 231180
rect 373868 231140 373874 231152
rect 429194 231140 429200 231152
rect 429252 231140 429258 231192
rect 365070 231072 365076 231124
rect 365128 231112 365134 231124
rect 421926 231112 421932 231124
rect 365128 231084 421932 231112
rect 365128 231072 365134 231084
rect 421926 231072 421932 231084
rect 421984 231072 421990 231124
rect 486970 231072 486976 231124
rect 487028 231112 487034 231124
rect 496814 231112 496820 231124
rect 487028 231084 496820 231112
rect 487028 231072 487034 231084
rect 496814 231072 496820 231084
rect 496872 231072 496878 231124
rect 44082 230732 44088 230784
rect 44140 230772 44146 230784
rect 46934 230772 46940 230784
rect 44140 230744 46940 230772
rect 44140 230732 44146 230744
rect 46934 230732 46940 230744
rect 46992 230732 46998 230784
rect 43898 230528 43904 230580
rect 43956 230568 43962 230580
rect 46014 230568 46020 230580
rect 43956 230540 46020 230568
rect 43956 230528 43962 230540
rect 46014 230528 46020 230540
rect 46072 230528 46078 230580
rect 35250 230460 35256 230512
rect 35308 230500 35314 230512
rect 45554 230500 45560 230512
rect 35308 230472 45560 230500
rect 35308 230460 35314 230472
rect 45554 230460 45560 230472
rect 45612 230460 45618 230512
rect 350442 230460 350448 230512
rect 350500 230500 350506 230512
rect 547322 230500 547328 230512
rect 350500 230472 547328 230500
rect 350500 230460 350506 230472
rect 547322 230460 547328 230472
rect 547380 230460 547386 230512
rect 376294 230392 376300 230444
rect 376352 230432 376358 230444
rect 540330 230432 540336 230444
rect 376352 230404 540336 230432
rect 376352 230392 376358 230404
rect 540330 230392 540336 230404
rect 540388 230392 540394 230444
rect 379330 230324 379336 230376
rect 379388 230364 379394 230376
rect 545850 230364 545856 230376
rect 379388 230336 545856 230364
rect 379388 230324 379394 230336
rect 545850 230324 545856 230336
rect 545908 230324 545914 230376
rect 380710 230256 380716 230308
rect 380768 230296 380774 230308
rect 548058 230296 548064 230308
rect 380768 230268 548064 230296
rect 380768 230256 380774 230268
rect 548058 230256 548064 230268
rect 548116 230256 548122 230308
rect 373166 230188 373172 230240
rect 373224 230228 373230 230240
rect 544654 230228 544660 230240
rect 373224 230200 544660 230228
rect 373224 230188 373230 230200
rect 544654 230188 544660 230200
rect 544712 230188 544718 230240
rect 370866 230120 370872 230172
rect 370924 230160 370930 230172
rect 541802 230160 541808 230172
rect 370924 230132 541808 230160
rect 370924 230120 370930 230132
rect 541802 230120 541808 230132
rect 541860 230120 541866 230172
rect 368290 230052 368296 230104
rect 368348 230092 368354 230104
rect 540514 230092 540520 230104
rect 368348 230064 540520 230092
rect 368348 230052 368354 230064
rect 540514 230052 540520 230064
rect 540572 230052 540578 230104
rect 367922 229984 367928 230036
rect 367980 230024 367986 230036
rect 543090 230024 543096 230036
rect 367980 229996 543096 230024
rect 367980 229984 367986 229996
rect 543090 229984 543096 229996
rect 543148 229984 543154 230036
rect 372246 229916 372252 229968
rect 372304 229956 372310 229968
rect 548242 229956 548248 229968
rect 372304 229928 548248 229956
rect 372304 229916 372310 229928
rect 548242 229916 548248 229928
rect 548300 229916 548306 229968
rect 399754 229848 399760 229900
rect 399812 229888 399818 229900
rect 576302 229888 576308 229900
rect 399812 229860 576308 229888
rect 399812 229848 399818 229860
rect 576302 229848 576308 229860
rect 576360 229848 576366 229900
rect 369762 229780 369768 229832
rect 369820 229820 369826 229832
rect 549346 229820 549352 229832
rect 369820 229792 549352 229820
rect 369820 229780 369826 229792
rect 549346 229780 549352 229792
rect 549404 229780 549410 229832
rect 46382 229712 46388 229764
rect 46440 229752 46446 229764
rect 46566 229752 46572 229764
rect 46440 229724 46572 229752
rect 46440 229712 46446 229724
rect 46566 229712 46572 229724
rect 46624 229712 46630 229764
rect 397270 229712 397276 229764
rect 397328 229752 397334 229764
rect 581822 229752 581828 229764
rect 397328 229724 581828 229752
rect 397328 229712 397334 229724
rect 581822 229712 581828 229724
rect 581880 229712 581886 229764
rect 396994 229644 397000 229696
rect 397052 229684 397058 229696
rect 545942 229684 545948 229696
rect 397052 229656 545948 229684
rect 397052 229644 397058 229656
rect 545942 229644 545948 229656
rect 546000 229644 546006 229696
rect 386874 229576 386880 229628
rect 386932 229616 386938 229628
rect 413554 229616 413560 229628
rect 386932 229588 413560 229616
rect 386932 229576 386938 229588
rect 413554 229576 413560 229588
rect 413612 229576 413618 229628
rect 509326 229576 509332 229628
rect 509384 229616 509390 229628
rect 572070 229616 572076 229628
rect 509384 229588 572076 229616
rect 509384 229576 509390 229588
rect 572070 229576 572076 229588
rect 572128 229576 572134 229628
rect 534718 229236 534724 229288
rect 534776 229276 534782 229288
rect 536834 229276 536840 229288
rect 534776 229248 536840 229276
rect 534776 229236 534782 229248
rect 536834 229236 536840 229248
rect 536892 229236 536898 229288
rect 350442 229100 350448 229152
rect 350500 229140 350506 229152
rect 358998 229140 359004 229152
rect 350500 229112 359004 229140
rect 350500 229100 350506 229112
rect 358998 229100 359004 229112
rect 359056 229100 359062 229152
rect 379422 228352 379428 228404
rect 379480 228392 379486 228404
rect 472066 228392 472072 228404
rect 379480 228364 472072 228392
rect 379480 228352 379486 228364
rect 472066 228352 472072 228364
rect 472124 228352 472130 228404
rect 32306 227740 32312 227792
rect 32364 227780 32370 227792
rect 45554 227780 45560 227792
rect 32364 227752 45560 227780
rect 32364 227740 32370 227752
rect 45554 227740 45560 227752
rect 45612 227740 45618 227792
rect 376478 227332 376484 227384
rect 376536 227372 376542 227384
rect 411622 227372 411628 227384
rect 376536 227344 411628 227372
rect 376536 227332 376542 227344
rect 411622 227332 411628 227344
rect 411680 227332 411686 227384
rect 390278 227264 390284 227316
rect 390336 227304 390342 227316
rect 448330 227304 448336 227316
rect 390336 227276 448336 227304
rect 390336 227264 390342 227276
rect 448330 227264 448336 227276
rect 448388 227264 448394 227316
rect 362218 227196 362224 227248
rect 362276 227236 362282 227248
rect 459922 227236 459928 227248
rect 362276 227208 459928 227236
rect 362276 227196 362282 227208
rect 459922 227196 459928 227208
rect 459980 227196 459986 227248
rect 508498 227196 508504 227248
rect 508556 227236 508562 227248
rect 543826 227236 543832 227248
rect 508556 227208 543832 227236
rect 508556 227196 508562 227208
rect 543826 227196 543832 227208
rect 543884 227196 543890 227248
rect 384758 227128 384764 227180
rect 384816 227168 384822 227180
rect 542998 227168 543004 227180
rect 384816 227140 543004 227168
rect 384816 227128 384822 227140
rect 542998 227128 543004 227140
rect 543056 227128 543062 227180
rect 403894 227060 403900 227112
rect 403952 227100 403958 227112
rect 580442 227100 580448 227112
rect 403952 227072 580448 227100
rect 403952 227060 403958 227072
rect 580442 227060 580448 227072
rect 580500 227060 580506 227112
rect 365254 226992 365260 227044
rect 365312 227032 365318 227044
rect 544102 227032 544108 227044
rect 365312 227004 544108 227032
rect 365312 226992 365318 227004
rect 544102 226992 544108 227004
rect 544160 226992 544166 227044
rect 379146 225700 379152 225752
rect 379204 225740 379210 225752
rect 435450 225740 435456 225752
rect 379204 225712 435456 225740
rect 379204 225700 379210 225712
rect 435450 225700 435456 225712
rect 435508 225700 435514 225752
rect 357158 225632 357164 225684
rect 357216 225672 357222 225684
rect 418062 225672 418068 225684
rect 357216 225644 418068 225672
rect 357216 225632 357222 225644
rect 418062 225632 418068 225644
rect 418120 225632 418126 225684
rect 383378 225564 383384 225616
rect 383436 225604 383442 225616
rect 525794 225604 525800 225616
rect 383436 225576 525800 225604
rect 383436 225564 383442 225576
rect 525794 225564 525800 225576
rect 525852 225564 525858 225616
rect 350350 224884 350356 224936
rect 350408 224924 350414 224936
rect 356422 224924 356428 224936
rect 350408 224896 356428 224924
rect 350408 224884 350414 224896
rect 356422 224884 356428 224896
rect 356480 224884 356486 224936
rect 357066 224340 357072 224392
rect 357124 224380 357130 224392
rect 400214 224380 400220 224392
rect 357124 224352 400220 224380
rect 357124 224340 357130 224352
rect 400214 224340 400220 224352
rect 400272 224340 400278 224392
rect 404722 224340 404728 224392
rect 404780 224380 404786 224392
rect 485038 224380 485044 224392
rect 404780 224352 485044 224380
rect 404780 224340 404786 224352
rect 485038 224340 485044 224352
rect 485096 224340 485102 224392
rect 363782 224272 363788 224324
rect 363840 224312 363846 224324
rect 476666 224312 476672 224324
rect 363840 224284 476672 224312
rect 363840 224272 363846 224284
rect 476666 224272 476672 224284
rect 476724 224272 476730 224324
rect 359642 224204 359648 224256
rect 359700 224244 359706 224256
rect 542446 224244 542452 224256
rect 359700 224216 542452 224244
rect 359700 224204 359706 224216
rect 542446 224204 542452 224216
rect 542504 224204 542510 224256
rect 31110 223592 31116 223644
rect 31168 223632 31174 223644
rect 46658 223632 46664 223644
rect 31168 223604 46664 223632
rect 31168 223592 31174 223604
rect 46658 223592 46664 223604
rect 46716 223592 46722 223644
rect 350442 223524 350448 223576
rect 350500 223564 350506 223576
rect 372338 223564 372344 223576
rect 350500 223536 372344 223564
rect 350500 223524 350506 223536
rect 372338 223524 372344 223536
rect 372396 223524 372402 223576
rect 358722 223456 358728 223508
rect 358780 223496 358786 223508
rect 359642 223496 359648 223508
rect 358780 223468 359648 223496
rect 358780 223456 358786 223468
rect 359642 223456 359648 223468
rect 359700 223456 359706 223508
rect 400674 222912 400680 222964
rect 400732 222952 400738 222964
rect 477954 222952 477960 222964
rect 400732 222924 477960 222952
rect 400732 222912 400738 222924
rect 477954 222912 477960 222924
rect 478012 222912 478018 222964
rect 356882 222844 356888 222896
rect 356940 222884 356946 222896
rect 445754 222884 445760 222896
rect 356940 222856 445760 222884
rect 356940 222844 356946 222856
rect 445754 222844 445760 222856
rect 445812 222844 445818 222896
rect 34790 222164 34796 222216
rect 34848 222204 34854 222216
rect 46658 222204 46664 222216
rect 34848 222176 46664 222204
rect 34848 222164 34854 222176
rect 46658 222164 46664 222176
rect 46716 222164 46722 222216
rect 46566 222096 46572 222148
rect 46624 222136 46630 222148
rect 47578 222136 47584 222148
rect 46624 222108 47584 222136
rect 46624 222096 46630 222108
rect 47578 222096 47584 222108
rect 47636 222096 47642 222148
rect 35342 221688 35348 221740
rect 35400 221728 35406 221740
rect 36354 221728 36360 221740
rect 35400 221700 36360 221728
rect 35400 221688 35406 221700
rect 36354 221688 36360 221700
rect 36412 221688 36418 221740
rect 39942 221688 39948 221740
rect 40000 221728 40006 221740
rect 42058 221728 42064 221740
rect 40000 221700 42064 221728
rect 40000 221688 40006 221700
rect 42058 221688 42064 221700
rect 42116 221688 42122 221740
rect 36998 221416 37004 221468
rect 37056 221456 37062 221468
rect 45922 221456 45928 221468
rect 37056 221428 45928 221456
rect 37056 221416 37062 221428
rect 45922 221416 45928 221428
rect 45980 221416 45986 221468
rect 398466 221416 398472 221468
rect 398524 221456 398530 221468
rect 521654 221456 521660 221468
rect 398524 221428 521660 221456
rect 398524 221416 398530 221428
rect 521654 221416 521660 221428
rect 521712 221416 521718 221468
rect 350442 221144 350448 221196
rect 350500 221184 350506 221196
rect 356514 221184 356520 221196
rect 350500 221156 356520 221184
rect 350500 221144 350506 221156
rect 356514 221144 356520 221156
rect 356572 221144 356578 221196
rect 31202 220804 31208 220856
rect 31260 220844 31266 220856
rect 46658 220844 46664 220856
rect 31260 220816 46664 220844
rect 31260 220804 31266 220816
rect 46658 220804 46664 220816
rect 46716 220804 46722 220856
rect 355410 220736 355416 220788
rect 355468 220776 355474 220788
rect 357618 220776 357624 220788
rect 355468 220748 357624 220776
rect 355468 220736 355474 220748
rect 357618 220736 357624 220748
rect 357676 220736 357682 220788
rect 37642 220260 37648 220312
rect 37700 220300 37706 220312
rect 39298 220300 39304 220312
rect 37700 220272 39304 220300
rect 37700 220260 37706 220272
rect 39298 220260 39304 220272
rect 39356 220260 39362 220312
rect 384114 220056 384120 220108
rect 384172 220096 384178 220108
rect 494054 220096 494060 220108
rect 384172 220068 494060 220096
rect 384172 220056 384178 220068
rect 494054 220056 494060 220068
rect 494112 220056 494118 220108
rect 42610 219444 42616 219496
rect 42668 219484 42674 219496
rect 45830 219484 45836 219496
rect 42668 219456 45836 219484
rect 42668 219444 42674 219456
rect 45830 219444 45836 219456
rect 45888 219444 45894 219496
rect 36906 218696 36912 218748
rect 36964 218736 36970 218748
rect 47670 218736 47676 218748
rect 36964 218708 47676 218736
rect 36964 218696 36970 218708
rect 47670 218696 47676 218708
rect 47728 218696 47734 218748
rect 365162 218696 365168 218748
rect 365220 218736 365226 218748
rect 481174 218736 481180 218748
rect 365220 218708 481180 218736
rect 365220 218696 365226 218708
rect 481174 218696 481180 218708
rect 481232 218696 481238 218748
rect 38102 218628 38108 218680
rect 38160 218668 38166 218680
rect 43622 218668 43628 218680
rect 38160 218640 43628 218668
rect 38160 218628 38166 218640
rect 43622 218628 43628 218640
rect 43680 218628 43686 218680
rect 43162 218560 43168 218612
rect 43220 218600 43226 218612
rect 46014 218600 46020 218612
rect 43220 218572 46020 218600
rect 43220 218560 43226 218572
rect 46014 218560 46020 218572
rect 46072 218560 46078 218612
rect 39298 218084 39304 218136
rect 39356 218124 39362 218136
rect 46658 218124 46664 218136
rect 39356 218096 46664 218124
rect 39356 218084 39362 218096
rect 46658 218084 46664 218096
rect 46716 218084 46722 218136
rect 35434 218016 35440 218068
rect 35492 218056 35498 218068
rect 46106 218056 46112 218068
rect 35492 218028 46112 218056
rect 35492 218016 35498 218028
rect 46106 218016 46112 218028
rect 46164 218016 46170 218068
rect 350442 218016 350448 218068
rect 350500 218056 350506 218068
rect 355042 218056 355048 218068
rect 350500 218028 355048 218056
rect 350500 218016 350506 218028
rect 355042 218016 355048 218028
rect 355100 218016 355106 218068
rect 350350 217948 350356 218000
rect 350408 217988 350414 218000
rect 354950 217988 354956 218000
rect 350408 217960 354956 217988
rect 350408 217948 350414 217960
rect 354950 217948 354956 217960
rect 355008 217948 355014 218000
rect 44082 217336 44088 217388
rect 44140 217376 44146 217388
rect 45738 217376 45744 217388
rect 44140 217348 45744 217376
rect 44140 217336 44146 217348
rect 45738 217336 45744 217348
rect 45796 217336 45802 217388
rect 438670 217336 438676 217388
rect 438728 217376 438734 217388
rect 477586 217376 477592 217388
rect 438728 217348 477592 217376
rect 438728 217336 438734 217348
rect 477586 217336 477592 217348
rect 477644 217336 477650 217388
rect 406654 217268 406660 217320
rect 406712 217308 406718 217320
rect 565998 217308 566004 217320
rect 406712 217280 566004 217308
rect 406712 217268 406718 217280
rect 565998 217268 566004 217280
rect 566056 217268 566062 217320
rect 350442 217200 350448 217252
rect 350500 217240 350506 217252
rect 355226 217240 355232 217252
rect 350500 217212 355232 217240
rect 350500 217200 350506 217212
rect 355226 217200 355232 217212
rect 355284 217200 355290 217252
rect 36906 216724 36912 216776
rect 36964 216764 36970 216776
rect 46290 216764 46296 216776
rect 36964 216736 46296 216764
rect 36964 216724 36970 216736
rect 46290 216724 46296 216736
rect 46348 216724 46354 216776
rect 36998 216656 37004 216708
rect 37056 216696 37062 216708
rect 46658 216696 46664 216708
rect 37056 216668 46664 216696
rect 37056 216656 37062 216668
rect 46658 216656 46664 216668
rect 46716 216656 46722 216708
rect 402422 215908 402428 215960
rect 402480 215948 402486 215960
rect 542814 215948 542820 215960
rect 402480 215920 542820 215948
rect 402480 215908 402486 215920
rect 542814 215908 542820 215920
rect 542872 215908 542878 215960
rect 37734 215296 37740 215348
rect 37792 215336 37798 215348
rect 46658 215336 46664 215348
rect 37792 215308 46664 215336
rect 37792 215296 37798 215308
rect 46658 215296 46664 215308
rect 46716 215296 46722 215348
rect 350442 215296 350448 215348
rect 350500 215336 350506 215348
rect 352742 215336 352748 215348
rect 350500 215308 352748 215336
rect 350500 215296 350506 215308
rect 352742 215296 352748 215308
rect 352800 215296 352806 215348
rect 380618 214548 380624 214600
rect 380676 214588 380682 214600
rect 512086 214588 512092 214600
rect 380676 214560 512092 214588
rect 380676 214548 380682 214560
rect 512086 214548 512092 214560
rect 512144 214548 512150 214600
rect 348602 213868 348608 213920
rect 348660 213908 348666 213920
rect 349338 213908 349344 213920
rect 348660 213880 349344 213908
rect 348660 213868 348666 213880
rect 349338 213868 349344 213880
rect 349396 213868 349402 213920
rect 352650 213868 352656 213920
rect 352708 213908 352714 213920
rect 355134 213908 355140 213920
rect 352708 213880 355140 213908
rect 352708 213868 352714 213880
rect 355134 213868 355140 213880
rect 355192 213868 355198 213920
rect 382642 213256 382648 213308
rect 382700 213296 382706 213308
rect 524966 213296 524972 213308
rect 382700 213268 524972 213296
rect 382700 213256 382706 213268
rect 524966 213256 524972 213268
rect 525024 213256 525030 213308
rect 384298 213188 384304 213240
rect 384356 213228 384362 213240
rect 535914 213228 535920 213240
rect 384356 213200 535920 213228
rect 384356 213188 384362 213200
rect 535914 213188 535920 213200
rect 535972 213188 535978 213240
rect 350442 212508 350448 212560
rect 350500 212548 350506 212560
rect 431218 212548 431224 212560
rect 350500 212520 431224 212548
rect 350500 212508 350506 212520
rect 431218 212508 431224 212520
rect 431276 212508 431282 212560
rect 433334 211760 433340 211812
rect 433392 211800 433398 211812
rect 581454 211800 581460 211812
rect 433392 211772 581460 211800
rect 433392 211760 433398 211772
rect 581454 211760 581460 211772
rect 581512 211760 581518 211812
rect 35066 211148 35072 211200
rect 35124 211188 35130 211200
rect 45554 211188 45560 211200
rect 35124 211160 45560 211188
rect 35124 211148 35130 211160
rect 45554 211148 45560 211160
rect 45612 211148 45618 211200
rect 44634 210536 44640 210588
rect 44692 210576 44698 210588
rect 47762 210576 47768 210588
rect 44692 210548 47768 210576
rect 44692 210536 44698 210548
rect 47762 210536 47768 210548
rect 47820 210536 47826 210588
rect 356790 210468 356796 210520
rect 356848 210508 356854 210520
rect 441614 210508 441620 210520
rect 356848 210480 441620 210508
rect 356848 210468 356854 210480
rect 441614 210468 441620 210480
rect 441672 210468 441678 210520
rect 44726 210400 44732 210452
rect 44784 210440 44790 210452
rect 45646 210440 45652 210452
rect 44784 210412 45652 210440
rect 44784 210400 44790 210412
rect 45646 210400 45652 210412
rect 45704 210400 45710 210452
rect 416958 210400 416964 210452
rect 417016 210440 417022 210452
rect 582926 210440 582932 210452
rect 417016 210412 582932 210440
rect 417016 210400 417022 210412
rect 582926 210400 582932 210412
rect 582984 210400 582990 210452
rect 350442 209856 350448 209908
rect 350500 209896 350506 209908
rect 356606 209896 356612 209908
rect 350500 209868 356612 209896
rect 350500 209856 350506 209868
rect 356606 209856 356612 209868
rect 356664 209856 356670 209908
rect 36354 209040 36360 209092
rect 36412 209080 36418 209092
rect 46290 209080 46296 209092
rect 36412 209052 46296 209080
rect 36412 209040 36418 209052
rect 46290 209040 46296 209052
rect 46348 209040 46354 209092
rect 350442 208360 350448 208412
rect 350500 208400 350506 208412
rect 545022 208400 545028 208412
rect 350500 208372 545028 208400
rect 350500 208360 350506 208372
rect 545022 208360 545028 208372
rect 545080 208360 545086 208412
rect 39574 208292 39580 208344
rect 39632 208332 39638 208344
rect 45554 208332 45560 208344
rect 39632 208304 45560 208332
rect 39632 208292 39638 208304
rect 45554 208292 45560 208304
rect 45612 208292 45618 208344
rect 46382 208292 46388 208344
rect 46440 208332 46446 208344
rect 47394 208332 47400 208344
rect 46440 208304 47400 208332
rect 46440 208292 46446 208304
rect 47394 208292 47400 208304
rect 47452 208292 47458 208344
rect 402606 207680 402612 207732
rect 402664 207720 402670 207732
rect 519170 207720 519176 207732
rect 402664 207692 519176 207720
rect 402664 207680 402670 207692
rect 519170 207680 519176 207692
rect 519228 207680 519234 207732
rect 370590 207612 370596 207664
rect 370648 207652 370654 207664
rect 497918 207652 497924 207664
rect 370648 207624 497924 207652
rect 370648 207612 370654 207624
rect 497918 207612 497924 207624
rect 497976 207612 497982 207664
rect 350442 207068 350448 207120
rect 350500 207108 350506 207120
rect 536098 207108 536104 207120
rect 350500 207080 536104 207108
rect 350500 207068 350506 207080
rect 536098 207068 536104 207080
rect 536156 207068 536162 207120
rect 350350 207000 350356 207052
rect 350408 207040 350414 207052
rect 544194 207040 544200 207052
rect 350408 207012 544200 207040
rect 350408 207000 350414 207012
rect 544194 207000 544200 207012
rect 544252 207000 544258 207052
rect 42426 206932 42432 206984
rect 42484 206972 42490 206984
rect 45646 206972 45652 206984
rect 42484 206944 45652 206972
rect 42484 206932 42490 206944
rect 45646 206932 45652 206944
rect 45704 206932 45710 206984
rect 350442 206932 350448 206984
rect 350500 206972 350506 206984
rect 399386 206972 399392 206984
rect 350500 206944 399392 206972
rect 350500 206932 350506 206944
rect 399386 206932 399392 206944
rect 399444 206932 399450 206984
rect 37182 205640 37188 205692
rect 37240 205680 37246 205692
rect 45646 205680 45652 205692
rect 37240 205652 45652 205680
rect 37240 205640 37246 205652
rect 45646 205640 45652 205652
rect 45704 205640 45710 205692
rect 410058 204892 410064 204944
rect 410116 204932 410122 204944
rect 500218 204932 500224 204944
rect 410116 204904 500224 204932
rect 410116 204892 410122 204904
rect 500218 204892 500224 204904
rect 500276 204892 500282 204944
rect 350350 204280 350356 204332
rect 350408 204320 350414 204332
rect 384298 204320 384304 204332
rect 350408 204292 384304 204320
rect 350408 204280 350414 204292
rect 384298 204280 384304 204292
rect 384356 204280 384362 204332
rect 350442 204212 350448 204264
rect 350500 204252 350506 204264
rect 418798 204252 418804 204264
rect 350500 204224 418804 204252
rect 350500 204212 350506 204224
rect 418798 204212 418804 204224
rect 418856 204212 418862 204264
rect 409874 203600 409880 203652
rect 409932 203640 409938 203652
rect 503714 203640 503720 203652
rect 409932 203612 503720 203640
rect 409932 203600 409938 203612
rect 503714 203600 503720 203612
rect 503772 203600 503778 203652
rect 350074 203532 350080 203584
rect 350132 203572 350138 203584
rect 537754 203572 537760 203584
rect 350132 203544 537760 203572
rect 350132 203532 350138 203544
rect 537754 203532 537760 203544
rect 537812 203532 537818 203584
rect 35710 202852 35716 202904
rect 35768 202892 35774 202904
rect 46658 202892 46664 202904
rect 35768 202864 46664 202892
rect 35768 202852 35774 202864
rect 46658 202852 46664 202864
rect 46716 202852 46722 202904
rect 350442 202852 350448 202904
rect 350500 202892 350506 202904
rect 414658 202892 414664 202904
rect 350500 202864 414664 202892
rect 350500 202852 350506 202864
rect 414658 202852 414664 202864
rect 414716 202852 414722 202904
rect 32950 202784 32956 202836
rect 33008 202824 33014 202836
rect 46382 202824 46388 202836
rect 33008 202796 46388 202824
rect 33008 202784 33014 202796
rect 46382 202784 46388 202796
rect 46440 202784 46446 202836
rect 411346 202104 411352 202156
rect 411404 202144 411410 202156
rect 476022 202144 476028 202156
rect 411404 202116 476028 202144
rect 411404 202104 411410 202116
rect 476022 202104 476028 202116
rect 476080 202104 476086 202156
rect 350442 201492 350448 201544
rect 350500 201532 350506 201544
rect 378686 201532 378692 201544
rect 350500 201504 378692 201532
rect 350500 201492 350506 201504
rect 378686 201492 378692 201504
rect 378744 201492 378750 201544
rect 378686 200812 378692 200864
rect 378744 200852 378750 200864
rect 386506 200852 386512 200864
rect 378744 200824 386512 200852
rect 378744 200812 378750 200824
rect 386506 200812 386512 200824
rect 386564 200812 386570 200864
rect 349890 200744 349896 200796
rect 349948 200784 349954 200796
rect 361758 200784 361764 200796
rect 349948 200756 361764 200784
rect 349948 200744 349954 200756
rect 361758 200744 361764 200756
rect 361816 200744 361822 200796
rect 363322 200744 363328 200796
rect 363380 200784 363386 200796
rect 507854 200784 507860 200796
rect 363380 200756 507860 200784
rect 363380 200744 363386 200756
rect 507854 200744 507860 200756
rect 507912 200744 507918 200796
rect 347774 200240 347780 200252
rect 347700 200212 347780 200240
rect 347700 200104 347728 200212
rect 347774 200200 347780 200212
rect 347832 200200 347838 200252
rect 347774 200104 347780 200116
rect 347700 200076 347780 200104
rect 347774 200064 347780 200076
rect 347832 200064 347838 200116
rect 346210 199860 346216 199912
rect 346268 199900 346274 199912
rect 353570 199900 353576 199912
rect 346268 199872 353576 199900
rect 346268 199860 346274 199872
rect 353570 199860 353576 199872
rect 353628 199860 353634 199912
rect 45002 199656 45008 199708
rect 45060 199696 45066 199708
rect 67082 199696 67088 199708
rect 45060 199668 67088 199696
rect 45060 199656 45066 199668
rect 67082 199656 67088 199668
rect 67140 199656 67146 199708
rect 47486 199588 47492 199640
rect 47544 199628 47550 199640
rect 75914 199628 75920 199640
rect 47544 199600 75920 199628
rect 47544 199588 47550 199600
rect 75914 199588 75920 199600
rect 75972 199588 75978 199640
rect 42610 199520 42616 199572
rect 42668 199560 42674 199572
rect 75454 199560 75460 199572
rect 42668 199532 75460 199560
rect 42668 199520 42674 199532
rect 75454 199520 75460 199532
rect 75512 199520 75518 199572
rect 347590 199520 347596 199572
rect 347648 199560 347654 199572
rect 380802 199560 380808 199572
rect 347648 199532 380808 199560
rect 347648 199520 347654 199532
rect 380802 199520 380808 199532
rect 380860 199520 380866 199572
rect 43898 199452 43904 199504
rect 43956 199492 43962 199504
rect 108942 199492 108948 199504
rect 43956 199464 108948 199492
rect 43956 199452 43962 199464
rect 108942 199452 108948 199464
rect 109000 199452 109006 199504
rect 347498 199452 347504 199504
rect 347556 199492 347562 199504
rect 349338 199492 349344 199504
rect 347556 199464 349344 199492
rect 347556 199452 347562 199464
rect 349338 199452 349344 199464
rect 349396 199452 349402 199504
rect 17402 199384 17408 199436
rect 17460 199424 17466 199436
rect 326982 199424 326988 199436
rect 17460 199396 326988 199424
rect 17460 199384 17466 199396
rect 326982 199384 326988 199396
rect 327040 199384 327046 199436
rect 342990 199384 342996 199436
rect 343048 199424 343054 199436
rect 361022 199424 361028 199436
rect 343048 199396 361028 199424
rect 343048 199384 343054 199396
rect 361022 199384 361028 199396
rect 361080 199384 361086 199436
rect 174262 199316 174268 199368
rect 174320 199356 174326 199368
rect 175090 199356 175096 199368
rect 174320 199328 175096 199356
rect 174320 199316 174326 199328
rect 175090 199316 175096 199328
rect 175148 199316 175154 199368
rect 317230 199316 317236 199368
rect 317288 199356 317294 199368
rect 348510 199356 348516 199368
rect 317288 199328 348516 199356
rect 317288 199316 317294 199328
rect 348510 199316 348516 199328
rect 348568 199316 348574 199368
rect 39666 199248 39672 199300
rect 39724 199288 39730 199300
rect 104618 199288 104624 199300
rect 39724 199260 104624 199288
rect 39724 199248 39730 199260
rect 104618 199248 104624 199260
rect 104676 199248 104682 199300
rect 328178 199248 328184 199300
rect 328236 199288 328242 199300
rect 361666 199288 361672 199300
rect 328236 199260 361672 199288
rect 328236 199248 328242 199260
rect 361666 199248 361672 199260
rect 361724 199248 361730 199300
rect 35526 199180 35532 199232
rect 35584 199220 35590 199232
rect 118786 199220 118792 199232
rect 35584 199192 118792 199220
rect 35584 199180 35590 199192
rect 118786 199180 118792 199192
rect 118844 199180 118850 199232
rect 187786 199180 187792 199232
rect 187844 199220 187850 199232
rect 257982 199220 257988 199232
rect 187844 199192 257988 199220
rect 187844 199180 187850 199192
rect 257982 199180 257988 199192
rect 258040 199180 258046 199232
rect 271506 199180 271512 199232
rect 271564 199220 271570 199232
rect 358446 199220 358452 199232
rect 271564 199192 358452 199220
rect 271564 199180 271570 199192
rect 358446 199180 358452 199192
rect 358504 199180 358510 199232
rect 27246 199112 27252 199164
rect 27304 199152 27310 199164
rect 160094 199152 160100 199164
rect 27304 199124 160100 199152
rect 27304 199112 27310 199124
rect 160094 199112 160100 199124
rect 160152 199112 160158 199164
rect 208394 199112 208400 199164
rect 208452 199152 208458 199164
rect 363690 199152 363696 199164
rect 208452 199124 363696 199152
rect 208452 199112 208458 199124
rect 363690 199112 363696 199124
rect 363748 199112 363754 199164
rect 25590 199044 25596 199096
rect 25648 199084 25654 199096
rect 127250 199084 127256 199096
rect 25648 199056 127256 199084
rect 25648 199044 25654 199056
rect 127250 199044 127256 199056
rect 127308 199044 127314 199096
rect 133046 199044 133052 199096
rect 133104 199084 133110 199096
rect 371326 199084 371332 199096
rect 133104 199056 371332 199084
rect 133104 199044 133110 199056
rect 371326 199044 371332 199056
rect 371384 199044 371390 199096
rect 104066 198976 104072 199028
rect 104124 199016 104130 199028
rect 361114 199016 361120 199028
rect 104124 198988 361120 199016
rect 104124 198976 104130 198988
rect 361114 198976 361120 198988
rect 361172 198976 361178 199028
rect 34054 198908 34060 198960
rect 34112 198948 34118 198960
rect 167822 198948 167828 198960
rect 34112 198920 167828 198948
rect 34112 198908 34118 198920
rect 167822 198908 167828 198920
rect 167880 198908 167886 198960
rect 170398 198908 170404 198960
rect 170456 198948 170462 198960
rect 296070 198948 296076 198960
rect 170456 198920 296076 198948
rect 170456 198908 170462 198920
rect 296070 198908 296076 198920
rect 296128 198908 296134 198960
rect 300486 198908 300492 198960
rect 300544 198948 300550 198960
rect 561030 198948 561036 198960
rect 300544 198920 561036 198948
rect 300544 198908 300550 198920
rect 561030 198908 561036 198920
rect 561088 198908 561094 198960
rect 39942 198840 39948 198892
rect 40000 198880 40006 198892
rect 221918 198880 221924 198892
rect 40000 198852 221924 198880
rect 40000 198840 40006 198852
rect 221918 198840 221924 198852
rect 221976 198840 221982 198892
rect 233510 198840 233516 198892
rect 233568 198880 233574 198892
rect 541894 198880 541900 198892
rect 233568 198852 541900 198880
rect 233568 198840 233574 198852
rect 541894 198840 541900 198852
rect 541952 198840 541958 198892
rect 46658 198772 46664 198824
rect 46716 198812 46722 198824
rect 50338 198812 50344 198824
rect 46716 198784 50344 198812
rect 46716 198772 46722 198784
rect 50338 198772 50344 198784
rect 50396 198772 50402 198824
rect 100846 198772 100852 198824
rect 100904 198812 100910 198824
rect 467926 198812 467932 198824
rect 100904 198784 467932 198812
rect 100904 198772 100910 198784
rect 467926 198772 467932 198784
rect 467984 198772 467990 198824
rect 31662 198704 31668 198756
rect 31720 198744 31726 198756
rect 174906 198744 174912 198756
rect 31720 198716 174912 198744
rect 31720 198704 31726 198716
rect 174906 198704 174912 198716
rect 174964 198704 174970 198756
rect 175090 198704 175096 198756
rect 175148 198744 175154 198756
rect 549530 198744 549536 198756
rect 175148 198716 549536 198744
rect 175148 198704 175154 198716
rect 549530 198704 549536 198716
rect 549588 198704 549594 198756
rect 21818 198636 21824 198688
rect 21876 198676 21882 198688
rect 48682 198676 48688 198688
rect 21876 198648 48688 198676
rect 21876 198636 21882 198648
rect 48682 198636 48688 198648
rect 48740 198636 48746 198688
rect 326982 198636 326988 198688
rect 327040 198676 327046 198688
rect 347590 198676 347596 198688
rect 327040 198648 347596 198676
rect 327040 198636 327046 198648
rect 347590 198636 347596 198648
rect 347648 198636 347654 198688
rect 28718 198568 28724 198620
rect 28776 198608 28782 198620
rect 105998 198608 106004 198620
rect 28776 198580 106004 198608
rect 28776 198568 28782 198580
rect 105998 198568 106004 198580
rect 106056 198568 106062 198620
rect 340414 198568 340420 198620
rect 340472 198608 340478 198620
rect 360194 198608 360200 198620
rect 340472 198580 360200 198608
rect 340472 198568 340478 198580
rect 360194 198568 360200 198580
rect 360252 198568 360258 198620
rect 29914 198500 29920 198552
rect 29972 198540 29978 198552
rect 101490 198540 101496 198552
rect 29972 198512 101496 198540
rect 29972 198500 29978 198512
rect 101490 198500 101496 198512
rect 101548 198500 101554 198552
rect 138198 198500 138204 198552
rect 138256 198540 138262 198552
rect 570782 198540 570788 198552
rect 138256 198512 570788 198540
rect 138256 198500 138262 198512
rect 570782 198500 570788 198512
rect 570840 198500 570846 198552
rect 39206 198432 39212 198484
rect 39264 198472 39270 198484
rect 73798 198472 73804 198484
rect 39264 198444 73804 198472
rect 39264 198432 39270 198444
rect 73798 198432 73804 198444
rect 73856 198432 73862 198484
rect 223850 198432 223856 198484
rect 223908 198472 223914 198484
rect 553854 198472 553860 198484
rect 223908 198444 553860 198472
rect 223908 198432 223914 198444
rect 553854 198432 553860 198444
rect 553912 198432 553918 198484
rect 32858 198364 32864 198416
rect 32916 198404 32922 198416
rect 67358 198404 67364 198416
rect 32916 198376 67364 198404
rect 32916 198364 32922 198376
rect 67358 198364 67364 198376
rect 67416 198364 67422 198416
rect 116302 198364 116308 198416
rect 116360 198404 116366 198416
rect 117958 198404 117964 198416
rect 116360 198376 117964 198404
rect 116360 198364 116366 198376
rect 117958 198364 117964 198376
rect 118016 198364 118022 198416
rect 201954 198364 201960 198416
rect 202012 198404 202018 198416
rect 491386 198404 491392 198416
rect 202012 198376 491392 198404
rect 202012 198364 202018 198376
rect 491386 198364 491392 198376
rect 491444 198364 491450 198416
rect 41138 198296 41144 198348
rect 41196 198336 41202 198348
rect 75638 198336 75644 198348
rect 41196 198308 75644 198336
rect 41196 198296 41202 198308
rect 75638 198296 75644 198308
rect 75696 198296 75702 198348
rect 147858 198296 147864 198348
rect 147916 198336 147922 198348
rect 200758 198336 200764 198348
rect 147916 198308 200764 198336
rect 147916 198296 147922 198308
rect 200758 198296 200764 198308
rect 200816 198296 200822 198348
rect 287606 198296 287612 198348
rect 287664 198336 287670 198348
rect 551186 198336 551192 198348
rect 287664 198308 551192 198336
rect 287664 198296 287670 198308
rect 551186 198296 551192 198308
rect 551244 198296 551250 198348
rect 22738 198228 22744 198280
rect 22796 198268 22802 198280
rect 55766 198268 55772 198280
rect 22796 198240 55772 198268
rect 22796 198228 22802 198240
rect 55766 198228 55772 198240
rect 55824 198228 55830 198280
rect 134334 198228 134340 198280
rect 134392 198268 134398 198280
rect 354766 198268 354772 198280
rect 134392 198240 354772 198268
rect 134392 198228 134398 198240
rect 354766 198228 354772 198240
rect 354824 198228 354830 198280
rect 31570 198160 31576 198212
rect 31628 198200 31634 198212
rect 64138 198200 64144 198212
rect 31628 198172 64144 198200
rect 31628 198160 31634 198172
rect 64138 198160 64144 198172
rect 64196 198160 64202 198212
rect 65058 198160 65064 198212
rect 65116 198200 65122 198212
rect 168466 198200 168472 198212
rect 65116 198172 168472 198200
rect 65116 198160 65122 198172
rect 168466 198160 168472 198172
rect 168524 198160 168530 198212
rect 190362 198160 190368 198212
rect 190420 198200 190426 198212
rect 367830 198200 367836 198212
rect 190420 198172 367836 198200
rect 190420 198160 190426 198172
rect 367830 198160 367836 198172
rect 367888 198160 367894 198212
rect 31478 198092 31484 198144
rect 31536 198132 31542 198144
rect 63586 198132 63592 198144
rect 31536 198104 63592 198132
rect 31536 198092 31542 198104
rect 63586 198092 63592 198104
rect 63644 198092 63650 198144
rect 65518 198092 65524 198144
rect 65576 198132 65582 198144
rect 113726 198132 113732 198144
rect 65576 198104 113732 198132
rect 65576 198092 65582 198104
rect 113726 198092 113732 198104
rect 113784 198092 113790 198144
rect 120718 198092 120724 198144
rect 120776 198132 120782 198144
rect 129826 198132 129832 198144
rect 120776 198104 129832 198132
rect 120776 198092 120782 198104
rect 129826 198092 129832 198104
rect 129884 198092 129890 198144
rect 156874 198092 156880 198144
rect 156932 198132 156938 198144
rect 283558 198132 283564 198144
rect 156932 198104 283564 198132
rect 156932 198092 156938 198104
rect 283558 198092 283564 198104
rect 283616 198092 283622 198144
rect 332042 198092 332048 198144
rect 332100 198132 332106 198144
rect 388346 198132 388352 198144
rect 332100 198104 388352 198132
rect 332100 198092 332106 198104
rect 388346 198092 388352 198104
rect 388404 198092 388410 198144
rect 44542 198024 44548 198076
rect 44600 198064 44606 198076
rect 90910 198064 90916 198076
rect 44600 198036 90916 198064
rect 44600 198024 44606 198036
rect 90910 198024 90916 198036
rect 90968 198024 90974 198076
rect 111150 198024 111156 198076
rect 111208 198064 111214 198076
rect 330478 198064 330484 198076
rect 111208 198036 330484 198064
rect 111208 198024 111214 198036
rect 330478 198024 330484 198036
rect 330536 198024 330542 198076
rect 44910 197956 44916 198008
rect 44968 197996 44974 198008
rect 158530 197996 158536 198008
rect 44968 197968 158536 197996
rect 44968 197956 44974 197968
rect 158530 197956 158536 197968
rect 158588 197956 158594 198008
rect 180058 197956 180064 198008
rect 180116 197996 180122 198008
rect 563882 197996 563888 198008
rect 180116 197968 563888 197996
rect 180116 197956 180122 197968
rect 563882 197956 563888 197968
rect 563940 197956 563946 198008
rect 25774 197888 25780 197940
rect 25832 197928 25838 197940
rect 48038 197928 48044 197940
rect 25832 197900 48044 197928
rect 25832 197888 25838 197900
rect 48038 197888 48044 197900
rect 48096 197888 48102 197940
rect 53282 197888 53288 197940
rect 53340 197928 53346 197940
rect 85298 197928 85304 197940
rect 53340 197900 85304 197928
rect 53340 197888 53346 197900
rect 85298 197888 85304 197900
rect 85356 197888 85362 197940
rect 262490 197888 262496 197940
rect 262548 197928 262554 197940
rect 265618 197928 265624 197940
rect 262548 197900 265624 197928
rect 262548 197888 262554 197900
rect 265618 197888 265624 197900
rect 265676 197888 265682 197940
rect 319806 197888 319812 197940
rect 319864 197928 319870 197940
rect 369118 197928 369124 197940
rect 319864 197900 369124 197928
rect 319864 197888 319870 197900
rect 369118 197888 369124 197900
rect 369176 197888 369182 197940
rect 49234 197820 49240 197872
rect 49292 197860 49298 197872
rect 79594 197860 79600 197872
rect 49292 197832 79600 197860
rect 49292 197820 49298 197832
rect 79594 197820 79600 197832
rect 79652 197820 79658 197872
rect 317874 197820 317880 197872
rect 317932 197860 317938 197872
rect 364978 197860 364984 197872
rect 317932 197832 364984 197860
rect 317932 197820 317938 197832
rect 364978 197820 364984 197832
rect 365036 197820 365042 197872
rect 52822 197752 52828 197804
rect 52880 197792 52886 197804
rect 72510 197792 72516 197804
rect 52880 197764 72516 197792
rect 52880 197752 52886 197764
rect 72510 197752 72516 197764
rect 72568 197752 72574 197804
rect 123386 197752 123392 197804
rect 123444 197792 123450 197804
rect 557074 197792 557080 197804
rect 123444 197764 557080 197792
rect 123444 197752 123450 197764
rect 557074 197752 557080 197764
rect 557132 197752 557138 197804
rect 36906 197684 36912 197736
rect 36964 197724 36970 197736
rect 487154 197724 487160 197736
rect 36964 197696 487160 197724
rect 36964 197684 36970 197696
rect 487154 197684 487160 197696
rect 487212 197684 487218 197736
rect 228450 197480 228456 197532
rect 228508 197520 228514 197532
rect 232866 197520 232872 197532
rect 228508 197492 232872 197520
rect 228508 197480 228514 197492
rect 232866 197480 232872 197492
rect 232924 197480 232930 197532
rect 49326 197344 49332 197396
rect 49384 197384 49390 197396
rect 53098 197384 53104 197396
rect 49384 197356 53104 197384
rect 49384 197344 49390 197356
rect 53098 197344 53104 197356
rect 53156 197344 53162 197396
rect 68278 197344 68284 197396
rect 68336 197384 68342 197396
rect 71130 197384 71136 197396
rect 68336 197356 71136 197384
rect 68336 197344 68342 197356
rect 71130 197344 71136 197356
rect 71188 197344 71194 197396
rect 310698 197344 310704 197396
rect 310756 197384 310762 197396
rect 338114 197384 338120 197396
rect 310756 197356 338120 197384
rect 310756 197344 310762 197356
rect 338114 197344 338120 197356
rect 338172 197344 338178 197396
rect 3418 197276 3424 197328
rect 3476 197316 3482 197328
rect 542354 197316 542360 197328
rect 3476 197288 542360 197316
rect 3476 197276 3482 197288
rect 542354 197276 542360 197288
rect 542412 197276 542418 197328
rect 28350 197208 28356 197260
rect 28408 197248 28414 197260
rect 550450 197248 550456 197260
rect 28408 197220 550456 197248
rect 28408 197208 28414 197220
rect 550450 197208 550456 197220
rect 550508 197208 550514 197260
rect 26970 197140 26976 197192
rect 27028 197180 27034 197192
rect 476206 197180 476212 197192
rect 27028 197152 476212 197180
rect 27028 197140 27034 197152
rect 476206 197140 476212 197152
rect 476264 197140 476270 197192
rect 35250 197072 35256 197124
rect 35308 197112 35314 197124
rect 463694 197112 463700 197124
rect 35308 197084 463700 197112
rect 35308 197072 35314 197084
rect 463694 197072 463700 197084
rect 463752 197072 463758 197124
rect 17310 197004 17316 197056
rect 17368 197044 17374 197056
rect 384206 197044 384212 197056
rect 17368 197016 384212 197044
rect 17368 197004 17374 197016
rect 384206 197004 384212 197016
rect 384264 197004 384270 197056
rect 42702 196936 42708 196988
rect 42760 196976 42766 196988
rect 196802 196976 196808 196988
rect 42760 196948 196808 196976
rect 42760 196936 42766 196948
rect 196802 196936 196808 196948
rect 196860 196936 196866 196988
rect 244458 196936 244464 196988
rect 244516 196976 244522 196988
rect 571886 196976 571892 196988
rect 244516 196948 571892 196976
rect 244516 196936 244522 196948
rect 571886 196936 571892 196948
rect 571944 196936 571950 196988
rect 44082 196868 44088 196920
rect 44140 196908 44146 196920
rect 65058 196908 65064 196920
rect 44140 196880 65064 196908
rect 44140 196868 44146 196880
rect 65058 196868 65064 196880
rect 65116 196868 65122 196920
rect 82170 196868 82176 196920
rect 82228 196908 82234 196920
rect 387426 196908 387432 196920
rect 82228 196880 387432 196908
rect 82228 196868 82234 196880
rect 387426 196868 387432 196880
rect 387484 196868 387490 196920
rect 21450 196800 21456 196852
rect 21508 196840 21514 196852
rect 310698 196840 310704 196852
rect 21508 196812 310704 196840
rect 21508 196800 21514 196812
rect 310698 196800 310704 196812
rect 310756 196800 310762 196852
rect 312722 196800 312728 196852
rect 312780 196840 312786 196852
rect 560846 196840 560852 196852
rect 312780 196812 560852 196840
rect 312780 196800 312786 196812
rect 560846 196800 560852 196812
rect 560904 196800 560910 196852
rect 37090 196732 37096 196784
rect 37148 196772 37154 196784
rect 121454 196772 121460 196784
rect 37148 196744 121460 196772
rect 37148 196732 37154 196744
rect 121454 196732 121460 196744
rect 121512 196732 121518 196784
rect 275370 196732 275376 196784
rect 275428 196772 275434 196784
rect 365806 196772 365812 196784
rect 275428 196744 365812 196772
rect 275428 196732 275434 196744
rect 365806 196732 365812 196744
rect 365864 196732 365870 196784
rect 42334 196664 42340 196716
rect 42392 196704 42398 196716
rect 141786 196704 141792 196716
rect 42392 196676 141792 196704
rect 42392 196664 42398 196676
rect 141786 196664 141792 196676
rect 141844 196664 141850 196716
rect 221642 196664 221648 196716
rect 221700 196704 221706 196716
rect 352374 196704 352380 196716
rect 221700 196676 352380 196704
rect 221700 196664 221706 196676
rect 352374 196664 352380 196676
rect 352432 196664 352438 196716
rect 40586 196596 40592 196648
rect 40644 196636 40650 196648
rect 183002 196636 183008 196648
rect 40644 196608 183008 196636
rect 40644 196596 40650 196608
rect 183002 196596 183008 196608
rect 183060 196596 183066 196648
rect 208118 196596 208124 196648
rect 208176 196636 208182 196648
rect 563422 196636 563428 196648
rect 208176 196608 563428 196636
rect 208176 196596 208182 196608
rect 563422 196596 563428 196608
rect 563480 196596 563486 196648
rect 258994 196528 259000 196580
rect 259052 196568 259058 196580
rect 349430 196568 349436 196580
rect 259052 196540 349436 196568
rect 259052 196528 259058 196540
rect 349430 196528 349436 196540
rect 349488 196528 349494 196580
rect 352006 196500 352012 196512
rect 287026 196472 352012 196500
rect 276014 196392 276020 196444
rect 276072 196432 276078 196444
rect 287026 196432 287054 196472
rect 352006 196460 352012 196472
rect 352064 196460 352070 196512
rect 276072 196404 287054 196432
rect 276072 196392 276078 196404
rect 338114 196392 338120 196444
rect 338172 196432 338178 196444
rect 390186 196432 390192 196444
rect 338172 196404 390192 196432
rect 338172 196392 338178 196404
rect 390186 196392 390192 196404
rect 390244 196392 390250 196444
rect 39758 195916 39764 195968
rect 39816 195956 39822 195968
rect 73522 195956 73528 195968
rect 39816 195928 73528 195956
rect 39816 195916 39822 195928
rect 73522 195916 73528 195928
rect 73580 195916 73586 195968
rect 120166 195916 120172 195968
rect 120224 195956 120230 195968
rect 560570 195956 560576 195968
rect 120224 195928 560576 195956
rect 120224 195916 120230 195928
rect 560570 195916 560576 195928
rect 560628 195916 560634 195968
rect 32214 195848 32220 195900
rect 32272 195888 32278 195900
rect 465074 195888 465080 195900
rect 32272 195860 465080 195888
rect 32272 195848 32278 195860
rect 465074 195848 465080 195860
rect 465132 195848 465138 195900
rect 49510 195780 49516 195832
rect 49568 195820 49574 195832
rect 189074 195820 189080 195832
rect 49568 195792 189080 195820
rect 49568 195780 49574 195792
rect 189074 195780 189080 195792
rect 189132 195780 189138 195832
rect 194226 195780 194232 195832
rect 194284 195820 194290 195832
rect 559466 195820 559472 195832
rect 194284 195792 559472 195820
rect 194284 195780 194290 195792
rect 559466 195780 559472 195792
rect 559524 195780 559530 195832
rect 32398 195712 32404 195764
rect 32456 195752 32462 195764
rect 369670 195752 369676 195764
rect 32456 195724 369676 195752
rect 32456 195712 32462 195724
rect 369670 195712 369676 195724
rect 369728 195712 369734 195764
rect 46750 195644 46756 195696
rect 46808 195684 46814 195696
rect 169110 195684 169116 195696
rect 46808 195656 169116 195684
rect 46808 195644 46814 195656
rect 169110 195644 169116 195656
rect 169168 195644 169174 195696
rect 182634 195644 182640 195696
rect 182692 195684 182698 195696
rect 348418 195684 348424 195696
rect 182692 195656 348424 195684
rect 182692 195644 182698 195656
rect 348418 195644 348424 195656
rect 348476 195644 348482 195696
rect 52270 195576 52276 195628
rect 52328 195616 52334 195628
rect 194870 195616 194876 195628
rect 52328 195588 194876 195616
rect 52328 195576 52334 195588
rect 194870 195576 194876 195588
rect 194928 195576 194934 195628
rect 249610 195576 249616 195628
rect 249668 195616 249674 195628
rect 368106 195616 368112 195628
rect 249668 195588 368112 195616
rect 249668 195576 249674 195588
rect 368106 195576 368112 195588
rect 368164 195576 368170 195628
rect 54846 195508 54852 195560
rect 54904 195548 54910 195560
rect 243078 195548 243084 195560
rect 54904 195520 243084 195548
rect 54904 195508 54910 195520
rect 243078 195508 243084 195520
rect 243136 195508 243142 195560
rect 276658 195508 276664 195560
rect 276716 195548 276722 195560
rect 349798 195548 349804 195560
rect 276716 195520 349804 195548
rect 276716 195508 276722 195520
rect 349798 195508 349804 195520
rect 349856 195508 349862 195560
rect 56042 195440 56048 195492
rect 56100 195480 56106 195492
rect 247678 195480 247684 195492
rect 56100 195452 247684 195480
rect 56100 195440 56106 195452
rect 247678 195440 247684 195452
rect 247736 195440 247742 195492
rect 304350 195440 304356 195492
rect 304408 195480 304414 195492
rect 364334 195480 364340 195492
rect 304408 195452 364340 195480
rect 304408 195440 304414 195452
rect 364334 195440 364340 195452
rect 364392 195440 364398 195492
rect 51534 195372 51540 195424
rect 51592 195412 51598 195424
rect 266906 195412 266912 195424
rect 51592 195384 266912 195412
rect 51592 195372 51598 195384
rect 266906 195372 266912 195384
rect 266964 195372 266970 195424
rect 285398 195372 285404 195424
rect 285456 195412 285462 195424
rect 359090 195412 359096 195424
rect 285456 195384 359096 195412
rect 285456 195372 285462 195384
rect 359090 195372 359096 195384
rect 359148 195372 359154 195424
rect 38286 195304 38292 195356
rect 38344 195344 38350 195356
rect 85574 195344 85580 195356
rect 38344 195316 85580 195344
rect 38344 195304 38350 195316
rect 85574 195304 85580 195316
rect 85632 195304 85638 195356
rect 127986 195304 127992 195356
rect 128044 195344 128050 195356
rect 383194 195344 383200 195356
rect 128044 195316 383200 195344
rect 128044 195304 128050 195316
rect 383194 195304 383200 195316
rect 383252 195304 383258 195356
rect 41966 195236 41972 195288
rect 42024 195276 42030 195288
rect 556614 195276 556620 195288
rect 42024 195248 214144 195276
rect 42024 195236 42030 195248
rect 51718 195168 51724 195220
rect 51776 195208 51782 195220
rect 165246 195208 165252 195220
rect 51776 195180 165252 195208
rect 51776 195168 51782 195180
rect 165246 195168 165252 195180
rect 165304 195168 165310 195220
rect 200114 195168 200120 195220
rect 200172 195208 200178 195220
rect 201310 195208 201316 195220
rect 200172 195180 201316 195208
rect 200172 195168 200178 195180
rect 201310 195168 201316 195180
rect 201368 195168 201374 195220
rect 208394 195168 208400 195220
rect 208452 195208 208458 195220
rect 209590 195208 209596 195220
rect 208452 195180 209596 195208
rect 208452 195168 208458 195180
rect 209590 195168 209596 195180
rect 209648 195168 209654 195220
rect 209774 195168 209780 195220
rect 209832 195208 209838 195220
rect 210970 195208 210976 195220
rect 209832 195180 210976 195208
rect 209832 195168 209838 195180
rect 210970 195168 210976 195180
rect 211028 195168 211034 195220
rect 214116 195152 214144 195248
rect 222304 195248 556620 195276
rect 222304 195152 222332 195248
rect 556614 195236 556620 195248
rect 556672 195236 556678 195288
rect 237374 195168 237380 195220
rect 237432 195208 237438 195220
rect 238570 195208 238576 195220
rect 237432 195180 238576 195208
rect 237432 195168 237438 195180
rect 238570 195168 238576 195180
rect 238628 195168 238634 195220
rect 238754 195168 238760 195220
rect 238812 195208 238818 195220
rect 239950 195208 239956 195220
rect 238812 195180 239956 195208
rect 238812 195168 238818 195180
rect 239950 195168 239956 195180
rect 240008 195168 240014 195220
rect 259454 195168 259460 195220
rect 259512 195208 259518 195220
rect 260558 195208 260564 195220
rect 259512 195180 260564 195208
rect 259512 195168 259518 195180
rect 260558 195168 260564 195180
rect 260616 195168 260622 195220
rect 315298 195168 315304 195220
rect 315356 195208 315362 195220
rect 353478 195208 353484 195220
rect 315356 195180 353484 195208
rect 315356 195168 315362 195180
rect 353478 195168 353484 195180
rect 353536 195168 353542 195220
rect 49418 195100 49424 195152
rect 49476 195140 49482 195152
rect 128446 195140 128452 195152
rect 49476 195112 128452 195140
rect 49476 195100 49482 195112
rect 128446 195100 128452 195112
rect 128504 195100 128510 195152
rect 150526 195100 150532 195152
rect 150584 195140 150590 195152
rect 151722 195140 151728 195152
rect 150584 195112 151728 195140
rect 150584 195100 150590 195112
rect 151722 195100 151728 195112
rect 151780 195100 151786 195152
rect 160186 195100 160192 195152
rect 160244 195140 160250 195152
rect 161382 195140 161388 195152
rect 160244 195112 161388 195140
rect 160244 195100 160250 195112
rect 161382 195100 161388 195112
rect 161440 195100 161446 195152
rect 214098 195100 214104 195152
rect 214156 195100 214162 195152
rect 222286 195100 222292 195152
rect 222344 195100 222350 195152
rect 304994 195100 305000 195152
rect 305052 195140 305058 195152
rect 305546 195140 305552 195152
rect 305052 195112 305552 195140
rect 305052 195100 305058 195112
rect 305546 195100 305552 195112
rect 305604 195100 305610 195152
rect 328454 195100 328460 195152
rect 328512 195140 328518 195152
rect 329374 195140 329380 195152
rect 328512 195112 329380 195140
rect 328512 195100 328518 195112
rect 329374 195100 329380 195112
rect 329432 195100 329438 195152
rect 333974 195100 333980 195152
rect 334032 195140 334038 195152
rect 335262 195140 335268 195152
rect 334032 195112 335268 195140
rect 334032 195100 334038 195112
rect 335262 195100 335268 195112
rect 335320 195100 335326 195152
rect 36262 195032 36268 195084
rect 36320 195072 36326 195084
rect 69014 195072 69020 195084
rect 36320 195044 69020 195072
rect 36320 195032 36326 195044
rect 69014 195032 69020 195044
rect 69072 195032 69078 195084
rect 73338 195032 73344 195084
rect 73396 195072 73402 195084
rect 74442 195072 74448 195084
rect 73396 195044 74448 195072
rect 73396 195032 73402 195044
rect 74442 195032 74448 195044
rect 74500 195032 74506 195084
rect 80054 195032 80060 195084
rect 80112 195072 80118 195084
rect 80790 195072 80796 195084
rect 80112 195044 80796 195072
rect 80112 195032 80118 195044
rect 80790 195032 80796 195044
rect 80848 195032 80854 195084
rect 85574 195032 85580 195084
rect 85632 195072 85638 195084
rect 86402 195072 86408 195084
rect 85632 195044 86408 195072
rect 85632 195032 85638 195044
rect 86402 195032 86408 195044
rect 86460 195032 86466 195084
rect 111794 195032 111800 195084
rect 111852 195072 111858 195084
rect 113082 195072 113088 195084
rect 111852 195044 113088 195072
rect 111852 195032 111858 195044
rect 113082 195032 113088 195044
rect 113140 195032 113146 195084
rect 40218 194828 40224 194880
rect 40276 194868 40282 194880
rect 45922 194868 45928 194880
rect 40276 194840 45928 194868
rect 40276 194828 40282 194840
rect 45922 194828 45928 194840
rect 45980 194828 45986 194880
rect 127066 194556 127072 194608
rect 127124 194596 127130 194608
rect 127986 194596 127992 194608
rect 127124 194568 127992 194596
rect 127124 194556 127130 194568
rect 127986 194556 127992 194568
rect 128044 194556 128050 194608
rect 20162 194488 20168 194540
rect 20220 194528 20226 194540
rect 573358 194528 573364 194540
rect 20220 194500 573364 194528
rect 20220 194488 20226 194500
rect 573358 194488 573364 194500
rect 573416 194488 573422 194540
rect 29546 194420 29552 194472
rect 29604 194460 29610 194472
rect 567562 194460 567568 194472
rect 29604 194432 567568 194460
rect 29604 194420 29610 194432
rect 567562 194420 567568 194432
rect 567620 194420 567626 194472
rect 33686 194352 33692 194404
rect 33744 194392 33750 194404
rect 519078 194392 519084 194404
rect 33744 194364 519084 194392
rect 33744 194352 33750 194364
rect 519078 194352 519084 194364
rect 519136 194352 519142 194404
rect 41230 194284 41236 194336
rect 41288 194324 41294 194336
rect 89254 194324 89260 194336
rect 41288 194296 89260 194324
rect 41288 194284 41294 194296
rect 89254 194284 89260 194296
rect 89312 194284 89318 194336
rect 205174 194284 205180 194336
rect 205232 194324 205238 194336
rect 574278 194324 574284 194336
rect 205232 194296 574284 194324
rect 205232 194284 205238 194296
rect 574278 194284 574284 194296
rect 574336 194284 574342 194336
rect 22646 194216 22652 194268
rect 22704 194256 22710 194268
rect 330754 194256 330760 194268
rect 22704 194228 330760 194256
rect 22704 194216 22710 194228
rect 330754 194216 330760 194228
rect 330812 194216 330818 194268
rect 342714 194216 342720 194268
rect 342772 194256 342778 194268
rect 354030 194256 354036 194268
rect 342772 194228 354036 194256
rect 342772 194216 342778 194228
rect 354030 194216 354036 194228
rect 354088 194216 354094 194268
rect 51258 194148 51264 194200
rect 51316 194188 51322 194200
rect 54570 194188 54576 194200
rect 51316 194160 54576 194188
rect 51316 194148 51322 194160
rect 54570 194148 54576 194160
rect 54628 194148 54634 194200
rect 116946 194148 116952 194200
rect 117004 194188 117010 194200
rect 399570 194188 399576 194200
rect 117004 194160 399576 194188
rect 117004 194148 117010 194160
rect 399570 194148 399576 194160
rect 399628 194148 399634 194200
rect 181346 194080 181352 194132
rect 181404 194120 181410 194132
rect 449894 194120 449900 194132
rect 181404 194092 449900 194120
rect 181404 194080 181410 194092
rect 449894 194080 449900 194092
rect 449952 194080 449958 194132
rect 102134 194012 102140 194064
rect 102192 194052 102198 194064
rect 366634 194052 366640 194064
rect 102192 194024 366640 194052
rect 102192 194012 102198 194024
rect 366634 194012 366640 194024
rect 366692 194012 366698 194064
rect 281166 193944 281172 193996
rect 281224 193984 281230 193996
rect 356146 193984 356152 193996
rect 281224 193956 356152 193984
rect 281224 193944 281230 193956
rect 356146 193944 356152 193956
rect 356204 193944 356210 193996
rect 241238 193876 241244 193928
rect 241296 193916 241302 193928
rect 362402 193916 362408 193928
rect 241296 193888 362408 193916
rect 241296 193876 241302 193888
rect 362402 193876 362408 193888
rect 362460 193876 362466 193928
rect 50430 193808 50436 193860
rect 50488 193848 50494 193860
rect 356514 193848 356520 193860
rect 50488 193820 356520 193848
rect 50488 193808 50494 193820
rect 356514 193808 356520 193820
rect 356572 193808 356578 193860
rect 169754 193740 169760 193792
rect 169812 193780 169818 193792
rect 352650 193780 352656 193792
rect 169812 193752 352656 193780
rect 169812 193740 169818 193752
rect 352650 193740 352656 193752
rect 352708 193740 352714 193792
rect 21726 193672 21732 193724
rect 21784 193712 21790 193724
rect 246390 193712 246396 193724
rect 21784 193684 246396 193712
rect 21784 193672 21790 193684
rect 246390 193672 246396 193684
rect 246448 193672 246454 193724
rect 248414 193672 248420 193724
rect 248472 193712 248478 193724
rect 358630 193712 358636 193724
rect 248472 193684 358636 193712
rect 248472 193672 248478 193684
rect 358630 193672 358636 193684
rect 358688 193672 358694 193724
rect 17218 193604 17224 193656
rect 17276 193644 17282 193656
rect 281718 193644 281724 193656
rect 17276 193616 281724 193644
rect 17276 193604 17282 193616
rect 281718 193604 281724 193616
rect 281776 193604 281782 193656
rect 295702 193604 295708 193656
rect 295760 193644 295766 193656
rect 350534 193644 350540 193656
rect 295760 193616 350540 193644
rect 295760 193604 295766 193616
rect 350534 193604 350540 193616
rect 350592 193604 350598 193656
rect 25314 193128 25320 193180
rect 25372 193168 25378 193180
rect 570414 193168 570420 193180
rect 25372 193140 570420 193168
rect 25372 193128 25378 193140
rect 570414 193128 570420 193140
rect 570472 193128 570478 193180
rect 571978 193128 571984 193180
rect 572036 193168 572042 193180
rect 580258 193168 580264 193180
rect 572036 193140 580264 193168
rect 572036 193128 572042 193140
rect 580258 193128 580264 193140
rect 580316 193128 580322 193180
rect 24026 193060 24032 193112
rect 24084 193100 24090 193112
rect 566458 193100 566464 193112
rect 24084 193072 566464 193100
rect 24084 193060 24090 193072
rect 566458 193060 566464 193072
rect 566516 193060 566522 193112
rect 26694 192992 26700 193044
rect 26752 193032 26758 193044
rect 478874 193032 478880 193044
rect 26752 193004 478880 193032
rect 26752 192992 26758 193004
rect 478874 192992 478880 193004
rect 478932 192992 478938 193044
rect 142062 192924 142068 192976
rect 142120 192964 142126 192976
rect 529934 192964 529940 192976
rect 142120 192936 529940 192964
rect 142120 192924 142126 192936
rect 529934 192924 529940 192936
rect 529992 192924 529998 192976
rect 30006 192856 30012 192908
rect 30064 192896 30070 192908
rect 337838 192896 337844 192908
rect 30064 192868 337844 192896
rect 30064 192856 30070 192868
rect 337838 192856 337844 192868
rect 337896 192856 337902 192908
rect 34054 192788 34060 192840
rect 34112 192828 34118 192840
rect 230934 192828 230940 192840
rect 34112 192800 230940 192828
rect 34112 192788 34118 192800
rect 230934 192788 230940 192800
rect 230992 192788 230998 192840
rect 278590 192788 278596 192840
rect 278648 192828 278654 192840
rect 351454 192828 351460 192840
rect 278648 192800 351460 192828
rect 278648 192788 278654 192800
rect 351454 192788 351460 192800
rect 351512 192788 351518 192840
rect 44634 192720 44640 192772
rect 44692 192760 44698 192772
rect 263778 192760 263784 192772
rect 44692 192732 263784 192760
rect 44692 192720 44698 192732
rect 263778 192720 263784 192732
rect 263836 192720 263842 192772
rect 280522 192720 280528 192772
rect 280580 192760 280586 192772
rect 353386 192760 353392 192772
rect 280580 192732 353392 192760
rect 280580 192720 280586 192732
rect 353386 192720 353392 192732
rect 353444 192720 353450 192772
rect 48038 192652 48044 192704
rect 48096 192692 48102 192704
rect 333330 192692 333336 192704
rect 48096 192664 333336 192692
rect 48096 192652 48102 192664
rect 333330 192652 333336 192664
rect 333388 192652 333394 192704
rect 36906 192584 36912 192636
rect 36964 192624 36970 192636
rect 326890 192624 326896 192636
rect 36964 192596 326896 192624
rect 36964 192584 36970 192596
rect 326890 192584 326896 192596
rect 326948 192584 326954 192636
rect 339494 192584 339500 192636
rect 339552 192624 339558 192636
rect 352558 192624 352564 192636
rect 339552 192596 352564 192624
rect 339552 192584 339558 192596
rect 352558 192584 352564 192596
rect 352616 192584 352622 192636
rect 52178 192516 52184 192568
rect 52236 192556 52242 192568
rect 360378 192556 360384 192568
rect 52236 192528 360384 192556
rect 52236 192516 52242 192528
rect 360378 192516 360384 192528
rect 360436 192516 360442 192568
rect 4798 192448 4804 192500
rect 4856 192488 4862 192500
rect 506474 192488 506480 192500
rect 4856 192460 506480 192488
rect 4856 192448 4862 192460
rect 506474 192448 506480 192460
rect 506532 192448 506538 192500
rect 31570 192380 31576 192432
rect 31628 192420 31634 192432
rect 216122 192420 216128 192432
rect 31628 192392 216128 192420
rect 31628 192380 31634 192392
rect 216122 192380 216128 192392
rect 216180 192380 216186 192432
rect 37090 192312 37096 192364
rect 37148 192352 37154 192364
rect 172974 192352 172980 192364
rect 37148 192324 172980 192352
rect 37148 192312 37154 192324
rect 172974 192312 172980 192324
rect 173032 192312 173038 192364
rect 192018 192312 192024 192364
rect 192076 192352 192082 192364
rect 359182 192352 359188 192364
rect 192076 192324 359188 192352
rect 192076 192312 192082 192324
rect 359182 192312 359188 192324
rect 359240 192312 359246 192364
rect 46290 192244 46296 192296
rect 46348 192284 46354 192296
rect 151814 192284 151820 192296
rect 46348 192256 151820 192284
rect 46348 192244 46354 192256
rect 151814 192244 151820 192256
rect 151872 192244 151878 192296
rect 204530 192244 204536 192296
rect 204588 192284 204594 192296
rect 354674 192284 354680 192296
rect 204588 192256 354680 192284
rect 204588 192244 204594 192256
rect 354674 192244 354680 192256
rect 354732 192244 354738 192296
rect 17494 191768 17500 191820
rect 17552 191808 17558 191820
rect 575934 191808 575940 191820
rect 17552 191780 575940 191808
rect 17552 191768 17558 191780
rect 575934 191768 575940 191780
rect 575992 191768 575998 191820
rect 56318 191700 56324 191752
rect 56376 191740 56382 191752
rect 180702 191740 180708 191752
rect 56376 191712 180708 191740
rect 56376 191700 56382 191712
rect 180702 191700 180708 191712
rect 180760 191700 180766 191752
rect 183922 191700 183928 191752
rect 183980 191740 183986 191752
rect 582650 191740 582656 191752
rect 183980 191712 582656 191740
rect 183980 191700 183986 191712
rect 582650 191700 582656 191712
rect 582708 191700 582714 191752
rect 146294 191632 146300 191684
rect 146352 191672 146358 191684
rect 356330 191672 356336 191684
rect 146352 191644 356336 191672
rect 146352 191632 146358 191644
rect 356330 191632 356336 191644
rect 356388 191632 356394 191684
rect 116670 191564 116676 191616
rect 116728 191604 116734 191616
rect 348234 191604 348240 191616
rect 116728 191576 348240 191604
rect 116728 191564 116734 191576
rect 348234 191564 348240 191576
rect 348292 191564 348298 191616
rect 297910 191496 297916 191548
rect 297968 191536 297974 191548
rect 358538 191536 358544 191548
rect 297968 191508 358544 191536
rect 297968 191496 297974 191508
rect 358538 191496 358544 191508
rect 358596 191496 358602 191548
rect 46842 191428 46848 191480
rect 46900 191468 46906 191480
rect 355686 191468 355692 191480
rect 46900 191440 355692 191468
rect 46900 191428 46906 191440
rect 355686 191428 355692 191440
rect 355744 191428 355750 191480
rect 50798 191360 50804 191412
rect 50856 191400 50862 191412
rect 361850 191400 361856 191412
rect 50856 191372 361856 191400
rect 50856 191360 50862 191372
rect 361850 191360 361856 191372
rect 361908 191360 361914 191412
rect 48222 191292 48228 191344
rect 48280 191332 48286 191344
rect 384482 191332 384488 191344
rect 48280 191304 384488 191332
rect 48280 191292 48286 191304
rect 384482 191292 384488 191304
rect 384540 191292 384546 191344
rect 3418 191224 3424 191276
rect 3476 191264 3482 191276
rect 365346 191264 365352 191276
rect 3476 191236 365352 191264
rect 3476 191224 3482 191236
rect 365346 191224 365352 191236
rect 365404 191224 365410 191276
rect 121454 191156 121460 191208
rect 121512 191196 121518 191208
rect 569310 191196 569316 191208
rect 121512 191168 569316 191196
rect 121512 191156 121518 191168
rect 569310 191156 569316 191168
rect 569368 191156 569374 191208
rect 35894 191088 35900 191140
rect 35952 191128 35958 191140
rect 555510 191128 555516 191140
rect 35952 191100 555516 191128
rect 35952 191088 35958 191100
rect 555510 191088 555516 191100
rect 555568 191088 555574 191140
rect 209406 191020 209412 191072
rect 209464 191060 209470 191072
rect 354858 191060 354864 191072
rect 209464 191032 354864 191060
rect 209464 191020 209470 191032
rect 354858 191020 354864 191032
rect 354916 191020 354922 191072
rect 58618 190952 58624 191004
rect 58676 190992 58682 191004
rect 314010 190992 314016 191004
rect 58676 190964 314016 190992
rect 58676 190952 58682 190964
rect 314010 190952 314016 190964
rect 314068 190952 314074 191004
rect 19978 190408 19984 190460
rect 20036 190448 20042 190460
rect 395706 190448 395712 190460
rect 20036 190420 395712 190448
rect 20036 190408 20042 190420
rect 395706 190408 395712 190420
rect 395764 190408 395770 190460
rect 173618 190340 173624 190392
rect 173676 190380 173682 190392
rect 359642 190380 359648 190392
rect 173676 190352 359648 190380
rect 173676 190340 173682 190352
rect 359642 190340 359648 190352
rect 359700 190340 359706 190392
rect 58710 190272 58716 190324
rect 58768 190312 58774 190324
rect 236730 190312 236736 190324
rect 58768 190284 236736 190312
rect 58768 190272 58774 190284
rect 236730 190272 236736 190284
rect 236788 190272 236794 190324
rect 242894 190272 242900 190324
rect 242952 190312 242958 190324
rect 367094 190312 367100 190324
rect 242952 190284 367100 190312
rect 242952 190272 242958 190284
rect 367094 190272 367100 190284
rect 367152 190272 367158 190324
rect 59630 190204 59636 190256
rect 59688 190244 59694 190256
rect 256050 190244 256056 190256
rect 59688 190216 256056 190244
rect 59688 190204 59694 190216
rect 256050 190204 256056 190216
rect 256108 190204 256114 190256
rect 287698 190204 287704 190256
rect 287756 190244 287762 190256
rect 480346 190244 480352 190256
rect 287756 190216 480352 190244
rect 287756 190204 287762 190216
rect 480346 190204 480352 190216
rect 480404 190204 480410 190256
rect 59906 190136 59912 190188
rect 59964 190176 59970 190188
rect 294690 190176 294696 190188
rect 59964 190148 294696 190176
rect 59964 190136 59970 190148
rect 294690 190136 294696 190148
rect 294748 190136 294754 190188
rect 322106 190136 322112 190188
rect 322164 190176 322170 190188
rect 558086 190176 558092 190188
rect 322164 190148 558092 190176
rect 322164 190136 322170 190148
rect 558086 190136 558092 190148
rect 558144 190136 558150 190188
rect 59170 190068 59176 190120
rect 59228 190108 59234 190120
rect 349154 190108 349160 190120
rect 59228 190080 349160 190108
rect 59228 190068 59234 190080
rect 349154 190068 349160 190080
rect 349212 190068 349218 190120
rect 58526 190000 58532 190052
rect 58584 190040 58590 190052
rect 355226 190040 355232 190052
rect 58584 190012 355232 190040
rect 58584 190000 58590 190012
rect 355226 190000 355232 190012
rect 355284 190000 355290 190052
rect 59814 189932 59820 189984
rect 59872 189972 59878 189984
rect 369946 189972 369952 189984
rect 59872 189944 369952 189972
rect 59872 189932 59878 189944
rect 369946 189932 369952 189944
rect 370004 189932 370010 189984
rect 35526 189864 35532 189916
rect 35584 189904 35590 189916
rect 370222 189904 370228 189916
rect 35584 189876 370228 189904
rect 35584 189864 35590 189876
rect 370222 189864 370228 189876
rect 370280 189864 370286 189916
rect 59538 189796 59544 189848
rect 59596 189836 59602 189848
rect 396074 189836 396080 189848
rect 59596 189808 396080 189836
rect 59596 189796 59602 189808
rect 396074 189796 396080 189808
rect 396132 189796 396138 189848
rect 31662 189728 31668 189780
rect 31720 189768 31726 189780
rect 373442 189768 373448 189780
rect 31720 189740 373448 189768
rect 31720 189728 31726 189740
rect 373442 189728 373448 189740
rect 373500 189728 373506 189780
rect 184566 189660 184572 189712
rect 184624 189700 184630 189712
rect 354122 189700 354128 189712
rect 184624 189672 354128 189700
rect 184624 189660 184630 189672
rect 354122 189660 354128 189672
rect 354180 189660 354186 189712
rect 198090 189592 198096 189644
rect 198148 189632 198154 189644
rect 302142 189632 302148 189644
rect 198148 189604 302148 189632
rect 198148 189592 198154 189604
rect 302142 189592 302148 189604
rect 302200 189592 302206 189644
rect 249978 189524 249984 189576
rect 250036 189564 250042 189576
rect 352282 189564 352288 189576
rect 250036 189536 352288 189564
rect 250036 189524 250042 189536
rect 352282 189524 352288 189536
rect 352340 189524 352346 189576
rect 21266 188980 21272 189032
rect 21324 189020 21330 189032
rect 581730 189020 581736 189032
rect 21324 188992 581736 189020
rect 21324 188980 21330 188992
rect 581730 188980 581736 188992
rect 581788 188980 581794 189032
rect 3510 188912 3516 188964
rect 3568 188952 3574 188964
rect 392670 188952 392676 188964
rect 3568 188924 392676 188952
rect 3568 188912 3574 188924
rect 392670 188912 392676 188924
rect 392728 188912 392734 188964
rect 195146 188844 195152 188896
rect 195204 188884 195210 188896
rect 201494 188884 201500 188896
rect 195204 188856 201500 188884
rect 195204 188844 195210 188856
rect 201494 188844 201500 188856
rect 201552 188844 201558 188896
rect 272518 188844 272524 188896
rect 272576 188884 272582 188896
rect 351086 188884 351092 188896
rect 272576 188856 351092 188884
rect 272576 188844 272582 188856
rect 351086 188844 351092 188856
rect 351144 188844 351150 188896
rect 226150 188776 226156 188828
rect 226208 188816 226214 188828
rect 324406 188816 324412 188828
rect 226208 188788 324412 188816
rect 226208 188776 226214 188788
rect 324406 188776 324412 188788
rect 324464 188776 324470 188828
rect 43162 188708 43168 188760
rect 43220 188748 43226 188760
rect 303706 188748 303712 188760
rect 43220 188720 303712 188748
rect 43220 188708 43226 188720
rect 303706 188708 303712 188720
rect 303764 188708 303770 188760
rect 255774 188640 255780 188692
rect 255832 188680 255838 188692
rect 555142 188680 555148 188692
rect 255832 188652 555148 188680
rect 255832 188640 255838 188652
rect 555142 188640 555148 188652
rect 555200 188640 555206 188692
rect 43254 188572 43260 188624
rect 43312 188612 43318 188624
rect 363138 188612 363144 188624
rect 43312 188584 363144 188612
rect 43312 188572 43318 188584
rect 363138 188572 363144 188584
rect 363196 188572 363202 188624
rect 41874 188504 41880 188556
rect 41932 188544 41938 188556
rect 363046 188544 363052 188556
rect 41932 188516 363052 188544
rect 41932 188504 41938 188516
rect 363046 188504 363052 188516
rect 363104 188504 363110 188556
rect 50614 188436 50620 188488
rect 50672 188476 50678 188488
rect 373994 188476 374000 188488
rect 50672 188448 374000 188476
rect 50672 188436 50678 188448
rect 373994 188436 374000 188448
rect 374052 188436 374058 188488
rect 34146 188368 34152 188420
rect 34204 188408 34210 188420
rect 371878 188408 371884 188420
rect 34204 188380 371884 188408
rect 34204 188368 34210 188380
rect 371878 188368 371884 188380
rect 371936 188368 371942 188420
rect 48958 188300 48964 188352
rect 49016 188340 49022 188352
rect 426526 188340 426532 188352
rect 49016 188312 426532 188340
rect 49016 188300 49022 188312
rect 426526 188300 426532 188312
rect 426584 188300 426590 188352
rect 384298 188164 384304 188216
rect 384356 188204 384362 188216
rect 389082 188204 389088 188216
rect 384356 188176 389088 188204
rect 384356 188164 384362 188176
rect 389082 188164 389088 188176
rect 389140 188164 389146 188216
rect 249334 187620 249340 187672
rect 249392 187660 249398 187672
rect 378226 187660 378232 187672
rect 249392 187632 378232 187660
rect 249392 187620 249398 187632
rect 378226 187620 378232 187632
rect 378284 187620 378290 187672
rect 187510 187552 187516 187604
rect 187568 187592 187574 187604
rect 353754 187592 353760 187604
rect 187568 187564 353760 187592
rect 187568 187552 187574 187564
rect 353754 187552 353760 187564
rect 353812 187552 353818 187604
rect 59078 187484 59084 187536
rect 59136 187524 59142 187536
rect 359274 187524 359280 187536
rect 59136 187496 359280 187524
rect 59136 187484 59142 187496
rect 359274 187484 359280 187496
rect 359332 187484 359338 187536
rect 58986 187416 58992 187468
rect 59044 187456 59050 187468
rect 362034 187456 362040 187468
rect 59044 187428 362040 187456
rect 59044 187416 59050 187428
rect 362034 187416 362040 187428
rect 362092 187416 362098 187468
rect 56410 187348 56416 187400
rect 56468 187388 56474 187400
rect 361942 187388 361948 187400
rect 56468 187360 361948 187388
rect 56468 187348 56474 187360
rect 361942 187348 361948 187360
rect 362000 187348 362006 187400
rect 40586 187280 40592 187332
rect 40644 187320 40650 187332
rect 376662 187320 376668 187332
rect 40644 187292 376668 187320
rect 40644 187280 40650 187292
rect 376662 187280 376668 187292
rect 376720 187280 376726 187332
rect 42426 187212 42432 187264
rect 42484 187252 42490 187264
rect 387334 187252 387340 187264
rect 42484 187224 387340 187252
rect 42484 187212 42490 187224
rect 387334 187212 387340 187224
rect 387392 187212 387398 187264
rect 44910 187144 44916 187196
rect 44968 187184 44974 187196
rect 409966 187184 409972 187196
rect 44968 187156 409972 187184
rect 44968 187144 44974 187156
rect 409966 187144 409972 187156
rect 410024 187144 410030 187196
rect 53650 187076 53656 187128
rect 53708 187116 53714 187128
rect 470594 187116 470600 187128
rect 53708 187088 470600 187116
rect 53708 187076 53714 187088
rect 470594 187076 470600 187088
rect 470652 187076 470658 187128
rect 116026 187008 116032 187060
rect 116084 187048 116090 187060
rect 552382 187048 552388 187060
rect 116084 187020 552388 187048
rect 116084 187008 116090 187020
rect 552382 187008 552388 187020
rect 552440 187008 552446 187060
rect 85758 186940 85764 186992
rect 85816 186980 85822 186992
rect 550082 186980 550088 186992
rect 85816 186952 550088 186980
rect 85816 186940 85822 186952
rect 550082 186940 550088 186952
rect 550140 186940 550146 186992
rect 239030 186872 239036 186924
rect 239088 186912 239094 186924
rect 352466 186912 352472 186924
rect 239088 186884 352472 186912
rect 239088 186872 239094 186884
rect 352466 186872 352472 186884
rect 352524 186872 352530 186924
rect 264146 186804 264152 186856
rect 264204 186844 264210 186856
rect 350810 186844 350816 186856
rect 264204 186816 350816 186844
rect 264204 186804 264210 186816
rect 350810 186804 350816 186816
rect 350868 186804 350874 186856
rect 351086 186804 351092 186856
rect 351144 186844 351150 186856
rect 392854 186844 392860 186856
rect 351144 186816 392860 186844
rect 351144 186804 351150 186816
rect 392854 186804 392860 186816
rect 392912 186804 392918 186856
rect 300854 186736 300860 186788
rect 300912 186776 300918 186788
rect 348142 186776 348148 186788
rect 300912 186748 348148 186776
rect 300912 186736 300918 186748
rect 348142 186736 348148 186748
rect 348200 186736 348206 186788
rect 266078 185988 266084 186040
rect 266136 186028 266142 186040
rect 348050 186028 348056 186040
rect 266136 186000 348056 186028
rect 266136 185988 266142 186000
rect 348050 185988 348056 186000
rect 348108 185988 348114 186040
rect 246114 185920 246120 185972
rect 246172 185960 246178 185972
rect 353662 185960 353668 185972
rect 246172 185932 353668 185960
rect 246172 185920 246178 185932
rect 353662 185920 353668 185932
rect 353720 185920 353726 185972
rect 43714 185852 43720 185904
rect 43772 185892 43778 185904
rect 154298 185892 154304 185904
rect 43772 185864 154304 185892
rect 43772 185852 43778 185864
rect 154298 185852 154304 185864
rect 154356 185852 154362 185904
rect 209866 185852 209872 185904
rect 209924 185892 209930 185904
rect 356238 185892 356244 185904
rect 209924 185864 356244 185892
rect 209924 185852 209930 185864
rect 356238 185852 356244 185864
rect 356296 185852 356302 185904
rect 52086 185784 52092 185836
rect 52144 185824 52150 185836
rect 356606 185824 356612 185836
rect 52144 185796 356612 185824
rect 52144 185784 52150 185796
rect 356606 185784 356612 185796
rect 356664 185784 356670 185836
rect 43530 185716 43536 185768
rect 43588 185756 43594 185768
rect 260834 185756 260840 185768
rect 43588 185728 260840 185756
rect 43588 185716 43594 185728
rect 260834 185716 260840 185728
rect 260892 185716 260898 185768
rect 268654 185716 268660 185768
rect 268712 185756 268718 185768
rect 580074 185756 580080 185768
rect 268712 185728 580080 185756
rect 268712 185716 268718 185728
rect 580074 185716 580080 185728
rect 580132 185716 580138 185768
rect 48866 185648 48872 185700
rect 48924 185688 48930 185700
rect 384574 185688 384580 185700
rect 48924 185660 384580 185688
rect 48924 185648 48930 185660
rect 384574 185648 384580 185660
rect 384632 185648 384638 185700
rect 46014 185580 46020 185632
rect 46072 185620 46078 185632
rect 581178 185620 581184 185632
rect 46072 185592 581184 185620
rect 46072 185580 46078 185592
rect 581178 185580 581184 185592
rect 581236 185580 581242 185632
rect 176654 184628 176660 184680
rect 176712 184668 176718 184680
rect 293954 184668 293960 184680
rect 176712 184640 293960 184668
rect 176712 184628 176718 184640
rect 293954 184628 293960 184640
rect 294012 184628 294018 184680
rect 318242 184628 318248 184680
rect 318300 184668 318306 184680
rect 328822 184668 328828 184680
rect 318300 184640 328828 184668
rect 318300 184628 318306 184640
rect 328822 184628 328828 184640
rect 328880 184628 328886 184680
rect 271874 184560 271880 184612
rect 271932 184600 271938 184612
rect 393038 184600 393044 184612
rect 271932 184572 393044 184600
rect 271932 184560 271938 184572
rect 393038 184560 393044 184572
rect 393096 184560 393102 184612
rect 33778 184492 33784 184544
rect 33836 184532 33842 184544
rect 135254 184532 135260 184544
rect 33836 184504 135260 184532
rect 33836 184492 33842 184504
rect 135254 184492 135260 184504
rect 135312 184492 135318 184544
rect 137278 184492 137284 184544
rect 137336 184532 137342 184544
rect 360286 184532 360292 184544
rect 137336 184504 360292 184532
rect 137336 184492 137342 184504
rect 360286 184492 360292 184504
rect 360344 184492 360350 184544
rect 58802 184424 58808 184476
rect 58860 184464 58866 184476
rect 349614 184464 349620 184476
rect 58860 184436 349620 184464
rect 58860 184424 58866 184436
rect 349614 184424 349620 184436
rect 349672 184424 349678 184476
rect 59446 184356 59452 184408
rect 59504 184396 59510 184408
rect 362954 184396 362960 184408
rect 59504 184368 362960 184396
rect 59504 184356 59510 184368
rect 362954 184356 362960 184368
rect 363012 184356 363018 184408
rect 59722 184288 59728 184340
rect 59780 184328 59786 184340
rect 370130 184328 370136 184340
rect 59780 184300 370136 184328
rect 59780 184288 59786 184300
rect 370130 184288 370136 184300
rect 370188 184288 370194 184340
rect 38102 184220 38108 184272
rect 38160 184260 38166 184272
rect 364518 184260 364524 184272
rect 38160 184232 364524 184260
rect 38160 184220 38166 184232
rect 364518 184220 364524 184232
rect 364576 184220 364582 184272
rect 38194 184152 38200 184204
rect 38252 184192 38258 184204
rect 367278 184192 367284 184204
rect 38252 184164 367284 184192
rect 38252 184152 38258 184164
rect 367278 184152 367284 184164
rect 367336 184152 367342 184204
rect 442994 184152 443000 184204
rect 443052 184192 443058 184204
rect 508222 184192 508228 184204
rect 443052 184164 508228 184192
rect 443052 184152 443058 184164
rect 508222 184152 508228 184164
rect 508280 184152 508286 184204
rect 108298 183540 108304 183592
rect 108356 183580 108362 183592
rect 382274 183580 382280 183592
rect 108356 183552 382280 183580
rect 108356 183540 108362 183552
rect 382274 183540 382280 183552
rect 382332 183540 382338 183592
rect 199746 183132 199752 183184
rect 199804 183172 199810 183184
rect 372062 183172 372068 183184
rect 199804 183144 372068 183172
rect 199804 183132 199810 183144
rect 372062 183132 372068 183144
rect 372120 183132 372126 183184
rect 40402 183064 40408 183116
rect 40460 183104 40466 183116
rect 220354 183104 220360 183116
rect 40460 183076 220360 183104
rect 40460 183064 40466 183076
rect 220354 183064 220360 183076
rect 220412 183064 220418 183116
rect 293126 183064 293132 183116
rect 293184 183104 293190 183116
rect 351270 183104 351276 183116
rect 293184 183076 351276 183104
rect 293184 183064 293190 183076
rect 351270 183064 351276 183076
rect 351328 183064 351334 183116
rect 46566 182996 46572 183048
rect 46624 183036 46630 183048
rect 369578 183036 369584 183048
rect 46624 183008 369584 183036
rect 46624 182996 46630 183008
rect 369578 182996 369584 183008
rect 369636 182996 369642 183048
rect 43530 182928 43536 182980
rect 43588 182968 43594 182980
rect 384850 182968 384856 182980
rect 43588 182940 384856 182968
rect 43588 182928 43594 182940
rect 384850 182928 384856 182940
rect 384908 182928 384914 182980
rect 80238 182860 80244 182912
rect 80296 182900 80302 182912
rect 550726 182900 550732 182912
rect 80296 182872 550732 182900
rect 80296 182860 80302 182872
rect 550726 182860 550732 182872
rect 550784 182860 550790 182912
rect 44818 182792 44824 182844
rect 44876 182832 44882 182844
rect 519814 182832 519820 182844
rect 44876 182804 519820 182832
rect 44876 182792 44882 182804
rect 519814 182792 519820 182804
rect 519872 182792 519878 182844
rect 284754 181976 284760 182028
rect 284812 182016 284818 182028
rect 364426 182016 364432 182028
rect 284812 181988 364432 182016
rect 284812 181976 284818 181988
rect 364426 181976 364432 181988
rect 364484 181976 364490 182028
rect 170766 181908 170772 181960
rect 170824 181948 170830 181960
rect 355502 181948 355508 181960
rect 170824 181920 355508 181948
rect 170824 181908 170830 181920
rect 355502 181908 355508 181920
rect 355560 181908 355566 181960
rect 33042 181840 33048 181892
rect 33100 181880 33106 181892
rect 353846 181880 353852 181892
rect 33100 181852 353852 181880
rect 33100 181840 33106 181852
rect 353846 181840 353852 181852
rect 353904 181840 353910 181892
rect 31386 181772 31392 181824
rect 31444 181812 31450 181824
rect 367186 181812 367192 181824
rect 31444 181784 367192 181812
rect 31444 181772 31450 181784
rect 367186 181772 367192 181784
rect 367244 181772 367250 181824
rect 33778 181704 33784 181756
rect 33836 181744 33842 181756
rect 370038 181744 370044 181756
rect 33836 181716 370044 181744
rect 33836 181704 33842 181716
rect 370038 181704 370044 181716
rect 370096 181704 370102 181756
rect 31478 181636 31484 181688
rect 31536 181676 31542 181688
rect 375006 181676 375012 181688
rect 31536 181648 375012 181676
rect 31536 181636 31542 181648
rect 375006 181636 375012 181648
rect 375064 181636 375070 181688
rect 34422 181568 34428 181620
rect 34480 181608 34486 181620
rect 380526 181608 380532 181620
rect 34480 181580 380532 181608
rect 34480 181568 34486 181580
rect 380526 181568 380532 181580
rect 380584 181568 380590 181620
rect 35250 181500 35256 181552
rect 35308 181540 35314 181552
rect 392946 181540 392952 181552
rect 35308 181512 392952 181540
rect 35308 181500 35314 181512
rect 392946 181500 392952 181512
rect 393004 181500 393010 181552
rect 174630 181432 174636 181484
rect 174688 181472 174694 181484
rect 581638 181472 581644 181484
rect 174688 181444 581644 181472
rect 174688 181432 174694 181444
rect 581638 181432 581644 181444
rect 581696 181432 581702 181484
rect 225506 180480 225512 180532
rect 225564 180520 225570 180532
rect 364058 180520 364064 180532
rect 225564 180492 364064 180520
rect 225564 180480 225570 180492
rect 364058 180480 364064 180492
rect 364116 180480 364122 180532
rect 217778 180412 217784 180464
rect 217836 180452 217842 180464
rect 372614 180452 372620 180464
rect 217836 180424 372620 180452
rect 217836 180412 217842 180424
rect 372614 180412 372620 180424
rect 372672 180412 372678 180464
rect 40494 180344 40500 180396
rect 40552 180384 40558 180396
rect 235166 180384 235172 180396
rect 40552 180356 235172 180384
rect 40552 180344 40558 180356
rect 235166 180344 235172 180356
rect 235224 180344 235230 180396
rect 99926 180276 99932 180328
rect 99984 180316 99990 180328
rect 373534 180316 373540 180328
rect 99984 180288 373540 180316
rect 99984 180276 99990 180288
rect 373534 180276 373540 180288
rect 373592 180276 373598 180328
rect 46106 180208 46112 180260
rect 46164 180248 46170 180260
rect 340874 180248 340880 180260
rect 46164 180220 340880 180248
rect 46164 180208 46170 180220
rect 340874 180208 340880 180220
rect 340932 180208 340938 180260
rect 53374 180140 53380 180192
rect 53432 180180 53438 180192
rect 369210 180180 369216 180192
rect 53432 180152 369216 180180
rect 53432 180140 53438 180152
rect 369210 180140 369216 180152
rect 369268 180140 369274 180192
rect 150526 180072 150532 180124
rect 150584 180112 150590 180124
rect 538950 180112 538956 180124
rect 150584 180084 538956 180112
rect 150584 180072 150590 180084
rect 538950 180072 538956 180084
rect 539008 180072 539014 180124
rect 301038 179324 301044 179376
rect 301096 179364 301102 179376
rect 468294 179364 468300 179376
rect 301096 179336 468300 179364
rect 301096 179324 301102 179336
rect 468294 179324 468300 179336
rect 468352 179324 468358 179376
rect 577498 179324 577504 179376
rect 577556 179364 577562 179376
rect 580074 179364 580080 179376
rect 577556 179336 580080 179364
rect 577556 179324 577562 179336
rect 580074 179324 580080 179336
rect 580132 179324 580138 179376
rect 66438 179256 66444 179308
rect 66496 179296 66502 179308
rect 348326 179296 348332 179308
rect 66496 179268 348332 179296
rect 66496 179256 66502 179268
rect 348326 179256 348332 179268
rect 348384 179256 348390 179308
rect 40862 179188 40868 179240
rect 40920 179228 40926 179240
rect 329190 179228 329196 179240
rect 40920 179200 329196 179228
rect 40920 179188 40926 179200
rect 329190 179188 329196 179200
rect 329248 179188 329254 179240
rect 55582 179120 55588 179172
rect 55640 179160 55646 179172
rect 347038 179160 347044 179172
rect 55640 179132 347044 179160
rect 55640 179120 55646 179132
rect 347038 179120 347044 179132
rect 347096 179120 347102 179172
rect 38654 179052 38660 179104
rect 38712 179092 38718 179104
rect 361206 179092 361212 179104
rect 38712 179064 361212 179092
rect 38712 179052 38718 179064
rect 361206 179052 361212 179064
rect 361264 179052 361270 179104
rect 42334 178984 42340 179036
rect 42392 179024 42398 179036
rect 368014 179024 368020 179036
rect 42392 178996 368020 179024
rect 42392 178984 42398 178996
rect 368014 178984 368020 178996
rect 368072 178984 368078 179036
rect 69658 178916 69664 178968
rect 69716 178956 69722 178968
rect 197354 178956 197360 178968
rect 69716 178928 197360 178956
rect 69716 178916 69722 178928
rect 197354 178916 197360 178928
rect 197412 178916 197418 178968
rect 234522 178916 234528 178968
rect 234580 178956 234586 178968
rect 560478 178956 560484 178968
rect 234580 178928 560484 178956
rect 234580 178916 234586 178928
rect 560478 178916 560484 178928
rect 560536 178916 560542 178968
rect 57606 178848 57612 178900
rect 57664 178888 57670 178900
rect 391474 178888 391480 178900
rect 57664 178860 391480 178888
rect 57664 178848 57670 178860
rect 391474 178848 391480 178860
rect 391532 178848 391538 178900
rect 54754 178780 54760 178832
rect 54812 178820 54818 178832
rect 392486 178820 392492 178832
rect 54812 178792 392492 178820
rect 54812 178780 54818 178792
rect 392486 178780 392492 178792
rect 392544 178780 392550 178832
rect 45002 178712 45008 178764
rect 45060 178752 45066 178764
rect 389910 178752 389916 178764
rect 45060 178724 389916 178752
rect 45060 178712 45066 178724
rect 389910 178712 389916 178724
rect 389968 178712 389974 178764
rect 166258 178644 166264 178696
rect 166316 178684 166322 178696
rect 552566 178684 552572 178696
rect 166316 178656 552572 178684
rect 166316 178644 166322 178656
rect 552566 178644 552572 178656
rect 552624 178644 552630 178696
rect 41046 178440 41052 178492
rect 41104 178480 41110 178492
rect 45554 178480 45560 178492
rect 41104 178452 45560 178480
rect 41104 178440 41110 178452
rect 45554 178440 45560 178452
rect 45612 178440 45618 178492
rect 285674 177828 285680 177880
rect 285732 177868 285738 177880
rect 364150 177868 364156 177880
rect 285732 177840 364156 177868
rect 285732 177828 285738 177840
rect 364150 177828 364156 177840
rect 364208 177828 364214 177880
rect 211982 177760 211988 177812
rect 212040 177800 212046 177812
rect 352098 177800 352104 177812
rect 212040 177772 352104 177800
rect 212040 177760 212046 177772
rect 352098 177760 352104 177772
rect 352156 177760 352162 177812
rect 119890 177692 119896 177744
rect 119948 177732 119954 177744
rect 358998 177732 359004 177744
rect 119948 177704 359004 177732
rect 119948 177692 119954 177704
rect 358998 177692 359004 177704
rect 359056 177692 359062 177744
rect 98638 177624 98644 177676
rect 98696 177664 98702 177676
rect 350994 177664 351000 177676
rect 98696 177636 351000 177664
rect 98696 177624 98702 177636
rect 350994 177624 351000 177636
rect 351052 177624 351058 177676
rect 56134 177556 56140 177608
rect 56192 177596 56198 177608
rect 349246 177596 349252 177608
rect 56192 177568 349252 177596
rect 56192 177556 56198 177568
rect 349246 177556 349252 177568
rect 349304 177556 349310 177608
rect 41138 177488 41144 177540
rect 41196 177528 41202 177540
rect 395246 177528 395252 177540
rect 41196 177500 395252 177528
rect 41196 177488 41202 177500
rect 395246 177488 395252 177500
rect 395304 177488 395310 177540
rect 34330 177420 34336 177472
rect 34388 177460 34394 177472
rect 401962 177460 401968 177472
rect 34388 177432 401968 177460
rect 34388 177420 34394 177432
rect 401962 177420 401968 177432
rect 402020 177420 402026 177472
rect 431218 177420 431224 177472
rect 431276 177460 431282 177472
rect 514018 177460 514024 177472
rect 431276 177432 514024 177460
rect 431276 177420 431282 177432
rect 514018 177420 514024 177432
rect 514076 177420 514082 177472
rect 77386 177352 77392 177404
rect 77444 177392 77450 177404
rect 539962 177392 539968 177404
rect 77444 177364 539968 177392
rect 77444 177352 77450 177364
rect 539962 177352 539968 177364
rect 540020 177352 540026 177404
rect 46198 177284 46204 177336
rect 46256 177324 46262 177336
rect 552290 177324 552296 177336
rect 46256 177296 552296 177324
rect 46256 177284 46262 177296
rect 552290 177284 552296 177296
rect 552348 177284 552354 177336
rect 44818 176604 44824 176656
rect 44876 176644 44882 176656
rect 45830 176644 45836 176656
rect 44876 176616 45836 176644
rect 44876 176604 44882 176616
rect 45830 176604 45836 176616
rect 45888 176604 45894 176656
rect 312446 176468 312452 176520
rect 312504 176508 312510 176520
rect 375374 176508 375380 176520
rect 312504 176480 375380 176508
rect 312504 176468 312510 176480
rect 375374 176468 375380 176480
rect 375432 176468 375438 176520
rect 188154 176400 188160 176452
rect 188212 176440 188218 176452
rect 381906 176440 381912 176452
rect 188212 176412 381912 176440
rect 188212 176400 188218 176412
rect 381906 176400 381912 176412
rect 381964 176400 381970 176452
rect 43438 176332 43444 176384
rect 43496 176372 43502 176384
rect 314378 176372 314384 176384
rect 43496 176344 314384 176372
rect 43496 176332 43502 176344
rect 314378 176332 314384 176344
rect 314436 176332 314442 176384
rect 53558 176264 53564 176316
rect 53616 176304 53622 176316
rect 386230 176304 386236 176316
rect 53616 176276 386236 176304
rect 53616 176264 53622 176276
rect 386230 176264 386236 176276
rect 386288 176264 386294 176316
rect 37182 176196 37188 176248
rect 37240 176236 37246 176248
rect 374822 176236 374828 176248
rect 37240 176208 374828 176236
rect 37240 176196 37246 176208
rect 374822 176196 374828 176208
rect 374880 176196 374886 176248
rect 41966 176128 41972 176180
rect 42024 176168 42030 176180
rect 385862 176168 385868 176180
rect 42024 176140 385868 176168
rect 42024 176128 42030 176140
rect 385862 176128 385868 176140
rect 385920 176128 385926 176180
rect 95234 176060 95240 176112
rect 95292 176100 95298 176112
rect 443178 176100 443184 176112
rect 95292 176072 443184 176100
rect 95292 176060 95298 176072
rect 443178 176060 443184 176072
rect 443236 176060 443242 176112
rect 40954 175992 40960 176044
rect 41012 176032 41018 176044
rect 389726 176032 389732 176044
rect 41012 176004 389732 176032
rect 41012 175992 41018 176004
rect 389726 175992 389732 176004
rect 389784 175992 389790 176044
rect 88334 175924 88340 175976
rect 88392 175964 88398 175976
rect 480530 175964 480536 175976
rect 88392 175936 480536 175964
rect 88392 175924 88398 175936
rect 480530 175924 480536 175936
rect 480588 175924 480594 175976
rect 254486 174904 254492 174956
rect 254544 174944 254550 174956
rect 377674 174944 377680 174956
rect 254544 174916 377680 174944
rect 254544 174904 254550 174916
rect 377674 174904 377680 174916
rect 377732 174904 377738 174956
rect 180794 174836 180800 174888
rect 180852 174876 180858 174888
rect 327074 174876 327080 174888
rect 180852 174848 327080 174876
rect 180852 174836 180858 174848
rect 327074 174836 327080 174848
rect 327132 174836 327138 174888
rect 205634 174768 205640 174820
rect 205692 174808 205698 174820
rect 384390 174808 384396 174820
rect 205692 174780 384396 174808
rect 205692 174768 205698 174780
rect 384390 174768 384396 174780
rect 384448 174768 384454 174820
rect 111978 174700 111984 174752
rect 112036 174740 112042 174752
rect 130194 174740 130200 174752
rect 112036 174712 130200 174740
rect 112036 174700 112042 174712
rect 130194 174700 130200 174712
rect 130252 174700 130258 174752
rect 318886 174700 318892 174752
rect 318944 174740 318950 174752
rect 562318 174740 562324 174752
rect 318944 174712 562324 174740
rect 318944 174700 318950 174712
rect 562318 174700 562324 174712
rect 562376 174700 562382 174752
rect 78030 174632 78036 174684
rect 78088 174672 78094 174684
rect 363966 174672 363972 174684
rect 78088 174644 363972 174672
rect 78088 174632 78094 174644
rect 363966 174632 363972 174644
rect 364024 174632 364030 174684
rect 46290 174564 46296 174616
rect 46348 174604 46354 174616
rect 364610 174604 364616 174616
rect 46348 174576 364616 174604
rect 46348 174564 46354 174576
rect 364610 174564 364616 174576
rect 364668 174564 364674 174616
rect 47946 174496 47952 174548
rect 48004 174536 48010 174548
rect 380894 174536 380900 174548
rect 48004 174508 380900 174536
rect 48004 174496 48010 174508
rect 380894 174496 380900 174508
rect 380952 174496 380958 174548
rect 568022 173816 568028 173868
rect 568080 173856 568086 173868
rect 570414 173856 570420 173868
rect 568080 173828 570420 173856
rect 568080 173816 568086 173828
rect 570414 173816 570420 173828
rect 570472 173816 570478 173868
rect 306466 173476 306472 173528
rect 306524 173516 306530 173528
rect 387058 173516 387064 173528
rect 306524 173488 387064 173516
rect 306524 173476 306530 173488
rect 387058 173476 387064 173488
rect 387116 173476 387122 173528
rect 241606 173408 241612 173460
rect 241664 173448 241670 173460
rect 347866 173448 347872 173460
rect 241664 173420 347872 173448
rect 241664 173408 241670 173420
rect 347866 173408 347872 173420
rect 347924 173408 347930 173460
rect 207474 173340 207480 173392
rect 207532 173380 207538 173392
rect 373258 173380 373264 173392
rect 207532 173352 373264 173380
rect 207532 173340 207538 173352
rect 373258 173340 373264 173352
rect 373316 173340 373322 173392
rect 38010 173272 38016 173324
rect 38068 173312 38074 173324
rect 175918 173312 175924 173324
rect 38068 173284 175924 173312
rect 38068 173272 38074 173284
rect 175918 173272 175924 173284
rect 175976 173272 175982 173324
rect 237374 173272 237380 173324
rect 237432 173312 237438 173324
rect 506934 173312 506940 173324
rect 237432 173284 506940 173312
rect 237432 173272 237438 173284
rect 506934 173272 506940 173284
rect 506992 173272 506998 173324
rect 79318 173204 79324 173256
rect 79376 173244 79382 173256
rect 355042 173244 355048 173256
rect 79376 173216 355048 173244
rect 79376 173204 79382 173216
rect 355042 173204 355048 173216
rect 355100 173204 355106 173256
rect 46474 173136 46480 173188
rect 46532 173176 46538 173188
rect 495434 173176 495440 173188
rect 46532 173148 495440 173176
rect 46532 173136 46538 173148
rect 495434 173136 495440 173148
rect 495492 173136 495498 173188
rect 96706 172320 96712 172372
rect 96764 172360 96770 172372
rect 242250 172360 242256 172372
rect 96764 172332 242256 172360
rect 96764 172320 96770 172332
rect 242250 172320 242256 172332
rect 242308 172320 242314 172372
rect 35158 172252 35164 172304
rect 35216 172292 35222 172304
rect 193214 172292 193220 172304
rect 35216 172264 193220 172292
rect 35216 172252 35222 172264
rect 193214 172252 193220 172264
rect 193272 172252 193278 172304
rect 283466 172252 283472 172304
rect 283524 172292 283530 172304
rect 368474 172292 368480 172304
rect 283524 172264 368480 172292
rect 283524 172252 283530 172264
rect 368474 172252 368480 172264
rect 368532 172252 368538 172304
rect 163038 172184 163044 172236
rect 163096 172224 163102 172236
rect 349706 172224 349712 172236
rect 163096 172196 349712 172224
rect 163096 172184 163102 172196
rect 349706 172184 349712 172196
rect 349764 172184 349770 172236
rect 146938 172116 146944 172168
rect 146996 172156 147002 172168
rect 351178 172156 351184 172168
rect 146996 172128 351184 172156
rect 146996 172116 147002 172128
rect 351178 172116 351184 172128
rect 351236 172116 351242 172168
rect 50522 172048 50528 172100
rect 50580 172088 50586 172100
rect 360470 172088 360476 172100
rect 50580 172060 360476 172088
rect 50580 172048 50586 172060
rect 360470 172048 360476 172060
rect 360528 172048 360534 172100
rect 46658 171980 46664 172032
rect 46716 172020 46722 172032
rect 359366 172020 359372 172032
rect 46716 171992 359372 172020
rect 46716 171980 46722 171992
rect 359366 171980 359372 171992
rect 359424 171980 359430 172032
rect 47762 171912 47768 171964
rect 47820 171952 47826 171964
rect 379606 171952 379612 171964
rect 47820 171924 379612 171952
rect 47820 171912 47826 171924
rect 379606 171912 379612 171924
rect 379664 171912 379670 171964
rect 43898 171844 43904 171896
rect 43956 171884 43962 171896
rect 379238 171884 379244 171896
rect 43956 171856 379244 171884
rect 43956 171844 43962 171856
rect 379238 171844 379244 171856
rect 379296 171844 379302 171896
rect 77386 171776 77392 171828
rect 77444 171816 77450 171828
rect 563514 171816 563520 171828
rect 77444 171788 563520 171816
rect 77444 171776 77450 171788
rect 563514 171776 563520 171788
rect 563572 171776 563578 171828
rect 259638 170756 259644 170808
rect 259696 170796 259702 170808
rect 309134 170796 309140 170808
rect 259696 170768 309140 170796
rect 259696 170756 259702 170768
rect 309134 170756 309140 170768
rect 309192 170756 309198 170808
rect 313734 170756 313740 170808
rect 313792 170796 313798 170808
rect 373902 170796 373908 170808
rect 313792 170768 373908 170796
rect 313792 170756 313798 170768
rect 373902 170756 373908 170768
rect 373960 170756 373966 170808
rect 195238 170688 195244 170740
rect 195296 170728 195302 170740
rect 352742 170728 352748 170740
rect 195296 170700 352748 170728
rect 195296 170688 195302 170700
rect 352742 170688 352748 170700
rect 352800 170688 352806 170740
rect 37918 170620 37924 170672
rect 37976 170660 37982 170672
rect 245470 170660 245476 170672
rect 37976 170632 245476 170660
rect 37976 170620 37982 170632
rect 245470 170620 245476 170632
rect 245528 170620 245534 170672
rect 279602 170620 279608 170672
rect 279660 170660 279666 170672
rect 356422 170660 356428 170672
rect 279660 170632 356428 170660
rect 279660 170620 279666 170632
rect 356422 170620 356428 170632
rect 356480 170620 356486 170672
rect 103790 170552 103796 170604
rect 103848 170592 103854 170604
rect 350718 170592 350724 170604
rect 103848 170564 350724 170592
rect 103848 170552 103854 170564
rect 350718 170552 350724 170564
rect 350776 170552 350782 170604
rect 369394 170552 369400 170604
rect 369452 170592 369458 170604
rect 400766 170592 400772 170604
rect 369452 170564 400772 170592
rect 369452 170552 369458 170564
rect 400766 170552 400772 170564
rect 400824 170552 400830 170604
rect 124398 170484 124404 170536
rect 124456 170524 124462 170536
rect 374086 170524 374092 170536
rect 124456 170496 374092 170524
rect 124456 170484 124462 170496
rect 374086 170484 374092 170496
rect 374144 170484 374150 170536
rect 84194 170416 84200 170468
rect 84252 170456 84258 170468
rect 371418 170456 371424 170468
rect 84252 170428 371424 170456
rect 84252 170416 84258 170428
rect 371418 170416 371424 170428
rect 371476 170416 371482 170468
rect 13814 170348 13820 170400
rect 13872 170388 13878 170400
rect 432046 170388 432052 170400
rect 13872 170360 432052 170388
rect 13872 170348 13878 170360
rect 432046 170348 432052 170360
rect 432104 170348 432110 170400
rect 462314 170348 462320 170400
rect 462372 170388 462378 170400
rect 552750 170388 552756 170400
rect 462372 170360 552756 170388
rect 462372 170348 462378 170360
rect 552750 170348 552756 170360
rect 552808 170348 552814 170400
rect 321462 169260 321468 169312
rect 321520 169300 321526 169312
rect 398098 169300 398104 169312
rect 321520 169272 398104 169300
rect 321520 169260 321526 169272
rect 398098 169260 398104 169272
rect 398156 169260 398162 169312
rect 354306 169192 354312 169244
rect 354364 169232 354370 169244
rect 467834 169232 467840 169244
rect 354364 169204 467840 169232
rect 354364 169192 354370 169204
rect 467834 169192 467840 169204
rect 467892 169192 467898 169244
rect 191834 169124 191840 169176
rect 191892 169164 191898 169176
rect 274450 169164 274456 169176
rect 191892 169136 274456 169164
rect 191892 169124 191898 169136
rect 274450 169124 274456 169136
rect 274508 169124 274514 169176
rect 292574 169124 292580 169176
rect 292632 169164 292638 169176
rect 439314 169164 439320 169176
rect 292632 169136 439320 169164
rect 292632 169124 292638 169136
rect 439314 169124 439320 169136
rect 439372 169124 439378 169176
rect 113174 169056 113180 169108
rect 113232 169096 113238 169108
rect 372430 169096 372436 169108
rect 113232 169068 372436 169096
rect 113232 169056 113238 169068
rect 372430 169056 372436 169068
rect 372488 169056 372494 169108
rect 397914 169056 397920 169108
rect 397972 169096 397978 169108
rect 407298 169096 407304 169108
rect 397972 169068 407304 169096
rect 397972 169056 397978 169068
rect 407298 169056 407304 169068
rect 407356 169056 407362 169108
rect 49694 168988 49700 169040
rect 49752 169028 49758 169040
rect 528830 169028 528836 169040
rect 49752 169000 528836 169028
rect 49752 168988 49758 169000
rect 528830 168988 528836 169000
rect 528888 168988 528894 169040
rect 271966 168104 271972 168156
rect 272024 168144 272030 168156
rect 309870 168144 309876 168156
rect 272024 168116 309876 168144
rect 272024 168104 272030 168116
rect 309870 168104 309876 168116
rect 309928 168104 309934 168156
rect 214006 168036 214012 168088
rect 214064 168076 214070 168088
rect 346578 168076 346584 168088
rect 214064 168048 346584 168076
rect 214064 168036 214070 168048
rect 346578 168036 346584 168048
rect 346636 168036 346642 168088
rect 228726 167968 228732 168020
rect 228784 168008 228790 168020
rect 378870 168008 378876 168020
rect 228784 167980 378876 168008
rect 228784 167968 228790 167980
rect 378870 167968 378876 167980
rect 378928 167968 378934 168020
rect 107746 167900 107752 167952
rect 107804 167940 107810 167952
rect 161750 167940 161756 167952
rect 107804 167912 161756 167940
rect 107804 167900 107810 167912
rect 161750 167900 161756 167912
rect 161808 167900 161814 167952
rect 250622 167900 250628 167952
rect 250680 167940 250686 167952
rect 547414 167940 547420 167952
rect 250680 167912 547420 167940
rect 250680 167900 250686 167912
rect 547414 167900 547420 167912
rect 547472 167900 547478 167952
rect 57514 167832 57520 167884
rect 57572 167872 57578 167884
rect 376570 167872 376576 167884
rect 57572 167844 376576 167872
rect 57572 167832 57578 167844
rect 376570 167832 376576 167844
rect 376628 167832 376634 167884
rect 407114 167832 407120 167884
rect 407172 167872 407178 167884
rect 438854 167872 438860 167884
rect 407172 167844 438860 167872
rect 407172 167832 407178 167844
rect 438854 167832 438860 167844
rect 438912 167832 438918 167884
rect 55950 167764 55956 167816
rect 56008 167804 56014 167816
rect 407850 167804 407856 167816
rect 56008 167776 407856 167804
rect 56008 167764 56014 167776
rect 407850 167764 407856 167776
rect 407908 167764 407914 167816
rect 145006 167696 145012 167748
rect 145064 167736 145070 167748
rect 552842 167736 552848 167748
rect 145064 167708 552848 167736
rect 145064 167696 145070 167708
rect 552842 167696 552848 167708
rect 552900 167696 552906 167748
rect 55030 167628 55036 167680
rect 55088 167668 55094 167680
rect 544470 167668 544476 167680
rect 55088 167640 544476 167668
rect 55088 167628 55094 167640
rect 544470 167628 544476 167640
rect 544528 167628 544534 167680
rect 41230 166540 41236 166592
rect 41288 166580 41294 166592
rect 77294 166580 77300 166592
rect 41288 166552 77300 166580
rect 41288 166540 41294 166552
rect 77294 166540 77300 166552
rect 77352 166540 77358 166592
rect 213270 166540 213276 166592
rect 213328 166580 213334 166592
rect 273254 166580 273260 166592
rect 213328 166552 273260 166580
rect 213328 166540 213334 166552
rect 273254 166540 273260 166552
rect 273312 166540 273318 166592
rect 278958 166540 278964 166592
rect 279016 166580 279022 166592
rect 366726 166580 366732 166592
rect 279016 166552 366732 166580
rect 279016 166540 279022 166552
rect 366726 166540 366732 166552
rect 366784 166540 366790 166592
rect 81894 166472 81900 166524
rect 81952 166512 81958 166524
rect 228358 166512 228364 166524
rect 81952 166484 228364 166512
rect 81952 166472 81958 166484
rect 228358 166472 228364 166484
rect 228416 166472 228422 166524
rect 233878 166472 233884 166524
rect 233936 166512 233942 166524
rect 385678 166512 385684 166524
rect 233936 166484 385684 166512
rect 233936 166472 233942 166484
rect 385678 166472 385684 166484
rect 385736 166472 385742 166524
rect 40770 166404 40776 166456
rect 40828 166444 40834 166456
rect 240134 166444 240140 166456
rect 40828 166416 240140 166444
rect 40828 166404 40834 166416
rect 240134 166404 240140 166416
rect 240192 166404 240198 166456
rect 271230 166404 271236 166456
rect 271288 166444 271294 166456
rect 402330 166444 402336 166456
rect 271288 166416 402336 166444
rect 271288 166404 271294 166416
rect 402330 166404 402336 166416
rect 402388 166404 402394 166456
rect 60826 166336 60832 166388
rect 60884 166376 60890 166388
rect 307938 166376 307944 166388
rect 60884 166348 307944 166376
rect 60884 166336 60890 166348
rect 307938 166336 307944 166348
rect 307996 166336 308002 166388
rect 342070 166336 342076 166388
rect 342128 166376 342134 166388
rect 347958 166376 347964 166388
rect 342128 166348 347964 166376
rect 342128 166336 342134 166348
rect 347958 166336 347964 166348
rect 348016 166336 348022 166388
rect 43346 166268 43352 166320
rect 43404 166308 43410 166320
rect 350442 166308 350448 166320
rect 43404 166280 350448 166308
rect 43404 166268 43410 166280
rect 350442 166268 350448 166280
rect 350500 166268 350506 166320
rect 251266 165180 251272 165232
rect 251324 165220 251330 165232
rect 402238 165220 402244 165232
rect 251324 165192 402244 165220
rect 251324 165180 251330 165192
rect 402238 165180 402244 165192
rect 402296 165180 402302 165232
rect 402698 165180 402704 165232
rect 402756 165220 402762 165232
rect 563422 165220 563428 165232
rect 402756 165192 563428 165220
rect 402756 165180 402762 165192
rect 563422 165180 563428 165192
rect 563480 165180 563486 165232
rect 142430 165112 142436 165164
rect 142488 165152 142494 165164
rect 361298 165152 361304 165164
rect 142488 165124 361304 165152
rect 142488 165112 142494 165124
rect 361298 165112 361304 165124
rect 361356 165112 361362 165164
rect 406562 165112 406568 165164
rect 406620 165152 406626 165164
rect 581638 165152 581644 165164
rect 406620 165124 581644 165152
rect 406620 165112 406626 165124
rect 581638 165112 581644 165124
rect 581696 165112 581702 165164
rect 328454 165044 328460 165096
rect 328512 165084 328518 165096
rect 560846 165084 560852 165096
rect 328512 165056 560852 165084
rect 328512 165044 328518 165056
rect 560846 165044 560852 165056
rect 560904 165044 560910 165096
rect 57422 164976 57428 165028
rect 57480 165016 57486 165028
rect 362310 165016 362316 165028
rect 57480 164988 362316 165016
rect 57480 164976 57486 164988
rect 362310 164976 362316 164988
rect 362368 164976 362374 165028
rect 377766 164976 377772 165028
rect 377824 165016 377830 165028
rect 574922 165016 574928 165028
rect 377824 164988 574928 165016
rect 377824 164976 377830 164988
rect 574922 164976 574928 164988
rect 574980 164976 574986 165028
rect 40678 164908 40684 164960
rect 40736 164948 40742 164960
rect 383930 164948 383936 164960
rect 40736 164920 383936 164948
rect 40736 164908 40742 164920
rect 383930 164908 383936 164920
rect 383988 164908 383994 164960
rect 391658 164908 391664 164960
rect 391716 164948 391722 164960
rect 581730 164948 581736 164960
rect 391716 164920 581736 164948
rect 391716 164908 391722 164920
rect 581730 164908 581736 164920
rect 581788 164908 581794 164960
rect 50154 164840 50160 164892
rect 50212 164880 50218 164892
rect 472158 164880 472164 164892
rect 50212 164852 472164 164880
rect 50212 164840 50218 164852
rect 472158 164840 472164 164852
rect 472216 164840 472222 164892
rect 277394 163752 277400 163804
rect 277452 163792 277458 163804
rect 371970 163792 371976 163804
rect 277452 163764 371976 163792
rect 277452 163752 277458 163764
rect 371970 163752 371976 163764
rect 372028 163752 372034 163804
rect 406286 163752 406292 163804
rect 406344 163792 406350 163804
rect 470226 163792 470232 163804
rect 406344 163764 470232 163792
rect 406344 163752 406350 163764
rect 470226 163752 470232 163764
rect 470284 163752 470290 163804
rect 200758 163684 200764 163736
rect 200816 163724 200822 163736
rect 369118 163724 369124 163736
rect 200816 163696 369124 163724
rect 200816 163684 200822 163696
rect 369118 163684 369124 163696
rect 369176 163684 369182 163736
rect 227714 163616 227720 163668
rect 227772 163656 227778 163668
rect 469214 163656 469220 163668
rect 227772 163628 469220 163656
rect 227772 163616 227778 163628
rect 469214 163616 469220 163628
rect 469272 163616 469278 163668
rect 42150 163548 42156 163600
rect 42208 163588 42214 163600
rect 345014 163588 345020 163600
rect 42208 163560 345020 163588
rect 42208 163548 42214 163560
rect 345014 163548 345020 163560
rect 345072 163548 345078 163600
rect 386966 163548 386972 163600
rect 387024 163588 387030 163600
rect 548334 163588 548340 163600
rect 387024 163560 548340 163588
rect 387024 163548 387030 163560
rect 548334 163548 548340 163560
rect 548392 163548 548398 163600
rect 224862 163480 224868 163532
rect 224920 163520 224926 163532
rect 563790 163520 563796 163532
rect 224920 163492 563796 163520
rect 224920 163480 224926 163492
rect 563790 163480 563796 163492
rect 563848 163480 563854 163532
rect 403342 162800 403348 162852
rect 403400 162840 403406 162852
rect 562318 162840 562324 162852
rect 403400 162812 562324 162840
rect 403400 162800 403406 162812
rect 562318 162800 562324 162812
rect 562376 162800 562382 162852
rect 392578 162732 392584 162784
rect 392636 162772 392642 162784
rect 550910 162772 550916 162784
rect 392636 162744 550916 162772
rect 392636 162732 392642 162744
rect 550910 162732 550916 162744
rect 550968 162732 550974 162784
rect 398558 162664 398564 162716
rect 398616 162704 398622 162716
rect 567286 162704 567292 162716
rect 398616 162676 567292 162704
rect 398616 162664 398622 162676
rect 567286 162664 567292 162676
rect 567344 162664 567350 162716
rect 406838 162596 406844 162648
rect 406896 162636 406902 162648
rect 582650 162636 582656 162648
rect 406896 162608 582656 162636
rect 406896 162596 406902 162608
rect 582650 162596 582656 162608
rect 582708 162596 582714 162648
rect 403710 162528 403716 162580
rect 403768 162568 403774 162580
rect 581178 162568 581184 162580
rect 403768 162540 581184 162568
rect 403768 162528 403774 162540
rect 581178 162528 581184 162540
rect 581236 162528 581242 162580
rect 358354 162460 358360 162512
rect 358412 162500 358418 162512
rect 537846 162500 537852 162512
rect 358412 162472 537852 162500
rect 358412 162460 358418 162472
rect 537846 162460 537852 162472
rect 537904 162460 537910 162512
rect 266354 162392 266360 162444
rect 266412 162432 266418 162444
rect 356238 162432 356244 162444
rect 266412 162404 356244 162432
rect 266412 162392 266418 162404
rect 356238 162392 356244 162404
rect 356296 162392 356302 162444
rect 392394 162392 392400 162444
rect 392452 162432 392458 162444
rect 580074 162432 580080 162444
rect 392452 162404 580080 162432
rect 392452 162392 392458 162404
rect 580074 162392 580080 162404
rect 580132 162392 580138 162444
rect 216490 162324 216496 162376
rect 216548 162364 216554 162376
rect 348694 162364 348700 162376
rect 216548 162336 348700 162364
rect 216548 162324 216554 162336
rect 348694 162324 348700 162336
rect 348752 162324 348758 162376
rect 377950 162324 377956 162376
rect 378008 162364 378014 162376
rect 574554 162364 574560 162376
rect 378008 162336 574560 162364
rect 378008 162324 378014 162336
rect 574554 162324 574560 162336
rect 574612 162324 574618 162376
rect 110874 162256 110880 162308
rect 110932 162296 110938 162308
rect 278774 162296 278780 162308
rect 110932 162268 278780 162296
rect 110932 162256 110938 162268
rect 278774 162256 278780 162268
rect 278832 162256 278838 162308
rect 282914 162256 282920 162308
rect 282972 162296 282978 162308
rect 549254 162296 549260 162308
rect 282972 162268 549260 162296
rect 282972 162256 282978 162268
rect 549254 162256 549260 162268
rect 549312 162256 549318 162308
rect 259546 162188 259552 162240
rect 259604 162228 259610 162240
rect 539042 162228 539048 162240
rect 259604 162200 539048 162228
rect 259604 162188 259610 162200
rect 539042 162188 539048 162200
rect 539100 162188 539106 162240
rect 25406 162120 25412 162172
rect 25464 162160 25470 162172
rect 568574 162160 568580 162172
rect 25464 162132 568580 162160
rect 25464 162120 25470 162132
rect 568574 162120 568580 162132
rect 568632 162120 568638 162172
rect 387518 162052 387524 162104
rect 387576 162092 387582 162104
rect 539226 162092 539232 162104
rect 387576 162064 539232 162092
rect 387576 162052 387582 162064
rect 539226 162052 539232 162064
rect 539284 162052 539290 162104
rect 410150 161984 410156 162036
rect 410208 162024 410214 162036
rect 539318 162024 539324 162036
rect 410208 161996 539324 162024
rect 410208 161984 410214 161996
rect 539318 161984 539324 161996
rect 539376 161984 539382 162036
rect 414658 161916 414664 161968
rect 414716 161956 414722 161968
rect 419994 161956 420000 161968
rect 414716 161928 420000 161956
rect 414716 161916 414722 161928
rect 419994 161916 420000 161928
rect 420052 161916 420058 161968
rect 328454 160964 328460 161016
rect 328512 161004 328518 161016
rect 391290 161004 391296 161016
rect 328512 160976 391296 161004
rect 328512 160964 328518 160976
rect 391290 160964 391296 160976
rect 391348 160964 391354 161016
rect 406378 160964 406384 161016
rect 406436 161004 406442 161016
rect 510154 161004 510160 161016
rect 406436 160976 510160 161004
rect 406436 160964 406442 160976
rect 510154 160964 510160 160976
rect 510212 160964 510218 161016
rect 320174 160896 320180 160948
rect 320232 160936 320238 160948
rect 578786 160936 578792 160948
rect 320232 160908 578792 160936
rect 320232 160896 320238 160908
rect 578786 160896 578792 160908
rect 578844 160896 578850 160948
rect 96706 160828 96712 160880
rect 96764 160868 96770 160880
rect 376018 160868 376024 160880
rect 96764 160840 376024 160868
rect 96764 160828 96770 160840
rect 376018 160828 376024 160840
rect 376076 160828 376082 160880
rect 378962 160828 378968 160880
rect 379020 160868 379026 160880
rect 549530 160868 549536 160880
rect 379020 160840 549536 160868
rect 379020 160828 379026 160840
rect 549530 160828 549536 160840
rect 549588 160828 549594 160880
rect 25958 160760 25964 160812
rect 26016 160800 26022 160812
rect 335630 160800 335636 160812
rect 26016 160772 335636 160800
rect 26016 160760 26022 160772
rect 335630 160760 335636 160772
rect 335688 160760 335694 160812
rect 380342 160760 380348 160812
rect 380400 160800 380406 160812
rect 552566 160800 552572 160812
rect 380400 160772 552572 160800
rect 380400 160760 380406 160772
rect 552566 160760 552572 160772
rect 552624 160760 552630 160812
rect 150434 160692 150440 160744
rect 150492 160732 150498 160744
rect 552382 160732 552388 160744
rect 150492 160704 552388 160732
rect 150492 160692 150498 160704
rect 552382 160692 552388 160704
rect 552440 160692 552446 160744
rect 408310 160012 408316 160064
rect 408368 160052 408374 160064
rect 559558 160052 559564 160064
rect 408368 160024 559564 160052
rect 408368 160012 408374 160024
rect 559558 160012 559564 160024
rect 559616 160012 559622 160064
rect 405182 159944 405188 159996
rect 405240 159984 405246 159996
rect 561030 159984 561036 159996
rect 405240 159956 561036 159984
rect 405240 159944 405246 159956
rect 561030 159944 561036 159956
rect 561088 159944 561094 159996
rect 386046 159876 386052 159928
rect 386104 159916 386110 159928
rect 545666 159916 545672 159928
rect 386104 159888 545672 159916
rect 386104 159876 386110 159888
rect 545666 159876 545672 159888
rect 545724 159876 545730 159928
rect 226794 159808 226800 159860
rect 226852 159848 226858 159860
rect 358170 159848 358176 159860
rect 226852 159820 358176 159848
rect 226852 159808 226858 159820
rect 358170 159808 358176 159820
rect 358228 159808 358234 159860
rect 374730 159808 374736 159860
rect 374788 159848 374794 159860
rect 536834 159848 536840 159860
rect 374788 159820 536840 159848
rect 374788 159808 374794 159820
rect 536834 159808 536840 159820
rect 536892 159808 536898 159860
rect 155310 159740 155316 159792
rect 155368 159780 155374 159792
rect 360930 159780 360936 159792
rect 155368 159752 360936 159780
rect 155368 159740 155374 159752
rect 360930 159740 360936 159752
rect 360988 159740 360994 159792
rect 373718 159740 373724 159792
rect 373776 159780 373782 159792
rect 546770 159780 546776 159792
rect 373776 159752 546776 159780
rect 373776 159740 373782 159752
rect 546770 159740 546776 159752
rect 546828 159740 546834 159792
rect 305086 159672 305092 159724
rect 305144 159712 305150 159724
rect 541066 159712 541072 159724
rect 305144 159684 541072 159712
rect 305144 159672 305150 159684
rect 541066 159672 541072 159684
rect 541124 159672 541130 159724
rect 201402 159604 201408 159656
rect 201460 159644 201466 159656
rect 454126 159644 454132 159656
rect 201460 159616 454132 159644
rect 201460 159604 201466 159616
rect 454126 159604 454132 159616
rect 454184 159604 454190 159656
rect 57330 159536 57336 159588
rect 57388 159576 57394 159588
rect 362494 159576 362500 159588
rect 57388 159548 362500 159576
rect 57388 159536 57394 159548
rect 362494 159536 362500 159548
rect 362552 159536 362558 159588
rect 372154 159536 372160 159588
rect 372212 159576 372218 159588
rect 562042 159576 562048 159588
rect 372212 159548 562048 159576
rect 372212 159536 372218 159548
rect 562042 159536 562048 159548
rect 562100 159536 562106 159588
rect 57698 159468 57704 159520
rect 57756 159508 57762 159520
rect 375190 159508 375196 159520
rect 57756 159480 375196 159508
rect 57756 159468 57762 159480
rect 375190 159468 375196 159480
rect 375248 159468 375254 159520
rect 409230 159468 409236 159520
rect 409288 159508 409294 159520
rect 571702 159508 571708 159520
rect 409288 159480 571708 159508
rect 409288 159468 409294 159480
rect 571702 159468 571708 159480
rect 571760 159468 571766 159520
rect 54938 159400 54944 159452
rect 54996 159440 55002 159452
rect 483106 159440 483112 159452
rect 54996 159412 483112 159440
rect 54996 159400 55002 159412
rect 483106 159400 483112 159412
rect 483164 159400 483170 159452
rect 31018 159332 31024 159384
rect 31076 159372 31082 159384
rect 559466 159372 559472 159384
rect 31076 159344 559472 159372
rect 31076 159332 31082 159344
rect 559466 159332 559472 159344
rect 559524 159332 559530 159384
rect 408218 159264 408224 159316
rect 408276 159304 408282 159316
rect 558270 159304 558276 159316
rect 408276 159276 558276 159304
rect 408276 159264 408282 159276
rect 558270 159264 558276 159276
rect 558328 159264 558334 159316
rect 282822 159196 282828 159248
rect 282880 159236 282886 159248
rect 426434 159236 426440 159248
rect 282880 159208 426440 159236
rect 282880 159196 282886 159208
rect 426434 159196 426440 159208
rect 426492 159196 426498 159248
rect 405090 159128 405096 159180
rect 405148 159168 405154 159180
rect 542906 159168 542912 159180
rect 405148 159140 542912 159168
rect 405148 159128 405154 159140
rect 542906 159128 542912 159140
rect 542964 159128 542970 159180
rect 265618 158448 265624 158500
rect 265676 158488 265682 158500
rect 406470 158488 406476 158500
rect 265676 158460 406476 158488
rect 265676 158448 265682 158460
rect 406470 158448 406476 158460
rect 406528 158448 406534 158500
rect 289262 158380 289268 158432
rect 289320 158420 289326 158432
rect 484394 158420 484400 158432
rect 289320 158392 484400 158420
rect 289320 158380 289326 158392
rect 484394 158380 484400 158392
rect 484452 158380 484458 158432
rect 150158 158312 150164 158364
rect 150216 158352 150222 158364
rect 358906 158352 358912 158364
rect 150216 158324 358912 158352
rect 150216 158312 150222 158324
rect 358906 158312 358912 158324
rect 358964 158312 358970 158364
rect 402514 158312 402520 158364
rect 402572 158352 402578 158364
rect 553854 158352 553860 158364
rect 402572 158324 553860 158352
rect 402572 158312 402578 158324
rect 553854 158312 553860 158324
rect 553912 158312 553918 158364
rect 92474 158244 92480 158296
rect 92532 158284 92538 158296
rect 320818 158284 320824 158296
rect 92532 158256 320824 158284
rect 92532 158244 92538 158256
rect 320818 158244 320824 158256
rect 320876 158244 320882 158296
rect 334066 158244 334072 158296
rect 334124 158284 334130 158296
rect 550082 158284 550088 158296
rect 334124 158256 550088 158284
rect 334124 158244 334130 158256
rect 550082 158244 550088 158256
rect 550140 158244 550146 158296
rect 56226 158176 56232 158228
rect 56284 158216 56290 158228
rect 349522 158216 349528 158228
rect 56284 158188 349528 158216
rect 56284 158176 56290 158188
rect 349522 158176 349528 158188
rect 349580 158176 349586 158228
rect 391750 158176 391756 158228
rect 391808 158216 391814 158228
rect 556430 158216 556436 158228
rect 391808 158188 556436 158216
rect 391808 158176 391814 158188
rect 556430 158176 556436 158188
rect 556488 158176 556494 158228
rect 57238 158108 57244 158160
rect 57296 158148 57302 158160
rect 353938 158148 353944 158160
rect 57296 158120 353944 158148
rect 57296 158108 57302 158120
rect 353938 158108 353944 158120
rect 353996 158108 354002 158160
rect 382090 158108 382096 158160
rect 382148 158148 382154 158160
rect 549806 158148 549812 158160
rect 382148 158120 549812 158148
rect 382148 158108 382154 158120
rect 549806 158108 549812 158120
rect 549864 158108 549870 158160
rect 47854 158040 47860 158092
rect 47912 158080 47918 158092
rect 204254 158080 204260 158092
rect 47912 158052 204260 158080
rect 47912 158040 47918 158052
rect 204254 158040 204260 158052
rect 204312 158040 204318 158092
rect 219710 158040 219716 158092
rect 219768 158080 219774 158092
rect 559190 158080 559196 158092
rect 219768 158052 559196 158080
rect 219768 158040 219774 158052
rect 559190 158040 559196 158052
rect 559248 158040 559254 158092
rect 33870 157972 33876 158024
rect 33928 158012 33934 158024
rect 529934 158012 529940 158024
rect 33928 157984 529940 158012
rect 33928 157972 33934 157984
rect 529934 157972 529940 157984
rect 529992 157972 529998 158024
rect 333974 157292 333980 157344
rect 334032 157332 334038 157344
rect 541342 157332 541348 157344
rect 334032 157304 541348 157332
rect 334032 157292 334038 157304
rect 541342 157292 541348 157304
rect 541400 157292 541406 157344
rect 117958 157224 117964 157276
rect 118016 157264 118022 157276
rect 343358 157264 343364 157276
rect 118016 157236 343364 157264
rect 118016 157224 118022 157236
rect 343358 157224 343364 157236
rect 343416 157224 343422 157276
rect 407942 157224 407948 157276
rect 408000 157264 408006 157276
rect 564618 157264 564624 157276
rect 408000 157236 564624 157264
rect 408000 157224 408006 157236
rect 564618 157224 564624 157236
rect 564676 157224 564682 157276
rect 78766 157156 78772 157208
rect 78824 157196 78830 157208
rect 323394 157196 323400 157208
rect 78824 157168 323400 157196
rect 78824 157156 78830 157168
rect 323394 157156 323400 157168
rect 323452 157156 323458 157208
rect 330478 157156 330484 157208
rect 330536 157196 330542 157208
rect 572162 157196 572168 157208
rect 330536 157168 572168 157196
rect 330536 157156 330542 157168
rect 572162 157156 572168 157168
rect 572220 157156 572226 157208
rect 106366 157088 106372 157140
rect 106424 157128 106430 157140
rect 370498 157128 370504 157140
rect 106424 157100 370504 157128
rect 106424 157088 106430 157100
rect 370498 157088 370504 157100
rect 370556 157088 370562 157140
rect 391014 157088 391020 157140
rect 391072 157128 391078 157140
rect 567654 157128 567660 157140
rect 391072 157100 567660 157128
rect 391072 157088 391078 157100
rect 567654 157088 567660 157100
rect 567712 157088 567718 157140
rect 80146 157020 80152 157072
rect 80204 157060 80210 157072
rect 281534 157060 281540 157072
rect 80204 157032 281540 157060
rect 80204 157020 80210 157032
rect 281534 157020 281540 157032
rect 281592 157020 281598 157072
rect 306374 157020 306380 157072
rect 306432 157060 306438 157072
rect 570690 157060 570696 157072
rect 306432 157032 570696 157060
rect 306432 157020 306438 157032
rect 570690 157020 570696 157032
rect 570748 157020 570754 157072
rect 253934 156952 253940 157004
rect 253992 156992 253998 157004
rect 555510 156992 555516 157004
rect 253992 156964 555516 156992
rect 253992 156952 253998 156964
rect 555510 156952 555516 156964
rect 555568 156952 555574 157004
rect 200114 156884 200120 156936
rect 200172 156924 200178 156936
rect 506290 156924 506296 156936
rect 200172 156896 506296 156924
rect 200172 156884 200178 156896
rect 506290 156884 506296 156896
rect 506348 156884 506354 156936
rect 231946 156816 231952 156868
rect 232004 156856 232010 156868
rect 567470 156856 567476 156868
rect 232004 156828 567476 156856
rect 232004 156816 232010 156828
rect 567470 156816 567476 156828
rect 567528 156816 567534 156868
rect 37826 156748 37832 156800
rect 37884 156788 37890 156800
rect 380710 156788 380716 156800
rect 37884 156760 380716 156788
rect 37884 156748 37890 156760
rect 380710 156748 380716 156760
rect 380768 156748 380774 156800
rect 381998 156748 382004 156800
rect 382056 156788 382062 156800
rect 577498 156788 577504 156800
rect 382056 156760 577504 156788
rect 382056 156748 382062 156760
rect 577498 156748 577504 156760
rect 577556 156748 577562 156800
rect 212534 156680 212540 156732
rect 212592 156720 212598 156732
rect 560478 156720 560484 156732
rect 212592 156692 560484 156720
rect 212592 156680 212598 156692
rect 560478 156680 560484 156692
rect 560536 156680 560542 156732
rect 184934 156612 184940 156664
rect 184992 156652 184998 156664
rect 568850 156652 568856 156664
rect 184992 156624 568856 156652
rect 184992 156612 184998 156624
rect 568850 156612 568856 156624
rect 568908 156612 568914 156664
rect 283558 156544 283564 156596
rect 283616 156584 283622 156596
rect 481818 156584 481824 156596
rect 283616 156556 481824 156584
rect 283616 156544 283622 156556
rect 481818 156544 481824 156556
rect 481876 156544 481882 156596
rect 388714 156476 388720 156528
rect 388772 156516 388778 156528
rect 542630 156516 542636 156528
rect 388772 156488 542636 156516
rect 388772 156476 388778 156488
rect 542630 156476 542636 156488
rect 542688 156476 542694 156528
rect 409782 156408 409788 156460
rect 409840 156448 409846 156460
rect 559190 156448 559196 156460
rect 409840 156420 559196 156448
rect 409840 156408 409846 156420
rect 559190 156408 559196 156420
rect 559248 156408 559254 156460
rect 47670 155864 47676 155916
rect 47728 155904 47734 155916
rect 141142 155904 141148 155916
rect 47728 155876 141148 155904
rect 47728 155864 47734 155876
rect 141142 155864 141148 155876
rect 141200 155864 141206 155916
rect 175274 155864 175280 155916
rect 175332 155904 175338 155916
rect 289814 155904 289820 155916
rect 175332 155876 289820 155904
rect 175332 155864 175338 155876
rect 289814 155864 289820 155876
rect 289872 155864 289878 155916
rect 407758 155864 407764 155916
rect 407816 155904 407822 155916
rect 540054 155904 540060 155916
rect 407816 155876 540060 155904
rect 407816 155864 407822 155876
rect 540054 155864 540060 155876
rect 540112 155864 540118 155916
rect 47854 155796 47860 155848
rect 47912 155836 47918 155848
rect 162854 155836 162860 155848
rect 47912 155808 162860 155836
rect 47912 155796 47918 155808
rect 162854 155796 162860 155808
rect 162912 155796 162918 155848
rect 232590 155796 232596 155848
rect 232648 155836 232654 155848
rect 348602 155836 348608 155848
rect 232648 155808 348608 155836
rect 232648 155796 232654 155808
rect 348602 155796 348608 155808
rect 348660 155796 348666 155848
rect 407390 155796 407396 155848
rect 407448 155836 407454 155848
rect 563054 155836 563060 155848
rect 407448 155808 563060 155836
rect 407448 155796 407454 155808
rect 563054 155796 563060 155808
rect 563112 155796 563118 155848
rect 39206 155728 39212 155780
rect 39264 155768 39270 155780
rect 160186 155768 160192 155780
rect 39264 155740 160192 155768
rect 39264 155728 39270 155740
rect 160186 155728 160192 155740
rect 160244 155728 160250 155780
rect 179414 155728 179420 155780
rect 179472 155768 179478 155780
rect 229370 155768 229376 155780
rect 179472 155740 229376 155768
rect 179472 155728 179478 155740
rect 229370 155728 229376 155740
rect 229428 155728 229434 155780
rect 230014 155728 230020 155780
rect 230072 155768 230078 155780
rect 354214 155768 354220 155780
rect 230072 155740 354220 155768
rect 230072 155728 230078 155740
rect 354214 155728 354220 155740
rect 354272 155728 354278 155780
rect 401410 155728 401416 155780
rect 401468 155768 401474 155780
rect 556522 155768 556528 155780
rect 401468 155740 556528 155768
rect 401468 155728 401474 155740
rect 556522 155728 556528 155740
rect 556580 155728 556586 155780
rect 46382 155660 46388 155712
rect 46440 155700 46446 155712
rect 204898 155700 204904 155712
rect 46440 155672 204904 155700
rect 46440 155660 46446 155672
rect 204898 155660 204904 155672
rect 204956 155660 204962 155712
rect 220814 155660 220820 155712
rect 220872 155700 220878 155712
rect 252646 155700 252652 155712
rect 220872 155672 252652 155700
rect 220872 155660 220878 155672
rect 252646 155660 252652 155672
rect 252704 155660 252710 155712
rect 291194 155660 291200 155712
rect 291252 155700 291258 155712
rect 340138 155700 340144 155712
rect 291252 155672 340144 155700
rect 291252 155660 291258 155672
rect 340138 155660 340144 155672
rect 340196 155660 340202 155712
rect 346394 155660 346400 155712
rect 346452 155700 346458 155712
rect 560754 155700 560760 155712
rect 346452 155672 560760 155700
rect 346452 155660 346458 155672
rect 560754 155660 560760 155672
rect 560812 155660 560818 155712
rect 28626 155592 28632 155644
rect 28684 155632 28690 155644
rect 240962 155632 240968 155644
rect 28684 155604 240968 155632
rect 28684 155592 28690 155604
rect 240962 155592 240968 155604
rect 241020 155592 241026 155644
rect 269114 155592 269120 155644
rect 269172 155632 269178 155644
rect 322750 155632 322756 155644
rect 269172 155604 322756 155632
rect 269172 155592 269178 155604
rect 322750 155592 322756 155604
rect 322808 155592 322814 155644
rect 338114 155592 338120 155644
rect 338172 155632 338178 155644
rect 562410 155632 562416 155644
rect 338172 155604 562416 155632
rect 338172 155592 338178 155604
rect 562410 155592 562416 155604
rect 562468 155592 562474 155644
rect 37734 155524 37740 155576
rect 37792 155564 37798 155576
rect 284110 155564 284116 155576
rect 37792 155536 284116 155564
rect 37792 155524 37798 155536
rect 284110 155524 284116 155536
rect 284168 155524 284174 155576
rect 302234 155524 302240 155576
rect 302292 155564 302298 155576
rect 560570 155564 560576 155576
rect 302292 155536 560576 155564
rect 302292 155524 302298 155536
rect 560570 155524 560576 155536
rect 560628 155524 560634 155576
rect 51994 155456 52000 155508
rect 52052 155496 52058 155508
rect 57974 155496 57980 155508
rect 52052 155468 57980 155496
rect 52052 155456 52058 155468
rect 57974 155456 57980 155468
rect 58032 155456 58038 155508
rect 74810 155456 74816 155508
rect 74868 155496 74874 155508
rect 376386 155496 376392 155508
rect 74868 155468 376392 155496
rect 74868 155456 74874 155468
rect 376386 155456 376392 155468
rect 376444 155456 376450 155508
rect 401226 155456 401232 155508
rect 401284 155496 401290 155508
rect 566458 155496 566464 155508
rect 401284 155468 566464 155496
rect 401284 155456 401290 155468
rect 566458 155456 566464 155468
rect 566516 155456 566522 155508
rect 55766 155388 55772 155440
rect 55824 155428 55830 155440
rect 365990 155428 365996 155440
rect 55824 155400 365996 155428
rect 55824 155388 55830 155400
rect 365990 155388 365996 155400
rect 366048 155388 366054 155440
rect 394418 155388 394424 155440
rect 394476 155428 394482 155440
rect 573450 155428 573456 155440
rect 394476 155400 573456 155428
rect 394476 155388 394482 155400
rect 573450 155388 573456 155400
rect 573508 155388 573514 155440
rect 50982 155320 50988 155372
rect 51040 155360 51046 155372
rect 371234 155360 371240 155372
rect 51040 155332 371240 155360
rect 51040 155320 51046 155332
rect 371234 155320 371240 155332
rect 371292 155320 371298 155372
rect 374914 155320 374920 155372
rect 374972 155360 374978 155372
rect 554038 155360 554044 155372
rect 374972 155332 554044 155360
rect 374972 155320 374978 155332
rect 554038 155320 554044 155332
rect 554096 155320 554102 155372
rect 40862 155252 40868 155304
rect 40920 155292 40926 155304
rect 365898 155292 365904 155304
rect 40920 155264 365904 155292
rect 40920 155252 40926 155264
rect 365898 155252 365904 155264
rect 365956 155252 365962 155304
rect 382182 155252 382188 155304
rect 382240 155292 382246 155304
rect 571886 155292 571892 155304
rect 382240 155264 571892 155292
rect 382240 155252 382246 155264
rect 571886 155252 571892 155264
rect 571944 155252 571950 155304
rect 38010 155184 38016 155236
rect 38068 155224 38074 155236
rect 208394 155224 208400 155236
rect 38068 155196 208400 155224
rect 38068 155184 38074 155196
rect 208394 155184 208400 155196
rect 208452 155184 208458 155236
rect 216674 155184 216680 155236
rect 216732 155224 216738 155236
rect 578234 155224 578240 155236
rect 216732 155196 578240 155224
rect 216732 155184 216738 155196
rect 578234 155184 578240 155196
rect 578292 155184 578298 155236
rect 49142 155116 49148 155168
rect 49200 155156 49206 155168
rect 136634 155156 136640 155168
rect 49200 155128 136640 155156
rect 49200 155116 49206 155128
rect 136634 155116 136640 155128
rect 136692 155116 136698 155168
rect 268010 155116 268016 155168
rect 268068 155156 268074 155168
rect 357618 155156 357624 155168
rect 268068 155128 357624 155156
rect 268068 155116 268074 155128
rect 357618 155116 357624 155128
rect 357676 155116 357682 155168
rect 251910 154776 251916 154828
rect 251968 154816 251974 154828
rect 259454 154816 259460 154828
rect 251968 154788 259460 154816
rect 251968 154776 251974 154788
rect 259454 154776 259460 154788
rect 259512 154776 259518 154828
rect 540606 154776 540612 154828
rect 540664 154776 540670 154828
rect 540624 154624 540652 154776
rect 540606 154572 540612 154624
rect 540664 154572 540670 154624
rect 401318 154504 401324 154556
rect 401376 154544 401382 154556
rect 540514 154544 540520 154556
rect 401376 154516 540520 154544
rect 401376 154504 401382 154516
rect 540514 154504 540520 154516
rect 540572 154504 540578 154556
rect 405274 154436 405280 154488
rect 405332 154476 405338 154488
rect 546310 154476 546316 154488
rect 405332 154448 546316 154476
rect 405332 154436 405338 154448
rect 546310 154436 546316 154448
rect 546368 154436 546374 154488
rect 404998 154368 405004 154420
rect 405056 154408 405062 154420
rect 557994 154408 558000 154420
rect 405056 154380 558000 154408
rect 405056 154368 405062 154380
rect 557994 154368 558000 154380
rect 558052 154368 558058 154420
rect 296346 154300 296352 154352
rect 296404 154340 296410 154352
rect 388806 154340 388812 154352
rect 296404 154312 388812 154340
rect 296404 154300 296410 154312
rect 388806 154300 388812 154312
rect 388864 154300 388870 154352
rect 391198 154300 391204 154352
rect 391256 154340 391262 154352
rect 546586 154340 546592 154352
rect 391256 154312 546592 154340
rect 391256 154300 391262 154312
rect 546586 154300 546592 154312
rect 546644 154300 546650 154352
rect 73430 154232 73436 154284
rect 73488 154272 73494 154284
rect 224218 154272 224224 154284
rect 73488 154244 224224 154272
rect 73488 154232 73494 154244
rect 224218 154232 224224 154244
rect 224276 154232 224282 154284
rect 382826 154232 382832 154284
rect 382884 154272 382890 154284
rect 542722 154272 542728 154284
rect 382884 154244 542728 154272
rect 382884 154232 382890 154244
rect 542722 154232 542728 154244
rect 542780 154232 542786 154284
rect 106274 154164 106280 154216
rect 106332 154204 106338 154216
rect 308582 154204 308588 154216
rect 106332 154176 308588 154204
rect 106332 154164 106338 154176
rect 308582 154164 308588 154176
rect 308640 154164 308646 154216
rect 395614 154164 395620 154216
rect 395672 154204 395678 154216
rect 565078 154204 565084 154216
rect 395672 154176 565084 154204
rect 395672 154164 395678 154176
rect 565078 154164 565084 154176
rect 565136 154164 565142 154216
rect 39574 154096 39580 154148
rect 39632 154136 39638 154148
rect 238754 154136 238760 154148
rect 39632 154108 238760 154136
rect 39632 154096 39638 154108
rect 238754 154096 238760 154108
rect 238812 154096 238818 154148
rect 260282 154096 260288 154148
rect 260340 154136 260346 154148
rect 299474 154136 299480 154148
rect 260340 154108 299480 154136
rect 260340 154096 260346 154108
rect 299474 154096 299480 154108
rect 299532 154096 299538 154148
rect 304994 154096 305000 154148
rect 305052 154136 305058 154148
rect 546862 154136 546868 154148
rect 305052 154108 546868 154136
rect 305052 154096 305058 154108
rect 546862 154096 546868 154108
rect 546920 154096 546926 154148
rect 58894 154028 58900 154080
rect 58952 154068 58958 154080
rect 359550 154068 359556 154080
rect 58952 154040 359556 154068
rect 58952 154028 58958 154040
rect 359550 154028 359556 154040
rect 359608 154028 359614 154080
rect 382918 154028 382924 154080
rect 382976 154068 382982 154080
rect 569218 154068 569224 154080
rect 382976 154040 569224 154068
rect 382976 154028 382982 154040
rect 569218 154028 569224 154040
rect 569276 154028 569282 154080
rect 91094 153960 91100 154012
rect 91152 154000 91158 154012
rect 166902 154000 166908 154012
rect 91152 153972 166908 154000
rect 91152 153960 91158 153972
rect 166902 153960 166908 153972
rect 166960 153960 166966 154012
rect 178034 153960 178040 154012
rect 178092 154000 178098 154012
rect 544930 154000 544936 154012
rect 178092 153972 544936 154000
rect 178092 153960 178098 153972
rect 544930 153960 544936 153972
rect 544988 153960 544994 154012
rect 124214 153892 124220 153944
rect 124272 153932 124278 153944
rect 548886 153932 548892 153944
rect 124272 153904 548892 153932
rect 124272 153892 124278 153904
rect 548886 153892 548892 153904
rect 548944 153892 548950 153944
rect 80054 153824 80060 153876
rect 80112 153864 80118 153876
rect 553026 153864 553032 153876
rect 80112 153836 553032 153864
rect 80112 153824 80118 153836
rect 553026 153824 553032 153836
rect 553084 153824 553090 153876
rect 408126 153756 408132 153808
rect 408184 153796 408190 153808
rect 540790 153796 540796 153808
rect 408184 153768 540796 153796
rect 408184 153756 408190 153768
rect 540790 153756 540796 153768
rect 540848 153756 540854 153808
rect 451274 153688 451280 153740
rect 451332 153728 451338 153740
rect 574278 153728 574284 153740
rect 451332 153700 574284 153728
rect 451332 153688 451338 153700
rect 574278 153688 574284 153700
rect 574336 153688 574342 153740
rect 518894 153620 518900 153672
rect 518952 153660 518958 153672
rect 568022 153660 568028 153672
rect 518952 153632 568028 153660
rect 518952 153620 518958 153632
rect 568022 153620 568028 153632
rect 568080 153620 568086 153672
rect 376938 153280 376944 153332
rect 376996 153320 377002 153332
rect 377214 153320 377220 153332
rect 376996 153292 377220 153320
rect 376996 153280 377002 153292
rect 377214 153280 377220 153292
rect 377272 153280 377278 153332
rect 29638 153144 29644 153196
rect 29696 153184 29702 153196
rect 88978 153184 88984 153196
rect 29696 153156 88984 153184
rect 29696 153144 29702 153156
rect 88978 153144 88984 153156
rect 89036 153144 89042 153196
rect 89806 153144 89812 153196
rect 89864 153184 89870 153196
rect 99282 153184 99288 153196
rect 89864 153156 99288 153184
rect 89864 153144 89870 153156
rect 99282 153144 99288 153156
rect 99340 153144 99346 153196
rect 347866 153144 347872 153196
rect 347924 153184 347930 153196
rect 347924 153156 369854 153184
rect 347924 153144 347930 153156
rect 24118 153076 24124 153128
rect 24176 153116 24182 153128
rect 107654 153116 107660 153128
rect 24176 153088 107660 153116
rect 24176 153076 24182 153088
rect 107654 153076 107660 153088
rect 107712 153076 107718 153128
rect 112162 153076 112168 153128
rect 112220 153116 112226 153128
rect 120718 153116 120724 153128
rect 112220 153088 120724 153116
rect 112220 153076 112226 153088
rect 120718 153076 120724 153088
rect 120776 153076 120782 153128
rect 135990 153076 135996 153128
rect 136048 153116 136054 153128
rect 166258 153116 166264 153128
rect 136048 153088 166264 153116
rect 136048 153076 136054 153088
rect 166258 153076 166264 153088
rect 166316 153076 166322 153128
rect 327258 153076 327264 153128
rect 327316 153116 327322 153128
rect 354858 153116 354864 153128
rect 327316 153088 354864 153116
rect 327316 153076 327322 153088
rect 354858 153076 354864 153088
rect 354916 153076 354922 153128
rect 354950 153076 354956 153128
rect 355008 153116 355014 153128
rect 358078 153116 358084 153128
rect 355008 153088 358084 153116
rect 355008 153076 355014 153088
rect 358078 153076 358084 153088
rect 358136 153076 358142 153128
rect 369826 153116 369854 153156
rect 374638 153144 374644 153196
rect 374696 153184 374702 153196
rect 383286 153184 383292 153196
rect 374696 153156 383292 153184
rect 374696 153144 374702 153156
rect 383286 153144 383292 153156
rect 383344 153144 383350 153196
rect 396718 153144 396724 153196
rect 396776 153184 396782 153196
rect 434162 153184 434168 153196
rect 396776 153156 434168 153184
rect 396776 153144 396782 153156
rect 434162 153144 434168 153156
rect 434220 153144 434226 153196
rect 500218 153144 500224 153196
rect 500276 153184 500282 153196
rect 507578 153184 507584 153196
rect 500276 153156 507584 153184
rect 500276 153144 500282 153156
rect 507578 153144 507584 153156
rect 507636 153144 507642 153196
rect 507670 153144 507676 153196
rect 507728 153184 507734 153196
rect 559650 153184 559656 153196
rect 507728 153156 559656 153184
rect 507728 153144 507734 153156
rect 559650 153144 559656 153156
rect 559708 153144 559714 153196
rect 376754 153116 376760 153128
rect 369826 153088 376760 153116
rect 376754 153076 376760 153088
rect 376812 153076 376818 153128
rect 380250 153076 380256 153128
rect 380308 153116 380314 153128
rect 425146 153116 425152 153128
rect 380308 153088 425152 153116
rect 380308 153076 380314 153088
rect 425146 153076 425152 153088
rect 425204 153076 425210 153128
rect 491294 153076 491300 153128
rect 491352 153116 491358 153128
rect 492122 153116 492128 153128
rect 491352 153088 492128 153116
rect 491352 153076 491358 153088
rect 492122 153076 492128 153088
rect 492180 153076 492186 153128
rect 498194 153076 498200 153128
rect 498252 153116 498258 153128
rect 572714 153116 572720 153128
rect 498252 153088 572720 153116
rect 498252 153076 498258 153088
rect 572714 153076 572720 153088
rect 572772 153076 572778 153128
rect 58250 153008 58256 153060
rect 58308 153048 58314 153060
rect 154574 153048 154580 153060
rect 58308 153020 154580 153048
rect 58308 153008 58314 153020
rect 154574 153008 154580 153020
rect 154632 153008 154638 153060
rect 160094 153008 160100 153060
rect 160152 153048 160158 153060
rect 188798 153048 188804 153060
rect 160152 153020 188804 153048
rect 160152 153008 160158 153020
rect 188798 153008 188804 153020
rect 188856 153008 188862 153060
rect 325050 153008 325056 153060
rect 325108 153048 325114 153060
rect 358814 153048 358820 153060
rect 325108 153020 358820 153048
rect 325108 153008 325114 153020
rect 358814 153008 358820 153020
rect 358872 153008 358878 153060
rect 394050 153008 394056 153060
rect 394108 153048 394114 153060
rect 448974 153048 448980 153060
rect 394108 153020 448980 153048
rect 394108 153008 394114 153020
rect 448974 153008 448980 153020
rect 449032 153008 449038 153060
rect 482922 153008 482928 153060
rect 482980 153048 482986 153060
rect 558086 153048 558092 153060
rect 482980 153020 558092 153048
rect 482980 153008 482986 153020
rect 558086 153008 558092 153020
rect 558144 153008 558150 153060
rect 30926 152940 30932 152992
rect 30984 152980 30990 152992
rect 93486 152980 93492 152992
rect 30984 152952 93492 152980
rect 30984 152940 30990 152952
rect 93486 152940 93492 152952
rect 93544 152940 93550 152992
rect 94774 152940 94780 152992
rect 94832 152980 94838 152992
rect 201402 152980 201408 152992
rect 94832 152952 201408 152980
rect 94832 152940 94838 152952
rect 201402 152940 201408 152952
rect 201460 152940 201466 152992
rect 316586 152940 316592 152992
rect 316644 152980 316650 152992
rect 356054 152980 356060 152992
rect 316644 152952 356060 152980
rect 316644 152940 316650 152952
rect 356054 152940 356060 152952
rect 356112 152940 356118 152992
rect 395338 152940 395344 152992
rect 395396 152980 395402 152992
rect 529198 152980 529204 152992
rect 395396 152952 529204 152980
rect 395396 152940 395402 152952
rect 529198 152940 529204 152952
rect 529256 152940 529262 152992
rect 531406 152940 531412 152992
rect 531464 152980 531470 152992
rect 534718 152980 534724 152992
rect 531464 152952 534724 152980
rect 531464 152940 531470 152952
rect 534718 152940 534724 152952
rect 534776 152940 534782 152992
rect 537570 152940 537576 152992
rect 537628 152980 537634 152992
rect 575934 152980 575940 152992
rect 537628 152952 575940 152980
rect 537628 152940 537634 152952
rect 575934 152940 575940 152952
rect 575992 152940 575998 152992
rect 55122 152872 55128 152924
rect 55180 152912 55186 152924
rect 198734 152912 198740 152924
rect 55180 152884 198740 152912
rect 55180 152872 55186 152884
rect 198734 152872 198740 152884
rect 198792 152872 198798 152924
rect 200390 152872 200396 152924
rect 200448 152912 200454 152924
rect 354766 152912 354772 152924
rect 200448 152884 354772 152912
rect 200448 152872 200454 152884
rect 354766 152872 354772 152884
rect 354824 152872 354830 152924
rect 354858 152872 354864 152924
rect 354916 152912 354922 152924
rect 361574 152912 361580 152924
rect 354916 152884 361580 152912
rect 354916 152872 354922 152884
rect 361574 152872 361580 152884
rect 361632 152872 361638 152924
rect 408034 152872 408040 152924
rect 408092 152912 408098 152924
rect 555142 152912 555148 152924
rect 408092 152884 555148 152912
rect 408092 152872 408098 152884
rect 555142 152872 555148 152884
rect 555200 152872 555206 152924
rect 26786 152804 26792 152856
rect 26844 152844 26850 152856
rect 125042 152844 125048 152856
rect 26844 152816 125048 152844
rect 26844 152804 26850 152816
rect 125042 152804 125048 152816
rect 125100 152804 125106 152856
rect 127618 152804 127624 152856
rect 127676 152844 127682 152856
rect 289262 152844 289268 152856
rect 127676 152816 289268 152844
rect 127676 152804 127682 152816
rect 289262 152804 289268 152816
rect 289320 152804 289326 152856
rect 334986 152804 334992 152856
rect 335044 152844 335050 152856
rect 378778 152844 378784 152856
rect 335044 152816 378784 152844
rect 335044 152804 335050 152816
rect 378778 152804 378784 152816
rect 378836 152804 378842 152856
rect 407022 152804 407028 152856
rect 407080 152844 407086 152856
rect 554130 152844 554136 152856
rect 407080 152816 554136 152844
rect 407080 152804 407086 152816
rect 554130 152804 554136 152816
rect 554188 152804 554194 152856
rect 32490 152736 32496 152788
rect 32548 152776 32554 152788
rect 202966 152776 202972 152788
rect 32548 152748 202972 152776
rect 32548 152736 32554 152748
rect 202966 152736 202972 152748
rect 203024 152736 203030 152788
rect 310514 152736 310520 152788
rect 310572 152776 310578 152788
rect 357434 152776 357440 152788
rect 310572 152748 357440 152776
rect 310572 152736 310578 152748
rect 357434 152736 357440 152748
rect 357492 152736 357498 152788
rect 381538 152736 381544 152788
rect 381596 152776 381602 152788
rect 391658 152776 391664 152788
rect 381596 152748 391664 152776
rect 381596 152736 381602 152748
rect 391658 152736 391664 152748
rect 391716 152736 391722 152788
rect 406930 152736 406936 152788
rect 406988 152776 406994 152788
rect 563882 152776 563888 152788
rect 406988 152748 563888 152776
rect 406988 152736 406994 152748
rect 563882 152736 563888 152748
rect 563940 152736 563946 152788
rect 37918 152668 37924 152720
rect 37976 152708 37982 152720
rect 209774 152708 209780 152720
rect 37976 152680 209780 152708
rect 37976 152668 37982 152680
rect 209774 152668 209780 152680
rect 209832 152668 209838 152720
rect 315022 152668 315028 152720
rect 315080 152708 315086 152720
rect 393958 152708 393964 152720
rect 315080 152680 393964 152708
rect 315080 152668 315086 152680
rect 393958 152668 393964 152680
rect 394016 152668 394022 152720
rect 409598 152668 409604 152720
rect 409656 152708 409662 152720
rect 566550 152708 566556 152720
rect 409656 152680 566556 152708
rect 409656 152668 409662 152680
rect 566550 152668 566556 152680
rect 566608 152668 566614 152720
rect 32306 152600 32312 152652
rect 32364 152640 32370 152652
rect 208762 152640 208768 152652
rect 32364 152612 208768 152640
rect 32364 152600 32370 152612
rect 208762 152600 208768 152612
rect 208820 152600 208826 152652
rect 287974 152600 287980 152652
rect 288032 152640 288038 152652
rect 377858 152640 377864 152652
rect 288032 152612 377864 152640
rect 288032 152600 288038 152612
rect 377858 152600 377864 152612
rect 377916 152600 377922 152652
rect 381630 152600 381636 152652
rect 381688 152640 381694 152652
rect 545114 152640 545120 152652
rect 381688 152612 545120 152640
rect 381688 152600 381694 152612
rect 545114 152600 545120 152612
rect 545172 152600 545178 152652
rect 36630 152532 36636 152584
rect 36688 152572 36694 152584
rect 297634 152572 297640 152584
rect 36688 152544 297640 152572
rect 36688 152532 36694 152544
rect 297634 152532 297640 152544
rect 297692 152532 297698 152584
rect 309226 152532 309232 152584
rect 309284 152572 309290 152584
rect 357526 152572 357532 152584
rect 309284 152544 357532 152572
rect 309284 152532 309290 152544
rect 357526 152532 357532 152544
rect 357584 152532 357590 152584
rect 376110 152532 376116 152584
rect 376168 152572 376174 152584
rect 542262 152572 542268 152584
rect 376168 152544 542268 152572
rect 376168 152532 376174 152544
rect 542262 152532 542268 152544
rect 542320 152532 542326 152584
rect 547322 152532 547328 152584
rect 547380 152572 547386 152584
rect 555326 152572 555332 152584
rect 547380 152544 555332 152572
rect 547380 152532 547386 152544
rect 555326 152532 555332 152544
rect 555384 152532 555390 152584
rect 36446 152464 36452 152516
rect 36504 152504 36510 152516
rect 326614 152504 326620 152516
rect 36504 152476 326620 152504
rect 36504 152464 36510 152476
rect 326614 152464 326620 152476
rect 326672 152464 326678 152516
rect 344002 152464 344008 152516
rect 344060 152504 344066 152516
rect 351914 152504 351920 152516
rect 344060 152476 351920 152504
rect 344060 152464 344066 152476
rect 351914 152464 351920 152476
rect 351972 152464 351978 152516
rect 354766 152464 354772 152516
rect 354824 152504 354830 152516
rect 360838 152504 360844 152516
rect 354824 152476 360844 152504
rect 354824 152464 354830 152476
rect 360838 152464 360844 152476
rect 360896 152464 360902 152516
rect 403250 152504 403256 152516
rect 361040 152476 403256 152504
rect 50338 152396 50344 152448
rect 50396 152436 50402 152448
rect 82538 152436 82544 152448
rect 50396 152408 82544 152436
rect 50396 152396 50402 152408
rect 82538 152396 82544 152408
rect 82596 152396 82602 152448
rect 341794 152396 341800 152448
rect 341852 152436 341858 152448
rect 341852 152408 354674 152436
rect 341852 152396 341858 152408
rect 54570 152328 54576 152380
rect 54628 152368 54634 152380
rect 65794 152368 65800 152380
rect 54628 152340 65800 152368
rect 54628 152328 54634 152340
rect 65794 152328 65800 152340
rect 65852 152328 65858 152380
rect 68738 152328 68744 152380
rect 68796 152368 68802 152380
rect 69658 152368 69664 152380
rect 68796 152340 69664 152368
rect 68796 152328 68802 152340
rect 69658 152328 69664 152340
rect 69716 152328 69722 152380
rect 61286 152260 61292 152312
rect 61344 152300 61350 152312
rect 68278 152300 68284 152312
rect 61344 152272 68284 152300
rect 61344 152260 61350 152272
rect 68278 152260 68284 152272
rect 68336 152260 68342 152312
rect 354646 152300 354674 152408
rect 355318 152328 355324 152380
rect 355376 152368 355382 152380
rect 361040 152368 361068 152476
rect 403250 152464 403256 152476
rect 403308 152464 403314 152516
rect 403802 152464 403808 152516
rect 403860 152504 403866 152516
rect 580258 152504 580264 152516
rect 403860 152476 580264 152504
rect 403860 152464 403866 152476
rect 580258 152464 580264 152476
rect 580316 152464 580322 152516
rect 367738 152436 367744 152448
rect 355376 152340 361068 152368
rect 364306 152408 367744 152436
rect 355376 152328 355382 152340
rect 364306 152300 364334 152408
rect 367738 152396 367744 152408
rect 367796 152396 367802 152448
rect 385770 152396 385776 152448
rect 385828 152436 385834 152448
rect 414842 152436 414848 152448
rect 385828 152408 414848 152436
rect 385828 152396 385834 152408
rect 414842 152396 414848 152408
rect 414900 152396 414906 152448
rect 457438 152396 457444 152448
rect 457496 152436 457502 152448
rect 499850 152436 499856 152448
rect 457496 152408 499856 152436
rect 457496 152396 457502 152408
rect 499850 152396 499856 152408
rect 499908 152396 499914 152448
rect 503070 152396 503076 152448
rect 503128 152436 503134 152448
rect 503128 152408 524414 152436
rect 503128 152396 503134 152408
rect 400858 152328 400864 152380
rect 400916 152368 400922 152380
rect 410334 152368 410340 152380
rect 400916 152340 410340 152368
rect 400916 152328 400922 152340
rect 410334 152328 410340 152340
rect 410392 152328 410398 152380
rect 499574 152328 499580 152380
rect 499632 152368 499638 152380
rect 507670 152368 507676 152380
rect 499632 152340 507676 152368
rect 499632 152328 499638 152340
rect 507670 152328 507676 152340
rect 507728 152328 507734 152380
rect 524386 152368 524414 152408
rect 529198 152396 529204 152448
rect 529256 152436 529262 152448
rect 534626 152436 534632 152448
rect 529256 152408 534632 152436
rect 529256 152396 529262 152408
rect 534626 152396 534632 152408
rect 534684 152396 534690 152448
rect 537478 152436 537484 152448
rect 535748 152408 537484 152436
rect 535748 152368 535776 152408
rect 537478 152396 537484 152408
rect 537536 152396 537542 152448
rect 537846 152396 537852 152448
rect 537904 152436 537910 152448
rect 540330 152436 540336 152448
rect 537904 152408 540336 152436
rect 537904 152396 537910 152408
rect 540330 152396 540336 152408
rect 540388 152396 540394 152448
rect 524386 152340 535776 152368
rect 536834 152328 536840 152380
rect 536892 152368 536898 152380
rect 541986 152368 541992 152380
rect 536892 152340 541992 152368
rect 536892 152328 536898 152340
rect 541986 152328 541992 152340
rect 542044 152328 542050 152380
rect 354646 152272 364334 152300
rect 409138 152260 409144 152312
rect 409196 152300 409202 152312
rect 419350 152300 419356 152312
rect 409196 152272 419356 152300
rect 409196 152260 409202 152272
rect 419350 152260 419356 152272
rect 419408 152260 419414 152312
rect 505646 152260 505652 152312
rect 505704 152300 505710 152312
rect 508498 152300 508504 152312
rect 505704 152272 508504 152300
rect 505704 152260 505710 152272
rect 508498 152260 508504 152272
rect 508556 152260 508562 152312
rect 199102 151784 199108 151836
rect 199160 151824 199166 151836
rect 360194 151824 360200 151836
rect 199160 151796 360200 151824
rect 199160 151784 199166 151796
rect 360194 151784 360200 151796
rect 360252 151784 360258 151836
rect 49050 151716 49056 151768
rect 49108 151756 49114 151768
rect 76006 151756 76012 151768
rect 49108 151728 76012 151756
rect 49108 151716 49114 151728
rect 76006 151716 76012 151728
rect 76064 151716 76070 151768
rect 398650 151716 398656 151768
rect 398708 151756 398714 151768
rect 563514 151756 563520 151768
rect 398708 151728 563520 151756
rect 398708 151716 398714 151728
rect 563514 151716 563520 151728
rect 563572 151716 563578 151768
rect 54202 151648 54208 151700
rect 54260 151688 54266 151700
rect 96614 151688 96620 151700
rect 54260 151660 96620 151688
rect 54260 151648 54266 151660
rect 96614 151648 96620 151660
rect 96672 151648 96678 151700
rect 324314 151648 324320 151700
rect 324372 151688 324378 151700
rect 543182 151688 543188 151700
rect 324372 151660 543188 151688
rect 324372 151648 324378 151660
rect 543182 151648 543188 151660
rect 543240 151648 543246 151700
rect 57882 151580 57888 151632
rect 57940 151620 57946 151632
rect 58894 151620 58900 151632
rect 57940 151592 58900 151620
rect 57940 151580 57946 151592
rect 58894 151580 58900 151592
rect 58952 151580 58958 151632
rect 59998 151580 60004 151632
rect 60056 151620 60062 151632
rect 226334 151620 226340 151632
rect 60056 151592 226340 151620
rect 60056 151580 60062 151592
rect 226334 151580 226340 151592
rect 226392 151580 226398 151632
rect 252554 151580 252560 151632
rect 252612 151620 252618 151632
rect 548426 151620 548432 151632
rect 252612 151592 548432 151620
rect 252612 151580 252618 151592
rect 548426 151580 548432 151592
rect 548484 151580 548490 151632
rect 30834 151512 30840 151564
rect 30892 151552 30898 151564
rect 360102 151552 360108 151564
rect 30892 151524 360108 151552
rect 30892 151512 30898 151524
rect 360102 151512 360108 151524
rect 360160 151512 360166 151564
rect 390094 151512 390100 151564
rect 390152 151552 390158 151564
rect 567746 151552 567752 151564
rect 390152 151524 567752 151552
rect 390152 151512 390158 151524
rect 567746 151512 567752 151524
rect 567804 151512 567810 151564
rect 53466 151444 53472 151496
rect 53524 151484 53530 151496
rect 113358 151484 113364 151496
rect 53524 151456 113364 151484
rect 53524 151444 53530 151456
rect 113358 151444 113364 151456
rect 113416 151444 113422 151496
rect 222194 151444 222200 151496
rect 222252 151484 222258 151496
rect 551738 151484 551744 151496
rect 222252 151456 551744 151484
rect 222252 151444 222258 151456
rect 551738 151444 551744 151456
rect 551796 151444 551802 151496
rect 44726 151376 44732 151428
rect 44784 151416 44790 151428
rect 375466 151416 375472 151428
rect 44784 151388 375472 151416
rect 44784 151376 44790 151388
rect 375466 151376 375472 151388
rect 375524 151376 375530 151428
rect 394234 151376 394240 151428
rect 394292 151416 394298 151428
rect 572806 151416 572812 151428
rect 394292 151388 572812 151416
rect 394292 151376 394298 151388
rect 572806 151376 572812 151388
rect 572864 151376 572870 151428
rect 46382 151308 46388 151360
rect 46440 151348 46446 151360
rect 414014 151348 414020 151360
rect 46440 151320 414020 151348
rect 46440 151308 46446 151320
rect 414014 151308 414020 151320
rect 414072 151308 414078 151360
rect 537662 151308 537668 151360
rect 537720 151348 537726 151360
rect 548150 151348 548156 151360
rect 537720 151320 548156 151348
rect 537720 151308 537726 151320
rect 548150 151308 548156 151320
rect 548208 151308 548214 151360
rect 51810 151240 51816 151292
rect 51868 151280 51874 151292
rect 126974 151280 126980 151292
rect 51868 151252 126980 151280
rect 51868 151240 51874 151252
rect 126974 151240 126980 151252
rect 127032 151240 127038 151292
rect 158714 151240 158720 151292
rect 158772 151280 158778 151292
rect 547046 151280 547052 151292
rect 158772 151252 547052 151280
rect 158772 151240 158778 151252
rect 547046 151240 547052 151252
rect 547104 151240 547110 151292
rect 547874 151240 547880 151292
rect 547932 151280 547938 151292
rect 559282 151280 559288 151292
rect 547932 151252 559288 151280
rect 547932 151240 547938 151252
rect 559282 151240 559288 151252
rect 559340 151240 559346 151292
rect 45922 151172 45928 151224
rect 45980 151212 45986 151224
rect 460934 151212 460940 151224
rect 45980 151184 460940 151212
rect 45980 151172 45986 151184
rect 460934 151172 460940 151184
rect 460992 151172 460998 151224
rect 536098 151172 536104 151224
rect 536156 151212 536162 151224
rect 552290 151212 552296 151224
rect 536156 151184 552296 151212
rect 536156 151172 536162 151184
rect 552290 151172 552296 151184
rect 552348 151172 552354 151224
rect 58158 151104 58164 151156
rect 58216 151144 58222 151156
rect 111794 151144 111800 151156
rect 58216 151116 111800 151144
rect 58216 151104 58222 151116
rect 111794 151104 111800 151116
rect 111852 151104 111858 151156
rect 111886 151104 111892 151156
rect 111944 151144 111950 151156
rect 545298 151144 545304 151156
rect 111944 151116 545304 151144
rect 111944 151104 111950 151116
rect 545298 151104 545304 151116
rect 545356 151104 545362 151156
rect 547230 151104 547236 151156
rect 547288 151144 547294 151156
rect 574830 151144 574836 151156
rect 547288 151116 574836 151144
rect 547288 151104 547294 151116
rect 574830 151104 574836 151116
rect 574888 151104 574894 151156
rect 35066 151036 35072 151088
rect 35124 151076 35130 151088
rect 551370 151076 551376 151088
rect 35124 151048 551376 151076
rect 35124 151036 35130 151048
rect 551370 151036 551376 151048
rect 551428 151036 551434 151088
rect 50706 150968 50712 151020
rect 50764 151008 50770 151020
rect 70486 151008 70492 151020
rect 50764 150980 70492 151008
rect 50764 150968 50770 150980
rect 70486 150968 70492 150980
rect 70544 150968 70550 151020
rect 380434 150968 380440 151020
rect 380492 151008 380498 151020
rect 541894 151008 541900 151020
rect 380492 150980 541900 151008
rect 380492 150968 380498 150980
rect 541894 150968 541900 150980
rect 541952 150968 541958 151020
rect 51902 150900 51908 150952
rect 51960 150940 51966 150952
rect 65518 150940 65524 150952
rect 51960 150912 65524 150940
rect 51960 150900 51966 150912
rect 65518 150900 65524 150912
rect 65576 150900 65582 150952
rect 408954 150900 408960 150952
rect 409012 150940 409018 150952
rect 562226 150940 562232 150952
rect 409012 150912 562232 150940
rect 409012 150900 409018 150912
rect 562226 150900 562232 150912
rect 562284 150900 562290 150952
rect 56502 150832 56508 150884
rect 56560 150872 56566 150884
rect 59998 150872 60004 150884
rect 56560 150844 60004 150872
rect 56560 150832 56566 150844
rect 59998 150832 60004 150844
rect 60056 150832 60062 150884
rect 406746 150832 406752 150884
rect 406804 150872 406810 150884
rect 553118 150872 553124 150884
rect 406804 150844 553124 150872
rect 406804 150832 406810 150844
rect 553118 150832 553124 150844
rect 553176 150832 553182 150884
rect 50062 150764 50068 150816
rect 50120 150804 50126 150816
rect 60734 150804 60740 150816
rect 50120 150776 60740 150804
rect 50120 150764 50126 150776
rect 60734 150764 60740 150776
rect 60792 150764 60798 150816
rect 549070 150628 549076 150680
rect 549128 150668 549134 150680
rect 556614 150668 556620 150680
rect 549128 150640 556620 150668
rect 549128 150628 549134 150640
rect 556614 150628 556620 150640
rect 556672 150628 556678 150680
rect 538858 150424 538864 150476
rect 538916 150464 538922 150476
rect 540974 150464 540980 150476
rect 538916 150436 540980 150464
rect 538916 150424 538922 150436
rect 540974 150424 540980 150436
rect 541032 150424 541038 150476
rect 539042 150356 539048 150408
rect 539100 150396 539106 150408
rect 549622 150396 549628 150408
rect 539100 150368 549628 150396
rect 539100 150356 539106 150368
rect 549622 150356 549628 150368
rect 549680 150356 549686 150408
rect 540606 150288 540612 150340
rect 540664 150328 540670 150340
rect 540664 150300 546632 150328
rect 540664 150288 540670 150300
rect 495434 150220 495440 150272
rect 495492 150260 495498 150272
rect 496630 150260 496636 150272
rect 495492 150232 496636 150260
rect 495492 150220 495498 150232
rect 496630 150220 496636 150232
rect 496688 150220 496694 150272
rect 539318 150084 539324 150136
rect 539376 150124 539382 150136
rect 546494 150124 546500 150136
rect 539376 150096 546500 150124
rect 539376 150084 539382 150096
rect 546494 150084 546500 150096
rect 546552 150084 546558 150136
rect 474642 150016 474648 150068
rect 474700 150056 474706 150068
rect 480070 150056 480076 150068
rect 474700 150028 480076 150056
rect 474700 150016 474706 150028
rect 480070 150016 480076 150028
rect 480128 150016 480134 150068
rect 515030 150016 515036 150068
rect 515088 150056 515094 150068
rect 515088 150028 524414 150056
rect 515088 150016 515094 150028
rect 54570 149948 54576 150000
rect 54628 149988 54634 150000
rect 59538 149988 59544 150000
rect 54628 149960 59544 149988
rect 54628 149948 54634 149960
rect 59538 149948 59544 149960
rect 59596 149948 59602 150000
rect 524386 149988 524414 150028
rect 537938 150016 537944 150068
rect 537996 150056 538002 150068
rect 540422 150056 540428 150068
rect 537996 150028 540428 150056
rect 537996 150016 538002 150028
rect 540422 150016 540428 150028
rect 540480 150016 540486 150068
rect 451246 149960 460934 149988
rect 51442 149880 51448 149932
rect 51500 149920 51506 149932
rect 349706 149920 349712 149932
rect 51500 149892 349712 149920
rect 51500 149880 51506 149892
rect 349706 149880 349712 149892
rect 349764 149880 349770 149932
rect 370958 149920 370964 149932
rect 354646 149892 370964 149920
rect 49602 149812 49608 149864
rect 49660 149852 49666 149864
rect 354646 149852 354674 149892
rect 370958 149880 370964 149892
rect 371016 149880 371022 149932
rect 403158 149880 403164 149932
rect 403216 149880 403222 149932
rect 49660 149824 354674 149852
rect 403176 149852 403204 149880
rect 451246 149852 451274 149960
rect 459554 149920 459560 149932
rect 403176 149824 451274 149852
rect 455432 149892 459560 149920
rect 49660 149812 49666 149824
rect 53006 149744 53012 149796
rect 53064 149784 53070 149796
rect 455432 149784 455460 149892
rect 459554 149880 459560 149892
rect 459612 149880 459618 149932
rect 460906 149852 460934 149960
rect 470566 149960 481634 149988
rect 470566 149852 470594 149960
rect 474642 149920 474648 149932
rect 460906 149824 470594 149852
rect 473326 149892 474648 149920
rect 53064 149756 455460 149784
rect 53064 149744 53070 149756
rect 3510 149676 3516 149728
rect 3568 149716 3574 149728
rect 473326 149716 473354 149892
rect 474642 149880 474648 149892
rect 474700 149880 474706 149932
rect 474734 149880 474740 149932
rect 474792 149880 474798 149932
rect 480070 149880 480076 149932
rect 480128 149880 480134 149932
rect 3568 149688 473354 149716
rect 3568 149676 3574 149688
rect 474752 149512 474780 149880
rect 480088 149784 480116 149880
rect 481606 149852 481634 149960
rect 500926 149960 515260 149988
rect 524386 149960 531314 149988
rect 487126 149892 495204 149920
rect 487126 149852 487154 149892
rect 495176 149852 495204 149892
rect 500926 149852 500954 149960
rect 515030 149920 515036 149932
rect 514956 149892 515036 149920
rect 481606 149824 487154 149852
rect 488506 149824 489914 149852
rect 495176 149824 500954 149852
rect 502306 149824 511994 149852
rect 488506 149784 488534 149824
rect 480088 149756 483014 149784
rect 482986 149716 483014 149756
rect 487126 149756 488534 149784
rect 482986 149688 484394 149716
rect 484366 149648 484394 149688
rect 484366 149620 485774 149648
rect 485746 149580 485774 149620
rect 487126 149580 487154 149756
rect 485746 149552 487154 149580
rect 474752 149484 483014 149512
rect 482986 149172 483014 149484
rect 489886 149444 489914 149824
rect 502306 149784 502334 149824
rect 500926 149756 502334 149784
rect 496786 149620 498194 149648
rect 491266 149484 492674 149512
rect 491266 149444 491294 149484
rect 489886 149416 491294 149444
rect 492646 149444 492674 149484
rect 494026 149484 495434 149512
rect 494026 149444 494054 149484
rect 492646 149416 494054 149444
rect 495406 149444 495434 149484
rect 496786 149444 496814 149620
rect 498166 149580 498194 149620
rect 498166 149552 499574 149580
rect 499546 149512 499574 149552
rect 500926 149512 500954 149756
rect 511966 149716 511994 149824
rect 513346 149756 514754 149784
rect 513346 149716 513374 149756
rect 511966 149688 513374 149716
rect 514726 149716 514754 149756
rect 514956 149716 514984 149892
rect 515030 149880 515036 149892
rect 515088 149880 515094 149932
rect 515232 149852 515260 149960
rect 531286 149920 531314 149960
rect 537754 149948 537760 150000
rect 537812 149988 537818 150000
rect 546604 149988 546632 150300
rect 552842 149988 552848 150000
rect 537812 149960 543734 149988
rect 546604 149960 552848 149988
rect 537812 149948 537818 149960
rect 538858 149920 538864 149932
rect 525766 149892 528554 149920
rect 531286 149892 538864 149920
rect 525766 149852 525794 149892
rect 515232 149824 525794 149852
rect 528526 149852 528554 149892
rect 538858 149880 538864 149892
rect 538916 149880 538922 149932
rect 538950 149880 538956 149932
rect 539008 149920 539014 149932
rect 540146 149920 540152 149932
rect 539008 149892 540152 149920
rect 539008 149880 539014 149892
rect 540146 149880 540152 149892
rect 540204 149880 540210 149932
rect 543706 149920 543734 149960
rect 552842 149948 552848 149960
rect 552900 149948 552906 150000
rect 551094 149920 551100 149932
rect 543706 149892 551100 149920
rect 551094 149880 551100 149892
rect 551152 149880 551158 149932
rect 565354 149852 565360 149864
rect 528526 149824 565360 149852
rect 565354 149812 565360 149824
rect 565412 149812 565418 149864
rect 546126 149784 546132 149796
rect 531286 149756 546132 149784
rect 514726 149688 514984 149716
rect 528526 149688 529934 149716
rect 528526 149580 528554 149688
rect 513346 149552 514754 149580
rect 513346 149512 513374 149552
rect 499546 149484 500954 149512
rect 502306 149484 513374 149512
rect 514726 149512 514754 149552
rect 527146 149552 528554 149580
rect 529906 149580 529934 149688
rect 531286 149580 531314 149756
rect 546126 149744 546132 149756
rect 546184 149744 546190 149796
rect 548518 149744 548524 149796
rect 548576 149784 548582 149796
rect 560294 149784 560300 149796
rect 548576 149756 560300 149784
rect 548576 149744 548582 149756
rect 560294 149744 560300 149756
rect 560352 149744 560358 149796
rect 544378 149676 544384 149728
rect 544436 149716 544442 149728
rect 550082 149716 550088 149728
rect 544436 149688 550088 149716
rect 544436 149676 544442 149688
rect 550082 149676 550088 149688
rect 550140 149676 550146 149728
rect 529906 149552 531314 149580
rect 527146 149512 527174 149552
rect 514726 149484 527174 149512
rect 502306 149444 502334 149484
rect 495406 149416 496814 149444
rect 499546 149416 502334 149444
rect 499546 149376 499574 149416
rect 489886 149348 491294 149376
rect 489886 149308 489914 149348
rect 485746 149280 489914 149308
rect 491266 149308 491294 149348
rect 495406 149348 496814 149376
rect 495406 149308 495434 149348
rect 491266 149280 495434 149308
rect 496786 149308 496814 149348
rect 498166 149348 499574 149376
rect 498166 149308 498194 149348
rect 496786 149280 498194 149308
rect 485746 149240 485774 149280
rect 484366 149212 485774 149240
rect 484366 149172 484394 149212
rect 482986 149144 484394 149172
rect 57146 149064 57152 149116
rect 57204 149104 57210 149116
rect 59630 149104 59636 149116
rect 57204 149076 59636 149104
rect 57204 149064 57210 149076
rect 59630 149064 59636 149076
rect 59688 149064 59694 149116
rect 543642 149064 543648 149116
rect 543700 149104 543706 149116
rect 545206 149104 545212 149116
rect 543700 149076 545212 149104
rect 543700 149064 543706 149076
rect 545206 149064 545212 149076
rect 545264 149064 545270 149116
rect 554130 149064 554136 149116
rect 554188 149104 554194 149116
rect 555418 149104 555424 149116
rect 554188 149076 555424 149104
rect 554188 149064 554194 149076
rect 555418 149064 555424 149076
rect 555476 149064 555482 149116
rect 546034 148996 546040 149048
rect 546092 149036 546098 149048
rect 547874 149036 547880 149048
rect 546092 149008 547880 149036
rect 546092 148996 546098 149008
rect 547874 148996 547880 149008
rect 547932 148996 547938 149048
rect 549898 148384 549904 148436
rect 549956 148424 549962 148436
rect 559006 148424 559012 148436
rect 549956 148396 559012 148424
rect 549956 148384 549962 148396
rect 559006 148384 559012 148396
rect 559064 148384 559070 148436
rect 549990 148316 549996 148368
rect 550048 148356 550054 148368
rect 567562 148356 567568 148368
rect 550048 148328 567568 148356
rect 550048 148316 550054 148328
rect 567562 148316 567568 148328
rect 567620 148316 567626 148368
rect 541710 147636 541716 147688
rect 541768 147676 541774 147688
rect 543734 147676 543740 147688
rect 541768 147648 543740 147676
rect 541768 147636 541774 147648
rect 543734 147636 543740 147648
rect 543792 147636 543798 147688
rect 543550 147568 543556 147620
rect 543608 147608 543614 147620
rect 561858 147608 561864 147620
rect 543608 147580 561864 147608
rect 543608 147568 543614 147580
rect 561858 147568 561864 147580
rect 561916 147568 561922 147620
rect 541526 147500 541532 147552
rect 541584 147540 541590 147552
rect 543918 147540 543924 147552
rect 541584 147512 543924 147540
rect 541584 147500 541590 147512
rect 543918 147500 543924 147512
rect 543976 147500 543982 147552
rect 50246 147296 50252 147348
rect 50304 147336 50310 147348
rect 55766 147336 55772 147348
rect 50304 147308 55772 147336
rect 50304 147296 50310 147308
rect 55766 147296 55772 147308
rect 55824 147296 55830 147348
rect 542906 147296 542912 147348
rect 542964 147296 542970 147348
rect 542924 147008 542952 147296
rect 54662 146956 54668 147008
rect 54720 146996 54726 147008
rect 58618 146996 58624 147008
rect 54720 146968 58624 146996
rect 54720 146956 54726 146968
rect 58618 146956 58624 146968
rect 58676 146956 58682 147008
rect 59078 146956 59084 147008
rect 59136 146996 59142 147008
rect 59538 146996 59544 147008
rect 59136 146968 59544 146996
rect 59136 146956 59142 146968
rect 59538 146956 59544 146968
rect 59596 146956 59602 147008
rect 542538 146956 542544 147008
rect 542596 146996 542602 147008
rect 542814 146996 542820 147008
rect 542596 146968 542820 146996
rect 542596 146956 542602 146968
rect 542814 146956 542820 146968
rect 542872 146956 542878 147008
rect 542906 146956 542912 147008
rect 542964 146956 542970 147008
rect 540698 146888 540704 146940
rect 540756 146928 540762 146940
rect 540756 146900 547874 146928
rect 540756 146888 540762 146900
rect 547846 146860 547874 146900
rect 549806 146860 549812 146872
rect 547846 146832 549812 146860
rect 549806 146820 549812 146832
rect 549864 146820 549870 146872
rect 549898 146820 549904 146872
rect 549956 146860 549962 146872
rect 550818 146860 550824 146872
rect 549956 146832 550824 146860
rect 549956 146820 549962 146832
rect 550818 146820 550824 146832
rect 550876 146820 550882 146872
rect 541250 146616 541256 146668
rect 541308 146656 541314 146668
rect 544654 146656 544660 146668
rect 541308 146628 544660 146656
rect 541308 146616 541314 146628
rect 544654 146616 544660 146628
rect 544712 146616 544718 146668
rect 59814 146316 59820 146328
rect 59280 146288 59820 146316
rect 52914 146208 52920 146260
rect 52972 146248 52978 146260
rect 56502 146248 56508 146260
rect 52972 146220 56508 146248
rect 52972 146208 52978 146220
rect 56502 146208 56508 146220
rect 56560 146208 56566 146260
rect 59280 146192 59308 146288
rect 59814 146276 59820 146288
rect 59872 146276 59878 146328
rect 541802 146276 541808 146328
rect 541860 146316 541866 146328
rect 543550 146316 543556 146328
rect 541860 146288 543556 146316
rect 541860 146276 541866 146288
rect 543550 146276 543556 146288
rect 543608 146276 543614 146328
rect 540698 146208 540704 146260
rect 540756 146248 540762 146260
rect 540974 146248 540980 146260
rect 540756 146220 540980 146248
rect 540756 146208 540762 146220
rect 540974 146208 540980 146220
rect 541032 146208 541038 146260
rect 542170 146208 542176 146260
rect 542228 146248 542234 146260
rect 544102 146248 544108 146260
rect 542228 146220 544108 146248
rect 542228 146208 542234 146220
rect 544102 146208 544108 146220
rect 544160 146208 544166 146260
rect 545942 146208 545948 146260
rect 546000 146248 546006 146260
rect 550358 146248 550364 146260
rect 546000 146220 550364 146248
rect 546000 146208 546006 146220
rect 550358 146208 550364 146220
rect 550416 146208 550422 146260
rect 59262 146140 59268 146192
rect 59320 146140 59326 146192
rect 543090 146140 543096 146192
rect 543148 146180 543154 146192
rect 545206 146180 545212 146192
rect 543148 146152 545212 146180
rect 543148 146140 543154 146152
rect 545206 146140 545212 146152
rect 545264 146140 545270 146192
rect 55766 146072 55772 146124
rect 55824 146112 55830 146124
rect 59446 146112 59452 146124
rect 55824 146084 59452 146112
rect 55824 146072 55830 146084
rect 59446 146072 59452 146084
rect 59504 146072 59510 146124
rect 540514 146072 540520 146124
rect 540572 146112 540578 146124
rect 543458 146112 543464 146124
rect 540572 146084 543464 146112
rect 540572 146072 540578 146084
rect 543458 146072 543464 146084
rect 543516 146072 543522 146124
rect 546402 146072 546408 146124
rect 546460 146112 546466 146124
rect 547966 146112 547972 146124
rect 546460 146084 547972 146112
rect 546460 146072 546466 146084
rect 547966 146072 547972 146084
rect 548024 146072 548030 146124
rect 546034 145596 546040 145648
rect 546092 145636 546098 145648
rect 549346 145636 549352 145648
rect 546092 145608 549352 145636
rect 546092 145596 546098 145608
rect 549346 145596 549352 145608
rect 549404 145596 549410 145648
rect 541710 145528 541716 145580
rect 541768 145568 541774 145580
rect 545758 145568 545764 145580
rect 541768 145540 545764 145568
rect 541768 145528 541774 145540
rect 545758 145528 545764 145540
rect 545816 145528 545822 145580
rect 545850 145460 545856 145512
rect 545908 145500 545914 145512
rect 549346 145500 549352 145512
rect 545908 145472 549352 145500
rect 545908 145460 545914 145472
rect 549346 145460 549352 145472
rect 549404 145460 549410 145512
rect 540146 144848 540152 144900
rect 540204 144888 540210 144900
rect 543274 144888 543280 144900
rect 540204 144860 543280 144888
rect 540204 144848 540210 144860
rect 543274 144848 543280 144860
rect 543332 144848 543338 144900
rect 543642 144848 543648 144900
rect 543700 144888 543706 144900
rect 544746 144888 544752 144900
rect 543700 144860 544752 144888
rect 543700 144848 543706 144860
rect 544746 144848 544752 144860
rect 544804 144848 544810 144900
rect 541618 144780 541624 144832
rect 541676 144820 541682 144832
rect 544378 144820 544384 144832
rect 541676 144792 544384 144820
rect 541676 144780 541682 144792
rect 544378 144780 544384 144792
rect 544436 144780 544442 144832
rect 543182 144712 543188 144764
rect 543240 144752 543246 144764
rect 544286 144752 544292 144764
rect 543240 144724 544292 144752
rect 543240 144712 543246 144724
rect 544286 144712 544292 144724
rect 544344 144712 544350 144764
rect 540514 144168 540520 144220
rect 540572 144208 540578 144220
rect 541158 144208 541164 144220
rect 540572 144180 541164 144208
rect 540572 144168 540578 144180
rect 541158 144168 541164 144180
rect 541216 144168 541222 144220
rect 544470 144100 544476 144152
rect 544528 144140 544534 144152
rect 549438 144140 549444 144152
rect 544528 144112 549444 144140
rect 544528 144100 544534 144112
rect 549438 144100 549444 144112
rect 549496 144100 549502 144152
rect 542078 143896 542084 143948
rect 542136 143936 542142 143948
rect 544010 143936 544016 143948
rect 542136 143908 544016 143936
rect 542136 143896 542142 143908
rect 544010 143896 544016 143908
rect 544068 143896 544074 143948
rect 542998 143556 543004 143608
rect 543056 143596 543062 143608
rect 543734 143596 543740 143608
rect 543056 143568 543740 143596
rect 543056 143556 543062 143568
rect 543734 143556 543740 143568
rect 543792 143556 543798 143608
rect 547966 143556 547972 143608
rect 548024 143596 548030 143608
rect 549254 143596 549260 143608
rect 548024 143568 549260 143596
rect 548024 143556 548030 143568
rect 549254 143556 549260 143568
rect 549312 143556 549318 143608
rect 55858 143488 55864 143540
rect 55916 143528 55922 143540
rect 56962 143528 56968 143540
rect 55916 143500 56968 143528
rect 55916 143488 55922 143500
rect 56962 143488 56968 143500
rect 57020 143488 57026 143540
rect 540882 143488 540888 143540
rect 540940 143528 540946 143540
rect 542814 143528 542820 143540
rect 540940 143500 542820 143528
rect 540940 143488 540946 143500
rect 542814 143488 542820 143500
rect 542872 143488 542878 143540
rect 543182 143488 543188 143540
rect 543240 143528 543246 143540
rect 563330 143528 563336 143540
rect 543240 143500 563336 143528
rect 543240 143488 543246 143500
rect 563330 143488 563336 143500
rect 563388 143488 563394 143540
rect 540790 143420 540796 143472
rect 540848 143460 540854 143472
rect 543918 143460 543924 143472
rect 540848 143432 543924 143460
rect 540848 143420 540854 143432
rect 543918 143420 543924 143432
rect 543976 143420 543982 143472
rect 540606 143352 540612 143404
rect 540664 143392 540670 143404
rect 542814 143392 542820 143404
rect 540664 143364 542820 143392
rect 540664 143352 540670 143364
rect 542814 143352 542820 143364
rect 542872 143352 542878 143404
rect 541986 143284 541992 143336
rect 542044 143324 542050 143336
rect 545482 143324 545488 143336
rect 542044 143296 545488 143324
rect 542044 143284 542050 143296
rect 545482 143284 545488 143296
rect 545540 143284 545546 143336
rect 543090 143148 543096 143200
rect 543148 143188 543154 143200
rect 545022 143188 545028 143200
rect 543148 143160 545028 143188
rect 543148 143148 543154 143160
rect 545022 143148 545028 143160
rect 545080 143148 545086 143200
rect 50798 142808 50804 142860
rect 50856 142848 50862 142860
rect 58618 142848 58624 142860
rect 50856 142820 58624 142848
rect 50856 142808 50862 142820
rect 58618 142808 58624 142820
rect 58676 142808 58682 142860
rect 49694 142196 49700 142248
rect 49752 142236 49758 142248
rect 57146 142236 57152 142248
rect 49752 142208 57152 142236
rect 49752 142196 49758 142208
rect 57146 142196 57152 142208
rect 57204 142196 57210 142248
rect 541158 142128 541164 142180
rect 541216 142168 541222 142180
rect 544194 142168 544200 142180
rect 541216 142140 544200 142168
rect 541216 142128 541222 142140
rect 544194 142128 544200 142140
rect 544252 142128 544258 142180
rect 55030 142060 55036 142112
rect 55088 142100 55094 142112
rect 57882 142100 57888 142112
rect 55088 142072 57888 142100
rect 55088 142060 55094 142072
rect 57882 142060 57888 142072
rect 57940 142060 57946 142112
rect 543642 142060 543648 142112
rect 543700 142100 543706 142112
rect 583570 142100 583576 142112
rect 543700 142072 583576 142100
rect 543700 142060 543706 142072
rect 583570 142060 583576 142072
rect 583628 142060 583634 142112
rect 550174 141992 550180 142044
rect 550232 142032 550238 142044
rect 554222 142032 554228 142044
rect 550232 142004 554228 142032
rect 550232 141992 550238 142004
rect 554222 141992 554228 142004
rect 554280 141992 554286 142044
rect 543182 141652 543188 141704
rect 543240 141692 543246 141704
rect 546586 141692 546592 141704
rect 543240 141664 546592 141692
rect 543240 141652 543246 141664
rect 546586 141652 546592 141664
rect 546644 141652 546650 141704
rect 53834 141380 53840 141432
rect 53892 141420 53898 141432
rect 58710 141420 58716 141432
rect 53892 141392 58716 141420
rect 53892 141380 53898 141392
rect 58710 141380 58716 141392
rect 58768 141380 58774 141432
rect 542170 141108 542176 141160
rect 542228 141148 542234 141160
rect 543274 141148 543280 141160
rect 542228 141120 543280 141148
rect 542228 141108 542234 141120
rect 543274 141108 543280 141120
rect 543332 141108 543338 141160
rect 56502 140836 56508 140888
rect 56560 140876 56566 140888
rect 59538 140876 59544 140888
rect 56560 140848 59544 140876
rect 56560 140836 56566 140848
rect 59538 140836 59544 140848
rect 59596 140836 59602 140888
rect 541526 140836 541532 140888
rect 541584 140876 541590 140888
rect 543826 140876 543832 140888
rect 541584 140848 543832 140876
rect 541584 140836 541590 140848
rect 543826 140836 543832 140848
rect 543884 140836 543890 140888
rect 57054 140768 57060 140820
rect 57112 140808 57118 140820
rect 59722 140808 59728 140820
rect 57112 140780 59728 140808
rect 57112 140768 57118 140780
rect 59722 140768 59728 140780
rect 59780 140768 59786 140820
rect 542262 140768 542268 140820
rect 542320 140808 542326 140820
rect 543550 140808 543556 140820
rect 542320 140780 543556 140808
rect 542320 140768 542326 140780
rect 543550 140768 543556 140780
rect 543608 140768 543614 140820
rect 563698 140768 563704 140820
rect 563756 140808 563762 140820
rect 565170 140808 565176 140820
rect 563756 140780 565176 140808
rect 563756 140768 563762 140780
rect 565170 140768 565176 140780
rect 565228 140768 565234 140820
rect 31294 140700 31300 140752
rect 31352 140740 31358 140752
rect 57882 140740 57888 140752
rect 31352 140712 57888 140740
rect 31352 140700 31358 140712
rect 57882 140700 57888 140712
rect 57940 140700 57946 140752
rect 40310 140632 40316 140684
rect 40368 140672 40374 140684
rect 57146 140672 57152 140684
rect 40368 140644 57152 140672
rect 40368 140632 40374 140644
rect 57146 140632 57152 140644
rect 57204 140632 57210 140684
rect 545114 140020 545120 140072
rect 545172 140060 545178 140072
rect 548058 140060 548064 140072
rect 545172 140032 548064 140060
rect 545172 140020 545178 140032
rect 548058 140020 548064 140032
rect 548116 140020 548122 140072
rect 540790 139544 540796 139596
rect 540848 139584 540854 139596
rect 541710 139584 541716 139596
rect 540848 139556 541716 139584
rect 540848 139544 540854 139556
rect 541710 139544 541716 139556
rect 541768 139544 541774 139596
rect 540606 139476 540612 139528
rect 540664 139516 540670 139528
rect 540882 139516 540888 139528
rect 540664 139488 540888 139516
rect 540664 139476 540670 139488
rect 540882 139476 540888 139488
rect 540940 139476 540946 139528
rect 541250 139476 541256 139528
rect 541308 139516 541314 139528
rect 545390 139516 545396 139528
rect 541308 139488 545396 139516
rect 541308 139476 541314 139488
rect 545390 139476 545396 139488
rect 545448 139476 545454 139528
rect 563790 139476 563796 139528
rect 563848 139516 563854 139528
rect 565170 139516 565176 139528
rect 563848 139488 565176 139516
rect 563848 139476 563854 139488
rect 565170 139476 565176 139488
rect 565228 139476 565234 139528
rect 565262 139476 565268 139528
rect 565320 139516 565326 139528
rect 566642 139516 566648 139528
rect 565320 139488 566648 139516
rect 565320 139476 565326 139488
rect 566642 139476 566648 139488
rect 566700 139476 566706 139528
rect 541158 139408 541164 139460
rect 541216 139448 541222 139460
rect 541802 139448 541808 139460
rect 541216 139420 541808 139448
rect 541216 139408 541222 139420
rect 541802 139408 541808 139420
rect 541860 139408 541866 139460
rect 565354 139408 565360 139460
rect 565412 139448 565418 139460
rect 565814 139448 565820 139460
rect 565412 139420 565820 139448
rect 565412 139408 565418 139420
rect 565814 139408 565820 139420
rect 565872 139408 565878 139460
rect 543550 139340 543556 139392
rect 543608 139380 543614 139392
rect 559466 139380 559472 139392
rect 543608 139352 559472 139380
rect 543608 139340 543614 139352
rect 559466 139340 559472 139352
rect 559524 139340 559530 139392
rect 567930 139340 567936 139392
rect 567988 139380 567994 139392
rect 580442 139380 580448 139392
rect 567988 139352 580448 139380
rect 567988 139340 567994 139352
rect 580442 139340 580448 139352
rect 580500 139340 580506 139392
rect 555602 138660 555608 138712
rect 555660 138700 555666 138712
rect 563790 138700 563796 138712
rect 555660 138672 563796 138700
rect 555660 138660 555666 138672
rect 563790 138660 563796 138672
rect 563848 138660 563854 138712
rect 542170 137980 542176 138032
rect 542228 138020 542234 138032
rect 545206 138020 545212 138032
rect 542228 137992 545212 138020
rect 542228 137980 542234 137992
rect 545206 137980 545212 137992
rect 545264 137980 545270 138032
rect 21542 137912 21548 137964
rect 21600 137952 21606 137964
rect 57882 137952 57888 137964
rect 21600 137924 57888 137952
rect 21600 137912 21606 137924
rect 57882 137912 57888 137924
rect 57940 137912 57946 137964
rect 3142 137844 3148 137896
rect 3200 137884 3206 137896
rect 32398 137884 32404 137896
rect 3200 137856 32404 137884
rect 3200 137844 3206 137856
rect 32398 137844 32404 137856
rect 32456 137844 32462 137896
rect 558178 137708 558184 137760
rect 558236 137748 558242 137760
rect 559466 137748 559472 137760
rect 558236 137720 559472 137748
rect 558236 137708 558242 137720
rect 559466 137708 559472 137720
rect 559524 137708 559530 137760
rect 544746 137504 544752 137556
rect 544804 137544 544810 137556
rect 545942 137544 545948 137556
rect 544804 137516 545948 137544
rect 544804 137504 544810 137516
rect 545942 137504 545948 137516
rect 546000 137504 546006 137556
rect 541986 137368 541992 137420
rect 542044 137408 542050 137420
rect 544746 137408 544752 137420
rect 542044 137380 544752 137408
rect 542044 137368 542050 137380
rect 544746 137368 544752 137380
rect 544804 137368 544810 137420
rect 540422 137300 540428 137352
rect 540480 137340 540486 137352
rect 540974 137340 540980 137352
rect 540480 137312 540980 137340
rect 540480 137300 540486 137312
rect 540974 137300 540980 137312
rect 541032 137300 541038 137352
rect 542814 137300 542820 137352
rect 542872 137340 542878 137352
rect 544654 137340 544660 137352
rect 542872 137312 544660 137340
rect 542872 137300 542878 137312
rect 544654 137300 544660 137312
rect 544712 137300 544718 137352
rect 558362 137300 558368 137352
rect 558420 137340 558426 137352
rect 559006 137340 559012 137352
rect 558420 137312 559012 137340
rect 558420 137300 558426 137312
rect 559006 137300 559012 137312
rect 559064 137300 559070 137352
rect 540238 137232 540244 137284
rect 540296 137272 540302 137284
rect 549806 137272 549812 137284
rect 540296 137244 549812 137272
rect 540296 137232 540302 137244
rect 549806 137232 549812 137244
rect 549864 137232 549870 137284
rect 51442 136552 51448 136604
rect 51500 136592 51506 136604
rect 53190 136592 53196 136604
rect 51500 136564 53196 136592
rect 51500 136552 51506 136564
rect 53190 136552 53196 136564
rect 53248 136552 53254 136604
rect 55122 136552 55128 136604
rect 55180 136592 55186 136604
rect 55858 136592 55864 136604
rect 55180 136564 55864 136592
rect 55180 136552 55186 136564
rect 55858 136552 55864 136564
rect 55916 136552 55922 136604
rect 543550 136552 543556 136604
rect 543608 136592 543614 136604
rect 572714 136592 572720 136604
rect 543608 136564 572720 136592
rect 543608 136552 543614 136564
rect 572714 136552 572720 136564
rect 572772 136552 572778 136604
rect 55766 136484 55772 136536
rect 55824 136524 55830 136536
rect 59630 136524 59636 136536
rect 55824 136496 59636 136524
rect 55824 136484 55830 136496
rect 59630 136484 59636 136496
rect 59688 136484 59694 136536
rect 543642 136484 543648 136536
rect 543700 136524 543706 136536
rect 564710 136524 564716 136536
rect 543700 136496 564716 136524
rect 543700 136484 543706 136496
rect 564710 136484 564716 136496
rect 564768 136484 564774 136536
rect 50982 136144 50988 136196
rect 51040 136184 51046 136196
rect 53006 136184 53012 136196
rect 51040 136156 53012 136184
rect 51040 136144 51046 136156
rect 53006 136144 53012 136156
rect 53064 136144 53070 136196
rect 54110 135872 54116 135924
rect 54168 135912 54174 135924
rect 59446 135912 59452 135924
rect 54168 135884 59452 135912
rect 54168 135872 54174 135884
rect 59446 135872 59452 135884
rect 59504 135872 59510 135924
rect 549438 135872 549444 135924
rect 549496 135912 549502 135924
rect 558178 135912 558184 135924
rect 549496 135884 558184 135912
rect 549496 135872 549502 135884
rect 558178 135872 558184 135884
rect 558236 135872 558242 135924
rect 543642 135396 543648 135448
rect 543700 135436 543706 135448
rect 546494 135436 546500 135448
rect 543700 135408 546500 135436
rect 543700 135396 543706 135408
rect 546494 135396 546500 135408
rect 546552 135396 546558 135448
rect 52362 135328 52368 135380
rect 52420 135368 52426 135380
rect 52914 135368 52920 135380
rect 52420 135340 52920 135368
rect 52420 135328 52426 135340
rect 52914 135328 52920 135340
rect 52972 135328 52978 135380
rect 545022 135260 545028 135312
rect 545080 135300 545086 135312
rect 549438 135300 549444 135312
rect 545080 135272 549444 135300
rect 545080 135260 545086 135272
rect 549438 135260 549444 135272
rect 549496 135260 549502 135312
rect 24670 135192 24676 135244
rect 24728 135232 24734 135244
rect 57882 135232 57888 135244
rect 24728 135204 57888 135232
rect 24728 135192 24734 135204
rect 57882 135192 57888 135204
rect 57940 135192 57946 135244
rect 543550 135192 543556 135244
rect 543608 135232 543614 135244
rect 568574 135232 568580 135244
rect 543608 135204 568580 135232
rect 543608 135192 543614 135204
rect 568574 135192 568580 135204
rect 568632 135192 568638 135244
rect 546034 135124 546040 135176
rect 546092 135164 546098 135176
rect 549254 135164 549260 135176
rect 546092 135136 549260 135164
rect 546092 135124 546098 135136
rect 549254 135124 549260 135136
rect 549312 135124 549318 135176
rect 58894 134716 58900 134768
rect 58952 134756 58958 134768
rect 59078 134756 59084 134768
rect 58952 134728 59084 134756
rect 58952 134716 58958 134728
rect 59078 134716 59084 134728
rect 59136 134716 59142 134768
rect 545114 133940 545120 133952
rect 542188 133912 545120 133940
rect 25866 133832 25872 133884
rect 25924 133872 25930 133884
rect 57882 133872 57888 133884
rect 25924 133844 57888 133872
rect 25924 133832 25930 133844
rect 57882 133832 57888 133844
rect 57940 133832 57946 133884
rect 542188 133736 542216 133912
rect 545114 133900 545120 133912
rect 545172 133900 545178 133952
rect 542262 133832 542268 133884
rect 542320 133872 542326 133884
rect 542538 133872 542544 133884
rect 542320 133844 542544 133872
rect 542320 133832 542326 133844
rect 542538 133832 542544 133844
rect 542596 133832 542602 133884
rect 543274 133832 543280 133884
rect 543332 133872 543338 133884
rect 545574 133872 545580 133884
rect 543332 133844 545580 133872
rect 543332 133832 543338 133844
rect 545574 133832 545580 133844
rect 545632 133832 545638 133884
rect 554222 133832 554228 133884
rect 554280 133872 554286 133884
rect 556982 133872 556988 133884
rect 554280 133844 556988 133872
rect 554280 133832 554286 133844
rect 556982 133832 556988 133844
rect 557040 133832 557046 133884
rect 542262 133736 542268 133748
rect 542188 133708 542268 133736
rect 542262 133696 542268 133708
rect 542320 133696 542326 133748
rect 546402 133152 546408 133204
rect 546460 133192 546466 133204
rect 548518 133192 548524 133204
rect 546460 133164 548524 133192
rect 546460 133152 546466 133164
rect 548518 133152 548524 133164
rect 548576 133152 548582 133204
rect 545942 133084 545948 133136
rect 546000 133124 546006 133136
rect 552014 133124 552020 133136
rect 546000 133096 552020 133124
rect 546000 133084 546006 133096
rect 552014 133084 552020 133096
rect 552072 133084 552078 133136
rect 546402 133016 546408 133068
rect 546460 133056 546466 133068
rect 547966 133056 547972 133068
rect 546460 133028 547972 133056
rect 546460 133016 546466 133028
rect 547966 133016 547972 133028
rect 548024 133016 548030 133068
rect 545850 132744 545856 132796
rect 545908 132784 545914 132796
rect 552106 132784 552112 132796
rect 545908 132756 552112 132784
rect 545908 132744 545914 132756
rect 552106 132744 552112 132756
rect 552164 132744 552170 132796
rect 57054 132676 57060 132728
rect 57112 132716 57118 132728
rect 57882 132716 57888 132728
rect 57112 132688 57888 132716
rect 57112 132676 57118 132688
rect 57882 132676 57888 132688
rect 57940 132676 57946 132728
rect 56502 132472 56508 132524
rect 56560 132512 56566 132524
rect 57146 132512 57152 132524
rect 56560 132484 57152 132512
rect 56560 132472 56566 132484
rect 57146 132472 57152 132484
rect 57204 132472 57210 132524
rect 32582 132404 32588 132456
rect 32640 132444 32646 132456
rect 57054 132444 57060 132456
rect 32640 132416 57060 132444
rect 32640 132404 32646 132416
rect 57054 132404 57060 132416
rect 57112 132404 57118 132456
rect 543550 132404 543556 132456
rect 543608 132444 543614 132456
rect 578786 132444 578792 132456
rect 543608 132416 578792 132444
rect 543608 132404 543614 132416
rect 578786 132404 578792 132416
rect 578844 132404 578850 132456
rect 56502 132336 56508 132388
rect 56560 132376 56566 132388
rect 59262 132376 59268 132388
rect 56560 132348 59268 132376
rect 56560 132336 56566 132348
rect 59262 132336 59268 132348
rect 59320 132336 59326 132388
rect 546126 132336 546132 132388
rect 546184 132376 546190 132388
rect 548978 132376 548984 132388
rect 546184 132348 548984 132376
rect 546184 132336 546190 132348
rect 548978 132336 548984 132348
rect 549036 132336 549042 132388
rect 543642 131452 543648 131504
rect 543700 131492 543706 131504
rect 548058 131492 548064 131504
rect 543700 131464 548064 131492
rect 543700 131452 543706 131464
rect 548058 131452 548064 131464
rect 548116 131452 548122 131504
rect 541710 131248 541716 131300
rect 541768 131288 541774 131300
rect 548242 131288 548248 131300
rect 541768 131260 548248 131288
rect 541768 131248 541774 131260
rect 548242 131248 548248 131260
rect 548300 131248 548306 131300
rect 541986 131180 541992 131232
rect 542044 131220 542050 131232
rect 546954 131220 546960 131232
rect 542044 131192 546960 131220
rect 542044 131180 542050 131192
rect 546954 131180 546960 131192
rect 547012 131180 547018 131232
rect 53374 131112 53380 131164
rect 53432 131152 53438 131164
rect 54570 131152 54576 131164
rect 53432 131124 54576 131152
rect 53432 131112 53438 131124
rect 54570 131112 54576 131124
rect 54628 131112 54634 131164
rect 58526 131112 58532 131164
rect 58584 131152 58590 131164
rect 59630 131152 59636 131164
rect 58584 131124 59636 131152
rect 58584 131112 58590 131124
rect 59630 131112 59636 131124
rect 59688 131112 59694 131164
rect 540974 131112 540980 131164
rect 541032 131112 541038 131164
rect 542170 131112 542176 131164
rect 542228 131152 542234 131164
rect 543734 131152 543740 131164
rect 542228 131124 543740 131152
rect 542228 131112 542234 131124
rect 543734 131112 543740 131124
rect 543792 131112 543798 131164
rect 540790 131044 540796 131096
rect 540848 131084 540854 131096
rect 540992 131084 541020 131112
rect 540848 131056 541020 131084
rect 540848 131044 540854 131056
rect 543550 131044 543556 131096
rect 543608 131084 543614 131096
rect 578234 131084 578240 131096
rect 543608 131056 578240 131084
rect 543608 131044 543614 131056
rect 578234 131044 578240 131056
rect 578292 131044 578298 131096
rect 545942 130976 545948 131028
rect 546000 131016 546006 131028
rect 546586 131016 546592 131028
rect 546000 130988 546592 131016
rect 546000 130976 546006 130988
rect 546586 130976 546592 130988
rect 546644 130976 546650 131028
rect 548610 130976 548616 131028
rect 548668 131016 548674 131028
rect 551278 131016 551284 131028
rect 548668 130988 551284 131016
rect 548668 130976 548674 130988
rect 551278 130976 551284 130988
rect 551336 130976 551342 131028
rect 544746 130908 544752 130960
rect 544804 130948 544810 130960
rect 545022 130948 545028 130960
rect 544804 130920 545028 130948
rect 544804 130908 544810 130920
rect 545022 130908 545028 130920
rect 545080 130908 545086 130960
rect 540698 130840 540704 130892
rect 540756 130880 540762 130892
rect 546954 130880 546960 130892
rect 540756 130852 546960 130880
rect 540756 130840 540762 130852
rect 546954 130840 546960 130852
rect 547012 130840 547018 130892
rect 544654 130772 544660 130824
rect 544712 130812 544718 130824
rect 547230 130812 547236 130824
rect 544712 130784 547236 130812
rect 544712 130772 544718 130784
rect 547230 130772 547236 130784
rect 547288 130772 547294 130824
rect 544470 130024 544476 130076
rect 544528 130064 544534 130076
rect 545390 130064 545396 130076
rect 544528 130036 545396 130064
rect 544528 130024 544534 130036
rect 545390 130024 545396 130036
rect 545448 130024 545454 130076
rect 54570 129684 54576 129736
rect 54628 129724 54634 129736
rect 55858 129724 55864 129736
rect 54628 129696 55864 129724
rect 54628 129684 54634 129696
rect 55858 129684 55864 129696
rect 55916 129684 55922 129736
rect 551462 129684 551468 129736
rect 551520 129724 551526 129736
rect 552106 129724 552112 129736
rect 551520 129696 552112 129724
rect 551520 129684 551526 129696
rect 552106 129684 552112 129696
rect 552164 129684 552170 129736
rect 54846 129616 54852 129668
rect 54904 129656 54910 129668
rect 57054 129656 57060 129668
rect 54904 129628 57060 129656
rect 54904 129616 54910 129628
rect 57054 129616 57060 129628
rect 57112 129616 57118 129668
rect 551278 129616 551284 129668
rect 551336 129656 551342 129668
rect 552014 129656 552020 129668
rect 551336 129628 552020 129656
rect 551336 129616 551342 129628
rect 552014 129616 552020 129628
rect 552072 129616 552078 129668
rect 55122 129548 55128 129600
rect 55180 129588 55186 129600
rect 56962 129588 56968 129600
rect 55180 129560 56968 129588
rect 55180 129548 55186 129560
rect 56962 129548 56968 129560
rect 57020 129548 57026 129600
rect 56410 128324 56416 128376
rect 56468 128364 56474 128376
rect 56870 128364 56876 128376
rect 56468 128336 56876 128364
rect 56468 128324 56474 128336
rect 56870 128324 56876 128336
rect 56928 128324 56934 128376
rect 39482 128256 39488 128308
rect 39540 128296 39546 128308
rect 57238 128296 57244 128308
rect 39540 128268 57244 128296
rect 39540 128256 39546 128268
rect 57238 128256 57244 128268
rect 57296 128256 57302 128308
rect 543550 128256 543556 128308
rect 543608 128296 543614 128308
rect 563054 128296 563060 128308
rect 543608 128268 563060 128296
rect 543608 128256 543614 128268
rect 563054 128256 563060 128268
rect 563112 128256 563118 128308
rect 542078 128188 542084 128240
rect 542136 128228 542142 128240
rect 544010 128228 544016 128240
rect 542136 128200 544016 128228
rect 542136 128188 542142 128200
rect 544010 128188 544016 128200
rect 544068 128188 544074 128240
rect 50982 127780 50988 127832
rect 51040 127820 51046 127832
rect 54386 127820 54392 127832
rect 51040 127792 54392 127820
rect 51040 127780 51046 127792
rect 54386 127780 54392 127792
rect 54444 127780 54450 127832
rect 53742 127576 53748 127628
rect 53800 127616 53806 127628
rect 58526 127616 58532 127628
rect 53800 127588 58532 127616
rect 53800 127576 53806 127588
rect 58526 127576 58532 127588
rect 58584 127576 58590 127628
rect 540974 127576 540980 127628
rect 541032 127616 541038 127628
rect 545022 127616 545028 127628
rect 541032 127588 545028 127616
rect 541032 127576 541038 127588
rect 545022 127576 545028 127588
rect 545080 127576 545086 127628
rect 49602 126896 49608 126948
rect 49660 126936 49666 126948
rect 50338 126936 50344 126948
rect 49660 126908 50344 126936
rect 49660 126896 49666 126908
rect 50338 126896 50344 126908
rect 50396 126896 50402 126948
rect 54754 126896 54760 126948
rect 54812 126936 54818 126948
rect 57238 126936 57244 126948
rect 54812 126908 57244 126936
rect 54812 126896 54818 126908
rect 57238 126896 57244 126908
rect 57296 126896 57302 126948
rect 58986 126896 58992 126948
rect 59044 126936 59050 126948
rect 59354 126936 59360 126948
rect 59044 126908 59360 126936
rect 59044 126896 59050 126908
rect 59354 126896 59360 126908
rect 59412 126896 59418 126948
rect 541894 126896 541900 126948
rect 541952 126936 541958 126948
rect 543182 126936 543188 126948
rect 541952 126908 543188 126936
rect 541952 126896 541958 126908
rect 543182 126896 543188 126908
rect 543240 126896 543246 126948
rect 541618 126828 541624 126880
rect 541676 126868 541682 126880
rect 543458 126868 543464 126880
rect 541676 126840 543464 126868
rect 541676 126828 541682 126840
rect 543458 126828 543464 126840
rect 543516 126828 543522 126880
rect 53742 126216 53748 126268
rect 53800 126256 53806 126268
rect 57146 126256 57152 126268
rect 53800 126228 57152 126256
rect 53800 126216 53806 126228
rect 57146 126216 57152 126228
rect 57204 126216 57210 126268
rect 540330 126216 540336 126268
rect 540388 126256 540394 126268
rect 556890 126256 556896 126268
rect 540388 126228 556896 126256
rect 540388 126216 540394 126228
rect 556890 126216 556896 126228
rect 556948 126216 556954 126268
rect 542262 125672 542268 125724
rect 542320 125712 542326 125724
rect 544562 125712 544568 125724
rect 542320 125684 544568 125712
rect 542320 125672 542326 125684
rect 544562 125672 544568 125684
rect 544620 125672 544626 125724
rect 540790 125604 540796 125656
rect 540848 125644 540854 125656
rect 541986 125644 541992 125656
rect 540848 125616 541992 125644
rect 540848 125604 540854 125616
rect 541986 125604 541992 125616
rect 542044 125604 542050 125656
rect 543734 125644 543740 125656
rect 543476 125616 543740 125644
rect 28902 125536 28908 125588
rect 28960 125576 28966 125588
rect 57238 125576 57244 125588
rect 28960 125548 57244 125576
rect 28960 125536 28966 125548
rect 57238 125536 57244 125548
rect 57296 125536 57302 125588
rect 542078 125536 542084 125588
rect 542136 125576 542142 125588
rect 543476 125576 543504 125616
rect 543734 125604 543740 125616
rect 543792 125604 543798 125656
rect 542136 125548 543504 125576
rect 542136 125536 542142 125548
rect 543550 125536 543556 125588
rect 543608 125576 543614 125588
rect 562318 125576 562324 125588
rect 543608 125548 562324 125576
rect 543608 125536 543614 125548
rect 562318 125536 562324 125548
rect 562376 125536 562382 125588
rect 52362 125468 52368 125520
rect 52420 125508 52426 125520
rect 55030 125508 55036 125520
rect 52420 125480 55036 125508
rect 52420 125468 52426 125480
rect 55030 125468 55036 125480
rect 55088 125468 55094 125520
rect 59262 124448 59268 124500
rect 59320 124488 59326 124500
rect 59814 124488 59820 124500
rect 59320 124460 59820 124488
rect 59320 124448 59326 124460
rect 59814 124448 59820 124460
rect 59872 124448 59878 124500
rect 22830 124108 22836 124160
rect 22888 124148 22894 124160
rect 57238 124148 57244 124160
rect 22888 124120 57244 124148
rect 22888 124108 22894 124120
rect 57238 124108 57244 124120
rect 57296 124108 57302 124160
rect 58894 124108 58900 124160
rect 58952 124148 58958 124160
rect 59446 124148 59452 124160
rect 58952 124120 59452 124148
rect 58952 124108 58958 124120
rect 59446 124108 59452 124120
rect 59504 124108 59510 124160
rect 544378 124108 544384 124160
rect 544436 124148 544442 124160
rect 545390 124148 545396 124160
rect 544436 124120 545396 124148
rect 544436 124108 544442 124120
rect 545390 124108 545396 124120
rect 545448 124108 545454 124160
rect 562318 124108 562324 124160
rect 562376 124148 562382 124160
rect 565262 124148 565268 124160
rect 562376 124120 565268 124148
rect 562376 124108 562382 124120
rect 565262 124108 565268 124120
rect 565320 124108 565326 124160
rect 56502 124040 56508 124092
rect 56560 124080 56566 124092
rect 58710 124080 58716 124092
rect 56560 124052 58716 124080
rect 56560 124040 56566 124052
rect 58710 124040 58716 124052
rect 58768 124040 58774 124092
rect 543366 123360 543372 123412
rect 543424 123400 543430 123412
rect 552474 123400 552480 123412
rect 543424 123372 552480 123400
rect 543424 123360 543430 123372
rect 552474 123360 552480 123372
rect 552532 123360 552538 123412
rect 55122 122884 55128 122936
rect 55180 122924 55186 122936
rect 55180 122884 55214 122924
rect 55186 122856 55214 122884
rect 55306 122856 55312 122868
rect 55186 122828 55312 122856
rect 55306 122816 55312 122828
rect 55364 122816 55370 122868
rect 544102 122816 544108 122868
rect 544160 122856 544166 122868
rect 546402 122856 546408 122868
rect 544160 122828 546408 122856
rect 544160 122816 544166 122828
rect 546402 122816 546408 122828
rect 546460 122816 546466 122868
rect 543550 122748 543556 122800
rect 543608 122788 543614 122800
rect 574922 122788 574928 122800
rect 543608 122760 574928 122788
rect 543608 122748 543614 122760
rect 574922 122748 574928 122760
rect 574980 122748 574986 122800
rect 546494 122680 546500 122732
rect 546552 122720 546558 122732
rect 549070 122720 549076 122732
rect 546552 122692 549076 122720
rect 546552 122680 546558 122692
rect 549070 122680 549076 122692
rect 549128 122680 549134 122732
rect 57146 121660 57152 121712
rect 57204 121700 57210 121712
rect 57882 121700 57888 121712
rect 57204 121672 57888 121700
rect 57204 121660 57210 121672
rect 57882 121660 57888 121672
rect 57940 121660 57946 121712
rect 58986 121592 58992 121644
rect 59044 121632 59050 121644
rect 59354 121632 59360 121644
rect 59044 121604 59360 121632
rect 59044 121592 59050 121604
rect 59354 121592 59360 121604
rect 59412 121592 59418 121644
rect 57330 121524 57336 121576
rect 57388 121564 57394 121576
rect 57882 121564 57888 121576
rect 57388 121536 57888 121564
rect 57388 121524 57394 121536
rect 57882 121524 57888 121536
rect 57940 121524 57946 121576
rect 545114 121456 545120 121508
rect 545172 121496 545178 121508
rect 548518 121496 548524 121508
rect 545172 121468 548524 121496
rect 545172 121456 545178 121468
rect 548518 121456 548524 121468
rect 548576 121456 548582 121508
rect 36170 121388 36176 121440
rect 36228 121428 36234 121440
rect 57330 121428 57336 121440
rect 36228 121400 57336 121428
rect 36228 121388 36234 121400
rect 57330 121388 57336 121400
rect 57388 121388 57394 121440
rect 543550 121388 543556 121440
rect 543608 121428 543614 121440
rect 560846 121428 560852 121440
rect 543608 121400 560852 121428
rect 543608 121388 543614 121400
rect 560846 121388 560852 121400
rect 560904 121388 560910 121440
rect 543182 121252 543188 121304
rect 543240 121292 543246 121304
rect 547874 121292 547880 121304
rect 543240 121264 547880 121292
rect 543240 121252 543246 121264
rect 547874 121252 547880 121264
rect 547932 121252 547938 121304
rect 54570 120708 54576 120760
rect 54628 120748 54634 120760
rect 55214 120748 55220 120760
rect 54628 120720 55220 120748
rect 54628 120708 54634 120720
rect 55214 120708 55220 120720
rect 55272 120708 55278 120760
rect 546034 120368 546040 120420
rect 546092 120408 546098 120420
rect 549254 120408 549260 120420
rect 546092 120380 549260 120408
rect 546092 120368 546098 120380
rect 549254 120368 549260 120380
rect 549312 120368 549318 120420
rect 59170 120164 59176 120216
rect 59228 120204 59234 120216
rect 59814 120204 59820 120216
rect 59228 120176 59820 120204
rect 59228 120164 59234 120176
rect 59814 120164 59820 120176
rect 59872 120164 59878 120216
rect 59262 120096 59268 120148
rect 59320 120136 59326 120148
rect 59446 120136 59452 120148
rect 59320 120108 59452 120136
rect 59320 120096 59326 120108
rect 59446 120096 59452 120108
rect 59504 120096 59510 120148
rect 540882 120096 540888 120148
rect 540940 120136 540946 120148
rect 543090 120136 543096 120148
rect 540940 120108 543096 120136
rect 540940 120096 540946 120108
rect 543090 120096 543096 120108
rect 543148 120096 543154 120148
rect 549990 120096 549996 120148
rect 550048 120136 550054 120148
rect 552106 120136 552112 120148
rect 550048 120108 552112 120136
rect 550048 120096 550054 120108
rect 552106 120096 552112 120108
rect 552164 120096 552170 120148
rect 40586 119960 40592 120012
rect 40644 120000 40650 120012
rect 57330 120000 57336 120012
rect 40644 119972 57336 120000
rect 40644 119960 40650 119972
rect 57330 119960 57336 119972
rect 57388 119960 57394 120012
rect 54754 119348 54760 119400
rect 54812 119388 54818 119400
rect 59630 119388 59636 119400
rect 54812 119360 59636 119388
rect 54812 119348 54818 119360
rect 59630 119348 59636 119360
rect 59688 119348 59694 119400
rect 548518 119348 548524 119400
rect 548576 119388 548582 119400
rect 565814 119388 565820 119400
rect 548576 119360 565820 119388
rect 548576 119348 548582 119360
rect 565814 119348 565820 119360
rect 565872 119348 565878 119400
rect 58710 118668 58716 118720
rect 58768 118708 58774 118720
rect 59538 118708 59544 118720
rect 58768 118680 59544 118708
rect 58768 118668 58774 118680
rect 59538 118668 59544 118680
rect 59596 118668 59602 118720
rect 54110 118600 54116 118652
rect 54168 118640 54174 118652
rect 56594 118640 56600 118652
rect 54168 118612 56600 118640
rect 54168 118600 54174 118612
rect 56594 118600 56600 118612
rect 56652 118600 56658 118652
rect 56502 118124 56508 118176
rect 56560 118164 56566 118176
rect 59722 118164 59728 118176
rect 56560 118136 59728 118164
rect 56560 118124 56566 118136
rect 59722 118124 59728 118136
rect 59780 118124 59786 118176
rect 57146 117988 57152 118040
rect 57204 118028 57210 118040
rect 59722 118028 59728 118040
rect 57204 118000 59728 118028
rect 57204 117988 57210 118000
rect 59722 117988 59728 118000
rect 59780 117988 59786 118040
rect 59170 117920 59176 117972
rect 59228 117960 59234 117972
rect 59354 117960 59360 117972
rect 59228 117932 59360 117960
rect 59228 117920 59234 117932
rect 59354 117920 59360 117932
rect 59412 117920 59418 117972
rect 540698 117512 540704 117564
rect 540756 117552 540762 117564
rect 546954 117552 546960 117564
rect 540756 117524 546960 117552
rect 540756 117512 540762 117524
rect 546954 117512 546960 117524
rect 547012 117512 547018 117564
rect 546126 117308 546132 117360
rect 546184 117348 546190 117360
rect 546586 117348 546592 117360
rect 546184 117320 546592 117348
rect 546184 117308 546190 117320
rect 546586 117308 546592 117320
rect 546644 117308 546650 117360
rect 22922 117240 22928 117292
rect 22980 117280 22986 117292
rect 57330 117280 57336 117292
rect 22980 117252 57336 117280
rect 22980 117240 22986 117252
rect 57330 117240 57336 117252
rect 57388 117240 57394 117292
rect 543550 117240 543556 117292
rect 543608 117280 543614 117292
rect 568022 117280 568028 117292
rect 543608 117252 568028 117280
rect 543608 117240 543614 117252
rect 568022 117240 568028 117252
rect 568080 117240 568086 117292
rect 545022 117172 545028 117224
rect 545080 117212 545086 117224
rect 546586 117212 546592 117224
rect 545080 117184 546592 117212
rect 545080 117172 545086 117184
rect 546586 117172 546592 117184
rect 546644 117172 546650 117224
rect 549070 117172 549076 117224
rect 549128 117212 549134 117224
rect 552106 117212 552112 117224
rect 549128 117184 552112 117212
rect 549128 117172 549134 117184
rect 552106 117172 552112 117184
rect 552164 117172 552170 117224
rect 547782 116628 547788 116680
rect 547840 116668 547846 116680
rect 548794 116668 548800 116680
rect 547840 116640 548800 116668
rect 547840 116628 547846 116640
rect 548794 116628 548800 116640
rect 548852 116628 548858 116680
rect 541802 116560 541808 116612
rect 541860 116600 541866 116612
rect 552198 116600 552204 116612
rect 541860 116572 552204 116600
rect 541860 116560 541866 116572
rect 552198 116560 552204 116572
rect 552256 116560 552262 116612
rect 54846 116424 54852 116476
rect 54904 116464 54910 116476
rect 56870 116464 56876 116476
rect 54904 116436 56876 116464
rect 54904 116424 54910 116436
rect 56870 116424 56876 116436
rect 56928 116424 56934 116476
rect 43162 115880 43168 115932
rect 43220 115920 43226 115932
rect 57330 115920 57336 115932
rect 43220 115892 57336 115920
rect 43220 115880 43226 115892
rect 57330 115880 57336 115892
rect 57388 115880 57394 115932
rect 541802 115880 541808 115932
rect 541860 115920 541866 115932
rect 542814 115920 542820 115932
rect 541860 115892 542820 115920
rect 541860 115880 541866 115892
rect 542814 115880 542820 115892
rect 542872 115880 542878 115932
rect 545758 115880 545764 115932
rect 545816 115920 545822 115932
rect 547230 115920 547236 115932
rect 545816 115892 547236 115920
rect 545816 115880 545822 115892
rect 547230 115880 547236 115892
rect 547288 115880 547294 115932
rect 558270 115920 558276 115932
rect 547846 115892 558276 115920
rect 543550 115812 543556 115864
rect 543608 115852 543614 115864
rect 547846 115852 547874 115892
rect 558270 115880 558276 115892
rect 558328 115880 558334 115932
rect 543608 115824 547874 115852
rect 543608 115812 543614 115824
rect 541986 115472 541992 115524
rect 542044 115512 542050 115524
rect 548794 115512 548800 115524
rect 542044 115484 548800 115512
rect 542044 115472 542050 115484
rect 548794 115472 548800 115484
rect 548852 115472 548858 115524
rect 541434 115404 541440 115456
rect 541492 115444 541498 115456
rect 542354 115444 542360 115456
rect 541492 115416 542360 115444
rect 541492 115404 541498 115416
rect 542354 115404 542360 115416
rect 542412 115404 542418 115456
rect 24302 115200 24308 115252
rect 24360 115240 24366 115252
rect 57146 115240 57152 115252
rect 24360 115212 57152 115240
rect 24360 115200 24366 115212
rect 57146 115200 57152 115212
rect 57204 115200 57210 115252
rect 544378 114996 544384 115048
rect 544436 115036 544442 115048
rect 545482 115036 545488 115048
rect 544436 115008 545488 115036
rect 544436 114996 544442 115008
rect 545482 114996 545488 115008
rect 545540 114996 545546 115048
rect 547782 114860 547788 114912
rect 547840 114900 547846 114912
rect 547966 114900 547972 114912
rect 547840 114872 547972 114900
rect 547840 114860 547846 114872
rect 547966 114860 547972 114872
rect 548024 114860 548030 114912
rect 545114 114588 545120 114640
rect 545172 114628 545178 114640
rect 547874 114628 547880 114640
rect 545172 114600 547880 114628
rect 545172 114588 545178 114600
rect 547874 114588 547880 114600
rect 547932 114588 547938 114640
rect 547322 114520 547328 114572
rect 547380 114560 547386 114572
rect 548058 114560 548064 114572
rect 547380 114532 548064 114560
rect 547380 114520 547386 114532
rect 548058 114520 548064 114532
rect 548116 114520 548122 114572
rect 542078 114452 542084 114504
rect 542136 114492 542142 114504
rect 542354 114492 542360 114504
rect 542136 114464 542360 114492
rect 542136 114452 542142 114464
rect 542354 114452 542360 114464
rect 542412 114452 542418 114504
rect 543550 114452 543556 114504
rect 543608 114492 543614 114504
rect 572162 114492 572168 114504
rect 543608 114464 572168 114492
rect 543608 114452 543614 114464
rect 572162 114452 572168 114464
rect 572220 114452 572226 114504
rect 543642 114384 543648 114436
rect 543700 114424 543706 114436
rect 559558 114424 559564 114436
rect 543700 114396 559564 114424
rect 543700 114384 543706 114396
rect 559558 114384 559564 114396
rect 559616 114384 559622 114436
rect 540514 114316 540520 114368
rect 540572 114356 540578 114368
rect 545482 114356 545488 114368
rect 540572 114328 545488 114356
rect 540572 114316 540578 114328
rect 545482 114316 545488 114328
rect 545540 114316 545546 114368
rect 540606 113976 540612 114028
rect 540664 114016 540670 114028
rect 546126 114016 546132 114028
rect 540664 113988 546132 114016
rect 540664 113976 540670 113988
rect 546126 113976 546132 113988
rect 546184 113976 546190 114028
rect 54662 113772 54668 113824
rect 54720 113812 54726 113824
rect 58710 113812 58716 113824
rect 54720 113784 58716 113812
rect 54720 113772 54726 113784
rect 58710 113772 58716 113784
rect 58768 113772 58774 113824
rect 542998 113500 543004 113552
rect 543056 113540 543062 113552
rect 547874 113540 547880 113552
rect 543056 113512 547880 113540
rect 543056 113500 543062 113512
rect 547874 113500 547880 113512
rect 547932 113500 547938 113552
rect 545114 113200 545120 113212
rect 542280 113172 545120 113200
rect 542280 113144 542308 113172
rect 545114 113160 545120 113172
rect 545172 113160 545178 113212
rect 547966 113160 547972 113212
rect 548024 113160 548030 113212
rect 557074 113160 557080 113212
rect 557132 113200 557138 113212
rect 558270 113200 558276 113212
rect 557132 113172 558276 113200
rect 557132 113160 557138 113172
rect 558270 113160 558276 113172
rect 558328 113160 558334 113212
rect 542262 113092 542268 113144
rect 542320 113092 542326 113144
rect 547984 113132 548012 113160
rect 549898 113132 549904 113144
rect 547984 113104 549904 113132
rect 549898 113092 549904 113104
rect 549956 113092 549962 113144
rect 576210 113092 576216 113144
rect 576268 113132 576274 113144
rect 580442 113132 580448 113144
rect 576268 113104 580448 113132
rect 576268 113092 576274 113104
rect 580442 113092 580448 113104
rect 580500 113092 580506 113144
rect 48866 112888 48872 112940
rect 48924 112928 48930 112940
rect 57330 112928 57336 112940
rect 48924 112900 57336 112928
rect 48924 112888 48930 112900
rect 57330 112888 57336 112900
rect 57388 112888 57394 112940
rect 59630 112072 59636 112124
rect 59688 112112 59694 112124
rect 59814 112112 59820 112124
rect 59688 112084 59820 112112
rect 59688 112072 59694 112084
rect 59814 112072 59820 112084
rect 59872 112072 59878 112124
rect 59262 111936 59268 111988
rect 59320 111976 59326 111988
rect 59814 111976 59820 111988
rect 59320 111948 59820 111976
rect 59320 111936 59326 111948
rect 59814 111936 59820 111948
rect 59872 111936 59878 111988
rect 558178 111868 558184 111920
rect 558236 111908 558242 111920
rect 565814 111908 565820 111920
rect 558236 111880 565820 111908
rect 558236 111868 558242 111880
rect 565814 111868 565820 111880
rect 565872 111868 565878 111920
rect 58894 111800 58900 111852
rect 58952 111840 58958 111852
rect 59538 111840 59544 111852
rect 58952 111812 59544 111840
rect 58952 111800 58958 111812
rect 59538 111800 59544 111812
rect 59596 111800 59602 111852
rect 546402 111800 546408 111852
rect 546460 111840 546466 111852
rect 549990 111840 549996 111852
rect 546460 111812 549996 111840
rect 546460 111800 546466 111812
rect 549990 111800 549996 111812
rect 550048 111800 550054 111852
rect 556982 111052 556988 111104
rect 557040 111092 557046 111104
rect 561674 111092 561680 111104
rect 557040 111064 561680 111092
rect 557040 111052 557046 111064
rect 561674 111052 561680 111064
rect 561732 111052 561738 111104
rect 543090 110576 543096 110628
rect 543148 110616 543154 110628
rect 543826 110616 543832 110628
rect 543148 110588 543832 110616
rect 543148 110576 543154 110588
rect 543826 110576 543832 110588
rect 543884 110576 543890 110628
rect 540882 110508 540888 110560
rect 540940 110548 540946 110560
rect 543366 110548 543372 110560
rect 540940 110520 543372 110548
rect 540940 110508 540946 110520
rect 543366 110508 543372 110520
rect 543424 110508 543430 110560
rect 56502 110440 56508 110492
rect 56560 110480 56566 110492
rect 59630 110480 59636 110492
rect 56560 110452 59636 110480
rect 56560 110440 56566 110452
rect 59630 110440 59636 110452
rect 59688 110440 59694 110492
rect 542998 110440 543004 110492
rect 543056 110480 543062 110492
rect 544010 110480 544016 110492
rect 543056 110452 544016 110480
rect 543056 110440 543062 110452
rect 544010 110440 544016 110452
rect 544068 110440 544074 110492
rect 543550 110372 543556 110424
rect 543608 110412 543614 110424
rect 551370 110412 551376 110424
rect 543608 110384 551376 110412
rect 543608 110372 543614 110384
rect 551370 110372 551376 110384
rect 551428 110372 551434 110424
rect 543182 109692 543188 109744
rect 543240 109732 543246 109744
rect 550726 109732 550732 109744
rect 543240 109704 550732 109732
rect 543240 109692 543246 109704
rect 550726 109692 550732 109704
rect 550784 109692 550790 109744
rect 43254 108944 43260 108996
rect 43312 108984 43318 108996
rect 57422 108984 57428 108996
rect 43312 108956 57428 108984
rect 43312 108944 43318 108956
rect 57422 108944 57428 108956
rect 57480 108944 57486 108996
rect 542262 108944 542268 108996
rect 542320 108984 542326 108996
rect 543090 108984 543096 108996
rect 542320 108956 543096 108984
rect 542320 108944 542326 108956
rect 543090 108944 543096 108956
rect 543148 108944 543154 108996
rect 44634 108876 44640 108928
rect 44692 108916 44698 108928
rect 57514 108916 57520 108928
rect 44692 108888 57520 108916
rect 44692 108876 44698 108888
rect 57514 108876 57520 108888
rect 57572 108876 57578 108928
rect 547874 108876 547880 108928
rect 547932 108916 547938 108928
rect 550082 108916 550088 108928
rect 547932 108888 550088 108916
rect 547932 108876 547938 108888
rect 550082 108876 550088 108888
rect 550140 108876 550146 108928
rect 543642 108808 543648 108860
rect 543700 108848 543706 108860
rect 544194 108848 544200 108860
rect 543700 108820 544200 108848
rect 543700 108808 543706 108820
rect 544194 108808 544200 108820
rect 544252 108808 544258 108860
rect 543734 108400 543740 108452
rect 543792 108440 543798 108452
rect 549622 108440 549628 108452
rect 543792 108412 549628 108440
rect 543792 108400 543798 108412
rect 549622 108400 549628 108412
rect 549680 108400 549686 108452
rect 542170 108332 542176 108384
rect 542228 108372 542234 108384
rect 542814 108372 542820 108384
rect 542228 108344 542820 108372
rect 542228 108332 542234 108344
rect 542814 108332 542820 108344
rect 542872 108332 542878 108384
rect 545022 108332 545028 108384
rect 545080 108372 545086 108384
rect 551278 108372 551284 108384
rect 545080 108344 551284 108372
rect 545080 108332 545086 108344
rect 551278 108332 551284 108344
rect 551336 108332 551342 108384
rect 546218 108264 546224 108316
rect 546276 108304 546282 108316
rect 550634 108304 550640 108316
rect 546276 108276 550640 108304
rect 546276 108264 546282 108276
rect 550634 108264 550640 108276
rect 550692 108264 550698 108316
rect 57882 108196 57888 108248
rect 57940 108236 57946 108248
rect 58802 108236 58808 108248
rect 57940 108208 58808 108236
rect 57940 108196 57946 108208
rect 58802 108196 58808 108208
rect 58860 108196 58866 108248
rect 542170 108196 542176 108248
rect 542228 108236 542234 108248
rect 544470 108236 544476 108248
rect 542228 108208 544476 108236
rect 542228 108196 542234 108208
rect 544470 108196 544476 108208
rect 544528 108196 544534 108248
rect 545942 108060 545948 108112
rect 546000 108100 546006 108112
rect 546586 108100 546592 108112
rect 546000 108072 546592 108100
rect 546000 108060 546006 108072
rect 546586 108060 546592 108072
rect 546644 108060 546650 108112
rect 543182 107856 543188 107908
rect 543240 107896 543246 107908
rect 548978 107896 548984 107908
rect 543240 107868 548984 107896
rect 543240 107856 543246 107868
rect 548978 107856 548984 107868
rect 549036 107856 549042 107908
rect 543826 107692 543832 107704
rect 541268 107664 543832 107692
rect 50246 107584 50252 107636
rect 50304 107624 50310 107636
rect 54662 107624 54668 107636
rect 50304 107596 54668 107624
rect 50304 107584 50310 107596
rect 54662 107584 54668 107596
rect 54720 107584 54726 107636
rect 540790 107584 540796 107636
rect 540848 107624 540854 107636
rect 541158 107624 541164 107636
rect 540848 107596 541164 107624
rect 540848 107584 540854 107596
rect 541158 107584 541164 107596
rect 541216 107584 541222 107636
rect 540790 107448 540796 107500
rect 540848 107488 540854 107500
rect 541268 107488 541296 107664
rect 543826 107652 543832 107664
rect 543884 107652 543890 107704
rect 543274 107584 543280 107636
rect 543332 107624 543338 107636
rect 562410 107624 562416 107636
rect 543332 107596 562416 107624
rect 543332 107584 543338 107596
rect 562410 107584 562416 107596
rect 562468 107584 562474 107636
rect 540848 107460 541296 107488
rect 540848 107448 540854 107460
rect 546034 106224 546040 106276
rect 546092 106264 546098 106276
rect 547414 106264 547420 106276
rect 546092 106236 547420 106264
rect 546092 106224 546098 106236
rect 547414 106224 547420 106236
rect 547472 106224 547478 106276
rect 548702 105884 548708 105936
rect 548760 105924 548766 105936
rect 552106 105924 552112 105936
rect 548760 105896 552112 105924
rect 548760 105884 548766 105896
rect 552106 105884 552112 105896
rect 552164 105884 552170 105936
rect 542354 104864 542360 104916
rect 542412 104864 542418 104916
rect 53282 104796 53288 104848
rect 53340 104836 53346 104848
rect 57422 104836 57428 104848
rect 53340 104808 57428 104836
rect 53340 104796 53346 104808
rect 57422 104796 57428 104808
rect 57480 104796 57486 104848
rect 542372 104836 542400 104864
rect 543826 104836 543832 104848
rect 542372 104808 543832 104836
rect 543826 104796 543832 104808
rect 543884 104796 543890 104848
rect 50430 104728 50436 104780
rect 50488 104768 50494 104780
rect 57514 104768 57520 104780
rect 50488 104740 57520 104768
rect 50488 104728 50494 104740
rect 57514 104728 57520 104740
rect 57572 104728 57578 104780
rect 541526 104728 541532 104780
rect 541584 104768 541590 104780
rect 544010 104768 544016 104780
rect 541584 104740 544016 104768
rect 541584 104728 541590 104740
rect 544010 104728 544016 104740
rect 544068 104728 544074 104780
rect 543458 104184 543464 104236
rect 543516 104224 543522 104236
rect 545022 104224 545028 104236
rect 543516 104196 545028 104224
rect 543516 104184 543522 104196
rect 545022 104184 545028 104196
rect 545080 104184 545086 104236
rect 558362 104224 558368 104236
rect 545132 104196 558368 104224
rect 541894 104116 541900 104168
rect 541952 104156 541958 104168
rect 545132 104156 545160 104196
rect 558362 104184 558368 104196
rect 558420 104184 558426 104236
rect 541952 104128 545160 104156
rect 541952 104116 541958 104128
rect 547230 104116 547236 104168
rect 547288 104156 547294 104168
rect 563790 104156 563796 104168
rect 547288 104128 563796 104156
rect 547288 104116 547294 104128
rect 563790 104116 563796 104128
rect 563848 104116 563854 104168
rect 24486 103436 24492 103488
rect 24544 103476 24550 103488
rect 57514 103476 57520 103488
rect 24544 103448 57520 103476
rect 24544 103436 24550 103448
rect 57514 103436 57520 103448
rect 57572 103436 57578 103488
rect 24394 103368 24400 103420
rect 24452 103408 24458 103420
rect 57422 103408 57428 103420
rect 24452 103380 57428 103408
rect 24452 103368 24458 103380
rect 57422 103368 57428 103380
rect 57480 103368 57486 103420
rect 549898 103096 549904 103148
rect 549956 103136 549962 103148
rect 552474 103136 552480 103148
rect 549956 103108 552480 103136
rect 549956 103096 549962 103108
rect 552474 103096 552480 103108
rect 552532 103096 552538 103148
rect 540882 102280 540888 102332
rect 540940 102320 540946 102332
rect 545022 102320 545028 102332
rect 540940 102292 545028 102320
rect 540940 102280 540946 102292
rect 545022 102280 545028 102292
rect 545080 102280 545086 102332
rect 542170 102212 542176 102264
rect 542228 102252 542234 102264
rect 543642 102252 543648 102264
rect 542228 102224 543648 102252
rect 542228 102212 542234 102224
rect 543642 102212 543648 102224
rect 543700 102212 543706 102264
rect 542262 102144 542268 102196
rect 542320 102184 542326 102196
rect 542814 102184 542820 102196
rect 542320 102156 542820 102184
rect 542320 102144 542326 102156
rect 542814 102144 542820 102156
rect 542872 102144 542878 102196
rect 563790 102144 563796 102196
rect 563848 102184 563854 102196
rect 565814 102184 565820 102196
rect 563848 102156 565820 102184
rect 563848 102144 563854 102156
rect 565814 102144 565820 102156
rect 565872 102144 565878 102196
rect 542170 102076 542176 102128
rect 542228 102116 542234 102128
rect 548794 102116 548800 102128
rect 542228 102088 548800 102116
rect 542228 102076 542234 102088
rect 548794 102076 548800 102088
rect 548852 102076 548858 102128
rect 53742 101940 53748 101992
rect 53800 101980 53806 101992
rect 55398 101980 55404 101992
rect 53800 101952 55404 101980
rect 53800 101940 53806 101952
rect 55398 101940 55404 101952
rect 55456 101940 55462 101992
rect 543090 101804 543096 101856
rect 543148 101844 543154 101856
rect 549622 101844 549628 101856
rect 543148 101816 549628 101844
rect 543148 101804 543154 101816
rect 549622 101804 549628 101816
rect 549680 101804 549686 101856
rect 544470 100716 544476 100768
rect 544528 100756 544534 100768
rect 545574 100756 545580 100768
rect 544528 100728 545580 100756
rect 544528 100716 544534 100728
rect 545574 100716 545580 100728
rect 545632 100716 545638 100768
rect 549990 100716 549996 100768
rect 550048 100756 550054 100768
rect 550726 100756 550732 100768
rect 550048 100728 550732 100756
rect 550048 100716 550054 100728
rect 550726 100716 550732 100728
rect 550784 100716 550790 100768
rect 560202 100716 560208 100768
rect 560260 100756 560266 100768
rect 560846 100756 560852 100768
rect 560260 100728 560852 100756
rect 560260 100716 560266 100728
rect 560846 100716 560852 100728
rect 560904 100716 560910 100768
rect 27338 100648 27344 100700
rect 27396 100688 27402 100700
rect 57514 100688 57520 100700
rect 27396 100660 57520 100688
rect 27396 100648 27402 100660
rect 57514 100648 57520 100660
rect 57572 100648 57578 100700
rect 540974 99968 540980 100020
rect 541032 100008 541038 100020
rect 570138 100008 570144 100020
rect 541032 99980 570144 100008
rect 541032 99968 541038 99980
rect 570138 99968 570144 99980
rect 570196 99968 570202 100020
rect 559558 99356 559564 99408
rect 559616 99396 559622 99408
rect 561674 99396 561680 99408
rect 559616 99368 561680 99396
rect 559616 99356 559622 99368
rect 561674 99356 561680 99368
rect 561732 99356 561738 99408
rect 540698 98812 540704 98864
rect 540756 98852 540762 98864
rect 542354 98852 542360 98864
rect 540756 98824 542360 98852
rect 540756 98812 540762 98824
rect 542354 98812 542360 98824
rect 542412 98812 542418 98864
rect 541434 98676 541440 98728
rect 541492 98716 541498 98728
rect 541986 98716 541992 98728
rect 541492 98688 541992 98716
rect 541492 98676 541498 98688
rect 541986 98676 541992 98688
rect 542044 98676 542050 98728
rect 543550 98608 543556 98660
rect 543608 98648 543614 98660
rect 551278 98648 551284 98660
rect 543608 98620 551284 98648
rect 543608 98608 543614 98620
rect 551278 98608 551284 98620
rect 551336 98608 551342 98660
rect 57974 97996 57980 98048
rect 58032 98036 58038 98048
rect 59722 98036 59728 98048
rect 58032 98008 59728 98036
rect 58032 97996 58038 98008
rect 59722 97996 59728 98008
rect 59780 97996 59786 98048
rect 540514 97996 540520 98048
rect 540572 98036 540578 98048
rect 542170 98036 542176 98048
rect 540572 98008 542176 98036
rect 540572 97996 540578 98008
rect 542170 97996 542176 98008
rect 542228 97996 542234 98048
rect 46106 97928 46112 97980
rect 46164 97968 46170 97980
rect 57514 97968 57520 97980
rect 46164 97940 57520 97968
rect 46164 97928 46170 97940
rect 57514 97928 57520 97940
rect 57572 97928 57578 97980
rect 57882 97928 57888 97980
rect 57940 97968 57946 97980
rect 58802 97968 58808 97980
rect 57940 97940 58808 97968
rect 57940 97928 57946 97940
rect 58802 97928 58808 97940
rect 58860 97928 58866 97980
rect 543550 97928 543556 97980
rect 543608 97968 543614 97980
rect 570046 97968 570052 97980
rect 543608 97940 570052 97968
rect 543608 97928 543614 97940
rect 570046 97928 570052 97940
rect 570104 97928 570110 97980
rect 53190 97860 53196 97912
rect 53248 97900 53254 97912
rect 55858 97900 55864 97912
rect 53248 97872 55864 97900
rect 53248 97860 53254 97872
rect 55858 97860 55864 97872
rect 55916 97860 55922 97912
rect 58526 97860 58532 97912
rect 58584 97900 58590 97912
rect 59722 97900 59728 97912
rect 58584 97872 59728 97900
rect 58584 97860 58590 97872
rect 59722 97860 59728 97872
rect 59780 97860 59786 97912
rect 2866 97724 2872 97776
rect 2924 97764 2930 97776
rect 4798 97764 4804 97776
rect 2924 97736 4804 97764
rect 2924 97724 2930 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 543090 97248 543096 97300
rect 543148 97288 543154 97300
rect 547322 97288 547328 97300
rect 543148 97260 547328 97288
rect 543148 97248 543154 97260
rect 547322 97248 547328 97260
rect 547380 97248 547386 97300
rect 543550 96568 543556 96620
rect 543608 96608 543614 96620
rect 575566 96608 575572 96620
rect 543608 96580 575572 96608
rect 543608 96568 543614 96580
rect 575566 96568 575572 96580
rect 575624 96568 575630 96620
rect 54754 96092 54760 96144
rect 54812 96132 54818 96144
rect 57422 96132 57428 96144
rect 54812 96104 57428 96132
rect 54812 96092 54818 96104
rect 57422 96092 57428 96104
rect 57480 96092 57486 96144
rect 547414 95276 547420 95328
rect 547472 95316 547478 95328
rect 547874 95316 547880 95328
rect 547472 95288 547880 95316
rect 547472 95276 547478 95288
rect 547874 95276 547880 95288
rect 547932 95276 547938 95328
rect 53282 95208 53288 95260
rect 53340 95248 53346 95260
rect 55306 95248 55312 95260
rect 53340 95220 55312 95248
rect 53340 95208 53346 95220
rect 55306 95208 55312 95220
rect 55364 95208 55370 95260
rect 547322 95208 547328 95260
rect 547380 95248 547386 95260
rect 547966 95248 547972 95260
rect 547380 95220 547972 95248
rect 547380 95208 547386 95220
rect 547966 95208 547972 95220
rect 548024 95208 548030 95260
rect 28166 95140 28172 95192
rect 28224 95180 28230 95192
rect 57514 95180 57520 95192
rect 28224 95152 57520 95180
rect 28224 95140 28230 95152
rect 57514 95140 57520 95152
rect 57572 95140 57578 95192
rect 542262 95140 542268 95192
rect 542320 95180 542326 95192
rect 543366 95180 543372 95192
rect 542320 95152 543372 95180
rect 542320 95140 542326 95152
rect 543366 95140 543372 95152
rect 543424 95140 543430 95192
rect 543550 95140 543556 95192
rect 543608 95180 543614 95192
rect 555510 95180 555516 95192
rect 543608 95152 555516 95180
rect 543608 95140 543614 95152
rect 555510 95140 555516 95152
rect 555568 95140 555574 95192
rect 548794 94188 548800 94240
rect 548852 94228 548858 94240
rect 554130 94228 554136 94240
rect 548852 94200 554136 94228
rect 548852 94188 548858 94200
rect 554130 94188 554136 94200
rect 554188 94188 554194 94240
rect 543274 94052 543280 94104
rect 543332 94092 543338 94104
rect 544562 94092 544568 94104
rect 543332 94064 544568 94092
rect 543332 94052 543338 94064
rect 544562 94052 544568 94064
rect 544620 94052 544626 94104
rect 57514 93916 57520 93968
rect 57572 93956 57578 93968
rect 57882 93956 57888 93968
rect 57572 93928 57888 93956
rect 57572 93916 57578 93928
rect 57882 93916 57888 93928
rect 57940 93916 57946 93968
rect 543550 93916 543556 93968
rect 543608 93956 543614 93968
rect 545114 93956 545120 93968
rect 543608 93928 545120 93956
rect 543608 93916 543614 93928
rect 545114 93916 545120 93928
rect 545172 93916 545178 93968
rect 51626 93780 51632 93832
rect 51684 93820 51690 93832
rect 57882 93820 57888 93832
rect 51684 93792 57888 93820
rect 51684 93780 51690 93792
rect 57882 93780 57888 93792
rect 57940 93780 57946 93832
rect 51626 92488 51632 92540
rect 51684 92528 51690 92540
rect 55398 92528 55404 92540
rect 51684 92500 55404 92528
rect 51684 92488 51690 92500
rect 55398 92488 55404 92500
rect 55456 92488 55462 92540
rect 543550 91196 543556 91248
rect 543608 91236 543614 91248
rect 549714 91236 549720 91248
rect 543608 91208 549720 91236
rect 543608 91196 543614 91208
rect 549714 91196 549720 91208
rect 549772 91196 549778 91248
rect 41230 90992 41236 91044
rect 41288 91032 41294 91044
rect 57882 91032 57888 91044
rect 41288 91004 57888 91032
rect 41288 90992 41294 91004
rect 57882 90992 57888 91004
rect 57940 90992 57946 91044
rect 542262 90856 542268 90908
rect 542320 90896 542326 90908
rect 549714 90896 549720 90908
rect 542320 90868 549720 90896
rect 542320 90856 542326 90868
rect 549714 90856 549720 90868
rect 549772 90856 549778 90908
rect 543458 90516 543464 90568
rect 543516 90556 543522 90568
rect 544102 90556 544108 90568
rect 543516 90528 544108 90556
rect 543516 90516 543522 90528
rect 544102 90516 544108 90528
rect 544160 90516 544166 90568
rect 540882 89768 540888 89820
rect 540940 89808 540946 89820
rect 543734 89808 543740 89820
rect 540940 89780 543740 89808
rect 540940 89768 540946 89780
rect 543734 89768 543740 89780
rect 543792 89768 543798 89820
rect 542630 89700 542636 89752
rect 542688 89740 542694 89752
rect 544194 89740 544200 89752
rect 542688 89712 544200 89740
rect 542688 89700 542694 89712
rect 544194 89700 544200 89712
rect 544252 89700 544258 89752
rect 30098 89632 30104 89684
rect 30156 89672 30162 89684
rect 57882 89672 57888 89684
rect 30156 89644 57888 89672
rect 30156 89632 30162 89644
rect 57882 89632 57888 89644
rect 57940 89632 57946 89684
rect 543550 89632 543556 89684
rect 543608 89672 543614 89684
rect 581730 89672 581736 89684
rect 543608 89644 581736 89672
rect 543608 89632 543614 89644
rect 581730 89632 581736 89644
rect 581788 89632 581794 89684
rect 546126 89564 546132 89616
rect 546184 89604 546190 89616
rect 547874 89604 547880 89616
rect 546184 89576 547880 89604
rect 546184 89564 546190 89576
rect 547874 89564 547880 89576
rect 547932 89564 547938 89616
rect 546402 89496 546408 89548
rect 546460 89536 546466 89548
rect 547966 89536 547972 89548
rect 546460 89508 547972 89536
rect 546460 89496 546466 89508
rect 547966 89496 547972 89508
rect 548024 89496 548030 89548
rect 547414 89428 547420 89480
rect 547472 89468 547478 89480
rect 549622 89468 549628 89480
rect 547472 89440 549628 89468
rect 547472 89428 547478 89440
rect 549622 89428 549628 89440
rect 549680 89428 549686 89480
rect 540606 88272 540612 88324
rect 540664 88312 540670 88324
rect 543826 88312 543832 88324
rect 540664 88284 543832 88312
rect 540664 88272 540670 88284
rect 543826 88272 543832 88284
rect 543884 88272 543890 88324
rect 545022 88272 545028 88324
rect 545080 88312 545086 88324
rect 545942 88312 545948 88324
rect 545080 88284 545948 88312
rect 545080 88272 545086 88284
rect 545942 88272 545948 88284
rect 546000 88272 546006 88324
rect 543458 87592 543464 87644
rect 543516 87632 543522 87644
rect 550634 87632 550640 87644
rect 543516 87604 550640 87632
rect 543516 87592 543522 87604
rect 550634 87592 550640 87604
rect 550692 87592 550698 87644
rect 540514 85756 540520 85808
rect 540572 85796 540578 85808
rect 543458 85796 543464 85808
rect 540572 85768 543464 85796
rect 540572 85756 540578 85768
rect 543458 85756 543464 85768
rect 543516 85756 543522 85808
rect 543826 85756 543832 85808
rect 543884 85796 543890 85808
rect 549254 85796 549260 85808
rect 543884 85768 549260 85796
rect 543884 85756 543890 85768
rect 549254 85756 549260 85768
rect 549312 85756 549318 85808
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 21358 85524 21364 85536
rect 3568 85496 21364 85524
rect 3568 85484 3574 85496
rect 21358 85484 21364 85496
rect 21416 85484 21422 85536
rect 540790 85484 540796 85536
rect 540848 85524 540854 85536
rect 547322 85524 547328 85536
rect 540848 85496 547328 85524
rect 540848 85484 540854 85496
rect 547322 85484 547328 85496
rect 547380 85484 547386 85536
rect 542354 84600 542360 84652
rect 542412 84640 542418 84652
rect 544930 84640 544936 84652
rect 542412 84612 544936 84640
rect 542412 84600 542418 84612
rect 544930 84600 544936 84612
rect 544988 84600 544994 84652
rect 543550 84124 543556 84176
rect 543608 84164 543614 84176
rect 552566 84164 552572 84176
rect 543608 84136 552572 84164
rect 543608 84124 543614 84136
rect 552566 84124 552572 84136
rect 552624 84124 552630 84176
rect 543734 83920 543740 83972
rect 543792 83960 543798 83972
rect 547874 83960 547880 83972
rect 543792 83932 547880 83960
rect 543792 83920 543798 83932
rect 547874 83920 547880 83932
rect 547932 83920 547938 83972
rect 545022 83852 545028 83904
rect 545080 83892 545086 83904
rect 546494 83892 546500 83904
rect 545080 83864 546500 83892
rect 545080 83852 545086 83864
rect 546494 83852 546500 83864
rect 546552 83852 546558 83904
rect 552934 83444 552940 83496
rect 552992 83484 552998 83496
rect 565170 83484 565176 83496
rect 552992 83456 565176 83484
rect 552992 83444 552998 83456
rect 565170 83444 565176 83456
rect 565228 83444 565234 83496
rect 544562 82968 544568 83020
rect 544620 83008 544626 83020
rect 547966 83008 547972 83020
rect 544620 82980 547972 83008
rect 544620 82968 544626 82980
rect 547966 82968 547972 82980
rect 548024 82968 548030 83020
rect 57054 82900 57060 82952
rect 57112 82940 57118 82952
rect 57606 82940 57612 82952
rect 57112 82912 57612 82940
rect 57112 82900 57118 82912
rect 57606 82900 57612 82912
rect 57664 82900 57670 82952
rect 540514 82900 540520 82952
rect 540572 82940 540578 82952
rect 546126 82940 546132 82952
rect 540572 82912 546132 82940
rect 540572 82900 540578 82912
rect 546126 82900 546132 82912
rect 546184 82900 546190 82952
rect 54754 82832 54760 82884
rect 54812 82872 54818 82884
rect 55214 82872 55220 82884
rect 54812 82844 55220 82872
rect 54812 82832 54818 82844
rect 55214 82832 55220 82844
rect 55272 82832 55278 82884
rect 546034 82832 546040 82884
rect 546092 82872 546098 82884
rect 547414 82872 547420 82884
rect 546092 82844 547420 82872
rect 546092 82832 546098 82844
rect 547414 82832 547420 82844
rect 547472 82832 547478 82884
rect 552842 82832 552848 82884
rect 552900 82872 552906 82884
rect 556614 82872 556620 82884
rect 552900 82844 556620 82872
rect 552900 82832 552906 82844
rect 556614 82832 556620 82844
rect 556672 82832 556678 82884
rect 23382 82764 23388 82816
rect 23440 82804 23446 82816
rect 57606 82804 57612 82816
rect 23440 82776 57612 82804
rect 23440 82764 23446 82776
rect 57606 82764 57612 82776
rect 57664 82764 57670 82816
rect 543550 82764 543556 82816
rect 543608 82804 543614 82816
rect 552382 82804 552388 82816
rect 543608 82776 552388 82804
rect 543608 82764 543614 82776
rect 552382 82764 552388 82776
rect 552440 82764 552446 82816
rect 47578 82696 47584 82748
rect 47636 82736 47642 82748
rect 57882 82736 57888 82748
rect 47636 82708 57888 82736
rect 47636 82696 47642 82708
rect 57882 82696 57888 82708
rect 57940 82696 57946 82748
rect 48958 82084 48964 82136
rect 49016 82124 49022 82136
rect 55950 82124 55956 82136
rect 49016 82096 55956 82124
rect 49016 82084 49022 82096
rect 55950 82084 55956 82096
rect 56008 82084 56014 82136
rect 551370 80044 551376 80096
rect 551428 80084 551434 80096
rect 552474 80084 552480 80096
rect 551428 80056 552480 80084
rect 551428 80044 551434 80056
rect 552474 80044 552480 80056
rect 552532 80044 552538 80096
rect 540146 79296 540152 79348
rect 540204 79336 540210 79348
rect 540422 79336 540428 79348
rect 540204 79308 540428 79336
rect 540204 79296 540210 79308
rect 540422 79296 540428 79308
rect 540480 79296 540486 79348
rect 543642 78616 543648 78668
rect 543700 78656 543706 78668
rect 563974 78656 563980 78668
rect 543700 78628 563980 78656
rect 543700 78616 543706 78628
rect 563974 78616 563980 78628
rect 564032 78616 564038 78668
rect 543550 78548 543556 78600
rect 543608 78588 543614 78600
rect 561030 78588 561036 78600
rect 543608 78560 561036 78588
rect 543608 78548 543614 78560
rect 561030 78548 561036 78560
rect 561088 78548 561094 78600
rect 543550 77188 543556 77240
rect 543608 77228 543614 77240
rect 559650 77228 559656 77240
rect 543608 77200 559656 77228
rect 543608 77188 543614 77200
rect 559650 77188 559656 77200
rect 559708 77188 559714 77240
rect 51718 75828 51724 75880
rect 51776 75868 51782 75880
rect 57606 75868 57612 75880
rect 51776 75840 57612 75868
rect 51776 75828 51782 75840
rect 57606 75828 57612 75840
rect 57664 75828 57670 75880
rect 540606 75828 540612 75880
rect 540664 75868 540670 75880
rect 542446 75868 542452 75880
rect 540664 75840 542452 75868
rect 540664 75828 540670 75840
rect 542446 75828 542452 75840
rect 542504 75828 542510 75880
rect 543550 75216 543556 75268
rect 543608 75256 543614 75268
rect 550266 75256 550272 75268
rect 543608 75228 550272 75256
rect 543608 75216 543614 75228
rect 550266 75216 550272 75228
rect 550324 75216 550330 75268
rect 545942 74536 545948 74588
rect 546000 74576 546006 74588
rect 549806 74576 549812 74588
rect 546000 74548 549812 74576
rect 546000 74536 546006 74548
rect 549806 74536 549812 74548
rect 549864 74536 549870 74588
rect 53282 73652 53288 73704
rect 53340 73692 53346 73704
rect 56962 73692 56968 73704
rect 53340 73664 56968 73692
rect 53340 73652 53346 73664
rect 56962 73652 56968 73664
rect 57020 73652 57026 73704
rect 542170 73176 542176 73228
rect 542228 73216 542234 73228
rect 544102 73216 544108 73228
rect 542228 73188 544108 73216
rect 542228 73176 542234 73188
rect 544102 73176 544108 73188
rect 544160 73176 544166 73228
rect 546034 73176 546040 73228
rect 546092 73176 546098 73228
rect 549898 73176 549904 73228
rect 549956 73216 549962 73228
rect 556890 73216 556896 73228
rect 549956 73188 556896 73216
rect 549956 73176 549962 73188
rect 556890 73176 556896 73188
rect 556948 73176 556954 73228
rect 546052 73148 546080 73176
rect 548242 73148 548248 73160
rect 546052 73120 548248 73148
rect 548242 73108 548248 73120
rect 548300 73108 548306 73160
rect 576118 73108 576124 73160
rect 576176 73148 576182 73160
rect 580258 73148 580264 73160
rect 576176 73120 580264 73148
rect 576176 73108 576182 73120
rect 580258 73108 580264 73120
rect 580316 73108 580322 73160
rect 543550 72428 543556 72480
rect 543608 72468 543614 72480
rect 562502 72468 562508 72480
rect 543608 72440 562508 72468
rect 543608 72428 543614 72440
rect 562502 72428 562508 72440
rect 562560 72428 562566 72480
rect 545114 72224 545120 72276
rect 545172 72264 545178 72276
rect 549990 72264 549996 72276
rect 545172 72236 549996 72264
rect 545172 72224 545178 72236
rect 549990 72224 549996 72236
rect 550048 72224 550054 72276
rect 547322 71680 547328 71732
rect 547380 71720 547386 71732
rect 549806 71720 549812 71732
rect 547380 71692 549812 71720
rect 547380 71680 547386 71692
rect 549806 71680 549812 71692
rect 549864 71680 549870 71732
rect 542814 71000 542820 71052
rect 542872 71040 542878 71052
rect 566734 71040 566740 71052
rect 542872 71012 566740 71040
rect 542872 71000 542878 71012
rect 566734 71000 566740 71012
rect 566792 71000 566798 71052
rect 542078 70592 542084 70644
rect 542136 70632 542142 70644
rect 546494 70632 546500 70644
rect 542136 70604 546500 70632
rect 542136 70592 542142 70604
rect 546494 70592 546500 70604
rect 546552 70592 546558 70644
rect 546494 70456 546500 70508
rect 546552 70496 546558 70508
rect 549254 70496 549260 70508
rect 546552 70468 549260 70496
rect 546552 70456 546558 70468
rect 549254 70456 549260 70468
rect 549312 70456 549318 70508
rect 543550 70320 543556 70372
rect 543608 70360 543614 70372
rect 552290 70360 552296 70372
rect 543608 70332 552296 70360
rect 543608 70320 543614 70332
rect 552290 70320 552296 70332
rect 552348 70320 552354 70372
rect 542630 69844 542636 69896
rect 542688 69884 542694 69896
rect 544102 69884 544108 69896
rect 542688 69856 544108 69884
rect 542688 69844 542694 69856
rect 544102 69844 544108 69856
rect 544160 69844 544166 69896
rect 45094 69640 45100 69692
rect 45152 69680 45158 69692
rect 57054 69680 57060 69692
rect 45152 69652 57060 69680
rect 45152 69640 45158 69652
rect 57054 69640 57060 69652
rect 57112 69640 57118 69692
rect 543734 69640 543740 69692
rect 543792 69680 543798 69692
rect 546954 69680 546960 69692
rect 543792 69652 546960 69680
rect 543792 69640 543798 69652
rect 546954 69640 546960 69652
rect 547012 69640 547018 69692
rect 18966 68960 18972 69012
rect 19024 69000 19030 69012
rect 57606 69000 57612 69012
rect 19024 68972 57612 69000
rect 19024 68960 19030 68972
rect 57606 68960 57612 68972
rect 57664 68960 57670 69012
rect 540882 68960 540888 69012
rect 540940 69000 540946 69012
rect 542630 69000 542636 69012
rect 540940 68972 542636 69000
rect 540940 68960 540946 68972
rect 542630 68960 542636 68972
rect 542688 68960 542694 69012
rect 56962 68076 56968 68128
rect 57020 68116 57026 68128
rect 57606 68116 57612 68128
rect 57020 68088 57612 68116
rect 57020 68076 57026 68088
rect 57606 68076 57612 68088
rect 57664 68076 57670 68128
rect 546034 67600 546040 67652
rect 546092 67640 546098 67652
rect 546494 67640 546500 67652
rect 546092 67612 546500 67640
rect 546092 67600 546098 67612
rect 546494 67600 546500 67612
rect 546552 67600 546558 67652
rect 50522 67124 50528 67176
rect 50580 67164 50586 67176
rect 56686 67164 56692 67176
rect 50580 67136 56692 67164
rect 50580 67124 50586 67136
rect 56686 67124 56692 67136
rect 56744 67124 56750 67176
rect 540606 66648 540612 66700
rect 540664 66688 540670 66700
rect 545114 66688 545120 66700
rect 540664 66660 545120 66688
rect 540664 66648 540670 66660
rect 545114 66648 545120 66660
rect 545172 66648 545178 66700
rect 543550 66172 543556 66224
rect 543608 66212 543614 66224
rect 577314 66212 577320 66224
rect 543608 66184 577320 66212
rect 543608 66172 543614 66184
rect 577314 66172 577320 66184
rect 577372 66172 577378 66224
rect 20438 64812 20444 64864
rect 20496 64852 20502 64864
rect 56962 64852 56968 64864
rect 20496 64824 56968 64852
rect 20496 64812 20502 64824
rect 56962 64812 56968 64824
rect 57020 64812 57026 64864
rect 46198 64744 46204 64796
rect 46256 64784 46262 64796
rect 57882 64784 57888 64796
rect 46256 64756 57888 64784
rect 46256 64744 46262 64756
rect 57882 64744 57888 64756
rect 57940 64744 57946 64796
rect 543550 63996 543556 64048
rect 543608 64036 543614 64048
rect 549530 64036 549536 64048
rect 543608 64008 549536 64036
rect 543608 63996 543614 64008
rect 549530 63996 549536 64008
rect 549588 63996 549594 64048
rect 57790 63656 57796 63708
rect 57848 63656 57854 63708
rect 57808 63504 57836 63656
rect 43530 63452 43536 63504
rect 43588 63492 43594 63504
rect 57698 63492 57704 63504
rect 43588 63464 57704 63492
rect 43588 63452 43594 63464
rect 57698 63452 57704 63464
rect 57756 63452 57762 63504
rect 57790 63452 57796 63504
rect 57848 63452 57854 63504
rect 41782 62024 41788 62076
rect 41840 62064 41846 62076
rect 57698 62064 57704 62076
rect 41840 62036 57704 62064
rect 41840 62024 41846 62036
rect 57698 62024 57704 62036
rect 57756 62024 57762 62076
rect 543550 62024 543556 62076
rect 543608 62064 543614 62076
rect 560754 62064 560760 62076
rect 543608 62036 560760 62064
rect 543608 62024 543614 62036
rect 560754 62024 560760 62036
rect 560812 62024 560818 62076
rect 543642 61956 543648 62008
rect 543700 61996 543706 62008
rect 560570 61996 560576 62008
rect 543700 61968 560576 61996
rect 543700 61956 543706 61968
rect 560570 61956 560576 61968
rect 560628 61956 560634 62008
rect 574738 60664 574744 60716
rect 574796 60704 574802 60716
rect 580258 60704 580264 60716
rect 574796 60676 580264 60704
rect 574796 60664 574802 60676
rect 580258 60664 580264 60676
rect 580316 60664 580322 60716
rect 26050 59304 26056 59356
rect 26108 59344 26114 59356
rect 57698 59344 57704 59356
rect 26108 59316 57704 59344
rect 26108 59304 26114 59316
rect 57698 59304 57704 59316
rect 57756 59304 57762 59356
rect 543550 57876 543556 57928
rect 543608 57916 543614 57928
rect 574094 57916 574100 57928
rect 543608 57888 574100 57916
rect 543608 57876 543614 57888
rect 574094 57876 574100 57888
rect 574152 57876 574158 57928
rect 54938 57264 54944 57316
rect 54996 57304 55002 57316
rect 57698 57304 57704 57316
rect 54996 57276 57704 57304
rect 54996 57264 55002 57276
rect 57698 57264 57704 57276
rect 57756 57264 57762 57316
rect 49234 53728 49240 53780
rect 49292 53768 49298 53780
rect 57698 53768 57704 53780
rect 49292 53740 57704 53768
rect 49292 53728 49298 53740
rect 57698 53728 57704 53740
rect 57756 53728 57762 53780
rect 543550 53728 543556 53780
rect 543608 53768 543614 53780
rect 569218 53768 569224 53780
rect 543608 53740 569224 53768
rect 543608 53728 543614 53740
rect 569218 53728 569224 53740
rect 569276 53728 569282 53780
rect 543458 50804 543464 50856
rect 543516 50844 543522 50856
rect 547046 50844 547052 50856
rect 543516 50816 547052 50844
rect 543516 50804 543522 50816
rect 547046 50804 547052 50816
rect 547104 50804 547110 50856
rect 543550 49648 543556 49700
rect 543608 49688 543614 49700
rect 551186 49688 551192 49700
rect 543608 49660 551192 49688
rect 543608 49648 543614 49660
rect 551186 49648 551192 49660
rect 551244 49648 551250 49700
rect 30190 48220 30196 48272
rect 30248 48260 30254 48272
rect 57698 48260 57704 48272
rect 30248 48232 57704 48260
rect 30248 48220 30254 48232
rect 57698 48220 57704 48232
rect 57756 48220 57762 48272
rect 543550 48220 543556 48272
rect 543608 48260 543614 48272
rect 575474 48260 575480 48272
rect 543608 48232 575480 48260
rect 543608 48220 543614 48232
rect 575474 48220 575480 48232
rect 575532 48220 575538 48272
rect 543550 45500 543556 45552
rect 543608 45540 543614 45552
rect 579890 45540 579896 45552
rect 543608 45512 579896 45540
rect 543608 45500 543614 45512
rect 579890 45500 579896 45512
rect 579948 45500 579954 45552
rect 543642 45432 543648 45484
rect 543700 45472 543706 45484
rect 563146 45472 563152 45484
rect 543700 45444 563152 45472
rect 543700 45432 543706 45444
rect 563146 45432 563152 45444
rect 563204 45432 563210 45484
rect 543550 44072 543556 44124
rect 543608 44112 543614 44124
rect 560478 44112 560484 44124
rect 543608 44084 560484 44112
rect 543608 44072 543614 44084
rect 560478 44072 560484 44084
rect 560536 44072 560542 44124
rect 542354 42304 542360 42356
rect 542412 42344 542418 42356
rect 544194 42344 544200 42356
rect 542412 42316 544200 42344
rect 542412 42304 542418 42316
rect 544194 42304 544200 42316
rect 544252 42304 544258 42356
rect 46290 41352 46296 41404
rect 46348 41392 46354 41404
rect 57698 41392 57704 41404
rect 46348 41364 57704 41392
rect 46348 41352 46354 41364
rect 57698 41352 57704 41364
rect 57756 41352 57762 41404
rect 543550 41352 543556 41404
rect 543608 41392 543614 41404
rect 563882 41392 563888 41404
rect 543608 41364 563888 41392
rect 543608 41352 543614 41364
rect 563882 41352 563888 41364
rect 563940 41352 563946 41404
rect 47026 39992 47032 40044
rect 47084 40032 47090 40044
rect 57698 40032 57704 40044
rect 47084 40004 57704 40032
rect 47084 39992 47090 40004
rect 57698 39992 57704 40004
rect 57756 39992 57762 40044
rect 543550 37204 543556 37256
rect 543608 37244 543614 37256
rect 562042 37244 562048 37256
rect 543608 37216 562048 37244
rect 543608 37204 543614 37216
rect 562042 37204 562048 37216
rect 562100 37204 562106 37256
rect 540882 36728 540888 36780
rect 540940 36768 540946 36780
rect 542538 36768 542544 36780
rect 540940 36740 542544 36768
rect 540940 36728 540946 36740
rect 542538 36728 542544 36740
rect 542596 36728 542602 36780
rect 543550 35844 543556 35896
rect 543608 35884 543614 35896
rect 581638 35884 581644 35896
rect 543608 35856 581644 35884
rect 543608 35844 543614 35856
rect 581638 35844 581644 35856
rect 581696 35844 581702 35896
rect 24578 34416 24584 34468
rect 24636 34456 24642 34468
rect 57698 34456 57704 34468
rect 24636 34428 57704 34456
rect 24636 34416 24642 34428
rect 57698 34416 57704 34428
rect 57756 34416 57762 34468
rect 33686 33056 33692 33108
rect 33744 33096 33750 33108
rect 57698 33096 57704 33108
rect 33744 33068 57704 33096
rect 33744 33056 33750 33068
rect 57698 33056 57704 33068
rect 57756 33056 57762 33108
rect 570598 33056 570604 33108
rect 570656 33096 570662 33108
rect 579798 33096 579804 33108
rect 570656 33068 579804 33096
rect 570656 33056 570662 33068
rect 579798 33056 579804 33068
rect 579856 33056 579862 33108
rect 34054 32988 34060 33040
rect 34112 33028 34118 33040
rect 57790 33028 57796 33040
rect 34112 33000 57796 33028
rect 34112 32988 34118 33000
rect 57790 32988 57796 33000
rect 57848 32988 57854 33040
rect 46566 31696 46572 31748
rect 46624 31736 46630 31748
rect 57698 31736 57704 31748
rect 46624 31708 57704 31736
rect 46624 31696 46630 31708
rect 57698 31696 57704 31708
rect 57756 31696 57762 31748
rect 543550 31696 543556 31748
rect 543608 31736 543614 31748
rect 583294 31736 583300 31748
rect 543608 31708 583300 31736
rect 543608 31696 543614 31708
rect 583294 31696 583300 31708
rect 583352 31696 583358 31748
rect 540882 31084 540888 31136
rect 540940 31124 540946 31136
rect 567746 31124 567752 31136
rect 540940 31096 567752 31124
rect 540940 31084 540946 31096
rect 567746 31084 567752 31096
rect 567804 31084 567810 31136
rect 540698 31016 540704 31068
rect 540756 31056 540762 31068
rect 568850 31056 568856 31068
rect 540756 31028 568856 31056
rect 540756 31016 540762 31028
rect 568850 31016 568856 31028
rect 568908 31016 568914 31068
rect 540606 30268 540612 30320
rect 540664 30308 540670 30320
rect 544470 30308 544476 30320
rect 540664 30280 544476 30308
rect 540664 30268 540670 30280
rect 544470 30268 544476 30280
rect 544528 30268 544534 30320
rect 168374 29860 168380 29912
rect 168432 29900 168438 29912
rect 169494 29900 169500 29912
rect 168432 29872 169500 29900
rect 168432 29860 168438 29872
rect 169494 29860 169500 29872
rect 169552 29860 169558 29912
rect 340874 29860 340880 29912
rect 340932 29900 340938 29912
rect 342086 29900 342092 29912
rect 340932 29872 342092 29900
rect 340932 29860 340938 29872
rect 342086 29860 342092 29872
rect 342144 29860 342150 29912
rect 361574 29860 361580 29912
rect 361632 29900 361638 29912
rect 362694 29900 362700 29912
rect 361632 29872 362700 29900
rect 361632 29860 361638 29872
rect 362694 29860 362700 29872
rect 362752 29860 362758 29912
rect 445846 29860 445852 29912
rect 445904 29900 445910 29912
rect 447058 29900 447064 29912
rect 445904 29872 447064 29900
rect 445904 29860 445910 29872
rect 447058 29860 447064 29872
rect 447116 29860 447122 29912
rect 458174 29860 458180 29912
rect 458232 29900 458238 29912
rect 459294 29900 459300 29912
rect 458232 29872 459300 29900
rect 458232 29860 458238 29872
rect 459294 29860 459300 29872
rect 459352 29860 459358 29912
rect 474734 29860 474740 29912
rect 474792 29900 474798 29912
rect 476038 29900 476044 29912
rect 474792 29872 476044 29900
rect 474792 29860 474798 29872
rect 476038 29860 476044 29872
rect 476096 29860 476102 29912
rect 525794 29860 525800 29912
rect 525852 29900 525858 29912
rect 526914 29900 526920 29912
rect 525852 29872 526920 29900
rect 525852 29860 525858 29872
rect 526914 29860 526920 29872
rect 526972 29860 526978 29912
rect 536834 29656 536840 29708
rect 536892 29696 536898 29708
rect 545850 29696 545856 29708
rect 536892 29668 545856 29696
rect 536892 29656 536898 29668
rect 545850 29656 545856 29668
rect 545908 29656 545914 29708
rect 45278 29588 45284 29640
rect 45336 29628 45342 29640
rect 69014 29628 69020 29640
rect 45336 29600 69020 29628
rect 45336 29588 45342 29600
rect 69014 29588 69020 29600
rect 69072 29588 69078 29640
rect 531406 29588 531412 29640
rect 531464 29628 531470 29640
rect 534810 29628 534816 29640
rect 531464 29600 534816 29628
rect 531464 29588 531470 29600
rect 534810 29588 534816 29600
rect 534868 29588 534874 29640
rect 535454 29588 535460 29640
rect 535512 29628 535518 29640
rect 581822 29628 581828 29640
rect 535512 29600 581828 29628
rect 535512 29588 535518 29600
rect 581822 29588 581828 29600
rect 581880 29588 581886 29640
rect 52822 29520 52828 29572
rect 52880 29560 52886 29572
rect 63218 29560 63224 29572
rect 52880 29532 63224 29560
rect 52880 29520 52886 29532
rect 63218 29520 63224 29532
rect 63276 29520 63282 29572
rect 474642 29520 474648 29572
rect 474700 29560 474706 29572
rect 474826 29560 474832 29572
rect 474700 29532 474832 29560
rect 474700 29520 474706 29532
rect 474826 29520 474832 29532
rect 474884 29520 474890 29572
rect 515950 29520 515956 29572
rect 516008 29560 516014 29572
rect 548150 29560 548156 29572
rect 516008 29532 548156 29560
rect 516008 29520 516014 29532
rect 548150 29520 548156 29532
rect 548208 29520 548214 29572
rect 43070 29452 43076 29504
rect 43128 29492 43134 29504
rect 69658 29492 69664 29504
rect 43128 29464 69664 29492
rect 43128 29452 43134 29464
rect 69658 29452 69664 29464
rect 69716 29452 69722 29504
rect 514018 29452 514024 29504
rect 514076 29492 514082 29504
rect 548334 29492 548340 29504
rect 514076 29464 548340 29492
rect 514076 29452 514082 29464
rect 548334 29452 548340 29464
rect 548392 29452 548398 29504
rect 33962 29384 33968 29436
rect 34020 29424 34026 29436
rect 71590 29424 71596 29436
rect 34020 29396 71596 29424
rect 34020 29384 34026 29396
rect 71590 29384 71596 29396
rect 71648 29384 71654 29436
rect 509510 29384 509516 29436
rect 509568 29424 509574 29436
rect 546770 29424 546776 29436
rect 509568 29396 546776 29424
rect 509568 29384 509574 29396
rect 546770 29384 546776 29396
rect 546828 29384 546834 29436
rect 42518 29316 42524 29368
rect 42576 29356 42582 29368
rect 159818 29356 159824 29368
rect 42576 29328 159824 29356
rect 42576 29316 42582 29328
rect 159818 29316 159824 29328
rect 159876 29316 159882 29368
rect 506934 29316 506940 29368
rect 506992 29356 506998 29368
rect 565906 29356 565912 29368
rect 506992 29328 565912 29356
rect 506992 29316 506998 29328
rect 565906 29316 565912 29328
rect 565964 29316 565970 29368
rect 51810 29248 51816 29300
rect 51868 29288 51874 29300
rect 170766 29288 170772 29300
rect 51868 29260 170772 29288
rect 51868 29248 51874 29260
rect 170766 29248 170772 29260
rect 170824 29248 170830 29300
rect 443178 29248 443184 29300
rect 443236 29288 443242 29300
rect 561950 29288 561956 29300
rect 443236 29260 561956 29288
rect 443236 29248 443242 29260
rect 561950 29248 561956 29260
rect 562008 29248 562014 29300
rect 47210 29180 47216 29232
rect 47268 29220 47274 29232
rect 199746 29220 199752 29232
rect 47268 29192 199752 29220
rect 47268 29180 47274 29192
rect 199746 29180 199752 29192
rect 199804 29180 199810 29232
rect 372982 29180 372988 29232
rect 373040 29220 373046 29232
rect 535454 29220 535460 29232
rect 373040 29192 535460 29220
rect 373040 29180 373046 29192
rect 535454 29180 535460 29192
rect 535512 29180 535518 29232
rect 537846 29180 537852 29232
rect 537904 29220 537910 29232
rect 546310 29220 546316 29232
rect 537904 29192 546316 29220
rect 537904 29180 537910 29192
rect 546310 29180 546316 29192
rect 546368 29180 546374 29232
rect 29730 29112 29736 29164
rect 29788 29152 29794 29164
rect 187510 29152 187516 29164
rect 29788 29124 187516 29152
rect 29788 29112 29794 29124
rect 187510 29112 187516 29124
rect 187568 29112 187574 29164
rect 356882 29112 356888 29164
rect 356940 29152 356946 29164
rect 560938 29152 560944 29164
rect 356940 29124 560944 29152
rect 356940 29112 356946 29124
rect 560938 29112 560944 29124
rect 560996 29112 561002 29164
rect 42242 29044 42248 29096
rect 42300 29084 42306 29096
rect 205542 29084 205548 29096
rect 42300 29056 205548 29084
rect 42300 29044 42306 29056
rect 205542 29044 205548 29056
rect 205600 29044 205606 29096
rect 287330 29044 287336 29096
rect 287388 29084 287394 29096
rect 287388 29056 533292 29084
rect 287388 29044 287394 29056
rect 31110 28976 31116 29028
rect 31168 29016 31174 29028
rect 109586 29016 109592 29028
rect 31168 28988 109592 29016
rect 31168 28976 31174 28988
rect 109586 28976 109592 28988
rect 109644 28976 109650 29028
rect 158530 28976 158536 29028
rect 158588 29016 158594 29028
rect 531222 29016 531228 29028
rect 158588 28988 531228 29016
rect 158588 28976 158594 28988
rect 531222 28976 531228 28988
rect 531280 28976 531286 29028
rect 533264 29016 533292 29056
rect 534810 29044 534816 29096
rect 534868 29084 534874 29096
rect 550910 29084 550916 29096
rect 534868 29056 550916 29084
rect 534868 29044 534874 29056
rect 550910 29044 550916 29056
rect 550968 29044 550974 29096
rect 539502 29016 539508 29028
rect 533264 28988 539508 29016
rect 539502 28976 539508 28988
rect 539560 28976 539566 29028
rect 52086 28908 52092 28960
rect 52144 28948 52150 28960
rect 70946 28948 70952 28960
rect 52144 28920 70952 28948
rect 52144 28908 52150 28920
rect 70946 28908 70952 28920
rect 71004 28908 71010 28960
rect 247402 28908 247408 28960
rect 247460 28948 247466 28960
rect 511258 28948 511264 28960
rect 247460 28920 511264 28948
rect 247460 28908 247466 28920
rect 511258 28908 511264 28920
rect 511316 28908 511322 28960
rect 49418 28840 49424 28892
rect 49476 28880 49482 28892
rect 67726 28880 67732 28892
rect 49476 28852 67732 28880
rect 49476 28840 49482 28852
rect 67726 28840 67732 28852
rect 67784 28840 67790 28892
rect 381354 28840 381360 28892
rect 381412 28880 381418 28892
rect 553946 28880 553952 28892
rect 381412 28852 553952 28880
rect 381412 28840 381418 28852
rect 553946 28840 553952 28852
rect 554004 28840 554010 28892
rect 39850 28772 39856 28824
rect 39908 28812 39914 28824
rect 82538 28812 82544 28824
rect 39908 28784 82544 28812
rect 39908 28772 39914 28784
rect 82538 28772 82544 28784
rect 82596 28772 82602 28824
rect 82814 28772 82820 28824
rect 82872 28812 82878 28824
rect 249978 28812 249984 28824
rect 82872 28784 249984 28812
rect 82872 28772 82878 28784
rect 249978 28772 249984 28784
rect 250036 28772 250042 28824
rect 451550 28772 451556 28824
rect 451608 28812 451614 28824
rect 561122 28812 561128 28824
rect 451608 28784 561128 28812
rect 451608 28772 451614 28784
rect 561122 28772 561128 28784
rect 561180 28772 561186 28824
rect 45462 28704 45468 28756
rect 45520 28744 45526 28756
rect 204898 28744 204904 28756
rect 45520 28716 204904 28744
rect 45520 28704 45526 28716
rect 204898 28704 204904 28716
rect 204956 28704 204962 28756
rect 275738 28704 275744 28756
rect 275796 28744 275802 28756
rect 387058 28744 387064 28756
rect 275796 28716 387064 28744
rect 275796 28704 275802 28716
rect 387058 28704 387064 28716
rect 387116 28704 387122 28756
rect 531222 28704 531228 28756
rect 531280 28744 531286 28756
rect 583386 28744 583392 28756
rect 531280 28716 583392 28744
rect 531280 28704 531286 28716
rect 583386 28704 583392 28716
rect 583444 28704 583450 28756
rect 41690 28636 41696 28688
rect 41748 28676 41754 28688
rect 195238 28676 195244 28688
rect 41748 28648 195244 28676
rect 41748 28636 41754 28648
rect 195238 28636 195244 28648
rect 195296 28636 195302 28688
rect 523034 28636 523040 28688
rect 523092 28676 523098 28688
rect 579706 28676 579712 28688
rect 523092 28648 579712 28676
rect 523092 28636 523098 28648
rect 579706 28636 579712 28648
rect 579764 28636 579770 28688
rect 34790 28568 34796 28620
rect 34848 28608 34854 28620
rect 103790 28608 103796 28620
rect 34848 28580 103796 28608
rect 34848 28568 34854 28580
rect 103790 28568 103796 28580
rect 103848 28568 103854 28620
rect 105630 28568 105636 28620
rect 105688 28608 105694 28620
rect 211338 28608 211344 28620
rect 105688 28580 211344 28608
rect 105688 28568 105694 28580
rect 211338 28568 211344 28580
rect 211396 28568 211402 28620
rect 322106 28568 322112 28620
rect 322164 28608 322170 28620
rect 504174 28608 504180 28620
rect 322164 28580 504180 28608
rect 322164 28568 322170 28580
rect 504174 28568 504180 28580
rect 504232 28568 504238 28620
rect 512086 28568 512092 28620
rect 512144 28608 512150 28620
rect 583202 28608 583208 28620
rect 512144 28580 583208 28608
rect 512144 28568 512150 28580
rect 583202 28568 583208 28580
rect 583260 28568 583266 28620
rect 35434 28500 35440 28552
rect 35492 28540 35498 28552
rect 73522 28540 73528 28552
rect 35492 28512 73528 28540
rect 35492 28500 35498 28512
rect 73522 28500 73528 28512
rect 73580 28500 73586 28552
rect 74626 28500 74632 28552
rect 74684 28540 74690 28552
rect 190730 28540 190736 28552
rect 74684 28512 190736 28540
rect 74684 28500 74690 28512
rect 190730 28500 190736 28512
rect 190788 28500 190794 28552
rect 271230 28500 271236 28552
rect 271288 28540 271294 28552
rect 473998 28540 474004 28552
rect 271288 28512 474004 28540
rect 271288 28500 271294 28512
rect 473998 28500 474004 28512
rect 474056 28500 474062 28552
rect 493410 28500 493416 28552
rect 493468 28540 493474 28552
rect 573174 28540 573180 28552
rect 493468 28512 573180 28540
rect 493468 28500 493474 28512
rect 573174 28500 573180 28512
rect 573232 28500 573238 28552
rect 46750 28432 46756 28484
rect 46808 28472 46814 28484
rect 105078 28472 105084 28484
rect 46808 28444 105084 28472
rect 46808 28432 46814 28444
rect 105078 28432 105084 28444
rect 105136 28432 105142 28484
rect 105538 28432 105544 28484
rect 105596 28472 105602 28484
rect 272518 28472 272524 28484
rect 105596 28444 272524 28472
rect 105596 28432 105602 28444
rect 272518 28432 272524 28444
rect 272576 28432 272582 28484
rect 295702 28432 295708 28484
rect 295760 28472 295766 28484
rect 527818 28472 527824 28484
rect 295760 28444 527824 28472
rect 295760 28432 295766 28444
rect 527818 28432 527824 28444
rect 527876 28432 527882 28484
rect 529474 28432 529480 28484
rect 529532 28472 529538 28484
rect 577406 28472 577412 28484
rect 529532 28444 577412 28472
rect 529532 28432 529538 28444
rect 577406 28432 577412 28444
rect 577464 28432 577470 28484
rect 41322 28364 41328 28416
rect 41380 28404 41386 28416
rect 89622 28404 89628 28416
rect 41380 28376 89628 28404
rect 41380 28364 41386 28376
rect 89622 28364 89628 28376
rect 89680 28364 89686 28416
rect 89714 28364 89720 28416
rect 89772 28404 89778 28416
rect 258994 28404 259000 28416
rect 89772 28376 259000 28404
rect 89772 28364 89778 28376
rect 258994 28364 259000 28376
rect 259052 28364 259058 28416
rect 266078 28364 266084 28416
rect 266136 28404 266142 28416
rect 522298 28404 522304 28416
rect 266136 28376 522304 28404
rect 266136 28364 266142 28376
rect 522298 28364 522304 28376
rect 522356 28364 522362 28416
rect 527174 28364 527180 28416
rect 527232 28404 527238 28416
rect 527232 28376 533384 28404
rect 527232 28364 527238 28376
rect 72510 28296 72516 28348
rect 72568 28336 72574 28348
rect 252554 28336 252560 28348
rect 72568 28308 252560 28336
rect 72568 28296 72574 28308
rect 252554 28296 252560 28308
rect 252612 28296 252618 28348
rect 268010 28296 268016 28348
rect 268068 28336 268074 28348
rect 528554 28336 528560 28348
rect 268068 28308 528560 28336
rect 268068 28296 268074 28308
rect 528554 28296 528560 28308
rect 528612 28296 528618 28348
rect 533356 28336 533384 28376
rect 537202 28364 537208 28416
rect 537260 28404 537266 28416
rect 546862 28404 546868 28416
rect 537260 28376 546868 28404
rect 537260 28364 537266 28376
rect 546862 28364 546868 28376
rect 546920 28364 546926 28416
rect 539502 28336 539508 28348
rect 533356 28308 539508 28336
rect 539502 28296 539508 28308
rect 539560 28296 539566 28348
rect 55582 28228 55588 28280
rect 55640 28268 55646 28280
rect 87690 28268 87696 28280
rect 55640 28240 87696 28268
rect 55640 28228 55646 28240
rect 87690 28228 87696 28240
rect 87748 28228 87754 28280
rect 89070 28228 89076 28280
rect 89128 28268 89134 28280
rect 213270 28268 213276 28280
rect 89128 28240 213276 28268
rect 89128 28228 89134 28240
rect 213270 28228 213276 28240
rect 213328 28228 213334 28280
rect 484394 28228 484400 28280
rect 484452 28268 484458 28280
rect 485038 28268 485044 28280
rect 484452 28240 485044 28268
rect 484452 28228 484458 28240
rect 485038 28228 485044 28240
rect 485096 28228 485102 28280
rect 505646 28228 505652 28280
rect 505704 28268 505710 28280
rect 548886 28268 548892 28280
rect 505704 28240 548892 28268
rect 505704 28228 505710 28240
rect 548886 28228 548892 28240
rect 548944 28228 548950 28280
rect 39114 28160 39120 28212
rect 39172 28200 39178 28212
rect 124398 28200 124404 28212
rect 39172 28172 124404 28200
rect 39172 28160 39178 28172
rect 124398 28160 124404 28172
rect 124456 28160 124462 28212
rect 147674 28160 147680 28212
rect 147732 28200 147738 28212
rect 148870 28200 148876 28212
rect 147732 28172 148876 28200
rect 147732 28160 147738 28172
rect 148870 28160 148876 28172
rect 148928 28160 148934 28212
rect 165614 28160 165620 28212
rect 165672 28200 165678 28212
rect 166258 28200 166264 28212
rect 165672 28172 166264 28200
rect 165672 28160 165678 28172
rect 166258 28160 166264 28172
rect 166316 28160 166322 28212
rect 166994 28160 167000 28212
rect 167052 28200 167058 28212
rect 168190 28200 168196 28212
rect 167052 28172 168196 28200
rect 167052 28160 167058 28172
rect 168190 28160 168196 28172
rect 168248 28160 168254 28212
rect 191834 28160 191840 28212
rect 191892 28200 191898 28212
rect 192662 28200 192668 28212
rect 191892 28172 192668 28200
rect 191892 28160 191898 28172
rect 192662 28160 192668 28172
rect 192720 28160 192726 28212
rect 194686 28160 194692 28212
rect 194744 28200 194750 28212
rect 195882 28200 195888 28212
rect 194744 28172 195888 28200
rect 194744 28160 194750 28172
rect 195882 28160 195888 28172
rect 195940 28160 195946 28212
rect 215294 28160 215300 28212
rect 215352 28200 215358 28212
rect 216490 28200 216496 28212
rect 215352 28172 216496 28200
rect 215352 28160 215358 28172
rect 216490 28160 216496 28172
rect 216548 28160 216554 28212
rect 300854 28160 300860 28212
rect 300912 28200 300918 28212
rect 302142 28200 302148 28212
rect 300912 28172 302148 28200
rect 300912 28160 300918 28172
rect 302142 28160 302148 28172
rect 302200 28160 302206 28212
rect 320174 28160 320180 28212
rect 320232 28200 320238 28212
rect 321462 28200 321468 28212
rect 320232 28172 321468 28200
rect 320232 28160 320238 28172
rect 321462 28160 321468 28172
rect 321520 28160 321526 28212
rect 321554 28160 321560 28212
rect 321612 28200 321618 28212
rect 322750 28200 322756 28212
rect 321612 28172 322756 28200
rect 321612 28160 321618 28172
rect 322750 28160 322756 28172
rect 322808 28160 322814 28212
rect 329834 28160 329840 28212
rect 329892 28200 329898 28212
rect 331122 28200 331128 28212
rect 329892 28172 331128 28200
rect 329892 28160 329898 28172
rect 331122 28160 331128 28172
rect 331180 28160 331186 28212
rect 347774 28160 347780 28212
rect 347832 28200 347838 28212
rect 348510 28200 348516 28212
rect 347832 28172 348516 28200
rect 347832 28160 347838 28172
rect 348510 28160 348516 28172
rect 348568 28160 348574 28212
rect 368474 28160 368480 28212
rect 368532 28200 368538 28212
rect 369762 28200 369768 28212
rect 368532 28172 369768 28200
rect 368532 28160 368538 28172
rect 369762 28160 369768 28172
rect 369820 28160 369826 28212
rect 426434 28160 426440 28212
rect 426492 28200 426498 28212
rect 427722 28200 427728 28212
rect 426492 28172 427728 28200
rect 426492 28160 426498 28172
rect 427722 28160 427728 28172
rect 427780 28160 427786 28212
rect 427814 28160 427820 28212
rect 427872 28200 427878 28212
rect 429010 28200 429016 28212
rect 427872 28172 429016 28200
rect 427872 28160 427878 28172
rect 429010 28160 429016 28172
rect 429068 28160 429074 28212
rect 436094 28160 436100 28212
rect 436152 28200 436158 28212
rect 437382 28200 437388 28212
rect 436152 28172 437388 28200
rect 436152 28160 436158 28172
rect 437382 28160 437388 28172
rect 437440 28160 437446 28212
rect 444374 28160 444380 28212
rect 444432 28200 444438 28212
rect 445110 28200 445116 28212
rect 444432 28172 445116 28200
rect 444432 28160 444438 28172
rect 445110 28160 445116 28172
rect 445168 28160 445174 28212
rect 447134 28160 447140 28212
rect 447192 28200 447198 28212
rect 448330 28200 448336 28212
rect 447192 28172 448336 28200
rect 447192 28160 447198 28172
rect 448330 28160 448336 28172
rect 448388 28160 448394 28212
rect 463694 28160 463700 28212
rect 463752 28200 463758 28212
rect 464430 28200 464436 28212
rect 463752 28172 464436 28200
rect 463752 28160 463758 28172
rect 464430 28160 464436 28172
rect 464488 28160 464494 28212
rect 474826 28160 474832 28212
rect 474884 28200 474890 28212
rect 552658 28200 552664 28212
rect 474884 28172 552664 28200
rect 474884 28160 474890 28172
rect 552658 28160 552664 28172
rect 552716 28160 552722 28212
rect 69750 28092 69756 28144
rect 69808 28132 69814 28144
rect 120534 28132 120540 28144
rect 69808 28104 120540 28132
rect 69808 28092 69814 28104
rect 120534 28092 120540 28104
rect 120592 28092 120598 28144
rect 155954 28092 155960 28144
rect 156012 28132 156018 28144
rect 157242 28132 157248 28144
rect 156012 28104 157248 28132
rect 156012 28092 156018 28104
rect 157242 28092 157248 28104
rect 157300 28092 157306 28144
rect 291194 28092 291200 28144
rect 291252 28132 291258 28144
rect 291838 28132 291844 28144
rect 291252 28104 291844 28132
rect 291252 28092 291258 28104
rect 291838 28092 291844 28104
rect 291896 28092 291902 28144
rect 378134 28092 378140 28144
rect 378192 28132 378198 28144
rect 379422 28132 379428 28144
rect 378192 28104 379428 28132
rect 378192 28092 378198 28104
rect 379422 28092 379428 28104
rect 379480 28092 379486 28144
rect 484486 28092 484492 28144
rect 484544 28132 484550 28144
rect 485682 28132 485688 28144
rect 484544 28104 485688 28132
rect 484544 28092 484550 28104
rect 485682 28092 485688 28104
rect 485740 28092 485746 28144
rect 505094 28092 505100 28144
rect 505152 28132 505158 28144
rect 506290 28132 506296 28144
rect 505152 28104 506296 28132
rect 505152 28092 505158 28104
rect 506290 28092 506296 28104
rect 506348 28092 506354 28144
rect 506382 28092 506388 28144
rect 506440 28132 506446 28144
rect 569954 28132 569960 28144
rect 506440 28104 569960 28132
rect 506440 28092 506446 28104
rect 569954 28092 569960 28104
rect 570012 28092 570018 28144
rect 39390 28024 39396 28076
rect 39448 28064 39454 28076
rect 128906 28064 128912 28076
rect 39448 28036 128912 28064
rect 39448 28024 39454 28036
rect 128906 28024 128912 28036
rect 128964 28024 128970 28076
rect 483106 28024 483112 28076
rect 483164 28064 483170 28076
rect 536834 28064 536840 28076
rect 483164 28036 536840 28064
rect 483164 28024 483170 28036
rect 536834 28024 536840 28036
rect 536892 28024 536898 28076
rect 43990 27956 43996 28008
rect 44048 27996 44054 28008
rect 217778 27996 217784 28008
rect 44048 27968 217784 27996
rect 44048 27956 44054 27968
rect 217778 27956 217784 27968
rect 217836 27956 217842 28008
rect 360102 27956 360108 28008
rect 360160 27996 360166 28008
rect 527174 27996 527180 28008
rect 360160 27968 527180 27996
rect 360160 27956 360166 27968
rect 527174 27956 527180 27968
rect 527232 27956 527238 28008
rect 43806 27888 43812 27940
rect 43864 27928 43870 27940
rect 92198 27928 92204 27940
rect 43864 27900 92204 27928
rect 43864 27888 43870 27900
rect 92198 27888 92204 27900
rect 92256 27888 92262 27940
rect 127618 27888 127624 27940
rect 127676 27928 127682 27940
rect 579982 27928 579988 27940
rect 127676 27900 579988 27928
rect 127676 27888 127682 27900
rect 579982 27888 579988 27900
rect 580040 27888 580046 27940
rect 389082 27820 389088 27872
rect 389140 27860 389146 27872
rect 534718 27860 534724 27872
rect 389140 27832 534724 27860
rect 389140 27820 389146 27832
rect 534718 27820 534724 27832
rect 534776 27820 534782 27872
rect 502334 27752 502340 27804
rect 502392 27792 502398 27804
rect 506382 27792 506388 27804
rect 502392 27764 506388 27792
rect 502392 27752 502398 27764
rect 506382 27752 506388 27764
rect 506440 27752 506446 27804
rect 88978 27616 88984 27668
rect 89036 27656 89042 27668
rect 89622 27656 89628 27668
rect 89036 27628 89628 27656
rect 89036 27616 89042 27628
rect 89622 27616 89628 27628
rect 89680 27616 89686 27668
rect 52178 27548 52184 27600
rect 52236 27588 52242 27600
rect 70302 27588 70308 27600
rect 52236 27560 70308 27588
rect 52236 27548 52242 27560
rect 70302 27548 70308 27560
rect 70360 27548 70366 27600
rect 528186 27548 528192 27600
rect 528244 27588 528250 27600
rect 553026 27588 553032 27600
rect 528244 27560 553032 27588
rect 528244 27548 528250 27560
rect 553026 27548 553032 27560
rect 553084 27548 553090 27600
rect 50890 27480 50896 27532
rect 50948 27520 50954 27532
rect 62574 27520 62580 27532
rect 50948 27492 62580 27520
rect 50948 27480 50954 27492
rect 62574 27480 62580 27492
rect 62632 27480 62638 27532
rect 492766 27480 492772 27532
rect 492824 27520 492830 27532
rect 555326 27520 555332 27532
rect 492824 27492 555332 27520
rect 492824 27480 492830 27492
rect 555326 27480 555332 27492
rect 555384 27480 555390 27532
rect 28810 27412 28816 27464
rect 28868 27452 28874 27464
rect 123754 27452 123760 27464
rect 28868 27424 123760 27452
rect 28868 27412 28874 27424
rect 123754 27412 123760 27424
rect 123812 27412 123818 27464
rect 174630 27412 174636 27464
rect 174688 27452 174694 27464
rect 578326 27452 578332 27464
rect 174688 27424 578332 27452
rect 174688 27412 174694 27424
rect 578326 27412 578332 27424
rect 578384 27412 578390 27464
rect 54478 27344 54484 27396
rect 54536 27384 54542 27396
rect 441246 27384 441252 27396
rect 54536 27356 441252 27384
rect 54536 27344 54542 27356
rect 441246 27344 441252 27356
rect 441304 27344 441310 27396
rect 511442 27344 511448 27396
rect 511500 27384 511506 27396
rect 545298 27384 545304 27396
rect 511500 27356 545304 27384
rect 511500 27344 511506 27356
rect 545298 27344 545304 27356
rect 545356 27344 545362 27396
rect 44450 27276 44456 27328
rect 44508 27316 44514 27328
rect 389726 27316 389732 27328
rect 44508 27288 389732 27316
rect 44508 27276 44514 27288
rect 389726 27276 389732 27288
rect 389784 27276 389790 27328
rect 398742 27276 398748 27328
rect 398800 27316 398806 27328
rect 582834 27316 582840 27328
rect 398800 27288 582840 27316
rect 398800 27276 398806 27288
rect 582834 27276 582840 27288
rect 582892 27276 582898 27328
rect 41874 27208 41880 27260
rect 41932 27248 41938 27260
rect 116670 27248 116676 27260
rect 41932 27220 116676 27248
rect 41932 27208 41938 27220
rect 116670 27208 116676 27220
rect 116728 27208 116734 27260
rect 224218 27208 224224 27260
rect 224276 27248 224282 27260
rect 548610 27248 548616 27260
rect 224276 27220 548616 27248
rect 224276 27208 224282 27220
rect 548610 27208 548616 27220
rect 548668 27208 548674 27260
rect 45186 27140 45192 27192
rect 45244 27180 45250 27192
rect 363966 27180 363972 27192
rect 45244 27152 363972 27180
rect 45244 27140 45250 27152
rect 363966 27140 363972 27152
rect 364024 27140 364030 27192
rect 365898 27140 365904 27192
rect 365956 27180 365962 27192
rect 579890 27180 579896 27192
rect 365956 27152 579896 27180
rect 365956 27140 365962 27152
rect 579890 27140 579896 27152
rect 579948 27140 579954 27192
rect 35618 27072 35624 27124
rect 35676 27112 35682 27124
rect 244182 27112 244188 27124
rect 35676 27084 244188 27112
rect 35676 27072 35682 27084
rect 244182 27072 244188 27084
rect 244240 27072 244246 27124
rect 268654 27072 268660 27124
rect 268712 27112 268718 27124
rect 578602 27112 578608 27124
rect 268712 27084 578608 27112
rect 268712 27072 268718 27084
rect 578602 27072 578608 27084
rect 578660 27072 578666 27124
rect 51994 27004 52000 27056
rect 52052 27044 52058 27056
rect 293126 27044 293132 27056
rect 52052 27016 293132 27044
rect 52052 27004 52058 27016
rect 293126 27004 293132 27016
rect 293184 27004 293190 27056
rect 327258 27004 327264 27056
rect 327316 27044 327322 27056
rect 560662 27044 560668 27056
rect 327316 27016 560668 27044
rect 327316 27004 327322 27016
rect 560662 27004 560668 27016
rect 560720 27004 560726 27056
rect 43622 26936 43628 26988
rect 43680 26976 43686 26988
rect 100570 26976 100576 26988
rect 43680 26948 100576 26976
rect 43680 26936 43686 26948
rect 100570 26936 100576 26948
rect 100628 26936 100634 26988
rect 344002 26936 344008 26988
rect 344060 26976 344066 26988
rect 562134 26976 562140 26988
rect 344060 26948 562140 26976
rect 344060 26936 344066 26948
rect 562134 26936 562140 26948
rect 562192 26936 562198 26988
rect 26878 26868 26884 26920
rect 26936 26908 26942 26920
rect 71774 26908 71780 26920
rect 26936 26880 71780 26908
rect 26936 26868 26942 26880
rect 71774 26868 71780 26880
rect 71832 26868 71838 26920
rect 410334 26868 410340 26920
rect 410392 26908 410398 26920
rect 556798 26908 556804 26920
rect 410392 26880 556804 26908
rect 410392 26868 410398 26880
rect 556798 26868 556804 26880
rect 556856 26868 556862 26920
rect 417418 26800 417424 26852
rect 417476 26840 417482 26852
rect 560386 26840 560392 26852
rect 417476 26812 560392 26840
rect 417476 26800 417482 26812
rect 560386 26800 560392 26812
rect 560444 26800 560450 26852
rect 409690 26732 409696 26784
rect 409748 26772 409754 26784
rect 540882 26772 540888 26784
rect 409748 26744 540888 26772
rect 409748 26732 409754 26744
rect 540882 26732 540888 26744
rect 540940 26732 540946 26784
rect 42058 26664 42064 26716
rect 42116 26704 42122 26716
rect 473446 26704 473452 26716
rect 42116 26676 473452 26704
rect 42116 26664 42122 26676
rect 473446 26664 473452 26676
rect 473504 26664 473510 26716
rect 516594 26664 516600 26716
rect 516652 26704 516658 26716
rect 574830 26704 574836 26716
rect 516652 26676 574836 26704
rect 516652 26664 516658 26676
rect 574830 26664 574836 26676
rect 574888 26664 574894 26716
rect 37642 26596 37648 26648
rect 37700 26636 37706 26648
rect 520458 26636 520464 26648
rect 37700 26608 520464 26636
rect 37700 26596 37706 26608
rect 520458 26596 520464 26608
rect 520516 26596 520522 26648
rect 27430 26188 27436 26240
rect 27488 26228 27494 26240
rect 523034 26228 523040 26240
rect 27488 26200 523040 26228
rect 27488 26188 27494 26200
rect 523034 26188 523040 26200
rect 523092 26188 523098 26240
rect 538214 26188 538220 26240
rect 538272 26228 538278 26240
rect 555694 26228 555700 26240
rect 538272 26200 555700 26228
rect 538272 26188 538278 26200
rect 555694 26188 555700 26200
rect 555752 26188 555758 26240
rect 35710 26120 35716 26172
rect 35768 26160 35774 26172
rect 494054 26160 494060 26172
rect 35768 26132 494060 26160
rect 35768 26120 35774 26132
rect 494054 26120 494060 26132
rect 494112 26120 494118 26172
rect 509234 26120 509240 26172
rect 509292 26160 509298 26172
rect 574554 26160 574560 26172
rect 509292 26132 574560 26160
rect 509292 26120 509298 26132
rect 574554 26120 574560 26132
rect 574612 26120 574618 26172
rect 29822 26052 29828 26104
rect 29880 26092 29886 26104
rect 470870 26092 470876 26104
rect 29880 26064 470876 26092
rect 29880 26052 29886 26064
rect 470870 26052 470876 26064
rect 470928 26052 470934 26104
rect 476206 26052 476212 26104
rect 476264 26092 476270 26104
rect 553118 26092 553124 26104
rect 476264 26064 553124 26092
rect 476264 26052 476270 26064
rect 553118 26052 553124 26064
rect 553176 26052 553182 26104
rect 20254 25984 20260 26036
rect 20312 26024 20318 26036
rect 391934 26024 391940 26036
rect 20312 25996 391940 26024
rect 20312 25984 20318 25996
rect 391934 25984 391940 25996
rect 391992 25984 391998 26036
rect 423674 25984 423680 26036
rect 423732 26024 423738 26036
rect 567654 26024 567660 26036
rect 423732 25996 567660 26024
rect 423732 25984 423738 25996
rect 567654 25984 567660 25996
rect 567712 25984 567718 26036
rect 40862 25916 40868 25968
rect 40920 25956 40926 25968
rect 387794 25956 387800 25968
rect 40920 25928 387800 25956
rect 40920 25916 40926 25928
rect 387794 25916 387800 25928
rect 387852 25916 387858 25968
rect 389266 25916 389272 25968
rect 389324 25956 389330 25968
rect 580074 25956 580080 25968
rect 389324 25928 580080 25956
rect 389324 25916 389330 25928
rect 580074 25916 580080 25928
rect 580132 25916 580138 25968
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 213914 25888 213920 25900
rect 23164 25860 213920 25888
rect 23164 25848 23170 25860
rect 213914 25848 213920 25860
rect 213972 25848 213978 25900
rect 280154 25848 280160 25900
rect 280212 25888 280218 25900
rect 575842 25888 575848 25900
rect 280212 25860 575848 25888
rect 280212 25848 280218 25860
rect 575842 25848 575848 25860
rect 575900 25848 575906 25900
rect 59722 25780 59728 25832
rect 59780 25820 59786 25832
rect 211246 25820 211252 25832
rect 59780 25792 211252 25820
rect 59780 25780 59786 25792
rect 211246 25780 211252 25792
rect 211304 25780 211310 25832
rect 322934 25780 322940 25832
rect 322992 25820 322998 25832
rect 578510 25820 578516 25832
rect 322992 25792 578516 25820
rect 322992 25780 322998 25792
rect 578510 25780 578516 25792
rect 578568 25780 578574 25832
rect 32122 25712 32128 25764
rect 32180 25752 32186 25764
rect 165706 25752 165712 25764
rect 32180 25724 165712 25752
rect 32180 25712 32186 25724
rect 165706 25712 165712 25724
rect 165764 25712 165770 25764
rect 325786 25712 325792 25764
rect 325844 25752 325850 25764
rect 578418 25752 578424 25764
rect 325844 25724 578424 25752
rect 325844 25712 325850 25724
rect 578418 25712 578424 25724
rect 578476 25712 578482 25764
rect 33594 25644 33600 25696
rect 33652 25684 33658 25696
rect 156046 25684 156052 25696
rect 33652 25656 156052 25684
rect 33652 25644 33658 25656
rect 156046 25644 156052 25656
rect 156104 25644 156110 25696
rect 430574 25644 430580 25696
rect 430632 25684 430638 25696
rect 540698 25684 540704 25696
rect 430632 25656 540704 25684
rect 430632 25644 430638 25656
rect 540698 25644 540704 25656
rect 540756 25644 540762 25696
rect 22554 25576 22560 25628
rect 22612 25616 22618 25628
rect 131206 25616 131212 25628
rect 22612 25588 131212 25616
rect 22612 25576 22618 25588
rect 131206 25576 131212 25588
rect 131264 25576 131270 25628
rect 477494 25576 477500 25628
rect 477552 25616 477558 25628
rect 572990 25616 572996 25628
rect 477552 25588 572996 25616
rect 477552 25576 477558 25588
rect 572990 25576 572996 25588
rect 573048 25576 573054 25628
rect 53558 25508 53564 25560
rect 53616 25548 53622 25560
rect 100754 25548 100760 25560
rect 53616 25520 100760 25548
rect 53616 25508 53622 25520
rect 100754 25508 100760 25520
rect 100812 25508 100818 25560
rect 396074 25508 396080 25560
rect 396132 25548 396138 25560
rect 547690 25548 547696 25560
rect 396132 25520 547696 25548
rect 396132 25508 396138 25520
rect 547690 25508 547696 25520
rect 547748 25508 547754 25560
rect 52270 25440 52276 25492
rect 52328 25480 52334 25492
rect 97994 25480 98000 25492
rect 52328 25452 98000 25480
rect 52328 25440 52334 25452
rect 97994 25440 98000 25452
rect 98052 25440 98058 25492
rect 513374 25440 513380 25492
rect 513432 25480 513438 25492
rect 569034 25480 569040 25492
rect 513432 25452 569040 25480
rect 513432 25440 513438 25452
rect 569034 25440 569040 25452
rect 569092 25440 569098 25492
rect 53650 25372 53656 25424
rect 53708 25412 53714 25424
rect 81434 25412 81440 25424
rect 53708 25384 81440 25412
rect 53708 25372 53714 25384
rect 81434 25372 81440 25384
rect 81492 25372 81498 25424
rect 520274 25372 520280 25424
rect 520332 25412 520338 25424
rect 571518 25412 571524 25424
rect 520332 25384 571524 25412
rect 520332 25372 520338 25384
rect 571518 25372 571524 25384
rect 571576 25372 571582 25424
rect 54294 25304 54300 25356
rect 54352 25344 54358 25356
rect 77294 25344 77300 25356
rect 54352 25316 77300 25344
rect 54352 25304 54358 25316
rect 77294 25304 77300 25316
rect 77352 25304 77358 25356
rect 516134 25304 516140 25356
rect 516192 25344 516198 25356
rect 568114 25344 568120 25356
rect 516192 25316 568120 25344
rect 516192 25304 516198 25316
rect 568114 25304 568120 25316
rect 568172 25304 568178 25356
rect 49050 24760 49056 24812
rect 49108 24800 49114 24812
rect 191926 24800 191932 24812
rect 49108 24772 191932 24800
rect 49108 24760 49114 24772
rect 191926 24760 191932 24772
rect 191984 24760 191990 24812
rect 534718 24760 534724 24812
rect 534776 24800 534782 24812
rect 544010 24800 544016 24812
rect 534776 24772 544016 24800
rect 534776 24760 534782 24772
rect 544010 24760 544016 24772
rect 544068 24760 544074 24812
rect 54202 24692 54208 24744
rect 54260 24732 54266 24744
rect 397454 24732 397460 24744
rect 54260 24704 397460 24732
rect 54260 24692 54266 24704
rect 397454 24692 397460 24704
rect 397512 24692 397518 24744
rect 409874 24692 409880 24744
rect 409932 24732 409938 24744
rect 555418 24732 555424 24744
rect 409932 24704 555424 24732
rect 409932 24692 409938 24704
rect 555418 24692 555424 24704
rect 555476 24692 555482 24744
rect 36998 24624 37004 24676
rect 37056 24664 37062 24676
rect 325694 24664 325700 24676
rect 37056 24636 325700 24664
rect 37056 24624 37062 24636
rect 325694 24624 325700 24636
rect 325752 24624 325758 24676
rect 385126 24624 385132 24676
rect 385184 24664 385190 24676
rect 580350 24664 580356 24676
rect 385184 24636 580356 24664
rect 385184 24624 385190 24636
rect 580350 24624 580356 24636
rect 580408 24624 580414 24676
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 285674 24596 285680 24608
rect 21968 24568 285680 24596
rect 21968 24556 21974 24568
rect 285674 24556 285680 24568
rect 285732 24556 285738 24608
rect 465166 24556 465172 24608
rect 465224 24596 465230 24608
rect 561766 24596 561772 24608
rect 465224 24568 561772 24596
rect 465224 24556 465230 24568
rect 561766 24556 561772 24568
rect 561824 24556 561830 24608
rect 47670 24488 47676 24540
rect 47728 24528 47734 24540
rect 291286 24528 291292 24540
rect 47728 24500 291292 24528
rect 47728 24488 47734 24500
rect 291286 24488 291292 24500
rect 291344 24488 291350 24540
rect 502518 24488 502524 24540
rect 502576 24528 502582 24540
rect 582650 24528 582656 24540
rect 502576 24500 582656 24528
rect 502576 24488 502582 24500
rect 582650 24488 582656 24500
rect 582708 24488 582714 24540
rect 24210 24420 24216 24472
rect 24268 24460 24274 24472
rect 266354 24460 266360 24472
rect 24268 24432 266360 24460
rect 24268 24420 24274 24432
rect 266354 24420 266360 24432
rect 266412 24420 266418 24472
rect 465258 24420 465264 24472
rect 465316 24460 465322 24472
rect 541066 24460 541072 24472
rect 465316 24432 541072 24460
rect 465316 24420 465322 24432
rect 541066 24420 541072 24432
rect 541124 24420 541130 24472
rect 31202 24352 31208 24404
rect 31260 24392 31266 24404
rect 256694 24392 256700 24404
rect 31260 24364 256700 24392
rect 31260 24352 31266 24364
rect 256694 24352 256700 24364
rect 256752 24352 256758 24404
rect 503714 24352 503720 24404
rect 503772 24392 503778 24404
rect 555234 24392 555240 24404
rect 503772 24364 555240 24392
rect 503772 24352 503778 24364
rect 555234 24352 555240 24364
rect 555292 24352 555298 24404
rect 33778 24284 33784 24336
rect 33836 24324 33842 24336
rect 219434 24324 219440 24336
rect 33836 24296 219440 24324
rect 33836 24284 33842 24296
rect 219434 24284 219440 24296
rect 219492 24284 219498 24336
rect 502426 24284 502432 24336
rect 502484 24324 502490 24336
rect 548426 24324 548432 24336
rect 502484 24296 548432 24324
rect 502484 24284 502490 24296
rect 548426 24284 548432 24296
rect 548484 24284 548490 24336
rect 44818 24216 44824 24268
rect 44876 24256 44882 24268
rect 219526 24256 219532 24268
rect 44876 24228 219532 24256
rect 44876 24216 44882 24228
rect 219526 24216 219532 24228
rect 219584 24216 219590 24268
rect 245654 24216 245660 24268
rect 245712 24256 245718 24268
rect 564894 24256 564900 24268
rect 245712 24228 564900 24256
rect 245712 24216 245718 24228
rect 564894 24216 564900 24228
rect 564952 24216 564958 24268
rect 51902 24148 51908 24200
rect 51960 24188 51966 24200
rect 209774 24188 209780 24200
rect 51960 24160 209780 24188
rect 51960 24148 51966 24160
rect 209774 24148 209780 24160
rect 209832 24148 209838 24200
rect 220814 24148 220820 24200
rect 220872 24188 220878 24200
rect 568666 24188 568672 24200
rect 220872 24160 568672 24188
rect 220872 24148 220878 24160
rect 568666 24148 568672 24160
rect 568724 24148 568730 24200
rect 55490 24080 55496 24132
rect 55548 24120 55554 24132
rect 197354 24120 197360 24132
rect 55548 24092 197360 24120
rect 55548 24080 55554 24092
rect 197354 24080 197360 24092
rect 197412 24080 197418 24132
rect 209866 24080 209872 24132
rect 209924 24120 209930 24132
rect 566182 24120 566188 24132
rect 209924 24092 566188 24120
rect 209924 24080 209930 24092
rect 566182 24080 566188 24092
rect 566240 24080 566246 24132
rect 47762 24012 47768 24064
rect 47820 24052 47826 24064
rect 161474 24052 161480 24064
rect 47820 24024 161480 24052
rect 47820 24012 47826 24024
rect 161474 24012 161480 24024
rect 161532 24012 161538 24064
rect 510614 24012 510620 24064
rect 510672 24052 510678 24064
rect 551646 24052 551652 24064
rect 510672 24024 551652 24052
rect 510672 24012 510678 24024
rect 551646 24012 551652 24024
rect 551704 24012 551710 24064
rect 53466 23944 53472 23996
rect 53524 23984 53530 23996
rect 142154 23984 142160 23996
rect 53524 23956 142160 23984
rect 53524 23944 53530 23956
rect 142154 23944 142160 23956
rect 142212 23944 142218 23996
rect 171134 23944 171140 23996
rect 171192 23984 171198 23996
rect 578234 23984 578240 23996
rect 171192 23956 578240 23984
rect 171192 23944 171198 23956
rect 578234 23944 578240 23956
rect 578292 23944 578298 23996
rect 51534 23876 51540 23928
rect 51592 23916 51598 23928
rect 95326 23916 95332 23928
rect 51592 23888 95332 23916
rect 51592 23876 51598 23888
rect 95326 23876 95332 23888
rect 95384 23876 95390 23928
rect 503714 23468 503720 23520
rect 503772 23508 503778 23520
rect 504358 23508 504364 23520
rect 503772 23480 504364 23508
rect 503772 23468 503778 23480
rect 504358 23468 504364 23480
rect 504416 23468 504422 23520
rect 48038 23400 48044 23452
rect 48096 23440 48102 23452
rect 69750 23440 69756 23452
rect 48096 23412 69756 23440
rect 48096 23400 48102 23412
rect 69750 23400 69756 23412
rect 69808 23400 69814 23452
rect 138014 23400 138020 23452
rect 138072 23440 138078 23452
rect 581086 23440 581092 23452
rect 138072 23412 581092 23440
rect 138072 23400 138078 23412
rect 581086 23400 581092 23412
rect 581144 23400 581150 23452
rect 185026 23332 185032 23384
rect 185084 23372 185090 23384
rect 581362 23372 581368 23384
rect 185084 23344 581368 23372
rect 185084 23332 185090 23344
rect 581362 23332 581368 23344
rect 581420 23332 581426 23384
rect 38470 23264 38476 23316
rect 38528 23304 38534 23316
rect 426526 23304 426532 23316
rect 38528 23276 426532 23304
rect 38528 23264 38534 23276
rect 426526 23264 426532 23276
rect 426584 23264 426590 23316
rect 434806 23264 434812 23316
rect 434864 23304 434870 23316
rect 564618 23304 564624 23316
rect 434864 23276 564624 23304
rect 434864 23264 434870 23276
rect 564618 23264 564624 23276
rect 564676 23264 564682 23316
rect 38562 23196 38568 23248
rect 38620 23236 38626 23248
rect 382274 23236 382280 23248
rect 38620 23208 382280 23236
rect 38620 23196 38626 23208
rect 382274 23196 382280 23208
rect 382332 23196 382338 23248
rect 383654 23196 383660 23248
rect 383712 23236 383718 23248
rect 574646 23236 574652 23248
rect 383712 23208 574652 23236
rect 383712 23196 383718 23208
rect 574646 23196 574652 23208
rect 574704 23196 574710 23248
rect 50062 23128 50068 23180
rect 50120 23168 50126 23180
rect 368474 23168 368480 23180
rect 50120 23140 368480 23168
rect 50120 23128 50126 23140
rect 368474 23128 368480 23140
rect 368532 23128 368538 23180
rect 376754 23128 376760 23180
rect 376812 23168 376818 23180
rect 576946 23168 576952 23180
rect 376812 23140 576952 23168
rect 376812 23128 376818 23140
rect 576946 23128 576952 23140
rect 577004 23128 577010 23180
rect 25682 23060 25688 23112
rect 25740 23100 25746 23112
rect 306374 23100 306380 23112
rect 25740 23072 306380 23100
rect 25740 23060 25746 23072
rect 306374 23060 306380 23072
rect 306432 23060 306438 23112
rect 361574 23060 361580 23112
rect 361632 23100 361638 23112
rect 552934 23100 552940 23112
rect 361632 23072 552940 23100
rect 361632 23060 361638 23072
rect 552934 23060 552940 23072
rect 552992 23060 552998 23112
rect 27154 22992 27160 23044
rect 27212 23032 27218 23044
rect 307754 23032 307760 23044
rect 27212 23004 307760 23032
rect 27212 22992 27218 23004
rect 307754 22992 307760 23004
rect 307812 22992 307818 23044
rect 447134 22992 447140 23044
rect 447192 23032 447198 23044
rect 565078 23032 565084 23044
rect 447192 23004 565084 23032
rect 447192 22992 447198 23004
rect 565078 22992 565084 23004
rect 565136 22992 565142 23044
rect 47302 22924 47308 22976
rect 47360 22964 47366 22976
rect 324314 22964 324320 22976
rect 47360 22936 324320 22964
rect 47360 22924 47366 22936
rect 324314 22924 324320 22936
rect 324372 22924 324378 22976
rect 484486 22924 484492 22976
rect 484544 22964 484550 22976
rect 563606 22964 563612 22976
rect 484544 22936 563612 22964
rect 484544 22924 484550 22936
rect 563606 22924 563612 22936
rect 563664 22924 563670 22976
rect 50706 22856 50712 22908
rect 50764 22896 50770 22908
rect 296714 22896 296720 22908
rect 50764 22868 296720 22896
rect 50764 22856 50770 22868
rect 296714 22856 296720 22868
rect 296772 22856 296778 22908
rect 434714 22856 434720 22908
rect 434772 22896 434778 22908
rect 559098 22896 559104 22908
rect 434772 22868 559104 22896
rect 434772 22856 434778 22868
rect 559098 22856 559104 22868
rect 559156 22856 559162 22908
rect 40954 22788 40960 22840
rect 41012 22828 41018 22840
rect 183554 22828 183560 22840
rect 41012 22800 183560 22828
rect 41012 22788 41018 22800
rect 183554 22788 183560 22800
rect 183612 22788 183618 22840
rect 389174 22788 389180 22840
rect 389232 22828 389238 22840
rect 556338 22828 556344 22840
rect 389232 22800 556344 22828
rect 389232 22788 389238 22800
rect 556338 22788 556344 22800
rect 556396 22788 556402 22840
rect 39666 22720 39672 22772
rect 39724 22760 39730 22772
rect 182174 22760 182180 22772
rect 39724 22732 182180 22760
rect 39724 22720 39730 22732
rect 182174 22720 182180 22732
rect 182232 22720 182238 22772
rect 360194 22720 360200 22772
rect 360252 22760 360258 22772
rect 547598 22760 547604 22772
rect 360252 22732 547604 22760
rect 360252 22720 360258 22732
rect 547598 22720 547604 22732
rect 547656 22720 547662 22772
rect 57238 22652 57244 22704
rect 57296 22692 57302 22704
rect 116026 22692 116032 22704
rect 57296 22664 116032 22692
rect 57296 22652 57302 22664
rect 116026 22652 116032 22664
rect 116084 22652 116090 22704
rect 498194 22652 498200 22704
rect 498252 22692 498258 22704
rect 545666 22692 545672 22704
rect 498252 22664 545672 22692
rect 498252 22652 498258 22664
rect 545666 22652 545672 22664
rect 545724 22652 545730 22704
rect 46842 22584 46848 22636
rect 46900 22624 46906 22636
rect 102134 22624 102140 22636
rect 46900 22596 102140 22624
rect 46900 22584 46906 22596
rect 102134 22584 102140 22596
rect 102192 22584 102198 22636
rect 31386 22516 31392 22568
rect 31444 22556 31450 22568
rect 131114 22556 131120 22568
rect 31444 22528 131120 22556
rect 31444 22516 31450 22528
rect 131114 22516 131120 22528
rect 131172 22516 131178 22568
rect 41046 22448 41052 22500
rect 41104 22488 41110 22500
rect 193214 22488 193220 22500
rect 41104 22460 193220 22488
rect 41104 22448 41110 22460
rect 193214 22448 193220 22460
rect 193272 22448 193278 22500
rect 56042 22040 56048 22092
rect 56100 22080 56106 22092
rect 69566 22080 69572 22092
rect 56100 22052 69572 22080
rect 56100 22040 56106 22052
rect 69566 22040 69572 22052
rect 69624 22040 69630 22092
rect 26142 21972 26148 22024
rect 26200 22012 26206 22024
rect 448606 22012 448612 22024
rect 26200 21984 448612 22012
rect 26200 21972 26206 21984
rect 448606 21972 448612 21984
rect 448664 21972 448670 22024
rect 488534 21972 488540 22024
rect 488592 22012 488598 22024
rect 577498 22012 577504 22024
rect 488592 21984 577504 22012
rect 488592 21972 488598 21984
rect 577498 21972 577504 21984
rect 577556 21972 577562 22024
rect 49142 21904 49148 21956
rect 49200 21944 49206 21956
rect 411254 21944 411260 21956
rect 49200 21916 411260 21944
rect 49200 21904 49206 21916
rect 411254 21904 411260 21916
rect 411312 21904 411318 21956
rect 420914 21904 420920 21956
rect 420972 21944 420978 21956
rect 552198 21944 552204 21956
rect 420972 21916 552204 21944
rect 420972 21904 420978 21916
rect 552198 21904 552204 21916
rect 552256 21904 552262 21956
rect 53098 21836 53104 21888
rect 53156 21876 53162 21888
rect 400214 21876 400220 21888
rect 53156 21848 400220 21876
rect 53156 21836 53162 21848
rect 400214 21836 400220 21848
rect 400272 21836 400278 21888
rect 419534 21836 419540 21888
rect 419592 21876 419598 21888
rect 543918 21876 543924 21888
rect 419592 21848 543924 21876
rect 419592 21836 419598 21848
rect 543918 21836 543924 21848
rect 543976 21836 543982 21888
rect 46474 21768 46480 21820
rect 46532 21808 46538 21820
rect 270494 21808 270500 21820
rect 46532 21780 270500 21808
rect 46532 21768 46538 21780
rect 270494 21768 270500 21780
rect 270552 21768 270558 21820
rect 523034 21768 523040 21820
rect 523092 21808 523098 21820
rect 575658 21808 575664 21820
rect 523092 21780 575664 21808
rect 523092 21768 523098 21780
rect 575658 21768 575664 21780
rect 575716 21768 575722 21820
rect 37918 21700 37924 21752
rect 37976 21740 37982 21752
rect 229094 21740 229100 21752
rect 37976 21712 229100 21740
rect 37976 21700 37982 21712
rect 229094 21700 229100 21712
rect 229152 21700 229158 21752
rect 470594 21700 470600 21752
rect 470652 21740 470658 21752
rect 556154 21740 556160 21752
rect 470652 21712 556160 21740
rect 470652 21700 470658 21712
rect 556154 21700 556160 21712
rect 556212 21700 556218 21752
rect 48866 21632 48872 21684
rect 48924 21672 48930 21684
rect 205634 21672 205640 21684
rect 48924 21644 205640 21672
rect 48924 21632 48930 21644
rect 205634 21632 205640 21644
rect 205692 21632 205698 21684
rect 416774 21632 416780 21684
rect 416832 21672 416838 21684
rect 557810 21672 557816 21684
rect 416832 21644 557816 21672
rect 416832 21632 416838 21644
rect 557810 21632 557816 21644
rect 557868 21632 557874 21684
rect 49510 21564 49516 21616
rect 49568 21604 49574 21616
rect 179414 21604 179420 21616
rect 49568 21576 179420 21604
rect 49568 21564 49574 21576
rect 179414 21564 179420 21576
rect 179472 21564 179478 21616
rect 407114 21564 407120 21616
rect 407172 21604 407178 21616
rect 555786 21604 555792 21616
rect 407172 21576 555792 21604
rect 407172 21564 407178 21576
rect 555786 21564 555792 21576
rect 555844 21564 555850 21616
rect 36906 21496 36912 21548
rect 36964 21536 36970 21548
rect 147674 21536 147680 21548
rect 36964 21508 147680 21536
rect 36964 21496 36970 21508
rect 147674 21496 147680 21508
rect 147732 21496 147738 21548
rect 249794 21496 249800 21548
rect 249852 21536 249858 21548
rect 568942 21536 568948 21548
rect 249852 21508 568948 21536
rect 249852 21496 249858 21508
rect 568942 21496 568948 21508
rect 569000 21496 569006 21548
rect 53374 21428 53380 21480
rect 53432 21468 53438 21480
rect 155954 21468 155960 21480
rect 53432 21440 155960 21468
rect 53432 21428 53438 21440
rect 155954 21428 155960 21440
rect 156012 21428 156018 21480
rect 229094 21428 229100 21480
rect 229152 21468 229158 21480
rect 574370 21468 574376 21480
rect 229152 21440 574376 21468
rect 229152 21428 229158 21440
rect 574370 21428 574376 21440
rect 574428 21428 574434 21480
rect 40218 21360 40224 21412
rect 40276 21400 40282 21412
rect 139394 21400 139400 21412
rect 40276 21372 139400 21400
rect 40276 21360 40282 21372
rect 139394 21360 139400 21372
rect 139452 21360 139458 21412
rect 176654 21360 176660 21412
rect 176712 21400 176718 21412
rect 572898 21400 572904 21412
rect 176712 21372 572904 21400
rect 176712 21360 176718 21372
rect 572898 21360 572904 21372
rect 572956 21360 572962 21412
rect 55858 21292 55864 21344
rect 55916 21332 55922 21344
rect 140774 21332 140780 21344
rect 55916 21304 140780 21332
rect 55916 21292 55922 21304
rect 140774 21292 140780 21304
rect 140832 21292 140838 21344
rect 58710 21224 58716 21276
rect 58768 21264 58774 21276
rect 128446 21264 128452 21276
rect 58768 21236 128452 21264
rect 58768 21224 58774 21236
rect 128446 21224 128452 21236
rect 128504 21224 128510 21276
rect 17770 21156 17776 21208
rect 17828 21196 17834 21208
rect 505094 21196 505100 21208
rect 17828 21168 505100 21196
rect 17828 21156 17834 21168
rect 505094 21156 505100 21168
rect 505152 21156 505158 21208
rect 179414 20816 179420 20868
rect 179472 20856 179478 20868
rect 569954 20856 569960 20868
rect 179472 20828 569960 20856
rect 179472 20816 179478 20828
rect 569954 20816 569960 20828
rect 570012 20816 570018 20868
rect 161474 20748 161480 20800
rect 161532 20788 161538 20800
rect 560294 20788 560300 20800
rect 161532 20760 560300 20788
rect 161532 20748 161538 20760
rect 560294 20748 560300 20760
rect 560352 20748 560358 20800
rect 135254 20680 135260 20732
rect 135312 20720 135318 20732
rect 571426 20720 571432 20732
rect 135312 20692 571432 20720
rect 135312 20680 135318 20692
rect 571426 20680 571432 20692
rect 571484 20680 571490 20732
rect 20346 20612 20352 20664
rect 20404 20652 20410 20664
rect 458174 20652 458180 20664
rect 20404 20624 458180 20652
rect 20404 20612 20410 20624
rect 458174 20612 458180 20624
rect 458232 20612 458238 20664
rect 527174 20612 527180 20664
rect 527232 20652 527238 20664
rect 547230 20652 547236 20664
rect 527232 20624 547236 20652
rect 527232 20612 527238 20624
rect 547230 20612 547236 20624
rect 547288 20612 547294 20664
rect 28534 20544 28540 20596
rect 28592 20584 28598 20596
rect 462314 20584 462320 20596
rect 28592 20556 462320 20584
rect 28592 20544 28598 20556
rect 462314 20544 462320 20556
rect 462372 20544 462378 20596
rect 469214 20544 469220 20596
rect 469272 20584 469278 20596
rect 567470 20584 567476 20596
rect 469272 20556 567476 20584
rect 469272 20544 469278 20556
rect 567470 20544 567476 20556
rect 567528 20544 567534 20596
rect 19058 20476 19064 20528
rect 19116 20516 19122 20528
rect 364426 20516 364432 20528
rect 19116 20488 364432 20516
rect 19116 20476 19122 20488
rect 364426 20476 364432 20488
rect 364484 20476 364490 20528
rect 449894 20476 449900 20528
rect 449952 20516 449958 20528
rect 558086 20516 558092 20528
rect 449952 20488 558092 20516
rect 449952 20476 449958 20488
rect 558086 20476 558092 20488
rect 558144 20476 558150 20528
rect 25498 20408 25504 20460
rect 25556 20448 25562 20460
rect 356054 20448 356060 20460
rect 25556 20420 356060 20448
rect 25556 20408 25562 20420
rect 356054 20408 356060 20420
rect 356112 20408 356118 20460
rect 459554 20408 459560 20460
rect 459612 20448 459618 20460
rect 544286 20448 544292 20460
rect 459612 20420 544292 20448
rect 459612 20408 459618 20420
rect 544286 20408 544292 20420
rect 544344 20408 544350 20460
rect 27522 20340 27528 20392
rect 27580 20380 27586 20392
rect 354674 20380 354680 20392
rect 27580 20352 354680 20380
rect 27580 20340 27586 20352
rect 354674 20340 354680 20352
rect 354732 20340 354738 20392
rect 477586 20340 477592 20392
rect 477644 20380 477650 20392
rect 554038 20380 554044 20392
rect 477644 20352 554044 20380
rect 477644 20340 477650 20352
rect 554038 20340 554044 20352
rect 554096 20340 554102 20392
rect 23014 20272 23020 20324
rect 23072 20312 23078 20324
rect 342254 20312 342260 20324
rect 23072 20284 342260 20312
rect 23072 20272 23078 20284
rect 342254 20272 342260 20284
rect 342312 20272 342318 20324
rect 463694 20272 463700 20324
rect 463752 20312 463758 20324
rect 540054 20312 540060 20324
rect 463752 20284 540060 20312
rect 463752 20272 463758 20284
rect 540054 20272 540060 20284
rect 540112 20272 540118 20324
rect 19150 20204 19156 20256
rect 19208 20244 19214 20256
rect 333974 20244 333980 20256
rect 19208 20216 333980 20244
rect 19208 20204 19214 20216
rect 333974 20204 333980 20216
rect 334032 20204 334038 20256
rect 474734 20204 474740 20256
rect 474792 20244 474798 20256
rect 551094 20244 551100 20256
rect 474792 20216 551100 20244
rect 474792 20204 474798 20216
rect 551094 20204 551100 20216
rect 551152 20204 551158 20256
rect 18874 20136 18880 20188
rect 18932 20176 18938 20188
rect 311894 20176 311900 20188
rect 18932 20148 311900 20176
rect 18932 20136 18938 20148
rect 311894 20136 311900 20148
rect 311952 20136 311958 20188
rect 452654 20136 452660 20188
rect 452712 20176 452718 20188
rect 557718 20176 557724 20188
rect 452712 20148 557724 20176
rect 452712 20136 452718 20148
rect 557718 20136 557724 20148
rect 557776 20136 557782 20188
rect 44726 20068 44732 20120
rect 44784 20108 44790 20120
rect 202874 20108 202880 20120
rect 44784 20080 202880 20108
rect 44784 20068 44790 20080
rect 202874 20068 202880 20080
rect 202932 20068 202938 20120
rect 427906 20068 427912 20120
rect 427964 20108 427970 20120
rect 543182 20108 543188 20120
rect 427964 20080 543188 20108
rect 427964 20068 427970 20080
rect 543182 20068 543188 20080
rect 543240 20068 543246 20120
rect 59814 20000 59820 20052
rect 59872 20040 59878 20052
rect 216766 20040 216772 20052
rect 59872 20012 216772 20040
rect 59872 20000 59878 20012
rect 216766 20000 216772 20012
rect 216824 20000 216830 20052
rect 296714 20000 296720 20052
rect 296772 20040 296778 20052
rect 563698 20040 563704 20052
rect 296772 20012 563704 20040
rect 296772 20000 296778 20012
rect 563698 20000 563704 20012
rect 563756 20000 563762 20052
rect 33042 19932 33048 19984
rect 33100 19972 33106 19984
rect 166994 19972 167000 19984
rect 33100 19944 167000 19972
rect 33100 19932 33106 19944
rect 166994 19932 167000 19944
rect 167052 19932 167058 19984
rect 271874 19932 271880 19984
rect 271932 19972 271938 19984
rect 556706 19972 556712 19984
rect 271932 19944 556712 19972
rect 271932 19932 271938 19944
rect 556706 19932 556712 19944
rect 556764 19932 556770 19984
rect 38102 19864 38108 19916
rect 38160 19904 38166 19916
rect 149054 19904 149060 19916
rect 38160 19876 149060 19904
rect 38160 19864 38166 19876
rect 149054 19864 149060 19876
rect 149112 19864 149118 19916
rect 504174 19864 504180 19916
rect 504232 19904 504238 19916
rect 544654 19904 544660 19916
rect 504232 19876 544660 19904
rect 504232 19864 504238 19876
rect 544654 19864 544660 19876
rect 544712 19864 544718 19916
rect 37090 19796 37096 19848
rect 37148 19836 37154 19848
rect 125594 19836 125600 19848
rect 37148 19808 125600 19836
rect 37148 19796 37154 19808
rect 125594 19796 125600 19808
rect 125652 19796 125658 19848
rect 533338 19796 533344 19848
rect 533396 19836 533402 19848
rect 550082 19836 550088 19848
rect 533396 19808 550088 19836
rect 533396 19796 533402 19808
rect 550082 19796 550088 19808
rect 550140 19796 550146 19848
rect 41138 19728 41144 19780
rect 41196 19768 41202 19780
rect 95234 19768 95240 19780
rect 41196 19740 95240 19768
rect 41196 19728 41202 19740
rect 95234 19728 95240 19740
rect 95292 19728 95298 19780
rect 461026 19728 461032 19780
rect 461084 19768 461090 19780
rect 562226 19768 562232 19780
rect 461084 19740 562232 19768
rect 461084 19728 461090 19740
rect 562226 19728 562232 19740
rect 562284 19728 562290 19780
rect 201586 19320 201592 19372
rect 201644 19360 201650 19372
rect 445846 19360 445852 19372
rect 201644 19332 445852 19360
rect 201644 19320 201650 19332
rect 445846 19320 445852 19332
rect 445904 19320 445910 19372
rect 58986 19252 58992 19304
rect 59044 19292 59050 19304
rect 88978 19292 88984 19304
rect 59044 19264 88984 19292
rect 59044 19252 59050 19264
rect 88978 19252 88984 19264
rect 89036 19252 89042 19304
rect 527818 19252 527824 19304
rect 527876 19292 527882 19304
rect 549806 19292 549812 19304
rect 527876 19264 549812 19292
rect 527876 19252 527882 19264
rect 549806 19252 549812 19264
rect 549864 19252 549870 19304
rect 57422 19184 57428 19236
rect 57480 19224 57486 19236
rect 72510 19224 72516 19236
rect 57480 19196 72516 19224
rect 57480 19184 57486 19196
rect 72510 19184 72516 19196
rect 72568 19184 72574 19236
rect 426434 19184 426440 19236
rect 426492 19224 426498 19236
rect 570690 19224 570696 19236
rect 426492 19196 570696 19224
rect 426492 19184 426498 19196
rect 570690 19184 570696 19196
rect 570748 19184 570754 19236
rect 54662 19116 54668 19168
rect 54720 19156 54726 19168
rect 336734 19156 336740 19168
rect 54720 19128 336740 19156
rect 54720 19116 54726 19128
rect 336734 19116 336740 19128
rect 336792 19116 336798 19168
rect 465074 19116 465080 19168
rect 465132 19156 465138 19168
rect 571978 19156 571984 19168
rect 465132 19128 571984 19156
rect 465132 19116 465138 19128
rect 571978 19116 571984 19128
rect 572036 19116 572042 19168
rect 57514 19048 57520 19100
rect 57572 19088 57578 19100
rect 215294 19088 215300 19100
rect 57572 19060 215300 19088
rect 57572 19048 57578 19060
rect 215294 19048 215300 19060
rect 215352 19048 215358 19100
rect 291194 19048 291200 19100
rect 291252 19088 291258 19100
rect 569126 19088 569132 19100
rect 291252 19060 569132 19088
rect 291252 19048 291258 19060
rect 569126 19048 569132 19060
rect 569184 19048 569190 19100
rect 54754 18980 54760 19032
rect 54812 19020 54818 19032
rect 293954 19020 293960 19032
rect 54812 18992 293960 19020
rect 54812 18980 54818 18992
rect 293954 18980 293960 18992
rect 294012 18980 294018 19032
rect 353294 18980 353300 19032
rect 353352 19020 353358 19032
rect 540330 19020 540336 19032
rect 353352 18992 540336 19020
rect 353352 18980 353358 18992
rect 540330 18980 540336 18992
rect 540388 18980 540394 19032
rect 38194 18912 38200 18964
rect 38252 18952 38258 18964
rect 194686 18952 194692 18964
rect 38252 18924 194692 18952
rect 38252 18912 38258 18924
rect 194686 18912 194692 18924
rect 194744 18912 194750 18964
rect 339586 18912 339592 18964
rect 339644 18952 339650 18964
rect 574186 18952 574192 18964
rect 339644 18924 574192 18952
rect 339644 18912 339650 18924
rect 574186 18912 574192 18924
rect 574244 18912 574250 18964
rect 39206 18844 39212 18896
rect 39264 18884 39270 18896
rect 189074 18884 189080 18896
rect 39264 18856 189080 18884
rect 39264 18844 39270 18856
rect 189074 18844 189080 18856
rect 189132 18844 189138 18896
rect 321554 18844 321560 18896
rect 321612 18884 321618 18896
rect 567378 18884 567384 18896
rect 321612 18856 567384 18884
rect 321612 18844 321618 18856
rect 567378 18844 567384 18856
rect 567436 18844 567442 18896
rect 39758 18776 39764 18828
rect 39816 18816 39822 18828
rect 150434 18816 150440 18828
rect 39816 18788 150440 18816
rect 39816 18776 39822 18788
rect 150434 18776 150440 18788
rect 150492 18776 150498 18828
rect 314746 18776 314752 18828
rect 314804 18816 314810 18828
rect 569402 18816 569408 18828
rect 314804 18788 569408 18816
rect 314804 18776 314810 18788
rect 569402 18776 569408 18788
rect 569460 18776 569466 18828
rect 43714 18708 43720 18760
rect 43772 18748 43778 18760
rect 146294 18748 146300 18760
rect 43772 18720 146300 18748
rect 43772 18708 43778 18720
rect 146294 18708 146300 18720
rect 146352 18708 146358 18760
rect 307754 18708 307760 18760
rect 307812 18748 307818 18760
rect 570322 18748 570328 18760
rect 307812 18720 570328 18748
rect 307812 18708 307818 18720
rect 570322 18708 570328 18720
rect 570380 18708 570386 18760
rect 55122 18640 55128 18692
rect 55180 18680 55186 18692
rect 154574 18680 154580 18692
rect 55180 18652 154580 18680
rect 55180 18640 55186 18652
rect 154574 18640 154580 18652
rect 154632 18640 154638 18692
rect 276106 18640 276112 18692
rect 276164 18680 276170 18692
rect 571518 18680 571524 18692
rect 276164 18652 571524 18680
rect 276164 18640 276170 18652
rect 571518 18640 571524 18652
rect 571576 18640 571582 18692
rect 56502 18572 56508 18624
rect 56560 18612 56566 18624
rect 105630 18612 105636 18624
rect 56560 18584 105636 18612
rect 56560 18572 56566 18584
rect 105630 18572 105636 18584
rect 105688 18572 105694 18624
rect 267734 18572 267740 18624
rect 267792 18612 267798 18624
rect 573542 18612 573548 18624
rect 267792 18584 573548 18612
rect 267792 18572 267798 18584
rect 573542 18572 573548 18584
rect 573600 18572 573606 18624
rect 58894 18504 58900 18556
rect 58952 18544 58958 18556
rect 89070 18544 89076 18556
rect 58952 18516 89076 18544
rect 58952 18504 58958 18516
rect 89070 18504 89076 18516
rect 89128 18504 89134 18556
rect 440326 18504 440332 18556
rect 440384 18544 440390 18556
rect 544102 18544 544108 18556
rect 440384 18516 544108 18544
rect 440384 18504 440390 18516
rect 544102 18504 544108 18516
rect 544160 18504 544166 18556
rect 47946 18436 47952 18488
rect 48004 18476 48010 18488
rect 164326 18476 164332 18488
rect 48004 18448 164332 18476
rect 48004 18436 48010 18448
rect 164326 18436 164332 18448
rect 164384 18436 164390 18488
rect 160094 18368 160100 18420
rect 160152 18408 160158 18420
rect 564986 18408 564992 18420
rect 160152 18380 564992 18408
rect 160152 18368 160158 18380
rect 564986 18368 564992 18380
rect 565044 18368 565050 18420
rect 38010 18300 38016 18352
rect 38068 18340 38074 18352
rect 364334 18340 364340 18352
rect 38068 18312 364340 18340
rect 38068 18300 38074 18312
rect 364334 18300 364340 18312
rect 364392 18300 364398 18352
rect 39298 17892 39304 17944
rect 39356 17932 39362 17944
rect 444374 17932 444380 17944
rect 39356 17904 444380 17932
rect 39356 17892 39362 17904
rect 444374 17892 444380 17904
rect 444432 17892 444438 17944
rect 445754 17892 445760 17944
rect 445812 17932 445818 17944
rect 577222 17932 577228 17944
rect 445812 17904 577228 17932
rect 445812 17892 445818 17904
rect 577222 17892 577228 17904
rect 577280 17892 577286 17944
rect 190546 17824 190552 17876
rect 190604 17864 190610 17876
rect 577590 17864 577596 17876
rect 190604 17836 577596 17864
rect 190604 17824 190610 17836
rect 577590 17824 577596 17836
rect 577648 17824 577654 17876
rect 47854 17756 47860 17808
rect 47912 17796 47918 17808
rect 427814 17796 427820 17808
rect 47912 17768 427820 17796
rect 47912 17756 47918 17768
rect 427814 17756 427820 17768
rect 427872 17756 427878 17808
rect 448514 17756 448520 17808
rect 448572 17796 448578 17808
rect 566550 17796 566556 17808
rect 448572 17768 566556 17796
rect 448572 17756 448578 17768
rect 566550 17756 566556 17768
rect 566608 17756 566614 17808
rect 235994 17688 236000 17740
rect 236052 17728 236058 17740
rect 582742 17728 582748 17740
rect 236052 17700 582748 17728
rect 236052 17688 236058 17700
rect 582742 17688 582748 17700
rect 582800 17688 582806 17740
rect 39574 17620 39580 17672
rect 39632 17660 39638 17672
rect 375374 17660 375380 17672
rect 39632 17632 375380 17660
rect 39632 17620 39638 17632
rect 375374 17620 375380 17632
rect 375432 17620 375438 17672
rect 438854 17620 438860 17672
rect 438912 17660 438918 17672
rect 541802 17660 541808 17672
rect 438912 17632 541808 17660
rect 438912 17620 438918 17632
rect 541802 17620 541808 17632
rect 541860 17620 541866 17672
rect 46658 17552 46664 17604
rect 46716 17592 46722 17604
rect 245746 17592 245752 17604
rect 46716 17564 245752 17592
rect 46716 17552 46722 17564
rect 245746 17552 245752 17564
rect 245804 17552 245810 17604
rect 251266 17552 251272 17604
rect 251324 17592 251330 17604
rect 583018 17592 583024 17604
rect 251324 17564 583024 17592
rect 251324 17552 251330 17564
rect 583018 17552 583024 17564
rect 583076 17552 583082 17604
rect 59630 17484 59636 17536
rect 59688 17524 59694 17536
rect 251174 17524 251180 17536
rect 59688 17496 251180 17524
rect 59688 17484 59694 17496
rect 251174 17484 251180 17496
rect 251232 17484 251238 17536
rect 260926 17484 260932 17536
rect 260984 17524 260990 17536
rect 581270 17524 581276 17536
rect 260984 17496 581276 17524
rect 260984 17484 260990 17496
rect 581270 17484 581276 17496
rect 581328 17484 581334 17536
rect 50338 17416 50344 17468
rect 50396 17456 50402 17468
rect 234614 17456 234620 17468
rect 50396 17428 234620 17456
rect 50396 17416 50402 17428
rect 234614 17416 234620 17428
rect 234672 17416 234678 17468
rect 299474 17416 299480 17468
rect 299532 17456 299538 17468
rect 543274 17456 543280 17468
rect 299532 17428 543280 17456
rect 299532 17416 299538 17428
rect 543274 17416 543280 17428
rect 543332 17416 543338 17468
rect 58802 17348 58808 17400
rect 58860 17388 58866 17400
rect 227714 17388 227720 17400
rect 58860 17360 227720 17388
rect 58860 17348 58866 17360
rect 227714 17348 227720 17360
rect 227772 17348 227778 17400
rect 259454 17348 259460 17400
rect 259512 17388 259518 17400
rect 542170 17388 542176 17400
rect 259512 17360 542176 17388
rect 259512 17348 259518 17360
rect 542170 17348 542176 17360
rect 542228 17348 542234 17400
rect 35526 17280 35532 17332
rect 35584 17320 35590 17332
rect 191834 17320 191840 17332
rect 35584 17292 191840 17320
rect 35584 17280 35590 17292
rect 191834 17280 191840 17292
rect 191892 17280 191898 17332
rect 256694 17280 256700 17332
rect 256752 17320 256758 17332
rect 543366 17320 543372 17332
rect 256752 17292 543372 17320
rect 256752 17280 256758 17292
rect 543366 17280 543372 17292
rect 543424 17280 543430 17332
rect 55950 17212 55956 17264
rect 56008 17252 56014 17264
rect 165614 17252 165620 17264
rect 56008 17224 165620 17252
rect 56008 17212 56014 17224
rect 165614 17212 165620 17224
rect 165672 17212 165678 17264
rect 234614 17212 234620 17264
rect 234672 17252 234678 17264
rect 553762 17252 553768 17264
rect 234672 17224 553768 17252
rect 234672 17212 234678 17224
rect 553762 17212 553768 17224
rect 553820 17212 553826 17264
rect 46382 17144 46388 17196
rect 46440 17184 46446 17196
rect 147674 17184 147680 17196
rect 46440 17156 147680 17184
rect 46440 17144 46446 17156
rect 147674 17144 147680 17156
rect 147732 17144 147738 17196
rect 460934 17144 460940 17196
rect 460992 17184 460998 17196
rect 542906 17184 542912 17196
rect 460992 17156 542912 17184
rect 460992 17144 460998 17156
rect 542906 17144 542912 17156
rect 542964 17144 542970 17196
rect 31478 17076 31484 17128
rect 31536 17116 31542 17128
rect 117314 17116 117320 17128
rect 31536 17088 117320 17116
rect 31536 17076 31542 17088
rect 117314 17076 117320 17088
rect 117372 17076 117378 17128
rect 511258 17076 511264 17128
rect 511316 17116 511322 17128
rect 580166 17116 580172 17128
rect 511316 17088 580172 17116
rect 511316 17076 511322 17088
rect 580166 17076 580172 17088
rect 580224 17076 580230 17128
rect 59262 17008 59268 17060
rect 59320 17048 59326 17060
rect 105538 17048 105544 17060
rect 59320 17020 105544 17048
rect 59320 17008 59326 17020
rect 105538 17008 105544 17020
rect 105596 17008 105602 17060
rect 31570 16940 31576 16992
rect 31628 16980 31634 16992
rect 201494 16980 201500 16992
rect 31628 16952 201500 16980
rect 31628 16940 31634 16952
rect 201494 16940 201500 16952
rect 201552 16940 201558 16992
rect 51626 16872 51632 16924
rect 51684 16912 51690 16924
rect 237374 16912 237380 16924
rect 51684 16884 237380 16912
rect 51684 16872 51690 16884
rect 237374 16872 237380 16884
rect 237432 16872 237438 16924
rect 522298 16532 522304 16584
rect 522356 16572 522362 16584
rect 549714 16572 549720 16584
rect 522356 16544 549720 16572
rect 522356 16532 522362 16544
rect 549714 16532 549720 16544
rect 549772 16532 549778 16584
rect 310606 16464 310612 16516
rect 310664 16504 310670 16516
rect 566274 16504 566280 16516
rect 310664 16476 566280 16504
rect 310664 16464 310670 16476
rect 566274 16464 566280 16476
rect 566332 16464 566338 16516
rect 403066 16396 403072 16448
rect 403124 16436 403130 16448
rect 582466 16436 582472 16448
rect 403124 16408 582472 16436
rect 403124 16396 403130 16408
rect 582466 16396 582472 16408
rect 582524 16396 582530 16448
rect 382366 16328 382372 16380
rect 382424 16368 382430 16380
rect 548518 16368 548524 16380
rect 382424 16340 548524 16368
rect 382424 16328 382430 16340
rect 548518 16328 548524 16340
rect 548576 16328 548582 16380
rect 364610 16260 364616 16312
rect 364668 16300 364674 16312
rect 541158 16300 541164 16312
rect 364668 16272 541164 16300
rect 364668 16260 364674 16272
rect 541158 16260 541164 16272
rect 541216 16260 541222 16312
rect 349154 16192 349160 16244
rect 349212 16232 349218 16244
rect 542998 16232 543004 16244
rect 349212 16204 543004 16232
rect 349212 16192 349218 16204
rect 542998 16192 543004 16204
rect 543056 16192 543062 16244
rect 357526 16124 357532 16176
rect 357584 16164 357590 16176
rect 562318 16164 562324 16176
rect 357584 16136 562324 16164
rect 357584 16124 357590 16136
rect 562318 16124 562324 16136
rect 562376 16124 562382 16176
rect 346946 16056 346952 16108
rect 347004 16096 347010 16108
rect 559466 16096 559472 16108
rect 347004 16068 559472 16096
rect 347004 16056 347010 16068
rect 559466 16056 559472 16068
rect 559524 16056 559530 16108
rect 342898 15988 342904 16040
rect 342956 16028 342962 16040
rect 575750 16028 575756 16040
rect 342956 16000 575756 16028
rect 342956 15988 342962 16000
rect 575750 15988 575756 16000
rect 575808 15988 575814 16040
rect 293218 15920 293224 15972
rect 293276 15960 293282 15972
rect 554958 15960 554964 15972
rect 293276 15932 554964 15960
rect 293276 15920 293282 15932
rect 554958 15920 554964 15932
rect 555016 15920 555022 15972
rect 120626 15852 120632 15904
rect 120684 15892 120690 15904
rect 576026 15892 576032 15904
rect 120684 15864 576032 15892
rect 120684 15852 120690 15864
rect 576026 15852 576032 15864
rect 576084 15852 576090 15904
rect 403618 15784 403624 15836
rect 403676 15824 403682 15836
rect 541894 15824 541900 15836
rect 403676 15796 541900 15824
rect 403676 15784 403682 15796
rect 541894 15784 541900 15796
rect 541952 15784 541958 15836
rect 433334 15716 433340 15768
rect 433392 15756 433398 15768
rect 551738 15756 551744 15768
rect 433392 15728 551744 15756
rect 433392 15716 433398 15728
rect 551738 15716 551744 15728
rect 551796 15716 551802 15768
rect 300854 15648 300860 15700
rect 300912 15688 300918 15700
rect 582374 15688 582380 15700
rect 300912 15660 582380 15688
rect 300912 15648 300918 15660
rect 582374 15648 582380 15660
rect 582432 15648 582438 15700
rect 220906 15104 220912 15156
rect 220964 15144 220970 15156
rect 564710 15144 564716 15156
rect 220964 15116 564716 15144
rect 220964 15104 220970 15116
rect 564710 15104 564716 15116
rect 564768 15104 564774 15156
rect 324406 15036 324412 15088
rect 324464 15076 324470 15088
rect 542078 15076 542084 15088
rect 324464 15048 542084 15076
rect 324464 15036 324470 15048
rect 542078 15036 542084 15048
rect 542136 15036 542142 15088
rect 380894 14968 380900 15020
rect 380952 15008 380958 15020
rect 567562 15008 567568 15020
rect 380952 14980 567568 15008
rect 380952 14968 380958 14980
rect 567562 14968 567568 14980
rect 567620 14968 567626 15020
rect 367738 14900 367744 14952
rect 367796 14940 367802 14952
rect 580994 14940 581000 14952
rect 367796 14912 581000 14940
rect 367796 14900 367802 14912
rect 580994 14900 581000 14912
rect 581052 14900 581058 14952
rect 254210 14832 254216 14884
rect 254268 14872 254274 14884
rect 540514 14872 540520 14884
rect 254268 14844 540520 14872
rect 254268 14832 254274 14844
rect 540514 14832 540520 14844
rect 540572 14832 540578 14884
rect 247586 14764 247592 14816
rect 247644 14804 247650 14816
rect 551370 14804 551376 14816
rect 247644 14776 551376 14804
rect 247644 14764 247650 14776
rect 551370 14764 551376 14776
rect 551428 14764 551434 14816
rect 264974 14696 264980 14748
rect 265032 14736 265038 14748
rect 570506 14736 570512 14748
rect 265032 14708 570512 14736
rect 265032 14696 265038 14708
rect 570506 14696 570512 14708
rect 570564 14696 570570 14748
rect 233418 14628 233424 14680
rect 233476 14668 233482 14680
rect 544562 14668 544568 14680
rect 233476 14640 544568 14668
rect 233476 14628 233482 14640
rect 544562 14628 544568 14640
rect 544620 14628 544626 14680
rect 253474 14560 253480 14612
rect 253532 14600 253538 14612
rect 576854 14600 576860 14612
rect 253532 14572 576860 14600
rect 253532 14560 253538 14572
rect 576854 14560 576860 14572
rect 576912 14560 576918 14612
rect 175458 14492 175464 14544
rect 175516 14532 175522 14544
rect 568758 14532 568764 14544
rect 175516 14504 568764 14532
rect 175516 14492 175522 14504
rect 568758 14492 568764 14504
rect 568816 14492 568822 14544
rect 171962 14424 171968 14476
rect 172020 14464 172026 14476
rect 564802 14464 564808 14476
rect 172020 14436 564808 14464
rect 172020 14424 172026 14436
rect 564802 14424 564808 14436
rect 564860 14424 564866 14476
rect 414290 14356 414296 14408
rect 414348 14396 414354 14408
rect 579246 14396 579252 14408
rect 414348 14368 579252 14396
rect 414348 14356 414354 14368
rect 579246 14356 579252 14368
rect 579304 14356 579310 14408
rect 473998 14288 474004 14340
rect 474056 14328 474062 14340
rect 540238 14328 540244 14340
rect 474056 14300 540244 14328
rect 474056 14288 474062 14300
rect 540238 14288 540244 14300
rect 540296 14288 540302 14340
rect 233234 13744 233240 13796
rect 233292 13784 233298 13796
rect 563790 13784 563796 13796
rect 233292 13756 563796 13784
rect 233292 13744 233298 13756
rect 563790 13744 563796 13756
rect 563848 13744 563854 13796
rect 320174 13676 320180 13728
rect 320232 13716 320238 13728
rect 544838 13716 544844 13728
rect 320232 13688 544844 13716
rect 320232 13676 320238 13688
rect 544838 13676 544844 13688
rect 544896 13676 544902 13728
rect 340874 13608 340880 13660
rect 340932 13648 340938 13660
rect 559558 13648 559564 13660
rect 340932 13620 559564 13648
rect 340932 13608 340938 13620
rect 559558 13608 559564 13620
rect 559616 13608 559622 13660
rect 351914 13540 351920 13592
rect 351972 13580 351978 13592
rect 551278 13580 551284 13592
rect 351972 13552 551284 13580
rect 351972 13540 351978 13552
rect 551278 13540 551284 13552
rect 551336 13540 551342 13592
rect 357434 13472 357440 13524
rect 357492 13512 357498 13524
rect 544378 13512 544384 13524
rect 357492 13484 544384 13512
rect 357492 13472 357498 13484
rect 544378 13472 544384 13484
rect 544436 13472 544442 13524
rect 363046 13404 363052 13456
rect 363104 13444 363110 13456
rect 545942 13444 545948 13456
rect 363104 13416 545948 13444
rect 363104 13404 363110 13416
rect 545942 13404 545948 13416
rect 546000 13404 546006 13456
rect 378134 13336 378140 13388
rect 378192 13376 378198 13388
rect 549438 13376 549444 13388
rect 378192 13348 549444 13376
rect 378192 13336 378198 13348
rect 549438 13336 549444 13348
rect 549496 13336 549502 13388
rect 404354 13268 404360 13320
rect 404412 13308 404418 13320
rect 560846 13308 560852 13320
rect 404412 13280 560852 13308
rect 404412 13268 404418 13280
rect 560846 13268 560852 13280
rect 560904 13268 560910 13320
rect 386414 13200 386420 13252
rect 386472 13240 386478 13252
rect 542446 13240 542452 13252
rect 386472 13212 542452 13240
rect 386472 13200 386478 13212
rect 542446 13200 542452 13212
rect 542504 13200 542510 13252
rect 398926 13132 398932 13184
rect 398984 13172 398990 13184
rect 576302 13172 576308 13184
rect 398984 13144 576308 13172
rect 398984 13132 398990 13144
rect 576302 13132 576308 13144
rect 576360 13132 576366 13184
rect 143534 13064 143540 13116
rect 143592 13104 143598 13116
rect 553394 13104 553400 13116
rect 143592 13076 553400 13104
rect 143592 13064 143598 13076
rect 553394 13064 553400 13076
rect 553452 13064 553458 13116
rect 393314 12996 393320 13048
rect 393372 13036 393378 13048
rect 548702 13036 548708 13048
rect 393372 13008 548708 13036
rect 393372 12996 393378 13008
rect 548702 12996 548708 13008
rect 548760 12996 548766 13048
rect 410794 12928 410800 12980
rect 410852 12968 410858 12980
rect 559742 12968 559748 12980
rect 410852 12940 559748 12968
rect 410852 12928 410858 12940
rect 559742 12928 559748 12940
rect 559800 12928 559806 12980
rect 456886 12860 456892 12912
rect 456944 12900 456950 12912
rect 551002 12900 551008 12912
rect 456944 12872 551008 12900
rect 456944 12860 456950 12872
rect 551002 12860 551008 12872
rect 551060 12860 551066 12912
rect 23198 12384 23204 12436
rect 23256 12424 23262 12436
rect 544194 12424 544200 12436
rect 23256 12396 544200 12424
rect 23256 12384 23262 12396
rect 544194 12384 544200 12396
rect 544252 12384 544258 12436
rect 313274 12316 313280 12368
rect 313332 12356 313338 12368
rect 542630 12356 542636 12368
rect 313332 12328 542636 12356
rect 313332 12316 313338 12328
rect 542630 12316 542636 12328
rect 542688 12316 542694 12368
rect 335446 12248 335452 12300
rect 335504 12288 335510 12300
rect 541986 12288 541992 12300
rect 335504 12260 541992 12288
rect 335504 12248 335510 12260
rect 541986 12248 541992 12260
rect 542044 12248 542050 12300
rect 347774 12180 347780 12232
rect 347832 12220 347838 12232
rect 549346 12220 549352 12232
rect 347832 12192 549352 12220
rect 347832 12180 347838 12192
rect 549346 12180 549352 12192
rect 549404 12180 549410 12232
rect 398834 12112 398840 12164
rect 398892 12152 398898 12164
rect 581178 12152 581184 12164
rect 398892 12124 581184 12152
rect 398892 12112 398898 12124
rect 581178 12112 581184 12124
rect 581236 12112 581242 12164
rect 467466 12044 467472 12096
rect 467524 12084 467530 12096
rect 545390 12084 545396 12096
rect 467524 12056 545396 12084
rect 467524 12044 467530 12056
rect 545390 12044 545396 12056
rect 545448 12044 545454 12096
rect 299474 11976 299480 12028
rect 299532 12016 299538 12028
rect 583662 12016 583668 12028
rect 299532 11988 583668 12016
rect 299532 11976 299538 11988
rect 583662 11976 583668 11988
rect 583720 11976 583726 12028
rect 228266 11908 228272 11960
rect 228324 11948 228330 11960
rect 545482 11948 545488 11960
rect 228324 11920 545488 11948
rect 228324 11908 228330 11920
rect 545482 11908 545488 11920
rect 545540 11908 545546 11960
rect 194410 11840 194416 11892
rect 194468 11880 194474 11892
rect 551554 11880 551560 11892
rect 194468 11852 551560 11880
rect 194468 11840 194474 11852
rect 551554 11840 551560 11852
rect 551612 11840 551618 11892
rect 36814 11772 36820 11824
rect 36872 11812 36878 11824
rect 132954 11812 132960 11824
rect 36872 11784 132960 11812
rect 36872 11772 36878 11784
rect 132954 11772 132960 11784
rect 133012 11812 133018 11824
rect 504358 11812 504364 11824
rect 133012 11784 504364 11812
rect 133012 11772 133018 11784
rect 504358 11772 504364 11784
rect 504416 11772 504422 11824
rect 56778 11704 56784 11756
rect 56836 11744 56842 11756
rect 574462 11744 574468 11756
rect 56836 11716 574468 11744
rect 56836 11704 56842 11716
rect 574462 11704 574468 11716
rect 574520 11704 574526 11756
rect 314654 10956 314660 11008
rect 314712 10996 314718 11008
rect 548242 10996 548248 11008
rect 314712 10968 548248 10996
rect 314712 10956 314718 10968
rect 548242 10956 548248 10968
rect 548300 10956 548306 11008
rect 328454 10888 328460 10940
rect 328512 10928 328518 10940
rect 546954 10928 546960 10940
rect 328512 10900 546960 10928
rect 328512 10888 328518 10900
rect 546954 10888 546960 10900
rect 547012 10888 547018 10940
rect 338114 10820 338120 10872
rect 338172 10860 338178 10872
rect 540606 10860 540612 10872
rect 338172 10832 540612 10860
rect 338172 10820 338178 10832
rect 540606 10820 540612 10832
rect 540664 10820 540670 10872
rect 339494 10752 339500 10804
rect 339552 10792 339558 10804
rect 540146 10792 540152 10804
rect 339552 10764 540152 10792
rect 339552 10752 339558 10764
rect 540146 10752 540152 10764
rect 540204 10752 540210 10804
rect 346394 10684 346400 10736
rect 346452 10724 346458 10736
rect 546034 10724 546040 10736
rect 346452 10696 546040 10724
rect 346452 10684 346458 10696
rect 546034 10684 546040 10696
rect 546092 10684 546098 10736
rect 387058 10616 387064 10668
rect 387116 10656 387122 10668
rect 540422 10656 540428 10668
rect 387116 10628 540428 10656
rect 387116 10616 387122 10628
rect 540422 10616 540428 10628
rect 540480 10616 540486 10668
rect 141234 10276 141240 10328
rect 141292 10316 141298 10328
rect 557902 10316 557908 10328
rect 141292 10288 557908 10316
rect 141292 10276 141298 10288
rect 557902 10276 557908 10288
rect 557960 10276 557966 10328
rect 371694 8984 371700 9036
rect 371752 9024 371758 9036
rect 553670 9024 553676 9036
rect 371752 8996 553676 9024
rect 371752 8984 371758 8996
rect 553670 8984 553676 8996
rect 553728 8984 553734 9036
rect 258258 8916 258264 8968
rect 258316 8956 258322 8968
rect 553486 8956 553492 8968
rect 258316 8928 553492 8956
rect 258316 8916 258322 8928
rect 553486 8916 553492 8928
rect 553544 8916 553550 8968
rect 421374 7556 421380 7608
rect 421432 7596 421438 7608
rect 559834 7596 559840 7608
rect 421432 7568 559840 7596
rect 421432 7556 421438 7568
rect 559834 7556 559840 7568
rect 559892 7556 559898 7608
rect 567838 7556 567844 7608
rect 567896 7596 567902 7608
rect 579798 7596 579804 7608
rect 567896 7568 579804 7596
rect 567896 7556 567902 7568
rect 579798 7556 579804 7568
rect 579856 7556 579862 7608
rect 506474 6808 506480 6860
rect 506532 6848 506538 6860
rect 566458 6848 566464 6860
rect 506532 6820 566464 6848
rect 506532 6808 506538 6820
rect 566458 6808 566464 6820
rect 566516 6808 566522 6860
rect 499390 6740 499396 6792
rect 499448 6780 499454 6792
rect 571886 6780 571892 6792
rect 499448 6752 571892 6780
rect 499448 6740 499454 6752
rect 571886 6740 571892 6752
rect 571944 6740 571950 6792
rect 460382 6672 460388 6724
rect 460440 6712 460446 6724
rect 541618 6712 541624 6724
rect 460440 6684 541624 6712
rect 460440 6672 460446 6684
rect 541618 6672 541624 6684
rect 541676 6672 541682 6724
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 485222 6604 485228 6656
rect 485280 6644 485286 6656
rect 567286 6644 567292 6656
rect 485280 6616 567292 6644
rect 485280 6604 485286 6616
rect 567286 6604 567292 6616
rect 567344 6604 567350 6656
rect 463970 6536 463976 6588
rect 464028 6576 464034 6588
rect 548794 6576 548800 6588
rect 464028 6548 548800 6576
rect 464028 6536 464034 6548
rect 548794 6536 548800 6548
rect 548852 6536 548858 6588
rect 446214 6468 446220 6520
rect 446272 6508 446278 6520
rect 543090 6508 543096 6520
rect 446272 6480 543096 6508
rect 446272 6468 446278 6480
rect 543090 6468 543096 6480
rect 543148 6468 543154 6520
rect 449802 6400 449808 6452
rect 449860 6440 449866 6452
rect 557994 6440 558000 6452
rect 449860 6412 558000 6440
rect 449860 6400 449866 6412
rect 557994 6400 558000 6412
rect 558052 6400 558058 6452
rect 442626 6332 442632 6384
rect 442684 6372 442690 6384
rect 559374 6372 559380 6384
rect 442684 6344 559380 6372
rect 442684 6332 442690 6344
rect 559374 6332 559380 6344
rect 559432 6332 559438 6384
rect 439130 6264 439136 6316
rect 439188 6304 439194 6316
rect 563514 6304 563520 6316
rect 439188 6276 563520 6304
rect 439188 6264 439194 6276
rect 563514 6264 563520 6276
rect 563572 6264 563578 6316
rect 432046 6196 432052 6248
rect 432104 6236 432110 6248
rect 573266 6236 573272 6248
rect 432104 6208 573272 6236
rect 432104 6196 432110 6208
rect 573266 6196 573272 6208
rect 573324 6196 573330 6248
rect 332686 6128 332692 6180
rect 332744 6168 332750 6180
rect 556246 6168 556252 6180
rect 332744 6140 556252 6168
rect 332744 6128 332750 6140
rect 556246 6128 556252 6140
rect 556304 6128 556310 6180
rect 288434 5448 288440 5500
rect 288492 5488 288498 5500
rect 550358 5488 550364 5500
rect 288492 5460 550364 5488
rect 288492 5448 288498 5460
rect 550358 5448 550364 5460
rect 550416 5448 550422 5500
rect 375282 4836 375288 4888
rect 375340 4876 375346 4888
rect 557534 4876 557540 4888
rect 375340 4848 557540 4876
rect 375340 4836 375346 4848
rect 557534 4836 557540 4848
rect 557592 4836 557598 4888
rect 318518 4768 318524 4820
rect 318576 4808 318582 4820
rect 547138 4808 547144 4820
rect 318576 4780 547144 4808
rect 318576 4768 318582 4780
rect 547138 4768 547144 4780
rect 547196 4768 547202 4820
rect 38286 4088 38292 4140
rect 38344 4128 38350 4140
rect 125870 4128 125876 4140
rect 38344 4100 125876 4128
rect 38344 4088 38350 4100
rect 125870 4088 125876 4100
rect 125928 4088 125934 4140
rect 492306 4088 492312 4140
rect 492364 4128 492370 4140
rect 553854 4128 553860 4140
rect 492364 4100 553860 4128
rect 492364 4088 492370 4100
rect 553854 4088 553860 4100
rect 553912 4088 553918 4140
rect 42334 4020 42340 4072
rect 42392 4060 42398 4072
rect 134150 4060 134156 4072
rect 42392 4032 134156 4060
rect 42392 4020 42398 4032
rect 134150 4020 134156 4032
rect 134208 4020 134214 4072
rect 488810 4020 488816 4072
rect 488868 4060 488874 4072
rect 566366 4060 566372 4072
rect 488868 4032 566372 4060
rect 488868 4020 488874 4032
rect 566366 4020 566372 4032
rect 566424 4020 566430 4072
rect 48774 3952 48780 4004
rect 48832 3992 48838 4004
rect 151814 3992 151820 4004
rect 48832 3964 151820 3992
rect 48832 3952 48838 3964
rect 151814 3952 151820 3964
rect 151872 3952 151878 4004
rect 424962 3952 424968 4004
rect 425020 3992 425026 4004
rect 555142 3992 555148 4004
rect 425020 3964 555148 3992
rect 425020 3952 425026 3964
rect 555142 3952 555148 3964
rect 555200 3952 555206 4004
rect 565814 3952 565820 4004
rect 565872 3992 565878 4004
rect 566090 3992 566096 4004
rect 565872 3964 566096 3992
rect 565872 3952 565878 3964
rect 566090 3952 566096 3964
rect 566148 3952 566154 4004
rect 43898 3884 43904 3936
rect 43956 3924 43962 3936
rect 158898 3924 158904 3936
rect 43956 3896 158904 3924
rect 43956 3884 43962 3896
rect 158898 3884 158904 3896
rect 158956 3884 158962 3936
rect 286594 3884 286600 3936
rect 286652 3924 286658 3936
rect 578694 3924 578700 3936
rect 286652 3896 578700 3924
rect 286652 3884 286658 3896
rect 578694 3884 578700 3896
rect 578752 3884 578758 3936
rect 48222 3816 48228 3868
rect 48280 3856 48286 3868
rect 173158 3856 173164 3868
rect 48280 3828 173164 3856
rect 48280 3816 48286 3828
rect 173158 3816 173164 3828
rect 173216 3816 173222 3868
rect 239306 3816 239312 3868
rect 239364 3856 239370 3868
rect 533338 3856 533344 3868
rect 239364 3828 533344 3856
rect 239364 3816 239370 3828
rect 533338 3816 533344 3828
rect 533396 3816 533402 3868
rect 534902 3816 534908 3868
rect 534960 3856 534966 3868
rect 573450 3856 573456 3868
rect 534960 3828 573456 3856
rect 534960 3816 534966 3828
rect 573450 3816 573456 3828
rect 573508 3816 573514 3868
rect 45002 3748 45008 3800
rect 45060 3788 45066 3800
rect 189718 3788 189724 3800
rect 45060 3760 189724 3788
rect 45060 3748 45066 3760
rect 189718 3748 189724 3760
rect 189776 3748 189782 3800
rect 244090 3748 244096 3800
rect 244148 3788 244154 3800
rect 545758 3788 545764 3800
rect 244148 3760 545764 3788
rect 244148 3748 244154 3760
rect 545758 3748 545764 3760
rect 545816 3748 545822 3800
rect 552658 3748 552664 3800
rect 552716 3788 552722 3800
rect 574278 3788 574284 3800
rect 552716 3760 574284 3788
rect 552716 3748 552722 3760
rect 574278 3748 574284 3760
rect 574336 3748 574342 3800
rect 34422 3680 34428 3732
rect 34480 3720 34486 3732
rect 193214 3720 193220 3732
rect 34480 3692 193220 3720
rect 34480 3680 34486 3692
rect 193214 3680 193220 3692
rect 193272 3680 193278 3732
rect 218146 3680 218152 3732
rect 218204 3720 218210 3732
rect 218204 3692 219388 3720
rect 218204 3680 218210 3692
rect 34146 3612 34152 3664
rect 34204 3652 34210 3664
rect 196802 3652 196808 3664
rect 34204 3624 196808 3652
rect 34204 3612 34210 3624
rect 196802 3612 196808 3624
rect 196860 3612 196866 3664
rect 219360 3652 219388 3692
rect 237006 3680 237012 3732
rect 237064 3720 237070 3732
rect 581546 3720 581552 3732
rect 237064 3692 581552 3720
rect 237064 3680 237070 3692
rect 581546 3680 581552 3692
rect 581604 3680 581610 3732
rect 571610 3652 571616 3664
rect 219360 3624 571616 3652
rect 571610 3612 571616 3624
rect 571668 3612 571674 3664
rect 31662 3544 31668 3596
rect 31720 3584 31726 3596
rect 212166 3584 212172 3596
rect 31720 3556 212172 3584
rect 31720 3544 31726 3556
rect 212166 3544 212172 3556
rect 212224 3544 212230 3596
rect 218054 3544 218060 3596
rect 218112 3584 218118 3596
rect 219250 3584 219256 3596
rect 218112 3556 219256 3584
rect 218112 3544 218118 3556
rect 219250 3544 219256 3556
rect 219308 3544 219314 3596
rect 219342 3544 219348 3596
rect 219400 3584 219406 3596
rect 573082 3584 573088 3596
rect 219400 3556 573088 3584
rect 219400 3544 219406 3556
rect 573082 3544 573088 3556
rect 573140 3544 573146 3596
rect 41966 3476 41972 3528
rect 42024 3516 42030 3528
rect 42024 3488 184796 3516
rect 42024 3476 42030 3488
rect 37182 3408 37188 3460
rect 37240 3448 37246 3460
rect 161290 3448 161296 3460
rect 37240 3420 161296 3448
rect 37240 3408 37246 3420
rect 161290 3408 161296 3420
rect 161348 3408 161354 3460
rect 168374 3408 168380 3460
rect 168432 3448 168438 3460
rect 168432 3420 180794 3448
rect 168432 3408 168438 3420
rect 42426 3340 42432 3392
rect 42484 3380 42490 3392
rect 130562 3380 130568 3392
rect 42484 3352 130568 3380
rect 42484 3340 42490 3352
rect 130562 3340 130568 3352
rect 130620 3340 130626 3392
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 136450 3380 136456 3392
rect 135312 3352 136456 3380
rect 135312 3340 135318 3352
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 50246 3272 50252 3324
rect 50304 3312 50310 3324
rect 110506 3312 110512 3324
rect 50304 3284 110512 3312
rect 50304 3272 50310 3284
rect 110506 3272 110512 3284
rect 110564 3272 110570 3324
rect 180766 3312 180794 3420
rect 184768 3380 184796 3488
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 186130 3516 186136 3528
rect 184992 3488 186136 3516
rect 184992 3476 184998 3488
rect 186130 3476 186136 3488
rect 186188 3476 186194 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 552842 3516 552848 3528
rect 190880 3488 552848 3516
rect 190880 3476 190886 3488
rect 552842 3476 552848 3488
rect 552900 3476 552906 3528
rect 572070 3476 572076 3528
rect 572128 3516 572134 3528
rect 573910 3516 573916 3528
rect 572128 3488 573916 3516
rect 572128 3476 572134 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 565814 3448 565820 3460
rect 190426 3420 565820 3448
rect 187326 3380 187332 3392
rect 184768 3352 187332 3380
rect 187326 3340 187332 3352
rect 187384 3340 187390 3392
rect 190426 3312 190454 3420
rect 565814 3408 565820 3420
rect 565872 3408 565878 3460
rect 215662 3340 215668 3392
rect 215720 3380 215726 3392
rect 219342 3380 219348 3392
rect 215720 3352 219348 3380
rect 215720 3340 215726 3352
rect 219342 3340 219348 3352
rect 219400 3340 219406 3392
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 235810 3380 235816 3392
rect 234672 3352 235816 3380
rect 234672 3340 234678 3352
rect 235810 3340 235816 3352
rect 235868 3340 235874 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260650 3380 260656 3392
rect 259512 3352 260656 3380
rect 259512 3340 259518 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 299474 3340 299480 3392
rect 299532 3380 299538 3392
rect 300762 3380 300768 3392
rect 299532 3352 300768 3380
rect 299532 3340 299538 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 495894 3340 495900 3392
rect 495952 3380 495958 3392
rect 556430 3380 556436 3392
rect 495952 3352 556436 3380
rect 495952 3340 495958 3352
rect 556430 3340 556436 3352
rect 556488 3340 556494 3392
rect 180766 3284 190454 3312
rect 510062 3272 510068 3324
rect 510120 3312 510126 3324
rect 563422 3312 563428 3324
rect 510120 3284 563428 3312
rect 510120 3272 510126 3284
rect 563422 3272 563428 3284
rect 563480 3272 563486 3324
rect 578970 3272 578976 3324
rect 579028 3312 579034 3324
rect 582190 3312 582196 3324
rect 579028 3284 582196 3312
rect 579028 3272 579034 3284
rect 582190 3272 582196 3284
rect 582248 3272 582254 3324
rect 545482 3204 545488 3256
rect 545540 3244 545546 3256
rect 571702 3244 571708 3256
rect 545540 3216 571708 3244
rect 545540 3204 545546 3216
rect 571702 3204 571708 3216
rect 571760 3204 571766 3256
rect 527818 3136 527824 3188
rect 527876 3176 527882 3188
rect 546678 3176 546684 3188
rect 527876 3148 546684 3176
rect 527876 3136 527882 3148
rect 546678 3136 546684 3148
rect 546736 3136 546742 3188
rect 552750 3000 552756 3052
rect 552808 3040 552814 3052
rect 556154 3040 556160 3052
rect 552808 3012 556160 3040
rect 552808 3000 552814 3012
rect 556154 3000 556160 3012
rect 556212 3000 556218 3052
rect 324314 2048 324320 2100
rect 324372 2088 324378 2100
rect 325602 2088 325608 2100
rect 324372 2060 325608 2088
rect 324372 2048 324378 2060
rect 325602 2048 325608 2060
rect 325660 2048 325666 2100
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 484400 700680 484452 700732
rect 543464 700680 543516 700732
rect 332508 700612 332560 700664
rect 398196 700612 398248 700664
rect 402888 700612 402940 700664
rect 527180 700612 527232 700664
rect 283840 700544 283892 700596
rect 399484 700544 399536 700596
rect 405004 700544 405056 700596
rect 559656 700544 559708 700596
rect 364984 700476 365036 700528
rect 551376 700476 551428 700528
rect 218980 700408 219032 700460
rect 342996 700408 343048 700460
rect 348792 700408 348844 700460
rect 566004 700408 566056 700460
rect 300124 700340 300176 700392
rect 551468 700340 551520 700392
rect 267648 700272 267700 700324
rect 566188 700272 566240 700324
rect 105452 698912 105504 698964
rect 399392 698912 399444 698964
rect 429844 698912 429896 698964
rect 550272 698912 550324 698964
rect 137836 697552 137888 697604
rect 389916 697552 389968 697604
rect 413652 697552 413704 697604
rect 552204 697552 552256 697604
rect 154120 696192 154172 696244
rect 552848 696192 552900 696244
rect 201500 694764 201552 694816
rect 498200 694764 498252 694816
rect 88340 693404 88392 693456
rect 551100 693404 551152 693456
rect 6920 692044 6972 692096
rect 550088 692044 550140 692096
rect 71780 690616 71832 690668
rect 383016 690616 383068 690668
rect 234620 687964 234672 688016
rect 538220 687964 538272 688016
rect 40040 687896 40092 687948
rect 373632 687896 373684 687948
rect 462320 687896 462372 687948
rect 550640 687896 550692 687948
rect 405096 687284 405148 687336
rect 457352 687284 457404 687336
rect 399760 687216 399812 687268
rect 554872 687216 554924 687268
rect 367744 686060 367796 686112
rect 476580 686060 476632 686112
rect 407764 685992 407816 686044
rect 554964 685992 555016 686044
rect 378784 685924 378836 685976
rect 528836 685924 528888 685976
rect 405188 685856 405240 685908
rect 580908 685856 580960 685908
rect 409144 685312 409196 685364
rect 470876 685312 470928 685364
rect 409052 685244 409104 685296
rect 454224 685244 454276 685296
rect 408408 685176 408460 685228
rect 436100 685176 436152 685228
rect 409696 685108 409748 685160
rect 450268 685108 450320 685160
rect 402428 685040 402480 685092
rect 490012 685040 490064 685092
rect 510528 685040 510580 685092
rect 581000 685040 581052 685092
rect 407948 684972 408000 685024
rect 456892 684972 456944 685024
rect 472808 684972 472860 685024
rect 582380 684972 582432 685024
rect 409236 684904 409288 684956
rect 523040 684904 523092 684956
rect 467012 684836 467064 684888
rect 582472 684836 582524 684888
rect 398748 684768 398800 684820
rect 521844 684768 521896 684820
rect 409512 684700 409564 684752
rect 535460 684700 535512 684752
rect 396816 684632 396868 684684
rect 539140 684632 539192 684684
rect 435456 684564 435508 684616
rect 576860 684564 576912 684616
rect 408040 684496 408092 684548
rect 555148 684496 555200 684548
rect 393964 684088 394016 684140
rect 470692 684088 470744 684140
rect 409788 684020 409840 684072
rect 449900 684020 449952 684072
rect 399852 683952 399904 684004
rect 468392 683952 468444 684004
rect 401508 683884 401560 683936
rect 476120 683884 476172 683936
rect 409328 683816 409380 683868
rect 497280 683816 497332 683868
rect 393228 683748 393280 683800
rect 499856 683748 499908 683800
rect 524880 683748 524932 683800
rect 582564 683748 582616 683800
rect 405372 683680 405424 683732
rect 437572 683680 437624 683732
rect 468300 683680 468352 683732
rect 579252 683680 579304 683732
rect 377404 683612 377456 683664
rect 422392 683612 422444 683664
rect 441252 683612 441304 683664
rect 554044 683612 554096 683664
rect 438676 683544 438728 683596
rect 567936 683544 567988 683596
rect 406476 683476 406528 683528
rect 552296 683476 552348 683528
rect 407856 683408 407908 683460
rect 553676 683408 553728 683460
rect 406568 683340 406620 683392
rect 553584 683340 553636 683392
rect 403808 683272 403860 683324
rect 555240 683272 555292 683324
rect 416688 683204 416740 683256
rect 571340 683204 571392 683256
rect 404084 683136 404136 683188
rect 580356 683136 580408 683188
rect 529664 682728 529716 682780
rect 551284 682728 551336 682780
rect 408132 682660 408184 682712
rect 553492 682660 553544 682712
rect 364248 682592 364300 682644
rect 546960 682592 547012 682644
rect 3424 682524 3476 682576
rect 550180 682524 550232 682576
rect 402336 682456 402388 682508
rect 441896 682456 441948 682508
rect 507584 682456 507636 682508
rect 553400 682456 553452 682508
rect 402244 682388 402296 682440
rect 458640 682388 458692 682440
rect 477500 682388 477552 682440
rect 566096 682388 566148 682440
rect 403716 682320 403768 682372
rect 463792 682320 463844 682372
rect 502248 682320 502300 682372
rect 560944 682320 560996 682372
rect 373264 682252 373316 682304
rect 439964 682252 440016 682304
rect 447140 682252 447192 682304
rect 509332 682252 509384 682304
rect 517244 682252 517296 682304
rect 574100 682252 574152 682304
rect 385684 682184 385736 682236
rect 480352 682184 480404 682236
rect 512736 682184 512788 682236
rect 575572 682184 575624 682236
rect 360844 682116 360896 682168
rect 429660 682116 429712 682168
rect 443000 682116 443052 682168
rect 458456 682116 458508 682168
rect 554780 682116 554832 682168
rect 398104 682048 398156 682100
rect 524972 682048 525024 682100
rect 549444 682048 549496 682100
rect 577044 682048 577096 682100
rect 549996 681980 550048 682032
rect 570144 681980 570196 682032
rect 387708 681912 387760 681964
rect 534080 681912 534132 681964
rect 535276 681912 535328 681964
rect 568764 681912 568816 681964
rect 403992 681844 404044 681896
rect 580448 681844 580500 681896
rect 537852 681776 537904 681828
rect 571616 681776 571668 681828
rect 499212 681708 499264 681760
rect 517520 681708 517572 681760
rect 541716 681708 541768 681760
rect 571984 681708 572036 681760
rect 400036 681300 400088 681352
rect 580724 681300 580776 681352
rect 517520 681232 517572 681284
rect 580264 681232 580316 681284
rect 174544 681164 174596 681216
rect 461216 681164 461268 681216
rect 501788 681164 501840 681216
rect 576124 681164 576176 681216
rect 407580 681096 407632 681148
rect 443000 681096 443052 681148
rect 496636 681096 496688 681148
rect 575480 681096 575532 681148
rect 408316 681028 408368 681080
rect 447140 681028 447192 681080
rect 484860 681028 484912 681080
rect 570052 681028 570104 681080
rect 342904 680960 342956 681012
rect 432052 680960 432104 681012
rect 434628 680960 434680 681012
rect 550732 680960 550784 681012
rect 409880 680892 409932 680944
rect 552940 680892 552992 680944
rect 408960 680824 409012 680876
rect 552112 680824 552164 680876
rect 406660 680756 406712 680808
rect 551192 680756 551244 680808
rect 406844 680688 406896 680740
rect 552756 680688 552808 680740
rect 406384 680620 406436 680672
rect 555056 680620 555108 680672
rect 399576 680552 399628 680604
rect 550916 680552 550968 680604
rect 400128 680484 400180 680536
rect 552664 680484 552716 680536
rect 409420 680416 409472 680468
rect 424508 680416 424560 680468
rect 399668 680348 399720 680400
rect 427912 680348 427964 680400
rect 439320 680348 439372 680400
rect 551008 680348 551060 680400
rect 437940 680076 437992 680128
rect 446220 680076 446272 680128
rect 441804 680008 441856 680060
rect 445760 680008 445812 680060
rect 435824 679940 435876 679992
rect 446956 679940 447008 679992
rect 441712 679872 441764 679924
rect 445944 679872 445996 679924
rect 465540 679872 465592 679924
rect 467104 679872 467156 679924
rect 411260 679804 411312 679856
rect 421472 679804 421524 679856
rect 413744 679736 413796 679788
rect 415216 679736 415268 679788
rect 409604 679668 409656 679720
rect 415492 679668 415544 679720
rect 442356 679736 442408 679788
rect 443920 679668 443972 679720
rect 406752 679464 406804 679516
rect 415354 679600 415406 679652
rect 411260 679464 411312 679516
rect 413744 679464 413796 679516
rect 405280 679396 405332 679448
rect 396724 679328 396776 679380
rect 399944 679260 399996 679312
rect 415216 679532 415268 679584
rect 358084 679192 358136 679244
rect 421472 679464 421524 679516
rect 432696 679532 432748 679584
rect 432788 679464 432840 679516
rect 432972 679464 433024 679516
rect 435824 679464 435876 679516
rect 437940 679464 437992 679516
rect 441712 679464 441764 679516
rect 441804 679464 441856 679516
rect 442356 679464 442408 679516
rect 443920 679464 443972 679516
rect 395528 679124 395580 679176
rect 9680 679056 9732 679108
rect 408868 679056 408920 679108
rect 3608 678988 3660 679040
rect 446220 679532 446272 679584
rect 466184 679804 466236 679856
rect 462412 679736 462464 679788
rect 467564 679736 467616 679788
rect 445760 679464 445812 679516
rect 445944 679464 445996 679516
rect 447094 679464 447146 679516
rect 462412 679464 462464 679516
rect 467196 679600 467248 679652
rect 473452 679600 473504 679652
rect 465540 679464 465592 679516
rect 466184 679464 466236 679516
rect 552020 679532 552072 679584
rect 467104 679464 467156 679516
rect 467472 679464 467524 679516
rect 467564 679464 467616 679516
rect 552388 679464 552440 679516
rect 557908 679396 557960 679448
rect 553768 679328 553820 679380
rect 580540 679260 580592 679312
rect 580816 679124 580868 679176
rect 579068 679056 579120 679108
rect 550824 678988 550876 679040
rect 552480 678988 552532 679040
rect 582656 678988 582708 679040
rect 552020 678920 552072 678972
rect 552480 678852 552532 678904
rect 407764 678512 407816 678564
rect 407764 678308 407816 678360
rect 165528 678240 165580 678292
rect 169760 678240 169812 678292
rect 337568 678240 337620 678292
rect 407948 678172 408000 678224
rect 408408 678172 408460 678224
rect 325056 677696 325108 677748
rect 343732 677696 343784 677748
rect 153108 677628 153160 677680
rect 171140 677628 171192 677680
rect 325792 677628 325844 677680
rect 353944 677628 353996 677680
rect 552112 677628 552164 677680
rect 572812 677628 572864 677680
rect 7564 677560 7616 677612
rect 407120 677560 407172 677612
rect 552020 677560 552072 677612
rect 579620 677560 579672 677612
rect 337568 676812 337620 676864
rect 400864 676812 400916 676864
rect 552020 674840 552072 674892
rect 574284 674840 574336 674892
rect 552572 674092 552624 674144
rect 552756 674092 552808 674144
rect 552020 672052 552072 672104
rect 571708 672052 571760 672104
rect 552112 671780 552164 671832
rect 552940 671780 552992 671832
rect 342996 670624 343048 670676
rect 407120 670624 407172 670676
rect 552756 669332 552808 669384
rect 563980 669332 564032 669384
rect 367836 667904 367888 667956
rect 407120 667904 407172 667956
rect 551284 667836 551336 667888
rect 552388 667836 552440 667888
rect 404912 666544 404964 666596
rect 407120 666544 407172 666596
rect 364984 665184 365036 665236
rect 407120 665184 407172 665236
rect 397460 663688 397512 663740
rect 407120 663688 407172 663740
rect 388536 661104 388588 661156
rect 407120 661104 407172 661156
rect 381544 661036 381596 661088
rect 407212 661036 407264 661088
rect 553308 656888 553360 656940
rect 563336 656888 563388 656940
rect 399392 655460 399444 655512
rect 407120 655460 407172 655512
rect 383568 654100 383620 654152
rect 407120 654100 407172 654152
rect 380164 652740 380216 652792
rect 407120 652740 407172 652792
rect 553308 652740 553360 652792
rect 560392 652740 560444 652792
rect 394608 651380 394660 651432
rect 407120 651380 407172 651432
rect 400864 651312 400916 651364
rect 407580 651312 407632 651364
rect 402520 648660 402572 648712
rect 407120 648660 407172 648712
rect 347044 648592 347096 648644
rect 407212 648592 407264 648644
rect 553308 648592 553360 648644
rect 561864 648592 561916 648644
rect 552940 646144 552992 646196
rect 556436 646144 556488 646196
rect 552940 644648 552992 644700
rect 556804 644648 556856 644700
rect 403440 644580 403492 644632
rect 407120 644580 407172 644632
rect 384948 644444 385000 644496
rect 407396 644444 407448 644496
rect 553308 644444 553360 644496
rect 565452 644444 565504 644496
rect 393136 643084 393188 643136
rect 407212 643084 407264 643136
rect 552020 642200 552072 642252
rect 555240 642200 555292 642252
rect 390468 641792 390520 641844
rect 407304 641792 407356 641844
rect 344284 641724 344336 641776
rect 407212 641724 407264 641776
rect 358176 640296 358228 640348
rect 407212 640296 407264 640348
rect 552480 637644 552532 637696
rect 563428 637644 563480 637696
rect 405648 637576 405700 637628
rect 407488 637576 407540 637628
rect 552020 637576 552072 637628
rect 564532 637576 564584 637628
rect 391848 636216 391900 636268
rect 407212 636216 407264 636268
rect 387064 633428 387116 633480
rect 407212 633428 407264 633480
rect 369124 632068 369176 632120
rect 407212 632068 407264 632120
rect 556804 632000 556856 632052
rect 580172 632000 580224 632052
rect 552020 631728 552072 631780
rect 556528 631728 556580 631780
rect 390376 630640 390428 630692
rect 407212 630640 407264 630692
rect 553308 629280 553360 629332
rect 571432 629280 571484 629332
rect 378968 627920 379020 627972
rect 407212 627920 407264 627972
rect 404728 625336 404780 625388
rect 407396 625336 407448 625388
rect 553308 623772 553360 623824
rect 562508 623772 562560 623824
rect 402612 622412 402664 622464
rect 407212 622412 407264 622464
rect 553308 619624 553360 619676
rect 577504 619624 577556 619676
rect 372068 618264 372120 618316
rect 407212 618264 407264 618316
rect 553308 616836 553360 616888
rect 577596 616836 577648 616888
rect 551284 615884 551336 615936
rect 552664 615884 552716 615936
rect 369308 615476 369360 615528
rect 407304 615476 407356 615528
rect 553308 614116 553360 614168
rect 581184 614116 581236 614168
rect 392860 612756 392912 612808
rect 407212 612756 407264 612808
rect 553308 612756 553360 612808
rect 578884 612756 578936 612808
rect 346308 611328 346360 611380
rect 371332 611328 371384 611380
rect 553308 611328 553360 611380
rect 569960 611328 570012 611380
rect 553308 609968 553360 610020
rect 570696 609968 570748 610020
rect 173808 608608 173860 608660
rect 202144 608608 202196 608660
rect 373356 608608 373408 608660
rect 407212 608608 407264 608660
rect 552480 608608 552532 608660
rect 555700 608608 555752 608660
rect 173808 607180 173860 607232
rect 199384 607180 199436 607232
rect 345112 607180 345164 607232
rect 364340 607180 364392 607232
rect 369216 607180 369268 607232
rect 407212 607180 407264 607232
rect 553308 607180 553360 607232
rect 562048 607180 562100 607232
rect 345572 605820 345624 605872
rect 365812 605820 365864 605872
rect 552020 603916 552072 603968
rect 554780 603916 554832 603968
rect 553308 603100 553360 603152
rect 563152 603100 563204 603152
rect 175924 601672 175976 601724
rect 203064 601672 203116 601724
rect 376024 601672 376076 601724
rect 407304 601672 407356 601724
rect 570604 600924 570656 600976
rect 580908 600924 580960 600976
rect 378876 598952 378928 599004
rect 407304 598952 407356 599004
rect 398656 596164 398708 596216
rect 407304 596164 407356 596216
rect 401416 594804 401468 594856
rect 407304 594804 407356 594856
rect 398564 592016 398616 592068
rect 407304 592016 407356 592068
rect 32680 591948 32732 592000
rect 204904 591948 204956 592000
rect 31576 591336 31628 591388
rect 32404 591336 32456 591388
rect 32864 591336 32916 591388
rect 78864 591336 78916 591388
rect 153660 591336 153712 591388
rect 171324 591336 171376 591388
rect 32772 591268 32824 591320
rect 306288 591268 306340 591320
rect 552020 590792 552072 590844
rect 555792 590792 555844 590844
rect 37004 590656 37056 590708
rect 407304 590656 407356 590708
rect 552480 590656 552532 590708
rect 581092 590656 581144 590708
rect 48964 590248 49016 590300
rect 60372 590248 60424 590300
rect 42616 590180 42668 590232
rect 50068 590180 50120 590232
rect 317420 590180 317472 590232
rect 343732 590180 343784 590232
rect 45284 590112 45336 590164
rect 77300 590112 77352 590164
rect 292764 590112 292816 590164
rect 406476 590112 406528 590164
rect 45100 590044 45152 590096
rect 78680 590044 78732 590096
rect 257344 590044 257396 590096
rect 406568 590044 406620 590096
rect 32864 589976 32916 590028
rect 69020 589976 69072 590028
rect 225144 589976 225196 590028
rect 400128 589976 400180 590028
rect 41236 589908 41288 589960
rect 171140 589908 171192 589960
rect 226432 589908 226484 589960
rect 405096 589908 405148 589960
rect 43720 589840 43772 589892
rect 92480 589840 92532 589892
rect 44640 589772 44692 589824
rect 127348 589772 127400 589824
rect 44732 589704 44784 589756
rect 129740 589704 129792 589756
rect 55864 589636 55916 589688
rect 227076 589636 227128 589688
rect 292120 589636 292172 589688
rect 348516 589636 348568 589688
rect 47584 589568 47636 589620
rect 241520 589568 241572 589620
rect 246672 589568 246724 589620
rect 351184 589568 351236 589620
rect 25780 589500 25832 589552
rect 223028 589500 223080 589552
rect 238392 589500 238444 589552
rect 355048 589500 355100 589552
rect 41144 589432 41196 589484
rect 99932 589432 99984 589484
rect 107568 589432 107620 589484
rect 308404 589432 308456 589484
rect 312084 589432 312136 589484
rect 354772 589432 354824 589484
rect 38384 589364 38436 589416
rect 251180 589364 251232 589416
rect 252376 589364 252428 589416
rect 355140 589364 355192 589416
rect 44916 589296 44968 589348
rect 259460 589296 259512 589348
rect 289544 589296 289596 589348
rect 350816 589296 350868 589348
rect 552020 588956 552072 589008
rect 554872 588956 554924 589008
rect 74816 588616 74868 588668
rect 295984 588616 296036 588668
rect 3516 588548 3568 588600
rect 371976 588548 372028 588600
rect 386328 587868 386380 587920
rect 407304 587868 407356 587920
rect 21824 587800 21876 587852
rect 122564 587800 122616 587852
rect 171692 587800 171744 587852
rect 236092 587800 236144 587852
rect 40960 587732 41012 587784
rect 203616 587732 203668 587784
rect 256056 587732 256108 587784
rect 359280 587732 359332 587784
rect 40868 587664 40920 587716
rect 203524 587664 203576 587716
rect 240600 587664 240652 587716
rect 354680 587664 354732 587716
rect 34888 587596 34940 587648
rect 225328 587596 225380 587648
rect 239312 587596 239364 587648
rect 399852 587596 399904 587648
rect 47032 587528 47084 587580
rect 345020 587528 345072 587580
rect 100852 587460 100904 587512
rect 405280 587460 405332 587512
rect 31576 587392 31628 587444
rect 78680 587392 78732 587444
rect 86040 587392 86092 587444
rect 396724 587392 396776 587444
rect 44088 587324 44140 587376
rect 399760 587324 399812 587376
rect 39948 587256 40000 587308
rect 399944 587256 399996 587308
rect 43996 587188 44048 587240
rect 406936 587188 406988 587240
rect 36728 587120 36780 587172
rect 402520 587120 402572 587172
rect 44824 587052 44876 587104
rect 137284 587052 137336 587104
rect 215484 587052 215536 587104
rect 278964 587052 279016 587104
rect 22744 586984 22796 587036
rect 104900 586984 104952 587036
rect 41972 586508 42024 586560
rect 407304 586508 407356 586560
rect 552020 586508 552072 586560
rect 578976 586508 579028 586560
rect 163320 585896 163372 585948
rect 231860 585896 231912 585948
rect 265072 585896 265124 585948
rect 293960 585896 294012 585948
rect 150440 585828 150492 585880
rect 171232 585828 171284 585880
rect 226616 585828 226668 585880
rect 351460 585828 351512 585880
rect 65432 585760 65484 585812
rect 351092 585760 351144 585812
rect 552020 585148 552072 585200
rect 577228 585148 577280 585200
rect 160100 584468 160152 584520
rect 254124 584468 254176 584520
rect 75736 584400 75788 584452
rect 132500 584400 132552 584452
rect 140780 584400 140832 584452
rect 345112 584400 345164 584452
rect 147220 583040 147272 583092
rect 271880 583040 271932 583092
rect 320456 583040 320508 583092
rect 381544 583040 381596 583092
rect 103428 582972 103480 583024
rect 349620 582972 349672 583024
rect 135628 581748 135680 581800
rect 248512 581748 248564 581800
rect 46664 581680 46716 581732
rect 172612 581680 172664 581732
rect 202880 581680 202932 581732
rect 242900 581680 242952 581732
rect 93768 581612 93820 581664
rect 222200 581612 222252 581664
rect 277308 581612 277360 581664
rect 350724 581612 350776 581664
rect 43904 580456 43956 580508
rect 117320 580456 117372 580508
rect 204904 580456 204956 580508
rect 250444 580456 250496 580508
rect 205548 580388 205600 580440
rect 278596 580388 278648 580440
rect 297916 580388 297968 580440
rect 347044 580388 347096 580440
rect 117320 580320 117372 580372
rect 233240 580320 233292 580372
rect 239956 580320 240008 580372
rect 350356 580320 350408 580372
rect 202144 580252 202196 580304
rect 349896 580252 349948 580304
rect 383292 579640 383344 579692
rect 407304 579640 407356 579692
rect 158628 578960 158680 579012
rect 270224 578960 270276 579012
rect 282828 578960 282880 579012
rect 350632 578960 350684 579012
rect 46388 578892 46440 578944
rect 299480 578892 299532 578944
rect 552020 578212 552072 578264
rect 563612 578212 563664 578264
rect 140688 577668 140740 577720
rect 163964 577668 164016 577720
rect 230296 577668 230348 577720
rect 306380 577668 306432 577720
rect 82636 577600 82688 577652
rect 147864 577600 147916 577652
rect 154580 577600 154632 577652
rect 251272 577600 251324 577652
rect 46848 577532 46900 577584
rect 236000 577532 236052 577584
rect 240048 577532 240100 577584
rect 349252 577532 349304 577584
rect 31392 577464 31444 577516
rect 348056 577464 348108 577516
rect 552020 577464 552072 577516
rect 556160 577464 556212 577516
rect 360936 576852 360988 576904
rect 407304 576852 407356 576904
rect 308404 576240 308456 576292
rect 330208 576240 330260 576292
rect 49056 576172 49108 576224
rect 220820 576172 220872 576224
rect 270408 576172 270460 576224
rect 307024 576172 307076 576224
rect 307760 576172 307812 576224
rect 343640 576172 343692 576224
rect 81348 576104 81400 576156
rect 347780 576104 347832 576156
rect 552020 575492 552072 575544
rect 560576 575492 560628 575544
rect 264796 574948 264848 575000
rect 354956 574948 355008 575000
rect 113088 574880 113140 574932
rect 211712 574880 211764 574932
rect 237288 574880 237340 574932
rect 347964 574880 348016 574932
rect 88248 574812 88300 574864
rect 349436 574812 349488 574864
rect 3608 574744 3660 574796
rect 384672 574744 384724 574796
rect 552020 574064 552072 574116
rect 563520 574064 563572 574116
rect 45376 573588 45428 573640
rect 223580 573588 223632 573640
rect 157248 573520 157300 573572
rect 347872 573520 347924 573572
rect 95148 573452 95200 573504
rect 331496 573452 331548 573504
rect 82728 573384 82780 573436
rect 349804 573384 349856 573436
rect 52736 573316 52788 573368
rect 405004 573316 405056 573368
rect 405372 572704 405424 572756
rect 407672 572704 407724 572756
rect 552020 572704 552072 572756
rect 582932 572704 582984 572756
rect 245844 572092 245896 572144
rect 344284 572092 344336 572144
rect 245568 572024 245620 572076
rect 353300 572024 353352 572076
rect 31484 571956 31536 572008
rect 349160 571956 349212 572008
rect 236184 571344 236236 571396
rect 363604 571344 363656 571396
rect 363696 571344 363748 571396
rect 407304 571344 407356 571396
rect 264888 571208 264940 571260
rect 350908 571208 350960 571260
rect 257896 571140 257948 571192
rect 349344 571140 349396 571192
rect 230204 571072 230256 571124
rect 361672 571072 361724 571124
rect 203892 571004 203944 571056
rect 352564 571004 352616 571056
rect 84108 570936 84160 570988
rect 237380 570936 237432 570988
rect 248328 570936 248380 570988
rect 349712 570936 349764 570988
rect 46572 570868 46624 570920
rect 260840 570868 260892 570920
rect 263508 570868 263560 570920
rect 360200 570868 360252 570920
rect 46204 570800 46256 570852
rect 296720 570800 296772 570852
rect 91008 570732 91060 570784
rect 348148 570732 348200 570784
rect 60648 570664 60700 570716
rect 352196 570664 352248 570716
rect 67548 570596 67600 570648
rect 378140 570596 378192 570648
rect 290924 569916 290976 569968
rect 368480 569916 368532 569968
rect 234528 569508 234580 569560
rect 348240 569508 348292 569560
rect 230388 569440 230440 569492
rect 352012 569440 352064 569492
rect 47676 569372 47728 569424
rect 133880 569372 133932 569424
rect 229008 569372 229060 569424
rect 356152 569372 356204 569424
rect 46480 569304 46532 569356
rect 249800 569304 249852 569356
rect 257988 569304 258040 569356
rect 353392 569304 353444 569356
rect 119988 569236 120040 569288
rect 352656 569236 352708 569288
rect 115848 569168 115900 569220
rect 353852 569168 353904 569220
rect 303988 568896 304040 568948
rect 366364 568896 366416 568948
rect 265164 568828 265216 568880
rect 357440 568828 357492 568880
rect 222016 568760 222068 568812
rect 371240 568760 371292 568812
rect 198188 568692 198240 568744
rect 357532 568692 357584 568744
rect 188528 568624 188580 568676
rect 377496 568624 377548 568676
rect 36544 568556 36596 568608
rect 407304 568556 407356 568608
rect 329656 568148 329708 568200
rect 363052 568148 363104 568200
rect 259276 568080 259328 568132
rect 348608 568080 348660 568132
rect 204168 568012 204220 568064
rect 351000 568012 351052 568064
rect 203800 567944 203852 567996
rect 356428 567944 356480 567996
rect 203984 567876 204036 567928
rect 359004 567876 359056 567928
rect 46296 567808 46348 567860
rect 234620 567808 234672 567860
rect 244188 567808 244240 567860
rect 352288 567808 352340 567860
rect 289176 567604 289228 567656
rect 374000 567604 374052 567656
rect 263232 567536 263284 567588
rect 351920 567536 351972 567588
rect 241336 567468 241388 567520
rect 358544 567468 358596 567520
rect 238668 567400 238720 567452
rect 356060 567400 356112 567452
rect 131212 567332 131264 567384
rect 354036 567332 354088 567384
rect 109960 567264 110012 567316
rect 368204 567264 368256 567316
rect 553124 567264 553176 567316
rect 559288 567264 559340 567316
rect 26056 567196 26108 567248
rect 352104 567196 352156 567248
rect 374920 567196 374972 567248
rect 407396 567196 407448 567248
rect 553308 567196 553360 567248
rect 560484 567196 560536 567248
rect 329748 566720 329800 566772
rect 353760 566720 353812 566772
rect 75644 566652 75696 566704
rect 225420 566652 225472 566704
rect 253848 566652 253900 566704
rect 349528 566652 349580 566704
rect 46756 566584 46808 566636
rect 175924 566584 175976 566636
rect 204076 566584 204128 566636
rect 353576 566584 353628 566636
rect 89628 566516 89680 566568
rect 253940 566516 253992 566568
rect 262128 566516 262180 566568
rect 348332 566516 348384 566568
rect 39580 566448 39632 566500
rect 62212 566448 62264 566500
rect 125508 566448 125560 566500
rect 353484 566448 353536 566500
rect 336280 566176 336332 566228
rect 382924 566176 382976 566228
rect 233792 566108 233844 566160
rect 347596 566108 347648 566160
rect 273168 566040 273220 566092
rect 387800 566040 387852 566092
rect 40776 565972 40828 566024
rect 372252 565972 372304 566024
rect 35624 565904 35676 565956
rect 370688 565904 370740 565956
rect 3240 565836 3292 565888
rect 17224 565836 17276 565888
rect 34428 565836 34480 565888
rect 380716 565836 380768 565888
rect 551468 565836 551520 565888
rect 552480 565836 552532 565888
rect 31208 565360 31260 565412
rect 405004 565360 405056 565412
rect 110328 565292 110380 565344
rect 219716 565292 219768 565344
rect 242808 565292 242860 565344
rect 281540 565292 281592 565344
rect 42156 565224 42208 565276
rect 172520 565224 172572 565276
rect 199384 565224 199436 565276
rect 243636 565224 243688 565276
rect 315948 565224 316000 565276
rect 376116 565224 376168 565276
rect 87696 565156 87748 565208
rect 244280 565156 244332 565208
rect 269856 565156 269908 565208
rect 387248 565156 387300 565208
rect 42432 565088 42484 565140
rect 51080 565088 51132 565140
rect 64788 565088 64840 565140
rect 247040 565088 247092 565140
rect 251824 565088 251876 565140
rect 369492 565088 369544 565140
rect 36912 565020 36964 565072
rect 111892 565020 111944 565072
rect 235080 565020 235132 565072
rect 355416 565020 355468 565072
rect 40684 564952 40736 565004
rect 162308 564952 162360 565004
rect 255136 564952 255188 565004
rect 388444 564952 388496 565004
rect 35348 564884 35400 564936
rect 168564 564884 168616 564936
rect 232504 564884 232556 564936
rect 369952 564884 370004 564936
rect 33968 564816 34020 564868
rect 244924 564816 244976 564868
rect 248328 564816 248380 564868
rect 391388 564816 391440 564868
rect 34980 564748 35032 564800
rect 124956 564748 125008 564800
rect 146208 564748 146260 564800
rect 358820 564748 358872 564800
rect 19248 564680 19300 564732
rect 301412 564680 301464 564732
rect 314936 564680 314988 564732
rect 377588 564680 377640 564732
rect 47860 564612 47912 564664
rect 58992 564612 59044 564664
rect 62488 564612 62540 564664
rect 400864 564612 400916 564664
rect 39856 564544 39908 564596
rect 381728 564544 381780 564596
rect 36636 564476 36688 564528
rect 405188 564476 405240 564528
rect 322112 564408 322164 564460
rect 356336 564408 356388 564460
rect 404636 564408 404688 564460
rect 407396 564408 407448 564460
rect 553308 564408 553360 564460
rect 563704 564408 563756 564460
rect 43444 564068 43496 564120
rect 407856 564068 407908 564120
rect 45192 564000 45244 564052
rect 89720 564000 89772 564052
rect 42064 563932 42116 563984
rect 86960 563932 87012 563984
rect 39672 563864 39724 563916
rect 85580 563864 85632 563916
rect 324688 563864 324740 563916
rect 354864 563864 354916 563916
rect 37096 563796 37148 563848
rect 84200 563796 84252 563848
rect 179696 563796 179748 563848
rect 258080 563796 258132 563848
rect 266268 563796 266320 563848
rect 346492 563796 346544 563848
rect 34152 563728 34204 563780
rect 81440 563728 81492 563780
rect 108304 563728 108356 563780
rect 230480 563728 230532 563780
rect 260748 563728 260800 563780
rect 343732 563728 343784 563780
rect 43628 563660 43680 563712
rect 91100 563660 91152 563712
rect 208032 563660 208084 563712
rect 354128 563660 354180 563712
rect 217784 563592 217836 563644
rect 370964 563592 371016 563644
rect 39304 563524 39356 563576
rect 86316 563524 86368 563576
rect 224224 563524 224276 563576
rect 390008 563524 390060 563576
rect 38108 563456 38160 563508
rect 191380 563456 191432 563508
rect 224776 563456 224828 563508
rect 395436 563456 395488 563508
rect 179144 563388 179196 563440
rect 381544 563388 381596 563440
rect 24768 563320 24820 563372
rect 255504 563320 255556 563372
rect 307760 563320 307812 563372
rect 308496 563320 308548 563372
rect 313096 563320 313148 563372
rect 361580 563320 361632 563372
rect 24492 563252 24544 563304
rect 255688 563252 255740 563304
rect 260748 563252 260800 563304
rect 372620 563252 372672 563304
rect 24308 563184 24360 563236
rect 325976 563184 326028 563236
rect 334992 563184 335044 563236
rect 367100 563184 367152 563236
rect 32496 563116 32548 563168
rect 395620 563116 395672 563168
rect 45008 563048 45060 563100
rect 181076 563048 181128 563100
rect 340144 563048 340196 563100
rect 354220 563048 354272 563100
rect 338028 562980 338080 563032
rect 342904 562980 342956 563032
rect 70308 562640 70360 562692
rect 91284 562640 91336 562692
rect 201408 562640 201460 562692
rect 379060 562640 379112 562692
rect 22928 562572 22980 562624
rect 65708 562572 65760 562624
rect 90824 562572 90876 562624
rect 171784 562572 171836 562624
rect 317972 562572 318024 562624
rect 365260 562572 365312 562624
rect 47216 562504 47268 562556
rect 74540 562504 74592 562556
rect 76656 562504 76708 562556
rect 174544 562504 174596 562556
rect 304080 562504 304132 562556
rect 363788 562504 363840 562556
rect 41880 562436 41932 562488
rect 50344 562436 50396 562488
rect 58992 562436 59044 562488
rect 164332 562436 164384 562488
rect 203156 562436 203208 562488
rect 340144 562436 340196 562488
rect 47308 562368 47360 562420
rect 75920 562368 75972 562420
rect 157800 562368 157852 562420
rect 303988 562368 304040 562420
rect 305920 562368 305972 562420
rect 365076 562368 365128 562420
rect 39764 562300 39816 562352
rect 81624 562300 81676 562352
rect 148784 562300 148836 562352
rect 336188 562300 336240 562352
rect 35808 562232 35860 562284
rect 83740 562232 83792 562284
rect 278320 562232 278372 562284
rect 347228 562232 347280 562284
rect 36268 562164 36320 562216
rect 94780 562164 94832 562216
rect 243544 562164 243596 562216
rect 363880 562164 363932 562216
rect 43352 562096 43404 562148
rect 50252 562096 50304 562148
rect 50344 562096 50396 562148
rect 99380 562096 99432 562148
rect 260288 562096 260340 562148
rect 387340 562096 387392 562148
rect 38292 562028 38344 562080
rect 45836 562028 45888 562080
rect 46020 562028 46072 562080
rect 105084 562028 105136 562080
rect 214472 562028 214524 562080
rect 347320 562028 347372 562080
rect 347688 562028 347740 562080
rect 391204 562028 391256 562080
rect 20628 561960 20680 562012
rect 43352 561960 43404 562012
rect 48228 561960 48280 562012
rect 49056 561960 49108 562012
rect 52828 561960 52880 562012
rect 138020 561960 138072 562012
rect 250444 561960 250496 562012
rect 403624 561960 403676 562012
rect 22836 561892 22888 561944
rect 113456 561892 113508 561944
rect 186872 561892 186924 561944
rect 340144 561892 340196 561944
rect 24400 561824 24452 561876
rect 51540 561824 51592 561876
rect 52000 561824 52052 561876
rect 181628 561824 181680 561876
rect 192576 561824 192628 561876
rect 365720 561824 365772 561876
rect 41328 561756 41380 561808
rect 193864 561756 193916 561808
rect 340052 561756 340104 561808
rect 358360 561756 358412 561808
rect 31484 561688 31536 561740
rect 138572 561688 138624 561740
rect 140504 561688 140556 561740
rect 319168 561688 319220 561740
rect 325608 561688 325660 561740
rect 355232 561688 355284 561740
rect 47124 561552 47176 561604
rect 66260 561552 66312 561604
rect 29920 561484 29972 561536
rect 51172 561484 51224 561536
rect 47492 561416 47544 561468
rect 73160 561416 73212 561468
rect 21732 561348 21784 561400
rect 53840 561348 53892 561400
rect 35532 561280 35584 561332
rect 67732 561280 67784 561332
rect 25596 561212 25648 561264
rect 58072 561212 58124 561264
rect 28724 561144 28776 561196
rect 62120 561144 62172 561196
rect 307668 561144 307720 561196
rect 355324 561144 355376 561196
rect 27252 561076 27304 561128
rect 60832 561076 60884 561128
rect 337568 561076 337620 561128
rect 405280 561076 405332 561128
rect 38200 561008 38252 561060
rect 71780 561008 71832 561060
rect 315672 561008 315724 561060
rect 395344 561008 395396 561060
rect 34060 560940 34112 560992
rect 67640 560940 67692 560992
rect 299388 560940 299440 560992
rect 380256 560940 380308 560992
rect 287888 560872 287940 560924
rect 374644 560872 374696 560924
rect 244832 560804 244884 560856
rect 376852 560804 376904 560856
rect 240968 560736 241020 560788
rect 376760 560736 376812 560788
rect 235816 560668 235868 560720
rect 396724 560668 396776 560720
rect 183008 560600 183060 560652
rect 394056 560600 394108 560652
rect 116584 560532 116636 560584
rect 358636 560532 358688 560584
rect 32772 560464 32824 560516
rect 381820 560464 381872 560516
rect 39488 560396 39540 560448
rect 395896 560396 395948 560448
rect 43536 560328 43588 560380
rect 405096 560328 405148 560380
rect 553308 560328 553360 560380
rect 566740 560328 566792 560380
rect 37832 560260 37884 560312
rect 407396 560260 407448 560312
rect 553124 560260 553176 560312
rect 568028 560260 568080 560312
rect 347596 560192 347648 560244
rect 351276 560192 351328 560244
rect 39396 559580 39448 559632
rect 52828 559988 52880 560040
rect 319168 559988 319220 560040
rect 45744 559920 45796 559972
rect 48872 559920 48924 559972
rect 52000 559920 52052 559972
rect 36820 559512 36872 559564
rect 41052 558900 41104 558952
rect 148968 559920 149020 559972
rect 327724 559920 327776 559972
rect 336648 559920 336700 559972
rect 340696 559920 340748 559972
rect 347228 559920 347280 559972
rect 347320 559920 347372 559972
rect 389180 559648 389232 559700
rect 407948 559580 408000 559632
rect 407672 559512 407724 559564
rect 349988 559444 350040 559496
rect 364432 559036 364484 559088
rect 356244 558968 356296 559020
rect 349988 558900 350040 558952
rect 380532 558900 380584 558952
rect 552940 557948 552992 558000
rect 556620 557948 556672 558000
rect 553308 557540 553360 557592
rect 568672 557540 568724 557592
rect 405280 557200 405332 557252
rect 407672 557200 407724 557252
rect 553308 556520 553360 556572
rect 559748 556520 559800 556572
rect 44548 556180 44600 556232
rect 46112 556180 46164 556232
rect 394516 556180 394568 556232
rect 407396 556180 407448 556232
rect 553308 556180 553360 556232
rect 573548 556180 573600 556232
rect 350448 554684 350500 554736
rect 353300 554684 353352 554736
rect 552020 553664 552072 553716
rect 555148 553664 555200 553716
rect 407856 552644 407908 552696
rect 408316 552644 408368 552696
rect 387616 552032 387668 552084
rect 407488 552032 407540 552084
rect 351368 551964 351420 552016
rect 407396 551964 407448 552016
rect 41788 551148 41840 551200
rect 46112 551148 46164 551200
rect 350448 551080 350500 551132
rect 356796 551080 356848 551132
rect 42340 550808 42392 550860
rect 46112 550808 46164 550860
rect 552020 550808 552072 550860
rect 555240 550808 555292 550860
rect 404176 550604 404228 550656
rect 407396 550604 407448 550656
rect 553308 550604 553360 550656
rect 562600 550604 562652 550656
rect 30196 549244 30248 549296
rect 46112 549244 46164 549296
rect 358452 549244 358504 549296
rect 407396 549244 407448 549296
rect 553308 549244 553360 549296
rect 574192 549244 574244 549296
rect 350172 549176 350224 549228
rect 352104 549176 352156 549228
rect 405188 549176 405240 549228
rect 407488 549176 407540 549228
rect 30288 547884 30340 547936
rect 46112 547884 46164 547936
rect 350448 546592 350500 546644
rect 384304 546592 384356 546644
rect 371884 546524 371936 546576
rect 407396 546524 407448 546576
rect 350264 546456 350316 546508
rect 385960 546456 386012 546508
rect 551376 546456 551428 546508
rect 552020 546456 552072 546508
rect 46112 545980 46164 546032
rect 46756 545980 46808 546032
rect 34336 545096 34388 545148
rect 46756 545096 46808 545148
rect 405188 543804 405240 543856
rect 407488 543804 407540 543856
rect 552572 543804 552624 543856
rect 555148 543804 555200 543856
rect 43076 543736 43128 543788
rect 46756 543736 46808 543788
rect 389824 543736 389876 543788
rect 407396 543736 407448 543788
rect 350448 542376 350500 542428
rect 398380 542376 398432 542428
rect 354036 542308 354088 542360
rect 407396 542308 407448 542360
rect 22008 540948 22060 541000
rect 46756 540948 46808 541000
rect 553308 539656 553360 539708
rect 562232 539656 562284 539708
rect 553124 539588 553176 539640
rect 567292 539588 567344 539640
rect 350448 538228 350500 538280
rect 365168 538228 365220 538280
rect 43444 538160 43496 538212
rect 46756 538160 46808 538212
rect 350448 536800 350500 536852
rect 386420 536800 386472 536852
rect 553308 535440 553360 535492
rect 560760 535440 560812 535492
rect 350448 534080 350500 534132
rect 362224 534080 362276 534132
rect 391296 534080 391348 534132
rect 407304 534080 407356 534132
rect 553308 534080 553360 534132
rect 581460 534080 581512 534132
rect 350264 532788 350316 532840
rect 358912 532788 358964 532840
rect 27436 532720 27488 532772
rect 46756 532720 46808 532772
rect 350448 532720 350500 532772
rect 386144 532720 386196 532772
rect 395712 532720 395764 532772
rect 407304 532720 407356 532772
rect 552388 532516 552440 532568
rect 553676 532516 553728 532568
rect 25872 531292 25924 531344
rect 46756 531292 46808 531344
rect 350448 531292 350500 531344
rect 353668 531292 353720 531344
rect 401324 531292 401376 531344
rect 407304 531292 407356 531344
rect 552388 530476 552440 530528
rect 553768 530476 553820 530528
rect 553308 530272 553360 530324
rect 558000 530272 558052 530324
rect 18972 529932 19024 529984
rect 46756 529932 46808 529984
rect 350448 529932 350500 529984
rect 380440 529932 380492 529984
rect 40408 528572 40460 528624
rect 46112 528572 46164 528624
rect 350448 527144 350500 527196
rect 366456 527144 366508 527196
rect 553308 527144 553360 527196
rect 566280 527144 566332 527196
rect 407120 526464 407172 526516
rect 407304 526464 407356 526516
rect 552388 526260 552440 526312
rect 553768 526260 553820 526312
rect 350448 525920 350500 525972
rect 356888 525920 356940 525972
rect 400128 525784 400180 525836
rect 407304 525784 407356 525836
rect 44088 525716 44140 525768
rect 46756 525716 46808 525768
rect 570696 525716 570748 525768
rect 580172 525716 580224 525768
rect 46020 524424 46072 524476
rect 47584 524424 47636 524476
rect 395988 524424 396040 524476
rect 407120 524424 407172 524476
rect 350264 524356 350316 524408
rect 353760 524356 353812 524408
rect 350448 522996 350500 523048
rect 369400 522996 369452 523048
rect 385868 522996 385920 523048
rect 407304 522996 407356 523048
rect 383016 522928 383068 522980
rect 407120 522928 407172 522980
rect 407488 522928 407540 522980
rect 409144 522928 409196 522980
rect 402704 521636 402756 521688
rect 407396 521636 407448 521688
rect 40960 521500 41012 521552
rect 46296 521500 46348 521552
rect 23296 520344 23348 520396
rect 45560 520344 45612 520396
rect 17868 520276 17920 520328
rect 45652 520276 45704 520328
rect 350172 520276 350224 520328
rect 352104 520276 352156 520328
rect 552020 520276 552072 520328
rect 571524 520276 571576 520328
rect 45836 519528 45888 519580
rect 46020 519528 46072 519580
rect 552020 519256 552072 519308
rect 553676 519256 553728 519308
rect 552020 518984 552072 519036
rect 564716 518984 564768 519036
rect 350448 517556 350500 517608
rect 381636 517556 381688 517608
rect 388260 517556 388312 517608
rect 407120 517556 407172 517608
rect 373448 517488 373500 517540
rect 407304 517488 407356 517540
rect 350264 516196 350316 516248
rect 387156 516196 387208 516248
rect 397368 516196 397420 516248
rect 407120 516196 407172 516248
rect 34244 516128 34296 516180
rect 45560 516128 45612 516180
rect 350448 516128 350500 516180
rect 361856 516128 361908 516180
rect 370504 516128 370556 516180
rect 407304 516128 407356 516180
rect 552020 516128 552072 516180
rect 570788 516128 570840 516180
rect 405096 516060 405148 516112
rect 407580 516060 407632 516112
rect 3424 514768 3476 514820
rect 26976 514768 27028 514820
rect 38568 514768 38620 514820
rect 45560 514768 45612 514820
rect 552020 514768 552072 514820
rect 564808 514768 564860 514820
rect 45836 514020 45888 514072
rect 46112 514020 46164 514072
rect 350264 513408 350316 513460
rect 353760 513408 353812 513460
rect 38016 513340 38068 513392
rect 46204 513340 46256 513392
rect 350448 513340 350500 513392
rect 394148 513340 394200 513392
rect 389916 513272 389968 513324
rect 407120 513272 407172 513324
rect 377680 511980 377732 512032
rect 407120 511980 407172 512032
rect 39856 510552 39908 510604
rect 46756 510552 46808 510604
rect 553308 509600 553360 509652
rect 559840 509600 559892 509652
rect 44916 509260 44968 509312
rect 46204 509260 46256 509312
rect 389916 509260 389968 509312
rect 407120 509260 407172 509312
rect 350448 509192 350500 509244
rect 406384 509192 406436 509244
rect 40684 508308 40736 508360
rect 44916 508308 44968 508360
rect 350448 506472 350500 506524
rect 375380 506472 375432 506524
rect 350264 506404 350316 506456
rect 399576 506404 399628 506456
rect 553308 506404 553360 506456
rect 570604 506404 570656 506456
rect 19156 505112 19208 505164
rect 46756 505112 46808 505164
rect 350448 505112 350500 505164
rect 383108 505112 383160 505164
rect 350448 503684 350500 503736
rect 360292 503684 360344 503736
rect 553308 503684 553360 503736
rect 574560 503684 574612 503736
rect 553308 502392 553360 502444
rect 557724 502392 557776 502444
rect 39948 502052 40000 502104
rect 45836 502052 45888 502104
rect 553308 501304 553360 501356
rect 559196 501304 559248 501356
rect 553308 500964 553360 501016
rect 574928 500964 574980 501016
rect 40868 500896 40920 500948
rect 46756 500896 46808 500948
rect 402428 500896 402480 500948
rect 407120 500896 407172 500948
rect 553308 499808 553360 499860
rect 557632 499808 557684 499860
rect 350448 499536 350500 499588
rect 384764 499536 384816 499588
rect 553308 498448 553360 498500
rect 557540 498448 557592 498500
rect 350448 498176 350500 498228
rect 354036 498176 354088 498228
rect 42524 498108 42576 498160
rect 45836 498108 45888 498160
rect 46020 497020 46072 497072
rect 46388 497020 46440 497072
rect 384488 496816 384540 496868
rect 407120 496816 407172 496868
rect 40776 496748 40828 496800
rect 46756 496748 46808 496800
rect 39120 495456 39172 495508
rect 46388 495456 46440 495508
rect 350448 495456 350500 495508
rect 386052 495456 386104 495508
rect 401140 495456 401192 495508
rect 407120 495456 407172 495508
rect 41972 495388 42024 495440
rect 46756 495388 46808 495440
rect 350448 493416 350500 493468
rect 351276 493416 351328 493468
rect 23204 492668 23256 492720
rect 46756 492668 46808 492720
rect 384396 492668 384448 492720
rect 407120 492668 407172 492720
rect 552664 492668 552716 492720
rect 563796 492668 563848 492720
rect 350264 491376 350316 491428
rect 359096 491376 359148 491428
rect 350448 491308 350500 491360
rect 367928 491308 367980 491360
rect 40868 489948 40920 490000
rect 46756 489948 46808 490000
rect 350448 489948 350500 490000
rect 379520 489948 379572 490000
rect 381912 489948 381964 490000
rect 407120 489948 407172 490000
rect 28632 489880 28684 489932
rect 46388 489880 46440 489932
rect 350264 489880 350316 489932
rect 392768 489880 392820 489932
rect 42616 489812 42668 489864
rect 46756 489812 46808 489864
rect 350172 489812 350224 489864
rect 352288 489812 352340 489864
rect 553308 488860 553360 488912
rect 559104 488860 559156 488912
rect 393044 488588 393096 488640
rect 407304 488588 407356 488640
rect 384580 488520 384632 488572
rect 407120 488520 407172 488572
rect 350264 488452 350316 488504
rect 372068 488452 372120 488504
rect 44640 488180 44692 488232
rect 46388 488180 46440 488232
rect 401232 487160 401284 487212
rect 407120 487160 407172 487212
rect 553308 487160 553360 487212
rect 572904 487160 572956 487212
rect 39856 485800 39908 485852
rect 46756 485800 46808 485852
rect 394332 485800 394384 485852
rect 407120 485800 407172 485852
rect 21640 484372 21692 484424
rect 46756 484372 46808 484424
rect 349988 484372 350040 484424
rect 352288 484372 352340 484424
rect 373540 484372 373592 484424
rect 407120 484372 407172 484424
rect 387432 483080 387484 483132
rect 407120 483080 407172 483132
rect 19064 483012 19116 483064
rect 46756 483012 46808 483064
rect 350264 483012 350316 483064
rect 377772 483012 377824 483064
rect 552664 483012 552716 483064
rect 574376 483012 574428 483064
rect 350448 481652 350500 481704
rect 370044 481652 370096 481704
rect 402796 481652 402848 481704
rect 407120 481652 407172 481704
rect 41880 480428 41932 480480
rect 45836 480428 45888 480480
rect 350264 480292 350316 480344
rect 366088 480292 366140 480344
rect 350448 480224 350500 480276
rect 370136 480224 370188 480276
rect 383016 478864 383068 478916
rect 407120 478864 407172 478916
rect 44732 478660 44784 478712
rect 46664 478660 46716 478712
rect 553308 477504 553360 477556
rect 562416 477504 562468 477556
rect 348516 476212 348568 476264
rect 349804 476212 349856 476264
rect 350172 476144 350224 476196
rect 361948 476144 362000 476196
rect 23112 476076 23164 476128
rect 46756 476076 46808 476128
rect 350264 476076 350316 476128
rect 370596 476076 370648 476128
rect 403348 474784 403400 474836
rect 407304 474784 407356 474836
rect 552572 474784 552624 474836
rect 561128 474784 561180 474836
rect 399576 474716 399628 474768
rect 407120 474716 407172 474768
rect 553308 474716 553360 474768
rect 561956 474716 562008 474768
rect 45100 474648 45152 474700
rect 46480 474648 46532 474700
rect 43536 474580 43588 474632
rect 46572 474580 46624 474632
rect 394424 473424 394476 473476
rect 407120 473424 407172 473476
rect 350264 473356 350316 473408
rect 352380 473356 352432 473408
rect 372068 473356 372120 473408
rect 407304 473356 407356 473408
rect 350448 471996 350500 472048
rect 353944 471996 353996 472048
rect 553308 470568 553360 470620
rect 567844 470568 567896 470620
rect 570696 470568 570748 470620
rect 580172 470568 580224 470620
rect 33600 469208 33652 469260
rect 46756 469208 46808 469260
rect 361028 469208 361080 469260
rect 407120 469208 407172 469260
rect 553308 469208 553360 469260
rect 577320 469208 577372 469260
rect 404084 469140 404136 469192
rect 407304 469140 407356 469192
rect 40776 467916 40828 467968
rect 46756 467916 46808 467968
rect 23020 467848 23072 467900
rect 46572 467848 46624 467900
rect 388904 467848 388956 467900
rect 407120 467848 407172 467900
rect 350448 466420 350500 466472
rect 392584 466420 392636 466472
rect 553308 466420 553360 466472
rect 567476 466420 567528 466472
rect 350264 466352 350316 466404
rect 403808 466352 403860 466404
rect 397276 465060 397328 465112
rect 407120 465060 407172 465112
rect 552020 465060 552072 465112
rect 575940 465060 575992 465112
rect 40592 464108 40644 464160
rect 46756 464108 46808 464160
rect 552020 463904 552072 463956
rect 556252 463904 556304 463956
rect 18880 463700 18932 463752
rect 45652 463700 45704 463752
rect 383200 463700 383252 463752
rect 407120 463700 407172 463752
rect 35624 463632 35676 463684
rect 46756 463632 46808 463684
rect 350448 462476 350500 462528
rect 395804 462476 395856 462528
rect 350264 462408 350316 462460
rect 376300 462408 376352 462460
rect 392676 462408 392728 462460
rect 407120 462408 407172 462460
rect 3516 462340 3568 462392
rect 19984 462340 20036 462392
rect 394240 462340 394292 462392
rect 407304 462340 407356 462392
rect 552020 462340 552072 462392
rect 573088 462340 573140 462392
rect 350448 461048 350500 461100
rect 362960 461048 363012 461100
rect 350264 460980 350316 461032
rect 364524 460980 364576 461032
rect 21916 460912 21968 460964
rect 46756 460912 46808 460964
rect 362316 460912 362368 460964
rect 407120 460912 407172 460964
rect 39488 460844 39540 460896
rect 46572 460844 46624 460896
rect 350448 459552 350500 459604
rect 396908 459552 396960 459604
rect 552020 459552 552072 459604
rect 560852 459552 560904 459604
rect 552020 459008 552072 459060
rect 553860 459008 553912 459060
rect 31392 458192 31444 458244
rect 46756 458192 46808 458244
rect 403900 458192 403952 458244
rect 407120 458192 407172 458244
rect 350448 456832 350500 456884
rect 367192 456832 367244 456884
rect 350264 456764 350316 456816
rect 375472 456764 375524 456816
rect 391480 456764 391532 456816
rect 407120 456764 407172 456816
rect 552020 456764 552072 456816
rect 576216 456764 576268 456816
rect 43996 456696 44048 456748
rect 46756 456696 46808 456748
rect 386052 456696 386104 456748
rect 407304 456696 407356 456748
rect 552020 456016 552072 456068
rect 553952 456016 554004 456068
rect 348976 455336 349028 455388
rect 350540 455336 350592 455388
rect 369492 455336 369544 455388
rect 407120 455336 407172 455388
rect 350448 454044 350500 454096
rect 380624 454044 380676 454096
rect 405280 454044 405332 454096
rect 407672 454044 407724 454096
rect 553308 454044 553360 454096
rect 565912 454044 565964 454096
rect 552848 452752 552900 452804
rect 556344 452752 556396 452804
rect 366548 452616 366600 452668
rect 407120 452616 407172 452668
rect 350448 451256 350500 451308
rect 386052 451256 386104 451308
rect 400956 451256 401008 451308
rect 407120 451256 407172 451308
rect 34428 451188 34480 451240
rect 46756 451188 46808 451240
rect 350448 449896 350500 449948
rect 362500 449896 362552 449948
rect 553308 449896 553360 449948
rect 578332 449896 578384 449948
rect 3148 448536 3200 448588
rect 17316 448536 17368 448588
rect 383476 448536 383528 448588
rect 407120 448536 407172 448588
rect 552572 448536 552624 448588
rect 575664 448536 575716 448588
rect 348884 447108 348936 447160
rect 349160 447108 349212 447160
rect 350448 447108 350500 447160
rect 367284 447108 367336 447160
rect 403532 447108 403584 447160
rect 407304 447108 407356 447160
rect 395620 447040 395672 447092
rect 407120 447040 407172 447092
rect 29644 445748 29696 445800
rect 46756 445748 46808 445800
rect 350264 445748 350316 445800
rect 370780 445748 370832 445800
rect 552572 445748 552624 445800
rect 566372 445748 566424 445800
rect 350448 445680 350500 445732
rect 399668 445680 399720 445732
rect 373632 445612 373684 445664
rect 407120 445612 407172 445664
rect 27068 444388 27120 444440
rect 46756 444388 46808 444440
rect 552572 444388 552624 444440
rect 581276 444388 581328 444440
rect 38476 442960 38528 443012
rect 46756 442960 46808 443012
rect 553308 442960 553360 443012
rect 569132 442960 569184 443012
rect 362408 441600 362460 441652
rect 407120 441600 407172 441652
rect 395896 441532 395948 441584
rect 407304 441532 407356 441584
rect 350448 440240 350500 440292
rect 395620 440240 395672 440292
rect 40684 438948 40736 439000
rect 46756 438948 46808 439000
rect 41696 438880 41748 438932
rect 46020 438880 46072 438932
rect 386236 438880 386288 438932
rect 407120 438880 407172 438932
rect 405004 438812 405056 438864
rect 407488 438812 407540 438864
rect 562416 437588 562468 437640
rect 563244 437588 563296 437640
rect 350264 437452 350316 437504
rect 398472 437452 398524 437504
rect 553308 437452 553360 437504
rect 562324 437452 562376 437504
rect 350448 437384 350500 437436
rect 403716 437384 403768 437436
rect 553032 437384 553084 437436
rect 556896 437384 556948 437436
rect 348884 436296 348936 436348
rect 349160 436296 349212 436348
rect 43536 436092 43588 436144
rect 46756 436092 46808 436144
rect 397184 436092 397236 436144
rect 407120 436092 407172 436144
rect 553308 436092 553360 436144
rect 577688 436092 577740 436144
rect 553032 435956 553084 436008
rect 553308 435956 553360 436008
rect 350448 434800 350500 434852
rect 370228 434800 370280 434852
rect 43996 434732 44048 434784
rect 46756 434732 46808 434784
rect 363972 434732 364024 434784
rect 407120 434732 407172 434784
rect 33876 433304 33928 433356
rect 46756 433304 46808 433356
rect 42524 431944 42576 431996
rect 46756 431944 46808 431996
rect 577596 431740 577648 431792
rect 579896 431740 579948 431792
rect 350448 430652 350500 430704
rect 373816 430652 373868 430704
rect 350264 430584 350316 430636
rect 397000 430584 397052 430636
rect 552204 430176 552256 430228
rect 555056 430176 555108 430228
rect 402612 429224 402664 429276
rect 407120 429224 407172 429276
rect 40500 427864 40552 427916
rect 46664 427864 46716 427916
rect 396632 427864 396684 427916
rect 407120 427864 407172 427916
rect 33784 427796 33836 427848
rect 46756 427796 46808 427848
rect 350448 427796 350500 427848
rect 375012 427796 375064 427848
rect 553032 427796 553084 427848
rect 563888 427796 563940 427848
rect 369492 426572 369544 426624
rect 407212 426572 407264 426624
rect 361120 426504 361172 426556
rect 407120 426504 407172 426556
rect 350448 426436 350500 426488
rect 399668 426436 399720 426488
rect 553032 426436 553084 426488
rect 577136 426436 577188 426488
rect 43444 425076 43496 425128
rect 45652 425076 45704 425128
rect 350448 425076 350500 425128
rect 359188 425076 359240 425128
rect 553032 425076 553084 425128
rect 569500 425076 569552 425128
rect 553032 423716 553084 423768
rect 570604 423716 570656 423768
rect 24124 423648 24176 423700
rect 46756 423648 46808 423700
rect 374828 423648 374880 423700
rect 407120 423648 407172 423700
rect 552940 423648 552992 423700
rect 574836 423648 574888 423700
rect 350448 422288 350500 422340
rect 376576 422288 376628 422340
rect 393872 422288 393924 422340
rect 407120 422288 407172 422340
rect 349988 420996 350040 421048
rect 352472 420996 352524 421048
rect 552204 420996 552256 421048
rect 554964 420996 555016 421048
rect 35164 420928 35216 420980
rect 45652 420928 45704 420980
rect 350448 420928 350500 420980
rect 383384 420928 383436 420980
rect 570788 420180 570840 420232
rect 580448 420180 580500 420232
rect 553032 420112 553084 420164
rect 559564 420112 559616 420164
rect 28356 419568 28408 419620
rect 45652 419568 45704 419620
rect 350448 419568 350500 419620
rect 368572 419568 368624 419620
rect 369584 419568 369636 419620
rect 407212 419568 407264 419620
rect 26792 419500 26844 419552
rect 45928 419500 45980 419552
rect 356980 419500 357032 419552
rect 407120 419500 407172 419552
rect 350448 418208 350500 418260
rect 382004 418208 382056 418260
rect 39488 418140 39540 418192
rect 45928 418140 45980 418192
rect 372344 418140 372396 418192
rect 407120 418140 407172 418192
rect 350448 416780 350500 416832
rect 379152 416780 379204 416832
rect 380716 416712 380768 416764
rect 407120 416712 407172 416764
rect 553032 416032 553084 416084
rect 559472 416032 559524 416084
rect 28816 415488 28868 415540
rect 45652 415488 45704 415540
rect 24216 415420 24268 415472
rect 45928 415420 45980 415472
rect 553032 415420 553084 415472
rect 579712 415420 579764 415472
rect 350448 414060 350500 414112
rect 374736 414060 374788 414112
rect 20168 413992 20220 414044
rect 46756 413992 46808 414044
rect 350264 413992 350316 414044
rect 376484 413992 376536 414044
rect 388996 413992 389048 414044
rect 407120 413992 407172 414044
rect 552388 412768 552440 412820
rect 555332 412768 555384 412820
rect 553032 412632 553084 412684
rect 580080 412632 580132 412684
rect 35624 411272 35676 411324
rect 46756 411272 46808 411324
rect 350448 411272 350500 411324
rect 375104 411272 375156 411324
rect 395896 411272 395948 411324
rect 407120 411272 407172 411324
rect 2964 411204 3016 411256
rect 32496 411204 32548 411256
rect 359556 409844 359608 409896
rect 407120 409844 407172 409896
rect 553032 409844 553084 409896
rect 570236 409844 570288 409896
rect 399944 408484 399996 408536
rect 407120 408484 407172 408536
rect 348976 407736 349028 407788
rect 350172 407736 350224 407788
rect 21456 407124 21508 407176
rect 46756 407124 46808 407176
rect 368020 405696 368072 405748
rect 407120 405696 407172 405748
rect 400036 405628 400088 405680
rect 407212 405628 407264 405680
rect 553032 405628 553084 405680
rect 579160 405628 579212 405680
rect 350264 404404 350316 404456
rect 364616 404404 364668 404456
rect 350448 404336 350500 404388
rect 368296 404336 368348 404388
rect 553032 403656 553084 403708
rect 557816 403656 557868 403708
rect 41972 402976 42024 403028
rect 46756 402976 46808 403028
rect 553032 402976 553084 403028
rect 579896 402976 579948 403028
rect 42156 402092 42208 402144
rect 44180 402092 44232 402144
rect 42156 400188 42208 400240
rect 46756 400188 46808 400240
rect 350448 400188 350500 400240
rect 372160 400188 372212 400240
rect 405004 400188 405056 400240
rect 407488 400188 407540 400240
rect 553032 400188 553084 400240
rect 582748 400188 582800 400240
rect 403992 400120 404044 400172
rect 407120 400120 407172 400172
rect 20444 398828 20496 398880
rect 46756 398828 46808 398880
rect 350448 398828 350500 398880
rect 360476 398828 360528 398880
rect 3516 397468 3568 397520
rect 17408 397468 17460 397520
rect 350448 397468 350500 397520
rect 388720 397468 388772 397520
rect 392952 397468 393004 397520
rect 407120 397468 407172 397520
rect 349804 396788 349856 396840
rect 352656 396788 352708 396840
rect 350448 396040 350500 396092
rect 382740 396040 382792 396092
rect 349896 395972 349948 396024
rect 351184 395972 351236 396024
rect 400036 394748 400088 394800
rect 407212 394748 407264 394800
rect 20536 394680 20588 394732
rect 46756 394680 46808 394732
rect 350264 394680 350316 394732
rect 352840 394680 352892 394732
rect 382188 394680 382240 394732
rect 407120 394680 407172 394732
rect 553032 394680 553084 394732
rect 581736 394680 581788 394732
rect 350448 394612 350500 394664
rect 392860 394612 392912 394664
rect 552204 393728 552256 393780
rect 554964 393728 555016 393780
rect 390100 393320 390152 393372
rect 407120 393320 407172 393372
rect 37924 392028 37976 392080
rect 46020 392028 46072 392080
rect 25688 391960 25740 392012
rect 46112 391960 46164 392012
rect 348884 391960 348936 392012
rect 349344 391960 349396 392012
rect 350448 391960 350500 392012
rect 402428 391960 402480 392012
rect 377864 390600 377916 390652
rect 407212 390600 407264 390652
rect 553032 390600 553084 390652
rect 581644 390600 581696 390652
rect 349620 390532 349672 390584
rect 351276 390532 351328 390584
rect 368112 390532 368164 390584
rect 407120 390532 407172 390584
rect 350448 390464 350500 390516
rect 395528 390464 395580 390516
rect 17776 389172 17828 389224
rect 46480 389172 46532 389224
rect 350264 389172 350316 389224
rect 373724 389172 373776 389224
rect 391756 389172 391808 389224
rect 407120 389172 407172 389224
rect 553032 389172 553084 389224
rect 570420 389172 570472 389224
rect 350448 387812 350500 387864
rect 377956 387812 378008 387864
rect 553032 387812 553084 387864
rect 579804 387812 579856 387864
rect 350264 387744 350316 387796
rect 400956 387744 401008 387796
rect 29828 386384 29880 386436
rect 46480 386384 46532 386436
rect 553032 386384 553084 386436
rect 561036 386384 561088 386436
rect 32404 386316 32456 386368
rect 46112 386316 46164 386368
rect 350448 386316 350500 386368
rect 352196 386316 352248 386368
rect 368204 386316 368256 386368
rect 407120 386316 407172 386368
rect 36176 385024 36228 385076
rect 46480 385024 46532 385076
rect 553032 385024 553084 385076
rect 562140 385024 562192 385076
rect 349068 384956 349120 385008
rect 352656 384956 352708 385008
rect 350448 384276 350500 384328
rect 359280 384276 359332 384328
rect 403164 383936 403216 383988
rect 407120 383936 407172 383988
rect 36728 383596 36780 383648
rect 46480 383596 46532 383648
rect 350264 382236 350316 382288
rect 400956 382236 401008 382288
rect 402520 382236 402572 382288
rect 407120 382236 407172 382288
rect 553032 381488 553084 381540
rect 558092 381488 558144 381540
rect 46480 381080 46532 381132
rect 46848 381080 46900 381132
rect 36452 380944 36504 380996
rect 45008 380944 45060 380996
rect 350080 380944 350132 380996
rect 380900 380944 380952 380996
rect 28448 380876 28500 380928
rect 46848 380876 46900 380928
rect 350264 380876 350316 380928
rect 385592 380876 385644 380928
rect 395528 380876 395580 380928
rect 407120 380876 407172 380928
rect 31300 379516 31352 379568
rect 46848 379516 46900 379568
rect 408132 378768 408184 378820
rect 409328 378768 409380 378820
rect 553032 378292 553084 378344
rect 557908 378292 557960 378344
rect 392860 378156 392912 378208
rect 407120 378156 407172 378208
rect 572076 378156 572128 378208
rect 580172 378156 580224 378208
rect 350080 378088 350132 378140
rect 352564 378088 352616 378140
rect 350264 376728 350316 376780
rect 408500 376728 408552 376780
rect 553032 376728 553084 376780
rect 582840 376728 582892 376780
rect 350080 375368 350132 375420
rect 403716 375368 403768 375420
rect 350264 375300 350316 375352
rect 374920 375300 374972 375352
rect 552204 372648 552256 372700
rect 555056 372648 555108 372700
rect 28264 372580 28316 372632
rect 46848 372580 46900 372632
rect 350264 372580 350316 372632
rect 374920 372580 374972 372632
rect 397092 372580 397144 372632
rect 407120 372580 407172 372632
rect 29736 371220 29788 371272
rect 46848 371220 46900 371272
rect 350264 371220 350316 371272
rect 380716 371220 380768 371272
rect 43812 371152 43864 371204
rect 45652 371152 45704 371204
rect 350080 371152 350132 371204
rect 356428 371152 356480 371204
rect 362500 371152 362552 371204
rect 407120 371152 407172 371204
rect 553032 369860 553084 369912
rect 560668 369860 560720 369912
rect 407672 369112 407724 369164
rect 408132 369112 408184 369164
rect 552204 368568 552256 368620
rect 555424 368568 555476 368620
rect 43812 368500 43864 368552
rect 46848 368500 46900 368552
rect 553032 368500 553084 368552
rect 572996 368500 573048 368552
rect 349068 368432 349120 368484
rect 349344 368432 349396 368484
rect 552020 367956 552072 368008
rect 553768 367956 553820 368008
rect 32128 367072 32180 367124
rect 46848 367072 46900 367124
rect 32772 367004 32824 367056
rect 46020 367004 46072 367056
rect 553032 365780 553084 365832
rect 567568 365780 567620 365832
rect 552940 365712 552992 365764
rect 578424 365712 578476 365764
rect 552020 365168 552072 365220
rect 554136 365168 554188 365220
rect 27160 362924 27212 362976
rect 46848 362924 46900 362976
rect 350080 362924 350132 362976
rect 352564 362924 352616 362976
rect 45284 361496 45336 361548
rect 46480 361496 46532 361548
rect 370780 361496 370832 361548
rect 407120 361496 407172 361548
rect 553032 360408 553084 360460
rect 557908 360408 557960 360460
rect 366640 360204 366692 360256
rect 407120 360204 407172 360256
rect 552940 360204 552992 360256
rect 574744 360204 574796 360256
rect 350264 358776 350316 358828
rect 363144 358776 363196 358828
rect 37832 358708 37884 358760
rect 46848 358708 46900 358760
rect 553032 358708 553084 358760
rect 572076 358708 572128 358760
rect 350264 357960 350316 358012
rect 355508 357960 355560 358012
rect 46480 357756 46532 357808
rect 46848 357756 46900 357808
rect 3148 357416 3200 357468
rect 28080 357416 28132 357468
rect 552940 357416 552992 357468
rect 573272 357416 573324 357468
rect 369676 356192 369728 356244
rect 407120 356192 407172 356244
rect 350264 356124 350316 356176
rect 378232 356124 378284 356176
rect 350264 355988 350316 356040
rect 396816 355988 396868 356040
rect 37832 354696 37884 354748
rect 46480 354696 46532 354748
rect 350264 354696 350316 354748
rect 359648 354696 359700 354748
rect 553032 354696 553084 354748
rect 568120 354696 568172 354748
rect 376392 353268 376444 353320
rect 407120 353268 407172 353320
rect 553032 353268 553084 353320
rect 575848 353268 575900 353320
rect 36544 353200 36596 353252
rect 46480 353200 46532 353252
rect 398840 351976 398892 352028
rect 407120 351976 407172 352028
rect 388812 351908 388864 351960
rect 407212 351908 407264 351960
rect 553124 350888 553176 350940
rect 558184 350888 558236 350940
rect 350264 350548 350316 350600
rect 362040 350548 362092 350600
rect 384856 350548 384908 350600
rect 407120 350548 407172 350600
rect 552848 350548 552900 350600
rect 583024 350548 583076 350600
rect 350080 349188 350132 349240
rect 364064 349188 364116 349240
rect 21548 349120 21600 349172
rect 46480 349120 46532 349172
rect 350264 349120 350316 349172
rect 365444 349120 365496 349172
rect 372436 349120 372488 349172
rect 407120 349120 407172 349172
rect 553124 349120 553176 349172
rect 583484 349120 583536 349172
rect 553124 346468 553176 346520
rect 575756 346468 575808 346520
rect 29552 346400 29604 346452
rect 46480 346400 46532 346452
rect 392400 346400 392452 346452
rect 407120 346400 407172 346452
rect 553032 346400 553084 346452
rect 578700 346400 578752 346452
rect 3516 345108 3568 345160
rect 29460 345108 29512 345160
rect 20352 345040 20404 345092
rect 46480 345040 46532 345092
rect 350264 345040 350316 345092
rect 379612 345040 379664 345092
rect 376576 344972 376628 345024
rect 407120 344972 407172 345024
rect 350264 343680 350316 343732
rect 361304 343680 361356 343732
rect 350080 343612 350132 343664
rect 382832 343612 382884 343664
rect 553032 343000 553084 343052
rect 556712 343000 556764 343052
rect 552020 342796 552072 342848
rect 553676 342796 553728 342848
rect 398012 342252 398064 342304
rect 407120 342252 407172 342304
rect 370780 339464 370832 339516
rect 407120 339464 407172 339516
rect 391664 338104 391716 338156
rect 407120 338104 407172 338156
rect 553124 338104 553176 338156
rect 569224 338104 569276 338156
rect 25412 336744 25464 336796
rect 46480 336744 46532 336796
rect 372252 336676 372304 336728
rect 407120 336676 407172 336728
rect 553032 335316 553084 335368
rect 566464 335316 566516 335368
rect 553124 335248 553176 335300
rect 566188 335248 566240 335300
rect 350356 334024 350408 334076
rect 357072 334024 357124 334076
rect 350356 332596 350408 332648
rect 359280 332596 359332 332648
rect 32680 331168 32732 331220
rect 46480 331168 46532 331220
rect 350356 329808 350408 329860
rect 374092 329808 374144 329860
rect 400772 329808 400824 329860
rect 407120 329808 407172 329860
rect 31024 328448 31076 328500
rect 46480 328448 46532 328500
rect 350356 328448 350408 328500
rect 370872 328448 370924 328500
rect 379244 328448 379296 328500
rect 407120 328448 407172 328500
rect 553032 327156 553084 327208
rect 570512 327156 570564 327208
rect 362500 327088 362552 327140
rect 407120 327088 407172 327140
rect 553124 327088 553176 327140
rect 578792 327088 578844 327140
rect 46296 327020 46348 327072
rect 46940 327020 46992 327072
rect 553032 325728 553084 325780
rect 581368 325728 581420 325780
rect 350356 325660 350408 325712
rect 364708 325660 364760 325712
rect 376576 325660 376628 325712
rect 407120 325660 407172 325712
rect 553124 325660 553176 325712
rect 583576 325660 583628 325712
rect 31208 325592 31260 325644
rect 46480 325592 46532 325644
rect 370688 325592 370740 325644
rect 407212 325592 407264 325644
rect 574928 325592 574980 325644
rect 580172 325592 580224 325644
rect 43352 323484 43404 323536
rect 44640 323484 44692 323536
rect 46296 323144 46348 323196
rect 46848 323144 46900 323196
rect 399852 323008 399904 323060
rect 407212 323008 407264 323060
rect 36544 322940 36596 322992
rect 46848 322940 46900 322992
rect 373908 322940 373960 322992
rect 407120 322940 407172 322992
rect 44916 322872 44968 322924
rect 45744 322872 45796 322924
rect 358636 322872 358688 322924
rect 407212 322872 407264 322924
rect 364708 322804 364760 322856
rect 407120 322804 407172 322856
rect 552020 322328 552072 322380
rect 553676 322328 553728 322380
rect 43352 321580 43404 321632
rect 46848 321580 46900 321632
rect 350356 321580 350408 321632
rect 373172 321580 373224 321632
rect 42248 321512 42300 321564
rect 46480 321512 46532 321564
rect 32404 320152 32456 320204
rect 46848 320152 46900 320204
rect 350356 320152 350408 320204
rect 379336 320152 379388 320204
rect 405096 320152 405148 320204
rect 407304 320152 407356 320204
rect 350264 320084 350316 320136
rect 383292 320084 383344 320136
rect 42248 318928 42300 318980
rect 46848 318928 46900 318980
rect 350356 318792 350408 318844
rect 382648 318792 382700 318844
rect 552756 317568 552808 317620
rect 559380 317568 559432 317620
rect 553124 317500 553176 317552
rect 566188 317500 566240 317552
rect 350356 317432 350408 317484
rect 370688 317432 370740 317484
rect 553032 317432 553084 317484
rect 579988 317432 580040 317484
rect 553124 316004 553176 316056
rect 576308 316004 576360 316056
rect 350356 315936 350408 315988
rect 390100 315936 390152 315988
rect 25504 314644 25556 314696
rect 46296 314644 46348 314696
rect 406200 314644 406252 314696
rect 407120 314644 407172 314696
rect 553124 314644 553176 314696
rect 571800 314644 571852 314696
rect 553032 313284 553084 313336
rect 583116 313284 583168 313336
rect 553124 313216 553176 313268
rect 566096 313216 566148 313268
rect 350356 311856 350408 311908
rect 390284 311856 390336 311908
rect 403808 310564 403860 310616
rect 407120 310564 407172 310616
rect 553124 310564 553176 310616
rect 572076 310564 572128 310616
rect 28540 310496 28592 310548
rect 46112 310496 46164 310548
rect 392492 310496 392544 310548
rect 407212 310496 407264 310548
rect 553032 310496 553084 310548
rect 573456 310496 573508 310548
rect 36636 310428 36688 310480
rect 46296 310428 46348 310480
rect 350172 310428 350224 310480
rect 350540 310428 350592 310480
rect 394148 310428 394200 310480
rect 407120 310428 407172 310480
rect 33692 309136 33744 309188
rect 46112 309136 46164 309188
rect 553124 309136 553176 309188
rect 577412 309136 577464 309188
rect 375196 307844 375248 307896
rect 407120 307844 407172 307896
rect 350356 307776 350408 307828
rect 390100 307776 390152 307828
rect 553124 307776 553176 307828
rect 575020 307776 575072 307828
rect 364064 307708 364116 307760
rect 407120 307708 407172 307760
rect 407580 307436 407632 307488
rect 407948 307436 408000 307488
rect 552020 307436 552072 307488
rect 553952 307436 554004 307488
rect 396540 307028 396592 307080
rect 409236 307028 409288 307080
rect 552204 305464 552256 305516
rect 555516 305464 555568 305516
rect 3516 304988 3568 305040
rect 26700 304988 26752 305040
rect 396816 304988 396868 305040
rect 407120 304988 407172 305040
rect 553124 304988 553176 305040
rect 583208 304988 583260 305040
rect 391572 304240 391624 304292
rect 407580 304240 407632 304292
rect 350448 303696 350500 303748
rect 369768 303696 369820 303748
rect 365352 303628 365404 303680
rect 407120 303628 407172 303680
rect 350172 302268 350224 302320
rect 350908 302268 350960 302320
rect 22560 302200 22612 302252
rect 46388 302200 46440 302252
rect 350448 302200 350500 302252
rect 382096 302200 382148 302252
rect 43720 302132 43772 302184
rect 46296 302132 46348 302184
rect 350448 300908 350500 300960
rect 372252 300908 372304 300960
rect 388352 300908 388404 300960
rect 407120 300908 407172 300960
rect 553032 300908 553084 300960
rect 566556 300908 566608 300960
rect 21272 300840 21324 300892
rect 46388 300840 46440 300892
rect 366732 300840 366784 300892
rect 407212 300840 407264 300892
rect 553124 300840 553176 300892
rect 574468 300840 574520 300892
rect 350448 299548 350500 299600
rect 379428 299548 379480 299600
rect 361212 299480 361264 299532
rect 407120 299480 407172 299532
rect 553124 299480 553176 299532
rect 574928 299480 574980 299532
rect 36636 298528 36688 298580
rect 39396 298528 39448 298580
rect 20260 298120 20312 298172
rect 46388 298120 46440 298172
rect 350448 298120 350500 298172
rect 384120 298120 384172 298172
rect 365260 297372 365312 297424
rect 375288 297372 375340 297424
rect 39396 296692 39448 296744
rect 46388 296692 46440 296744
rect 553124 296692 553176 296744
rect 573364 296692 573416 296744
rect 350448 296624 350500 296676
rect 363052 296624 363104 296676
rect 349252 295740 349304 295792
rect 350816 295740 350868 295792
rect 406108 295400 406160 295452
rect 407856 295400 407908 295452
rect 350448 295332 350500 295384
rect 365260 295332 365312 295384
rect 399760 295332 399812 295384
rect 407120 295332 407172 295384
rect 350356 294040 350408 294092
rect 350816 294040 350868 294092
rect 43260 293972 43312 294024
rect 44180 293972 44232 294024
rect 350448 293972 350500 294024
rect 363052 293972 363104 294024
rect 35256 293904 35308 293956
rect 46112 293904 46164 293956
rect 552020 293088 552072 293140
rect 553768 293088 553820 293140
rect 3516 292544 3568 292596
rect 17500 292544 17552 292596
rect 32496 292544 32548 292596
rect 46388 292544 46440 292596
rect 364064 292544 364116 292596
rect 407212 292544 407264 292596
rect 371976 292476 372028 292528
rect 407120 292476 407172 292528
rect 402704 292408 402756 292460
rect 407212 292408 407264 292460
rect 552020 291728 552072 291780
rect 554044 291728 554096 291780
rect 43720 291184 43772 291236
rect 46388 291184 46440 291236
rect 553124 291184 553176 291236
rect 583300 291184 583352 291236
rect 373632 290436 373684 290488
rect 403532 290436 403584 290488
rect 553124 289824 553176 289876
rect 566096 289824 566148 289876
rect 402152 288464 402204 288516
rect 407120 288464 407172 288516
rect 553032 288464 553084 288516
rect 564992 288464 565044 288516
rect 350448 288396 350500 288448
rect 403532 288396 403584 288448
rect 404912 288396 404964 288448
rect 407304 288396 407356 288448
rect 553124 288396 553176 288448
rect 578516 288396 578568 288448
rect 401140 288328 401192 288380
rect 402704 288328 402756 288380
rect 350448 287104 350500 287156
rect 357164 287104 357216 287156
rect 401140 287104 401192 287156
rect 407120 287104 407172 287156
rect 380808 287036 380860 287088
rect 407212 287036 407264 287088
rect 553124 287036 553176 287088
rect 570328 287036 570380 287088
rect 390192 285744 390244 285796
rect 407120 285744 407172 285796
rect 28172 285676 28224 285728
rect 46388 285676 46440 285728
rect 350448 285676 350500 285728
rect 401048 285676 401100 285728
rect 350356 285608 350408 285660
rect 400772 285608 400824 285660
rect 393044 284928 393096 284980
rect 394148 284928 394200 284980
rect 43628 284656 43680 284708
rect 45652 284656 45704 284708
rect 384212 284316 384264 284368
rect 407120 284316 407172 284368
rect 365444 284248 365496 284300
rect 407212 284248 407264 284300
rect 553124 283568 553176 283620
rect 566188 283568 566240 283620
rect 393044 282888 393096 282940
rect 407120 282888 407172 282940
rect 566188 282888 566240 282940
rect 566648 282888 566700 282940
rect 553124 282820 553176 282872
rect 566004 282820 566056 282872
rect 348516 281936 348568 281988
rect 350172 281936 350224 281988
rect 39212 281664 39264 281716
rect 44824 281664 44876 281716
rect 32588 281596 32640 281648
rect 46848 281596 46900 281648
rect 24032 281528 24084 281580
rect 45652 281528 45704 281580
rect 387524 281460 387576 281512
rect 387800 281460 387852 281512
rect 553124 280236 553176 280288
rect 566832 280236 566884 280288
rect 553032 280168 553084 280220
rect 571892 280168 571944 280220
rect 553124 280100 553176 280152
rect 566280 280100 566332 280152
rect 349068 279012 349120 279064
rect 350816 279012 350868 279064
rect 400772 278808 400824 278860
rect 407120 278808 407172 278860
rect 553124 278808 553176 278860
rect 557080 278808 557132 278860
rect 388168 278740 388220 278792
rect 407212 278740 407264 278792
rect 25320 277380 25372 277432
rect 46848 277380 46900 277432
rect 350448 277380 350500 277432
rect 381452 277380 381504 277432
rect 553124 277380 553176 277432
rect 567384 277380 567436 277432
rect 380532 277312 380584 277364
rect 407120 277312 407172 277364
rect 408408 276768 408460 276820
rect 409144 276768 409196 276820
rect 553032 276088 553084 276140
rect 556804 276088 556856 276140
rect 46480 276020 46532 276072
rect 47584 276020 47636 276072
rect 350448 275952 350500 276004
rect 388536 275952 388588 276004
rect 384672 275884 384724 275936
rect 407120 275884 407172 275936
rect 46480 274660 46532 274712
rect 47308 274660 47360 274712
rect 351368 274660 351420 274712
rect 354128 274660 354180 274712
rect 376668 274660 376720 274712
rect 379520 274660 379572 274712
rect 553124 274660 553176 274712
rect 565084 274660 565136 274712
rect 350448 273300 350500 273352
rect 364708 273300 364760 273352
rect 32680 273232 32732 273284
rect 46848 273232 46900 273284
rect 350356 273232 350408 273284
rect 393780 273232 393832 273284
rect 553124 273232 553176 273284
rect 576032 273232 576084 273284
rect 575020 273164 575072 273216
rect 580172 273164 580224 273216
rect 46480 272552 46532 272604
rect 46848 272552 46900 272604
rect 407488 272552 407540 272604
rect 407764 272552 407816 272604
rect 405372 271804 405424 271856
rect 407120 271804 407172 271856
rect 553124 270512 553176 270564
rect 578608 270512 578660 270564
rect 350448 270444 350500 270496
rect 378968 270444 379020 270496
rect 36820 269764 36872 269816
rect 45560 269764 45612 269816
rect 358636 269084 358688 269136
rect 407120 269084 407172 269136
rect 350448 269016 350500 269068
rect 378140 269016 378192 269068
rect 33968 268336 34020 268388
rect 47124 268336 47176 268388
rect 36820 267792 36872 267844
rect 46388 267792 46440 267844
rect 30932 267724 30984 267776
rect 46480 267724 46532 267776
rect 401968 267724 402020 267776
rect 407120 267724 407172 267776
rect 45468 266364 45520 266416
rect 46940 266364 46992 266416
rect 350448 266364 350500 266416
rect 378968 266364 379020 266416
rect 405372 266364 405424 266416
rect 407764 266364 407816 266416
rect 553124 266364 553176 266416
rect 574652 266364 574704 266416
rect 552020 265208 552072 265260
rect 554228 265208 554280 265260
rect 350448 263644 350500 263696
rect 371424 263644 371476 263696
rect 360384 263576 360436 263628
rect 407120 263576 407172 263628
rect 553124 263576 553176 263628
rect 564440 263576 564492 263628
rect 552020 263168 552072 263220
rect 554780 263168 554832 263220
rect 394148 262896 394200 262948
rect 395160 262896 395212 262948
rect 389088 262624 389140 262676
rect 392400 262624 392452 262676
rect 364156 262216 364208 262268
rect 407120 262216 407172 262268
rect 349068 262148 349120 262200
rect 349988 262148 350040 262200
rect 350448 262148 350500 262200
rect 360384 262148 360436 262200
rect 394148 261536 394200 261588
rect 395712 261536 395764 261588
rect 351828 261400 351880 261452
rect 355140 261400 355192 261452
rect 404820 261128 404872 261180
rect 407488 261128 407540 261180
rect 407580 261128 407632 261180
rect 407580 260924 407632 260976
rect 380532 260856 380584 260908
rect 407120 260856 407172 260908
rect 552020 260856 552072 260908
rect 568580 260856 568632 260908
rect 552848 260380 552900 260432
rect 553032 260380 553084 260432
rect 552112 259496 552164 259548
rect 569040 259496 569092 259548
rect 395712 259428 395764 259480
rect 407120 259428 407172 259480
rect 552020 259428 552072 259480
rect 583392 259428 583444 259480
rect 552112 258136 552164 258188
rect 560300 258136 560352 258188
rect 44456 258068 44508 258120
rect 46020 258068 46072 258120
rect 350448 258068 350500 258120
rect 386972 258068 387024 258120
rect 552020 258068 552072 258120
rect 568948 258068 569000 258120
rect 37188 257320 37240 257372
rect 45652 257320 45704 257372
rect 402520 257320 402572 257372
rect 406568 257320 406620 257372
rect 46848 257184 46900 257236
rect 47400 257184 47452 257236
rect 399392 256776 399444 256828
rect 407120 256776 407172 256828
rect 45468 256708 45520 256760
rect 46020 256708 46072 256760
rect 371976 256708 372028 256760
rect 407212 256708 407264 256760
rect 552020 256708 552072 256760
rect 565820 256708 565872 256760
rect 35072 255960 35124 256012
rect 36636 255960 36688 256012
rect 375012 255960 375064 256012
rect 384672 255960 384724 256012
rect 387340 255960 387392 256012
rect 391112 255960 391164 256012
rect 402060 255960 402112 256012
rect 407488 255960 407540 256012
rect 349896 255416 349948 255468
rect 350540 255416 350592 255468
rect 350356 255348 350408 255400
rect 391020 255348 391072 255400
rect 350448 255280 350500 255332
rect 397920 255280 397972 255332
rect 3148 255212 3200 255264
rect 26884 255212 26936 255264
rect 405188 255212 405240 255264
rect 407488 255212 407540 255264
rect 406752 253988 406804 254040
rect 407304 253988 407356 254040
rect 552112 253988 552164 254040
rect 566188 253988 566240 254040
rect 36636 253920 36688 253972
rect 46848 253920 46900 253972
rect 350448 253920 350500 253972
rect 355692 253920 355744 253972
rect 387340 253920 387392 253972
rect 407120 253920 407172 253972
rect 552020 253920 552072 253972
rect 573180 253920 573232 253972
rect 36452 253648 36504 253700
rect 43168 253648 43220 253700
rect 43628 253648 43680 253700
rect 44824 253648 44876 253700
rect 354128 253444 354180 253496
rect 355048 253444 355100 253496
rect 402152 253172 402204 253224
rect 409236 253172 409288 253224
rect 553124 252560 553176 252612
rect 570788 252560 570840 252612
rect 552664 252492 552716 252544
rect 553952 252492 554004 252544
rect 361304 251812 361356 251864
rect 378692 251812 378744 251864
rect 402520 251200 402572 251252
rect 407120 251200 407172 251252
rect 553124 251200 553176 251252
rect 561680 251200 561732 251252
rect 402888 251132 402940 251184
rect 407212 251132 407264 251184
rect 361304 249840 361356 249892
rect 407120 249840 407172 249892
rect 552664 249840 552716 249892
rect 553400 249840 553452 249892
rect 350448 249772 350500 249824
rect 400680 249772 400732 249824
rect 552020 249772 552072 249824
rect 553400 249704 553452 249756
rect 405556 248752 405608 248804
rect 407764 248752 407816 248804
rect 350448 248412 350500 248464
rect 402152 248412 402204 248464
rect 349528 248140 349580 248192
rect 351460 248140 351512 248192
rect 37188 247664 37240 247716
rect 45560 247664 45612 247716
rect 552940 247664 552992 247716
rect 567200 247664 567252 247716
rect 36452 247052 36504 247104
rect 46848 247052 46900 247104
rect 351460 247052 351512 247104
rect 353852 247052 353904 247104
rect 404268 247052 404320 247104
rect 404820 247052 404872 247104
rect 405004 247052 405056 247104
rect 406292 247052 406344 247104
rect 553124 247052 553176 247104
rect 561680 247052 561732 247104
rect 405004 245828 405056 245880
rect 406384 245828 406436 245880
rect 405188 245760 405240 245812
rect 406476 245760 406528 245812
rect 406752 245760 406804 245812
rect 407580 245760 407632 245812
rect 395252 245692 395304 245744
rect 407120 245692 407172 245744
rect 552204 245692 552256 245744
rect 564900 245692 564952 245744
rect 350448 245624 350500 245676
rect 359372 245624 359424 245676
rect 375012 245624 375064 245676
rect 407212 245624 407264 245676
rect 553124 245624 553176 245676
rect 572260 245624 572312 245676
rect 45468 245556 45520 245608
rect 46020 245556 46072 245608
rect 382924 245556 382976 245608
rect 385500 245556 385552 245608
rect 400128 245556 400180 245608
rect 408960 245556 409012 245608
rect 44824 245488 44876 245540
rect 45928 245488 45980 245540
rect 44640 245420 44692 245472
rect 45652 245420 45704 245472
rect 44640 245284 44692 245336
rect 45744 245284 45796 245336
rect 45652 245216 45704 245268
rect 45652 245012 45704 245064
rect 349988 244876 350040 244928
rect 358728 244876 358780 244928
rect 404912 244672 404964 244724
rect 406384 244672 406436 244724
rect 389732 244332 389784 244384
rect 407120 244332 407172 244384
rect 350448 244264 350500 244316
rect 392400 244264 392452 244316
rect 405464 244264 405516 244316
rect 407304 244264 407356 244316
rect 407764 244264 407816 244316
rect 408500 244264 408552 244316
rect 409052 244264 409104 244316
rect 409420 244264 409472 244316
rect 553124 244264 553176 244316
rect 577596 244264 577648 244316
rect 351828 244196 351880 244248
rect 355140 244196 355192 244248
rect 395896 243516 395948 243568
rect 408868 243516 408920 243568
rect 350448 242904 350500 242956
rect 382924 242904 382976 242956
rect 375104 242836 375156 242888
rect 407120 242836 407172 242888
rect 550364 241476 550416 241528
rect 552112 241476 552164 241528
rect 378692 241272 378744 241324
rect 581460 241272 581512 241324
rect 381728 241204 381780 241256
rect 576308 241204 576360 241256
rect 405372 241136 405424 241188
rect 569132 241136 569184 241188
rect 409512 241068 409564 241120
rect 571708 241068 571760 241120
rect 401968 240728 402020 240780
rect 409512 240592 409564 240644
rect 410156 240592 410208 240644
rect 537668 240592 537720 240644
rect 550548 240524 550600 240576
rect 560300 240728 560352 240780
rect 549996 240252 550048 240304
rect 550456 240252 550508 240304
rect 549260 240184 549312 240236
rect 552480 240184 552532 240236
rect 3056 240116 3108 240168
rect 32220 240116 32272 240168
rect 549536 240116 549588 240168
rect 550272 240116 550324 240168
rect 550456 240116 550508 240168
rect 554136 240116 554188 240168
rect 391572 240048 391624 240100
rect 566372 240048 566424 240100
rect 395528 239980 395580 240032
rect 396080 239980 396132 240032
rect 400956 239980 401008 240032
rect 573456 239980 573508 240032
rect 397368 239912 397420 239964
rect 568580 239912 568632 239964
rect 396908 239844 396960 239896
rect 564440 239844 564492 239896
rect 402152 239776 402204 239828
rect 567476 239776 567528 239828
rect 349068 239708 349120 239760
rect 349896 239708 349948 239760
rect 408960 239708 409012 239760
rect 566648 239708 566700 239760
rect 409052 239640 409104 239692
rect 552020 239640 552072 239692
rect 409420 239572 409472 239624
rect 550456 239572 550508 239624
rect 552756 239572 552808 239624
rect 561680 239572 561732 239624
rect 549076 239504 549128 239556
rect 568764 239504 568816 239556
rect 382740 239436 382792 239488
rect 547788 239436 547840 239488
rect 552848 239436 552900 239488
rect 577688 239436 577740 239488
rect 350264 239368 350316 239420
rect 547236 239368 547288 239420
rect 547420 239368 547472 239420
rect 569316 239368 569368 239420
rect 571800 239368 571852 239420
rect 574928 239300 574980 239352
rect 350448 238960 350500 239012
rect 457444 238960 457496 239012
rect 535276 238960 535328 239012
rect 551376 238960 551428 239012
rect 381452 238892 381504 238944
rect 463148 238892 463200 238944
rect 506664 238892 506716 238944
rect 555332 238892 555384 238944
rect 350356 238824 350408 238876
rect 355232 238824 355284 238876
rect 405556 238824 405608 238876
rect 504364 238824 504416 238876
rect 505652 238824 505704 238876
rect 570696 238824 570748 238876
rect 350448 238756 350500 238808
rect 386880 238756 386932 238808
rect 398196 238756 398248 238808
rect 427820 238756 427872 238808
rect 436744 238756 436796 238808
rect 551100 238756 551152 238808
rect 37004 238688 37056 238740
rect 46664 238688 46716 238740
rect 403532 238688 403584 238740
rect 545580 238688 545632 238740
rect 547788 238688 547840 238740
rect 564808 238688 564860 238740
rect 390008 238620 390060 238672
rect 528836 238620 528888 238672
rect 532056 238620 532108 238672
rect 558184 238620 558236 238672
rect 399668 238552 399720 238604
rect 440240 238552 440292 238604
rect 447048 238552 447100 238604
rect 570512 238552 570564 238604
rect 395436 238484 395488 238536
rect 416688 238484 416740 238536
rect 497924 238484 497976 238536
rect 556896 238484 556948 238536
rect 398748 238416 398800 238468
rect 432236 238416 432288 238468
rect 445116 238416 445168 238468
rect 554228 238416 554280 238468
rect 392768 238348 392820 238400
rect 454132 238348 454184 238400
rect 457352 238348 457404 238400
rect 551284 238348 551336 238400
rect 409328 238280 409380 238332
rect 442540 238280 442592 238332
rect 470600 238280 470652 238332
rect 556436 238280 556488 238332
rect 401048 238212 401100 238264
rect 428372 238212 428424 238264
rect 472624 238212 472676 238264
rect 550824 238212 550876 238264
rect 403624 238144 403676 238196
rect 422576 238144 422628 238196
rect 423588 238144 423640 238196
rect 476396 238144 476448 238196
rect 554780 238144 554832 238196
rect 421288 238076 421340 238128
rect 543924 238076 543976 238128
rect 37004 238008 37056 238060
rect 45744 238008 45796 238060
rect 414848 238008 414900 238060
rect 541164 238008 541216 238060
rect 549168 238008 549220 238060
rect 583668 238008 583720 238060
rect 416688 237940 416740 237992
rect 490564 237940 490616 237992
rect 491116 237940 491168 237992
rect 501788 237940 501840 237992
rect 547604 237940 547656 237992
rect 423588 237872 423640 237924
rect 482928 237872 482980 237924
rect 528192 237872 528244 237924
rect 560392 237872 560444 237924
rect 391388 237804 391440 237856
rect 515312 237804 515364 237856
rect 544200 237736 544252 237788
rect 560300 237736 560352 237788
rect 529848 237600 529900 237652
rect 547696 237600 547748 237652
rect 541900 237464 541952 237516
rect 549628 237464 549680 237516
rect 413560 237396 413612 237448
rect 414020 237396 414072 237448
rect 482928 237396 482980 237448
rect 483756 237396 483808 237448
rect 547144 237396 547196 237448
rect 547880 237396 547932 237448
rect 560944 237396 560996 237448
rect 561772 237396 561824 237448
rect 350448 237328 350500 237380
rect 370780 237328 370832 237380
rect 391112 237328 391164 237380
rect 583484 237328 583536 237380
rect 385592 237260 385644 237312
rect 573088 237260 573140 237312
rect 394516 237192 394568 237244
rect 580448 237192 580500 237244
rect 395160 237124 395212 237176
rect 578700 237124 578752 237176
rect 384672 237056 384724 237108
rect 567200 237056 567252 237108
rect 389088 236988 389140 237040
rect 569224 236988 569276 237040
rect 405464 236920 405516 236972
rect 582932 236920 582984 236972
rect 402060 236852 402112 236904
rect 574560 236852 574612 236904
rect 398380 236784 398432 236836
rect 552204 236784 552256 236836
rect 560300 236784 560352 236836
rect 560944 236784 560996 236836
rect 395804 236716 395856 236768
rect 532700 236716 532752 236768
rect 547512 236716 547564 236768
rect 567292 236716 567344 236768
rect 417424 236648 417476 236700
rect 550640 236648 550692 236700
rect 404636 236580 404688 236632
rect 514760 236580 514812 236632
rect 478604 236512 478656 236564
rect 550916 236512 550968 236564
rect 499212 236444 499264 236496
rect 555424 236444 555476 236496
rect 42708 235968 42760 236020
rect 43260 235968 43312 236020
rect 396540 235900 396592 235952
rect 580356 235900 580408 235952
rect 404268 235832 404320 235884
rect 549996 235832 550048 235884
rect 474648 235764 474700 235816
rect 541624 235764 541676 235816
rect 481548 235696 481600 235748
rect 570512 235696 570564 235748
rect 393780 235628 393832 235680
rect 527548 235628 527600 235680
rect 528744 235628 528796 235680
rect 568764 235628 568816 235680
rect 370688 235560 370740 235612
rect 511448 235560 511500 235612
rect 524328 235560 524380 235612
rect 564992 235560 565044 235612
rect 430304 235492 430356 235544
rect 573272 235492 573324 235544
rect 395988 235424 396040 235476
rect 565176 235424 565228 235476
rect 385040 235356 385092 235408
rect 556528 235356 556580 235408
rect 376944 235288 376996 235340
rect 555240 235288 555292 235340
rect 378140 235220 378192 235272
rect 559564 235220 559616 235272
rect 493416 235152 493468 235204
rect 558000 235152 558052 235204
rect 488632 235084 488684 235136
rect 551284 235084 551336 235136
rect 491208 235016 491260 235068
rect 552112 235016 552164 235068
rect 44088 234812 44140 234864
rect 45928 234812 45980 234864
rect 30840 234608 30892 234660
rect 46664 234608 46716 234660
rect 350448 234608 350500 234660
rect 360384 234608 360436 234660
rect 453488 234540 453540 234592
rect 571616 234540 571668 234592
rect 436744 234472 436796 234524
rect 559288 234472 559340 234524
rect 456708 234404 456760 234456
rect 580448 234404 580500 234456
rect 401140 234336 401192 234388
rect 541716 234336 541768 234388
rect 400772 234268 400824 234320
rect 545212 234268 545264 234320
rect 393872 234200 393924 234252
rect 544844 234200 544896 234252
rect 394240 234132 394292 234184
rect 544384 234132 544436 234184
rect 388168 234064 388220 234116
rect 552480 234064 552532 234116
rect 43904 233996 43956 234048
rect 45928 233996 45980 234048
rect 398012 233996 398064 234048
rect 578700 233996 578752 234048
rect 349988 233928 350040 233980
rect 541440 233928 541492 233980
rect 543832 233928 543884 233980
rect 544292 233928 544344 233980
rect 355600 233860 355652 233912
rect 554044 233860 554096 233912
rect 409972 233792 410024 233844
rect 410340 233792 410392 233844
rect 418804 233792 418856 233844
rect 420000 233792 420052 233844
rect 461216 233792 461268 233844
rect 562232 233792 562284 233844
rect 409696 233724 409748 233776
rect 491300 233724 491352 233776
rect 406200 233656 406252 233708
rect 472808 233656 472860 233708
rect 45468 233384 45520 233436
rect 45744 233384 45796 233436
rect 349068 233180 349120 233232
rect 349712 233180 349764 233232
rect 390376 233180 390428 233232
rect 580172 233180 580224 233232
rect 401508 233112 401560 233164
rect 540428 233112 540480 233164
rect 407580 233044 407632 233096
rect 548524 233044 548576 233096
rect 400036 232976 400088 233028
rect 542544 232976 542596 233028
rect 387616 232908 387668 232960
rect 538864 232908 538916 232960
rect 399852 232840 399904 232892
rect 555608 232840 555660 232892
rect 394608 232772 394660 232824
rect 556988 232772 557040 232824
rect 394332 232704 394384 232756
rect 558184 232704 558236 232756
rect 383568 232636 383620 232688
rect 549904 232636 549956 232688
rect 396816 232568 396868 232620
rect 566648 232568 566700 232620
rect 383476 232500 383528 232552
rect 580356 232500 580408 232552
rect 403440 232432 403492 232484
rect 416780 232432 416832 232484
rect 452568 232432 452620 232484
rect 569132 232432 569184 232484
rect 460940 232364 460992 232416
rect 564808 232364 564860 232416
rect 491116 232296 491168 232348
rect 566280 232296 566332 232348
rect 580172 232228 580224 232280
rect 580448 232228 580500 232280
rect 33968 231820 34020 231872
rect 45560 231820 45612 231872
rect 350448 231820 350500 231872
rect 353852 231820 353904 231872
rect 358544 231752 358596 231804
rect 359004 231752 359056 231804
rect 405648 231208 405700 231260
rect 444472 231208 444524 231260
rect 373816 231140 373868 231192
rect 429200 231140 429252 231192
rect 365076 231072 365128 231124
rect 421932 231072 421984 231124
rect 486976 231072 487028 231124
rect 496820 231072 496872 231124
rect 44088 230732 44140 230784
rect 46940 230732 46992 230784
rect 43904 230528 43956 230580
rect 46020 230528 46072 230580
rect 35256 230460 35308 230512
rect 45560 230460 45612 230512
rect 350448 230460 350500 230512
rect 547328 230460 547380 230512
rect 376300 230392 376352 230444
rect 540336 230392 540388 230444
rect 379336 230324 379388 230376
rect 545856 230324 545908 230376
rect 380716 230256 380768 230308
rect 548064 230256 548116 230308
rect 373172 230188 373224 230240
rect 544660 230188 544712 230240
rect 370872 230120 370924 230172
rect 541808 230120 541860 230172
rect 368296 230052 368348 230104
rect 540520 230052 540572 230104
rect 367928 229984 367980 230036
rect 543096 229984 543148 230036
rect 372252 229916 372304 229968
rect 548248 229916 548300 229968
rect 399760 229848 399812 229900
rect 576308 229848 576360 229900
rect 369768 229780 369820 229832
rect 549352 229780 549404 229832
rect 46388 229712 46440 229764
rect 46572 229712 46624 229764
rect 397276 229712 397328 229764
rect 581828 229712 581880 229764
rect 397000 229644 397052 229696
rect 545948 229644 546000 229696
rect 386880 229576 386932 229628
rect 413560 229576 413612 229628
rect 509332 229576 509384 229628
rect 572076 229576 572128 229628
rect 534724 229236 534776 229288
rect 536840 229236 536892 229288
rect 350448 229100 350500 229152
rect 359004 229100 359056 229152
rect 379428 228352 379480 228404
rect 472072 228352 472124 228404
rect 32312 227740 32364 227792
rect 45560 227740 45612 227792
rect 376484 227332 376536 227384
rect 411628 227332 411680 227384
rect 390284 227264 390336 227316
rect 448336 227264 448388 227316
rect 362224 227196 362276 227248
rect 459928 227196 459980 227248
rect 508504 227196 508556 227248
rect 543832 227196 543884 227248
rect 384764 227128 384816 227180
rect 543004 227128 543056 227180
rect 403900 227060 403952 227112
rect 580448 227060 580500 227112
rect 365260 226992 365312 227044
rect 544108 226992 544160 227044
rect 379152 225700 379204 225752
rect 435456 225700 435508 225752
rect 357164 225632 357216 225684
rect 418068 225632 418120 225684
rect 383384 225564 383436 225616
rect 525800 225564 525852 225616
rect 350356 224884 350408 224936
rect 356428 224884 356480 224936
rect 357072 224340 357124 224392
rect 400220 224340 400272 224392
rect 404728 224340 404780 224392
rect 485044 224340 485096 224392
rect 363788 224272 363840 224324
rect 476672 224272 476724 224324
rect 359648 224204 359700 224256
rect 542452 224204 542504 224256
rect 31116 223592 31168 223644
rect 46664 223592 46716 223644
rect 350448 223524 350500 223576
rect 372344 223524 372396 223576
rect 358728 223456 358780 223508
rect 359648 223456 359700 223508
rect 400680 222912 400732 222964
rect 477960 222912 478012 222964
rect 356888 222844 356940 222896
rect 445760 222844 445812 222896
rect 34796 222164 34848 222216
rect 46664 222164 46716 222216
rect 46572 222096 46624 222148
rect 47584 222096 47636 222148
rect 35348 221688 35400 221740
rect 36360 221688 36412 221740
rect 39948 221688 40000 221740
rect 42064 221688 42116 221740
rect 37004 221416 37056 221468
rect 45928 221416 45980 221468
rect 398472 221416 398524 221468
rect 521660 221416 521712 221468
rect 350448 221144 350500 221196
rect 356520 221144 356572 221196
rect 31208 220804 31260 220856
rect 46664 220804 46716 220856
rect 355416 220736 355468 220788
rect 357624 220736 357676 220788
rect 37648 220260 37700 220312
rect 39304 220260 39356 220312
rect 384120 220056 384172 220108
rect 494060 220056 494112 220108
rect 42616 219444 42668 219496
rect 45836 219444 45888 219496
rect 36912 218696 36964 218748
rect 47676 218696 47728 218748
rect 365168 218696 365220 218748
rect 481180 218696 481232 218748
rect 38108 218628 38160 218680
rect 43628 218628 43680 218680
rect 43168 218560 43220 218612
rect 46020 218560 46072 218612
rect 39304 218084 39356 218136
rect 46664 218084 46716 218136
rect 35440 218016 35492 218068
rect 46112 218016 46164 218068
rect 350448 218016 350500 218068
rect 355048 218016 355100 218068
rect 350356 217948 350408 218000
rect 354956 217948 355008 218000
rect 44088 217336 44140 217388
rect 45744 217336 45796 217388
rect 438676 217336 438728 217388
rect 477592 217336 477644 217388
rect 406660 217268 406712 217320
rect 566004 217268 566056 217320
rect 350448 217200 350500 217252
rect 355232 217200 355284 217252
rect 36912 216724 36964 216776
rect 46296 216724 46348 216776
rect 37004 216656 37056 216708
rect 46664 216656 46716 216708
rect 402428 215908 402480 215960
rect 542820 215908 542872 215960
rect 37740 215296 37792 215348
rect 46664 215296 46716 215348
rect 350448 215296 350500 215348
rect 352748 215296 352800 215348
rect 380624 214548 380676 214600
rect 512092 214548 512144 214600
rect 348608 213868 348660 213920
rect 349344 213868 349396 213920
rect 352656 213868 352708 213920
rect 355140 213868 355192 213920
rect 382648 213256 382700 213308
rect 524972 213256 525024 213308
rect 384304 213188 384356 213240
rect 535920 213188 535972 213240
rect 350448 212508 350500 212560
rect 431224 212508 431276 212560
rect 433340 211760 433392 211812
rect 581460 211760 581512 211812
rect 35072 211148 35124 211200
rect 45560 211148 45612 211200
rect 44640 210536 44692 210588
rect 47768 210536 47820 210588
rect 356796 210468 356848 210520
rect 441620 210468 441672 210520
rect 44732 210400 44784 210452
rect 45652 210400 45704 210452
rect 416964 210400 417016 210452
rect 582932 210400 582984 210452
rect 350448 209856 350500 209908
rect 356612 209856 356664 209908
rect 36360 209040 36412 209092
rect 46296 209040 46348 209092
rect 350448 208360 350500 208412
rect 545028 208360 545080 208412
rect 39580 208292 39632 208344
rect 45560 208292 45612 208344
rect 46388 208292 46440 208344
rect 47400 208292 47452 208344
rect 402612 207680 402664 207732
rect 519176 207680 519228 207732
rect 370596 207612 370648 207664
rect 497924 207612 497976 207664
rect 350448 207068 350500 207120
rect 536104 207068 536156 207120
rect 350356 207000 350408 207052
rect 544200 207000 544252 207052
rect 42432 206932 42484 206984
rect 45652 206932 45704 206984
rect 350448 206932 350500 206984
rect 399392 206932 399444 206984
rect 37188 205640 37240 205692
rect 45652 205640 45704 205692
rect 410064 204892 410116 204944
rect 500224 204892 500276 204944
rect 350356 204280 350408 204332
rect 384304 204280 384356 204332
rect 350448 204212 350500 204264
rect 418804 204212 418856 204264
rect 409880 203600 409932 203652
rect 503720 203600 503772 203652
rect 350080 203532 350132 203584
rect 537760 203532 537812 203584
rect 35716 202852 35768 202904
rect 46664 202852 46716 202904
rect 350448 202852 350500 202904
rect 414664 202852 414716 202904
rect 32956 202784 33008 202836
rect 46388 202784 46440 202836
rect 411352 202104 411404 202156
rect 476028 202104 476080 202156
rect 350448 201492 350500 201544
rect 378692 201492 378744 201544
rect 378692 200812 378744 200864
rect 386512 200812 386564 200864
rect 349896 200744 349948 200796
rect 361764 200744 361816 200796
rect 363328 200744 363380 200796
rect 507860 200744 507912 200796
rect 347780 200200 347832 200252
rect 347780 200064 347832 200116
rect 346216 199860 346268 199912
rect 353576 199860 353628 199912
rect 45008 199656 45060 199708
rect 67088 199656 67140 199708
rect 47492 199588 47544 199640
rect 75920 199588 75972 199640
rect 42616 199520 42668 199572
rect 75460 199520 75512 199572
rect 347596 199520 347648 199572
rect 380808 199520 380860 199572
rect 43904 199452 43956 199504
rect 108948 199452 109000 199504
rect 347504 199452 347556 199504
rect 349344 199452 349396 199504
rect 17408 199384 17460 199436
rect 326988 199384 327040 199436
rect 342996 199384 343048 199436
rect 361028 199384 361080 199436
rect 174268 199316 174320 199368
rect 175096 199316 175148 199368
rect 317236 199316 317288 199368
rect 348516 199316 348568 199368
rect 39672 199248 39724 199300
rect 104624 199248 104676 199300
rect 328184 199248 328236 199300
rect 361672 199248 361724 199300
rect 35532 199180 35584 199232
rect 118792 199180 118844 199232
rect 187792 199180 187844 199232
rect 257988 199180 258040 199232
rect 271512 199180 271564 199232
rect 358452 199180 358504 199232
rect 27252 199112 27304 199164
rect 160100 199112 160152 199164
rect 208400 199112 208452 199164
rect 363696 199112 363748 199164
rect 25596 199044 25648 199096
rect 127256 199044 127308 199096
rect 133052 199044 133104 199096
rect 371332 199044 371384 199096
rect 104072 198976 104124 199028
rect 361120 198976 361172 199028
rect 34060 198908 34112 198960
rect 167828 198908 167880 198960
rect 170404 198908 170456 198960
rect 296076 198908 296128 198960
rect 300492 198908 300544 198960
rect 561036 198908 561088 198960
rect 39948 198840 40000 198892
rect 221924 198840 221976 198892
rect 233516 198840 233568 198892
rect 541900 198840 541952 198892
rect 46664 198772 46716 198824
rect 50344 198772 50396 198824
rect 100852 198772 100904 198824
rect 467932 198772 467984 198824
rect 31668 198704 31720 198756
rect 174912 198704 174964 198756
rect 175096 198704 175148 198756
rect 549536 198704 549588 198756
rect 21824 198636 21876 198688
rect 48688 198636 48740 198688
rect 326988 198636 327040 198688
rect 347596 198636 347648 198688
rect 28724 198568 28776 198620
rect 106004 198568 106056 198620
rect 340420 198568 340472 198620
rect 360200 198568 360252 198620
rect 29920 198500 29972 198552
rect 101496 198500 101548 198552
rect 138204 198500 138256 198552
rect 570788 198500 570840 198552
rect 39212 198432 39264 198484
rect 73804 198432 73856 198484
rect 223856 198432 223908 198484
rect 553860 198432 553912 198484
rect 32864 198364 32916 198416
rect 67364 198364 67416 198416
rect 116308 198364 116360 198416
rect 117964 198364 118016 198416
rect 201960 198364 202012 198416
rect 491392 198364 491444 198416
rect 41144 198296 41196 198348
rect 75644 198296 75696 198348
rect 147864 198296 147916 198348
rect 200764 198296 200816 198348
rect 287612 198296 287664 198348
rect 551192 198296 551244 198348
rect 22744 198228 22796 198280
rect 55772 198228 55824 198280
rect 134340 198228 134392 198280
rect 354772 198228 354824 198280
rect 31576 198160 31628 198212
rect 64144 198160 64196 198212
rect 65064 198160 65116 198212
rect 168472 198160 168524 198212
rect 190368 198160 190420 198212
rect 367836 198160 367888 198212
rect 31484 198092 31536 198144
rect 63592 198092 63644 198144
rect 65524 198092 65576 198144
rect 113732 198092 113784 198144
rect 120724 198092 120776 198144
rect 129832 198092 129884 198144
rect 156880 198092 156932 198144
rect 283564 198092 283616 198144
rect 332048 198092 332100 198144
rect 388352 198092 388404 198144
rect 44548 198024 44600 198076
rect 90916 198024 90968 198076
rect 111156 198024 111208 198076
rect 330484 198024 330536 198076
rect 44916 197956 44968 198008
rect 158536 197956 158588 198008
rect 180064 197956 180116 198008
rect 563888 197956 563940 198008
rect 25780 197888 25832 197940
rect 48044 197888 48096 197940
rect 53288 197888 53340 197940
rect 85304 197888 85356 197940
rect 262496 197888 262548 197940
rect 265624 197888 265676 197940
rect 319812 197888 319864 197940
rect 369124 197888 369176 197940
rect 49240 197820 49292 197872
rect 79600 197820 79652 197872
rect 317880 197820 317932 197872
rect 364984 197820 365036 197872
rect 52828 197752 52880 197804
rect 72516 197752 72568 197804
rect 123392 197752 123444 197804
rect 557080 197752 557132 197804
rect 36912 197684 36964 197736
rect 487160 197684 487212 197736
rect 228456 197480 228508 197532
rect 232872 197480 232924 197532
rect 49332 197344 49384 197396
rect 53104 197344 53156 197396
rect 68284 197344 68336 197396
rect 71136 197344 71188 197396
rect 310704 197344 310756 197396
rect 338120 197344 338172 197396
rect 3424 197276 3476 197328
rect 542360 197276 542412 197328
rect 28356 197208 28408 197260
rect 550456 197208 550508 197260
rect 26976 197140 27028 197192
rect 476212 197140 476264 197192
rect 35256 197072 35308 197124
rect 463700 197072 463752 197124
rect 17316 197004 17368 197056
rect 384212 197004 384264 197056
rect 42708 196936 42760 196988
rect 196808 196936 196860 196988
rect 244464 196936 244516 196988
rect 571892 196936 571944 196988
rect 44088 196868 44140 196920
rect 65064 196868 65116 196920
rect 82176 196868 82228 196920
rect 387432 196868 387484 196920
rect 21456 196800 21508 196852
rect 310704 196800 310756 196852
rect 312728 196800 312780 196852
rect 560852 196800 560904 196852
rect 37096 196732 37148 196784
rect 121460 196732 121512 196784
rect 275376 196732 275428 196784
rect 365812 196732 365864 196784
rect 42340 196664 42392 196716
rect 141792 196664 141844 196716
rect 221648 196664 221700 196716
rect 352380 196664 352432 196716
rect 40592 196596 40644 196648
rect 183008 196596 183060 196648
rect 208124 196596 208176 196648
rect 563428 196596 563480 196648
rect 259000 196528 259052 196580
rect 349436 196528 349488 196580
rect 276020 196392 276072 196444
rect 352012 196460 352064 196512
rect 338120 196392 338172 196444
rect 390192 196392 390244 196444
rect 39764 195916 39816 195968
rect 73528 195916 73580 195968
rect 120172 195916 120224 195968
rect 560576 195916 560628 195968
rect 32220 195848 32272 195900
rect 465080 195848 465132 195900
rect 49516 195780 49568 195832
rect 189080 195780 189132 195832
rect 194232 195780 194284 195832
rect 559472 195780 559524 195832
rect 32404 195712 32456 195764
rect 369676 195712 369728 195764
rect 46756 195644 46808 195696
rect 169116 195644 169168 195696
rect 182640 195644 182692 195696
rect 348424 195644 348476 195696
rect 52276 195576 52328 195628
rect 194876 195576 194928 195628
rect 249616 195576 249668 195628
rect 368112 195576 368164 195628
rect 54852 195508 54904 195560
rect 243084 195508 243136 195560
rect 276664 195508 276716 195560
rect 349804 195508 349856 195560
rect 56048 195440 56100 195492
rect 247684 195440 247736 195492
rect 304356 195440 304408 195492
rect 364340 195440 364392 195492
rect 51540 195372 51592 195424
rect 266912 195372 266964 195424
rect 285404 195372 285456 195424
rect 359096 195372 359148 195424
rect 38292 195304 38344 195356
rect 85580 195304 85632 195356
rect 127992 195304 128044 195356
rect 383200 195304 383252 195356
rect 41972 195236 42024 195288
rect 51724 195168 51776 195220
rect 165252 195168 165304 195220
rect 200120 195168 200172 195220
rect 201316 195168 201368 195220
rect 208400 195168 208452 195220
rect 209596 195168 209648 195220
rect 209780 195168 209832 195220
rect 210976 195168 211028 195220
rect 556620 195236 556672 195288
rect 237380 195168 237432 195220
rect 238576 195168 238628 195220
rect 238760 195168 238812 195220
rect 239956 195168 240008 195220
rect 259460 195168 259512 195220
rect 260564 195168 260616 195220
rect 315304 195168 315356 195220
rect 353484 195168 353536 195220
rect 49424 195100 49476 195152
rect 128452 195100 128504 195152
rect 150532 195100 150584 195152
rect 151728 195100 151780 195152
rect 160192 195100 160244 195152
rect 161388 195100 161440 195152
rect 214104 195100 214156 195152
rect 222292 195100 222344 195152
rect 305000 195100 305052 195152
rect 305552 195100 305604 195152
rect 328460 195100 328512 195152
rect 329380 195100 329432 195152
rect 333980 195100 334032 195152
rect 335268 195100 335320 195152
rect 36268 195032 36320 195084
rect 69020 195032 69072 195084
rect 73344 195032 73396 195084
rect 74448 195032 74500 195084
rect 80060 195032 80112 195084
rect 80796 195032 80848 195084
rect 85580 195032 85632 195084
rect 86408 195032 86460 195084
rect 111800 195032 111852 195084
rect 113088 195032 113140 195084
rect 40224 194828 40276 194880
rect 45928 194828 45980 194880
rect 127072 194556 127124 194608
rect 127992 194556 128044 194608
rect 20168 194488 20220 194540
rect 573364 194488 573416 194540
rect 29552 194420 29604 194472
rect 567568 194420 567620 194472
rect 33692 194352 33744 194404
rect 519084 194352 519136 194404
rect 41236 194284 41288 194336
rect 89260 194284 89312 194336
rect 205180 194284 205232 194336
rect 574284 194284 574336 194336
rect 22652 194216 22704 194268
rect 330760 194216 330812 194268
rect 342720 194216 342772 194268
rect 354036 194216 354088 194268
rect 51264 194148 51316 194200
rect 54576 194148 54628 194200
rect 116952 194148 117004 194200
rect 399576 194148 399628 194200
rect 181352 194080 181404 194132
rect 449900 194080 449952 194132
rect 102140 194012 102192 194064
rect 366640 194012 366692 194064
rect 281172 193944 281224 193996
rect 356152 193944 356204 193996
rect 241244 193876 241296 193928
rect 362408 193876 362460 193928
rect 50436 193808 50488 193860
rect 356520 193808 356572 193860
rect 169760 193740 169812 193792
rect 352656 193740 352708 193792
rect 21732 193672 21784 193724
rect 246396 193672 246448 193724
rect 248420 193672 248472 193724
rect 358636 193672 358688 193724
rect 17224 193604 17276 193656
rect 281724 193604 281776 193656
rect 295708 193604 295760 193656
rect 350540 193604 350592 193656
rect 25320 193128 25372 193180
rect 570420 193128 570472 193180
rect 571984 193128 572036 193180
rect 580264 193128 580316 193180
rect 24032 193060 24084 193112
rect 566464 193060 566516 193112
rect 26700 192992 26752 193044
rect 478880 192992 478932 193044
rect 142068 192924 142120 192976
rect 529940 192924 529992 192976
rect 30012 192856 30064 192908
rect 337844 192856 337896 192908
rect 34060 192788 34112 192840
rect 230940 192788 230992 192840
rect 278596 192788 278648 192840
rect 351460 192788 351512 192840
rect 44640 192720 44692 192772
rect 263784 192720 263836 192772
rect 280528 192720 280580 192772
rect 353392 192720 353444 192772
rect 48044 192652 48096 192704
rect 333336 192652 333388 192704
rect 36912 192584 36964 192636
rect 326896 192584 326948 192636
rect 339500 192584 339552 192636
rect 352564 192584 352616 192636
rect 52184 192516 52236 192568
rect 360384 192516 360436 192568
rect 4804 192448 4856 192500
rect 506480 192448 506532 192500
rect 31576 192380 31628 192432
rect 216128 192380 216180 192432
rect 37096 192312 37148 192364
rect 172980 192312 173032 192364
rect 192024 192312 192076 192364
rect 359188 192312 359240 192364
rect 46296 192244 46348 192296
rect 151820 192244 151872 192296
rect 204536 192244 204588 192296
rect 354680 192244 354732 192296
rect 17500 191768 17552 191820
rect 575940 191768 575992 191820
rect 56324 191700 56376 191752
rect 180708 191700 180760 191752
rect 183928 191700 183980 191752
rect 582656 191700 582708 191752
rect 146300 191632 146352 191684
rect 356336 191632 356388 191684
rect 116676 191564 116728 191616
rect 348240 191564 348292 191616
rect 297916 191496 297968 191548
rect 358544 191496 358596 191548
rect 46848 191428 46900 191480
rect 355692 191428 355744 191480
rect 50804 191360 50856 191412
rect 361856 191360 361908 191412
rect 48228 191292 48280 191344
rect 384488 191292 384540 191344
rect 3424 191224 3476 191276
rect 365352 191224 365404 191276
rect 121460 191156 121512 191208
rect 569316 191156 569368 191208
rect 35900 191088 35952 191140
rect 555516 191088 555568 191140
rect 209412 191020 209464 191072
rect 354864 191020 354916 191072
rect 58624 190952 58676 191004
rect 314016 190952 314068 191004
rect 19984 190408 20036 190460
rect 395712 190408 395764 190460
rect 173624 190340 173676 190392
rect 359648 190340 359700 190392
rect 58716 190272 58768 190324
rect 236736 190272 236788 190324
rect 242900 190272 242952 190324
rect 367100 190272 367152 190324
rect 59636 190204 59688 190256
rect 256056 190204 256108 190256
rect 287704 190204 287756 190256
rect 480352 190204 480404 190256
rect 59912 190136 59964 190188
rect 294696 190136 294748 190188
rect 322112 190136 322164 190188
rect 558092 190136 558144 190188
rect 59176 190068 59228 190120
rect 349160 190068 349212 190120
rect 58532 190000 58584 190052
rect 355232 190000 355284 190052
rect 59820 189932 59872 189984
rect 369952 189932 370004 189984
rect 35532 189864 35584 189916
rect 370228 189864 370280 189916
rect 59544 189796 59596 189848
rect 396080 189796 396132 189848
rect 31668 189728 31720 189780
rect 373448 189728 373500 189780
rect 184572 189660 184624 189712
rect 354128 189660 354180 189712
rect 198096 189592 198148 189644
rect 302148 189592 302200 189644
rect 249984 189524 250036 189576
rect 352288 189524 352340 189576
rect 21272 188980 21324 189032
rect 581736 188980 581788 189032
rect 3516 188912 3568 188964
rect 392676 188912 392728 188964
rect 195152 188844 195204 188896
rect 201500 188844 201552 188896
rect 272524 188844 272576 188896
rect 351092 188844 351144 188896
rect 226156 188776 226208 188828
rect 324412 188776 324464 188828
rect 43168 188708 43220 188760
rect 303712 188708 303764 188760
rect 255780 188640 255832 188692
rect 555148 188640 555200 188692
rect 43260 188572 43312 188624
rect 363144 188572 363196 188624
rect 41880 188504 41932 188556
rect 363052 188504 363104 188556
rect 50620 188436 50672 188488
rect 374000 188436 374052 188488
rect 34152 188368 34204 188420
rect 371884 188368 371936 188420
rect 48964 188300 49016 188352
rect 426532 188300 426584 188352
rect 384304 188164 384356 188216
rect 389088 188164 389140 188216
rect 249340 187620 249392 187672
rect 378232 187620 378284 187672
rect 187516 187552 187568 187604
rect 353760 187552 353812 187604
rect 59084 187484 59136 187536
rect 359280 187484 359332 187536
rect 58992 187416 59044 187468
rect 362040 187416 362092 187468
rect 56416 187348 56468 187400
rect 361948 187348 362000 187400
rect 40592 187280 40644 187332
rect 376668 187280 376720 187332
rect 42432 187212 42484 187264
rect 387340 187212 387392 187264
rect 44916 187144 44968 187196
rect 409972 187144 410024 187196
rect 53656 187076 53708 187128
rect 470600 187076 470652 187128
rect 116032 187008 116084 187060
rect 552388 187008 552440 187060
rect 85764 186940 85816 186992
rect 550088 186940 550140 186992
rect 239036 186872 239088 186924
rect 352472 186872 352524 186924
rect 264152 186804 264204 186856
rect 350816 186804 350868 186856
rect 351092 186804 351144 186856
rect 392860 186804 392912 186856
rect 300860 186736 300912 186788
rect 348148 186736 348200 186788
rect 266084 185988 266136 186040
rect 348056 185988 348108 186040
rect 246120 185920 246172 185972
rect 353668 185920 353720 185972
rect 43720 185852 43772 185904
rect 154304 185852 154356 185904
rect 209872 185852 209924 185904
rect 356244 185852 356296 185904
rect 52092 185784 52144 185836
rect 356612 185784 356664 185836
rect 43536 185716 43588 185768
rect 260840 185716 260892 185768
rect 268660 185716 268712 185768
rect 580080 185716 580132 185768
rect 48872 185648 48924 185700
rect 384580 185648 384632 185700
rect 46020 185580 46072 185632
rect 581184 185580 581236 185632
rect 176660 184628 176712 184680
rect 293960 184628 294012 184680
rect 318248 184628 318300 184680
rect 328828 184628 328880 184680
rect 271880 184560 271932 184612
rect 393044 184560 393096 184612
rect 33784 184492 33836 184544
rect 135260 184492 135312 184544
rect 137284 184492 137336 184544
rect 360292 184492 360344 184544
rect 58808 184424 58860 184476
rect 349620 184424 349672 184476
rect 59452 184356 59504 184408
rect 362960 184356 363012 184408
rect 59728 184288 59780 184340
rect 370136 184288 370188 184340
rect 38108 184220 38160 184272
rect 364524 184220 364576 184272
rect 38200 184152 38252 184204
rect 367284 184152 367336 184204
rect 443000 184152 443052 184204
rect 508228 184152 508280 184204
rect 108304 183540 108356 183592
rect 382280 183540 382332 183592
rect 199752 183132 199804 183184
rect 372068 183132 372120 183184
rect 40408 183064 40460 183116
rect 220360 183064 220412 183116
rect 293132 183064 293184 183116
rect 351276 183064 351328 183116
rect 46572 182996 46624 183048
rect 369584 182996 369636 183048
rect 43536 182928 43588 182980
rect 384856 182928 384908 182980
rect 80244 182860 80296 182912
rect 550732 182860 550784 182912
rect 44824 182792 44876 182844
rect 519820 182792 519872 182844
rect 284760 181976 284812 182028
rect 364432 181976 364484 182028
rect 170772 181908 170824 181960
rect 355508 181908 355560 181960
rect 33048 181840 33100 181892
rect 353852 181840 353904 181892
rect 31392 181772 31444 181824
rect 367192 181772 367244 181824
rect 33784 181704 33836 181756
rect 370044 181704 370096 181756
rect 31484 181636 31536 181688
rect 375012 181636 375064 181688
rect 34428 181568 34480 181620
rect 380532 181568 380584 181620
rect 35256 181500 35308 181552
rect 392952 181500 393004 181552
rect 174636 181432 174688 181484
rect 581644 181432 581696 181484
rect 225512 180480 225564 180532
rect 364064 180480 364116 180532
rect 217784 180412 217836 180464
rect 372620 180412 372672 180464
rect 40500 180344 40552 180396
rect 235172 180344 235224 180396
rect 99932 180276 99984 180328
rect 373540 180276 373592 180328
rect 46112 180208 46164 180260
rect 340880 180208 340932 180260
rect 53380 180140 53432 180192
rect 369216 180140 369268 180192
rect 150532 180072 150584 180124
rect 538956 180072 539008 180124
rect 301044 179324 301096 179376
rect 468300 179324 468352 179376
rect 577504 179324 577556 179376
rect 580080 179324 580132 179376
rect 66444 179256 66496 179308
rect 348332 179256 348384 179308
rect 40868 179188 40920 179240
rect 329196 179188 329248 179240
rect 55588 179120 55640 179172
rect 347044 179120 347096 179172
rect 38660 179052 38712 179104
rect 361212 179052 361264 179104
rect 42340 178984 42392 179036
rect 368020 178984 368072 179036
rect 69664 178916 69716 178968
rect 197360 178916 197412 178968
rect 234528 178916 234580 178968
rect 560484 178916 560536 178968
rect 57612 178848 57664 178900
rect 391480 178848 391532 178900
rect 54760 178780 54812 178832
rect 392492 178780 392544 178832
rect 45008 178712 45060 178764
rect 389916 178712 389968 178764
rect 166264 178644 166316 178696
rect 552572 178644 552624 178696
rect 41052 178440 41104 178492
rect 45560 178440 45612 178492
rect 285680 177828 285732 177880
rect 364156 177828 364208 177880
rect 211988 177760 212040 177812
rect 352104 177760 352156 177812
rect 119896 177692 119948 177744
rect 359004 177692 359056 177744
rect 98644 177624 98696 177676
rect 351000 177624 351052 177676
rect 56140 177556 56192 177608
rect 349252 177556 349304 177608
rect 41144 177488 41196 177540
rect 395252 177488 395304 177540
rect 34336 177420 34388 177472
rect 401968 177420 402020 177472
rect 431224 177420 431276 177472
rect 514024 177420 514076 177472
rect 77392 177352 77444 177404
rect 539968 177352 540020 177404
rect 46204 177284 46256 177336
rect 552296 177284 552348 177336
rect 44824 176604 44876 176656
rect 45836 176604 45888 176656
rect 312452 176468 312504 176520
rect 375380 176468 375432 176520
rect 188160 176400 188212 176452
rect 381912 176400 381964 176452
rect 43444 176332 43496 176384
rect 314384 176332 314436 176384
rect 53564 176264 53616 176316
rect 386236 176264 386288 176316
rect 37188 176196 37240 176248
rect 374828 176196 374880 176248
rect 41972 176128 42024 176180
rect 385868 176128 385920 176180
rect 95240 176060 95292 176112
rect 443184 176060 443236 176112
rect 40960 175992 41012 176044
rect 389732 175992 389784 176044
rect 88340 175924 88392 175976
rect 480536 175924 480588 175976
rect 254492 174904 254544 174956
rect 377680 174904 377732 174956
rect 180800 174836 180852 174888
rect 327080 174836 327132 174888
rect 205640 174768 205692 174820
rect 384396 174768 384448 174820
rect 111984 174700 112036 174752
rect 130200 174700 130252 174752
rect 318892 174700 318944 174752
rect 562324 174700 562376 174752
rect 78036 174632 78088 174684
rect 363972 174632 364024 174684
rect 46296 174564 46348 174616
rect 364616 174564 364668 174616
rect 47952 174496 48004 174548
rect 380900 174496 380952 174548
rect 568028 173816 568080 173868
rect 570420 173816 570472 173868
rect 306472 173476 306524 173528
rect 387064 173476 387116 173528
rect 241612 173408 241664 173460
rect 347872 173408 347924 173460
rect 207480 173340 207532 173392
rect 373264 173340 373316 173392
rect 38016 173272 38068 173324
rect 175924 173272 175976 173324
rect 237380 173272 237432 173324
rect 506940 173272 506992 173324
rect 79324 173204 79376 173256
rect 355048 173204 355100 173256
rect 46480 173136 46532 173188
rect 495440 173136 495492 173188
rect 96712 172320 96764 172372
rect 242256 172320 242308 172372
rect 35164 172252 35216 172304
rect 193220 172252 193272 172304
rect 283472 172252 283524 172304
rect 368480 172252 368532 172304
rect 163044 172184 163096 172236
rect 349712 172184 349764 172236
rect 146944 172116 146996 172168
rect 351184 172116 351236 172168
rect 50528 172048 50580 172100
rect 360476 172048 360528 172100
rect 46664 171980 46716 172032
rect 359372 171980 359424 172032
rect 47768 171912 47820 171964
rect 379612 171912 379664 171964
rect 43904 171844 43956 171896
rect 379244 171844 379296 171896
rect 77392 171776 77444 171828
rect 563520 171776 563572 171828
rect 259644 170756 259696 170808
rect 309140 170756 309192 170808
rect 313740 170756 313792 170808
rect 373908 170756 373960 170808
rect 195244 170688 195296 170740
rect 352748 170688 352800 170740
rect 37924 170620 37976 170672
rect 245476 170620 245528 170672
rect 279608 170620 279660 170672
rect 356428 170620 356480 170672
rect 103796 170552 103848 170604
rect 350724 170552 350776 170604
rect 369400 170552 369452 170604
rect 400772 170552 400824 170604
rect 124404 170484 124456 170536
rect 374092 170484 374144 170536
rect 84200 170416 84252 170468
rect 371424 170416 371476 170468
rect 13820 170348 13872 170400
rect 432052 170348 432104 170400
rect 462320 170348 462372 170400
rect 552756 170348 552808 170400
rect 321468 169260 321520 169312
rect 398104 169260 398156 169312
rect 354312 169192 354364 169244
rect 467840 169192 467892 169244
rect 191840 169124 191892 169176
rect 274456 169124 274508 169176
rect 292580 169124 292632 169176
rect 439320 169124 439372 169176
rect 113180 169056 113232 169108
rect 372436 169056 372488 169108
rect 397920 169056 397972 169108
rect 407304 169056 407356 169108
rect 49700 168988 49752 169040
rect 528836 168988 528888 169040
rect 271972 168104 272024 168156
rect 309876 168104 309928 168156
rect 214012 168036 214064 168088
rect 346584 168036 346636 168088
rect 228732 167968 228784 168020
rect 378876 167968 378928 168020
rect 107752 167900 107804 167952
rect 161756 167900 161808 167952
rect 250628 167900 250680 167952
rect 547420 167900 547472 167952
rect 57520 167832 57572 167884
rect 376576 167832 376628 167884
rect 407120 167832 407172 167884
rect 438860 167832 438912 167884
rect 55956 167764 56008 167816
rect 407856 167764 407908 167816
rect 145012 167696 145064 167748
rect 552848 167696 552900 167748
rect 55036 167628 55088 167680
rect 544476 167628 544528 167680
rect 41236 166540 41288 166592
rect 77300 166540 77352 166592
rect 213276 166540 213328 166592
rect 273260 166540 273312 166592
rect 278964 166540 279016 166592
rect 366732 166540 366784 166592
rect 81900 166472 81952 166524
rect 228364 166472 228416 166524
rect 233884 166472 233936 166524
rect 385684 166472 385736 166524
rect 40776 166404 40828 166456
rect 240140 166404 240192 166456
rect 271236 166404 271288 166456
rect 402336 166404 402388 166456
rect 60832 166336 60884 166388
rect 307944 166336 307996 166388
rect 342076 166336 342128 166388
rect 347964 166336 348016 166388
rect 43352 166268 43404 166320
rect 350448 166268 350500 166320
rect 251272 165180 251324 165232
rect 402244 165180 402296 165232
rect 402704 165180 402756 165232
rect 563428 165180 563480 165232
rect 142436 165112 142488 165164
rect 361304 165112 361356 165164
rect 406568 165112 406620 165164
rect 581644 165112 581696 165164
rect 328460 165044 328512 165096
rect 560852 165044 560904 165096
rect 57428 164976 57480 165028
rect 362316 164976 362368 165028
rect 377772 164976 377824 165028
rect 574928 164976 574980 165028
rect 40684 164908 40736 164960
rect 383936 164908 383988 164960
rect 391664 164908 391716 164960
rect 581736 164908 581788 164960
rect 50160 164840 50212 164892
rect 472164 164840 472216 164892
rect 277400 163752 277452 163804
rect 371976 163752 372028 163804
rect 406292 163752 406344 163804
rect 470232 163752 470284 163804
rect 200764 163684 200816 163736
rect 369124 163684 369176 163736
rect 227720 163616 227772 163668
rect 469220 163616 469272 163668
rect 42156 163548 42208 163600
rect 345020 163548 345072 163600
rect 386972 163548 387024 163600
rect 548340 163548 548392 163600
rect 224868 163480 224920 163532
rect 563796 163480 563848 163532
rect 403348 162800 403400 162852
rect 562324 162800 562376 162852
rect 392584 162732 392636 162784
rect 550916 162732 550968 162784
rect 398564 162664 398616 162716
rect 567292 162664 567344 162716
rect 406844 162596 406896 162648
rect 582656 162596 582708 162648
rect 403716 162528 403768 162580
rect 581184 162528 581236 162580
rect 358360 162460 358412 162512
rect 537852 162460 537904 162512
rect 266360 162392 266412 162444
rect 356244 162392 356296 162444
rect 392400 162392 392452 162444
rect 580080 162392 580132 162444
rect 216496 162324 216548 162376
rect 348700 162324 348752 162376
rect 377956 162324 378008 162376
rect 574560 162324 574612 162376
rect 110880 162256 110932 162308
rect 278780 162256 278832 162308
rect 282920 162256 282972 162308
rect 549260 162256 549312 162308
rect 259552 162188 259604 162240
rect 539048 162188 539100 162240
rect 25412 162120 25464 162172
rect 568580 162120 568632 162172
rect 387524 162052 387576 162104
rect 539232 162052 539284 162104
rect 410156 161984 410208 162036
rect 539324 161984 539376 162036
rect 414664 161916 414716 161968
rect 420000 161916 420052 161968
rect 328460 160964 328512 161016
rect 391296 160964 391348 161016
rect 406384 160964 406436 161016
rect 510160 160964 510212 161016
rect 320180 160896 320232 160948
rect 578792 160896 578844 160948
rect 96712 160828 96764 160880
rect 376024 160828 376076 160880
rect 378968 160828 379020 160880
rect 549536 160828 549588 160880
rect 25964 160760 26016 160812
rect 335636 160760 335688 160812
rect 380348 160760 380400 160812
rect 552572 160760 552624 160812
rect 150440 160692 150492 160744
rect 552388 160692 552440 160744
rect 408316 160012 408368 160064
rect 559564 160012 559616 160064
rect 405188 159944 405240 159996
rect 561036 159944 561088 159996
rect 386052 159876 386104 159928
rect 545672 159876 545724 159928
rect 226800 159808 226852 159860
rect 358176 159808 358228 159860
rect 374736 159808 374788 159860
rect 536840 159808 536892 159860
rect 155316 159740 155368 159792
rect 360936 159740 360988 159792
rect 373724 159740 373776 159792
rect 546776 159740 546828 159792
rect 305092 159672 305144 159724
rect 541072 159672 541124 159724
rect 201408 159604 201460 159656
rect 454132 159604 454184 159656
rect 57336 159536 57388 159588
rect 362500 159536 362552 159588
rect 372160 159536 372212 159588
rect 562048 159536 562100 159588
rect 57704 159468 57756 159520
rect 375196 159468 375248 159520
rect 409236 159468 409288 159520
rect 571708 159468 571760 159520
rect 54944 159400 54996 159452
rect 483112 159400 483164 159452
rect 31024 159332 31076 159384
rect 559472 159332 559524 159384
rect 408224 159264 408276 159316
rect 558276 159264 558328 159316
rect 282828 159196 282880 159248
rect 426440 159196 426492 159248
rect 405096 159128 405148 159180
rect 542912 159128 542964 159180
rect 265624 158448 265676 158500
rect 406476 158448 406528 158500
rect 289268 158380 289320 158432
rect 484400 158380 484452 158432
rect 150164 158312 150216 158364
rect 358912 158312 358964 158364
rect 402520 158312 402572 158364
rect 553860 158312 553912 158364
rect 92480 158244 92532 158296
rect 320824 158244 320876 158296
rect 334072 158244 334124 158296
rect 550088 158244 550140 158296
rect 56232 158176 56284 158228
rect 349528 158176 349580 158228
rect 391756 158176 391808 158228
rect 556436 158176 556488 158228
rect 57244 158108 57296 158160
rect 353944 158108 353996 158160
rect 382096 158108 382148 158160
rect 549812 158108 549864 158160
rect 47860 158040 47912 158092
rect 204260 158040 204312 158092
rect 219716 158040 219768 158092
rect 559196 158040 559248 158092
rect 33876 157972 33928 158024
rect 529940 157972 529992 158024
rect 333980 157292 334032 157344
rect 541348 157292 541400 157344
rect 117964 157224 118016 157276
rect 343364 157224 343416 157276
rect 407948 157224 408000 157276
rect 564624 157224 564676 157276
rect 78772 157156 78824 157208
rect 323400 157156 323452 157208
rect 330484 157156 330536 157208
rect 572168 157156 572220 157208
rect 106372 157088 106424 157140
rect 370504 157088 370556 157140
rect 391020 157088 391072 157140
rect 567660 157088 567712 157140
rect 80152 157020 80204 157072
rect 281540 157020 281592 157072
rect 306380 157020 306432 157072
rect 570696 157020 570748 157072
rect 253940 156952 253992 157004
rect 555516 156952 555568 157004
rect 200120 156884 200172 156936
rect 506296 156884 506348 156936
rect 231952 156816 232004 156868
rect 567476 156816 567528 156868
rect 37832 156748 37884 156800
rect 380716 156748 380768 156800
rect 382004 156748 382056 156800
rect 577504 156748 577556 156800
rect 212540 156680 212592 156732
rect 560484 156680 560536 156732
rect 184940 156612 184992 156664
rect 568856 156612 568908 156664
rect 283564 156544 283616 156596
rect 481824 156544 481876 156596
rect 388720 156476 388772 156528
rect 542636 156476 542688 156528
rect 409788 156408 409840 156460
rect 559196 156408 559248 156460
rect 47676 155864 47728 155916
rect 141148 155864 141200 155916
rect 175280 155864 175332 155916
rect 289820 155864 289872 155916
rect 407764 155864 407816 155916
rect 540060 155864 540112 155916
rect 47860 155796 47912 155848
rect 162860 155796 162912 155848
rect 232596 155796 232648 155848
rect 348608 155796 348660 155848
rect 407396 155796 407448 155848
rect 563060 155796 563112 155848
rect 39212 155728 39264 155780
rect 160192 155728 160244 155780
rect 179420 155728 179472 155780
rect 229376 155728 229428 155780
rect 230020 155728 230072 155780
rect 354220 155728 354272 155780
rect 401416 155728 401468 155780
rect 556528 155728 556580 155780
rect 46388 155660 46440 155712
rect 204904 155660 204956 155712
rect 220820 155660 220872 155712
rect 252652 155660 252704 155712
rect 291200 155660 291252 155712
rect 340144 155660 340196 155712
rect 346400 155660 346452 155712
rect 560760 155660 560812 155712
rect 28632 155592 28684 155644
rect 240968 155592 241020 155644
rect 269120 155592 269172 155644
rect 322756 155592 322808 155644
rect 338120 155592 338172 155644
rect 562416 155592 562468 155644
rect 37740 155524 37792 155576
rect 284116 155524 284168 155576
rect 302240 155524 302292 155576
rect 560576 155524 560628 155576
rect 52000 155456 52052 155508
rect 57980 155456 58032 155508
rect 74816 155456 74868 155508
rect 376392 155456 376444 155508
rect 401232 155456 401284 155508
rect 566464 155456 566516 155508
rect 55772 155388 55824 155440
rect 365996 155388 366048 155440
rect 394424 155388 394476 155440
rect 573456 155388 573508 155440
rect 50988 155320 51040 155372
rect 371240 155320 371292 155372
rect 374920 155320 374972 155372
rect 554044 155320 554096 155372
rect 40868 155252 40920 155304
rect 365904 155252 365956 155304
rect 382188 155252 382240 155304
rect 571892 155252 571944 155304
rect 38016 155184 38068 155236
rect 208400 155184 208452 155236
rect 216680 155184 216732 155236
rect 578240 155184 578292 155236
rect 49148 155116 49200 155168
rect 136640 155116 136692 155168
rect 268016 155116 268068 155168
rect 357624 155116 357676 155168
rect 251916 154776 251968 154828
rect 259460 154776 259512 154828
rect 540612 154776 540664 154828
rect 540612 154572 540664 154624
rect 401324 154504 401376 154556
rect 540520 154504 540572 154556
rect 405280 154436 405332 154488
rect 546316 154436 546368 154488
rect 405004 154368 405056 154420
rect 558000 154368 558052 154420
rect 296352 154300 296404 154352
rect 388812 154300 388864 154352
rect 391204 154300 391256 154352
rect 546592 154300 546644 154352
rect 73436 154232 73488 154284
rect 224224 154232 224276 154284
rect 382832 154232 382884 154284
rect 542728 154232 542780 154284
rect 106280 154164 106332 154216
rect 308588 154164 308640 154216
rect 395620 154164 395672 154216
rect 565084 154164 565136 154216
rect 39580 154096 39632 154148
rect 238760 154096 238812 154148
rect 260288 154096 260340 154148
rect 299480 154096 299532 154148
rect 305000 154096 305052 154148
rect 546868 154096 546920 154148
rect 58900 154028 58952 154080
rect 359556 154028 359608 154080
rect 382924 154028 382976 154080
rect 569224 154028 569276 154080
rect 91100 153960 91152 154012
rect 166908 153960 166960 154012
rect 178040 153960 178092 154012
rect 544936 153960 544988 154012
rect 124220 153892 124272 153944
rect 548892 153892 548944 153944
rect 80060 153824 80112 153876
rect 553032 153824 553084 153876
rect 408132 153756 408184 153808
rect 540796 153756 540848 153808
rect 451280 153688 451332 153740
rect 574284 153688 574336 153740
rect 518900 153620 518952 153672
rect 568028 153620 568080 153672
rect 376944 153280 376996 153332
rect 377220 153280 377272 153332
rect 29644 153144 29696 153196
rect 88984 153144 89036 153196
rect 89812 153144 89864 153196
rect 99288 153144 99340 153196
rect 347872 153144 347924 153196
rect 24124 153076 24176 153128
rect 107660 153076 107712 153128
rect 112168 153076 112220 153128
rect 120724 153076 120776 153128
rect 135996 153076 136048 153128
rect 166264 153076 166316 153128
rect 327264 153076 327316 153128
rect 354864 153076 354916 153128
rect 354956 153076 355008 153128
rect 358084 153076 358136 153128
rect 374644 153144 374696 153196
rect 383292 153144 383344 153196
rect 396724 153144 396776 153196
rect 434168 153144 434220 153196
rect 500224 153144 500276 153196
rect 507584 153144 507636 153196
rect 507676 153144 507728 153196
rect 559656 153144 559708 153196
rect 376760 153076 376812 153128
rect 380256 153076 380308 153128
rect 425152 153076 425204 153128
rect 491300 153076 491352 153128
rect 492128 153076 492180 153128
rect 498200 153076 498252 153128
rect 572720 153076 572772 153128
rect 58256 153008 58308 153060
rect 154580 153008 154632 153060
rect 160100 153008 160152 153060
rect 188804 153008 188856 153060
rect 325056 153008 325108 153060
rect 358820 153008 358872 153060
rect 394056 153008 394108 153060
rect 448980 153008 449032 153060
rect 482928 153008 482980 153060
rect 558092 153008 558144 153060
rect 30932 152940 30984 152992
rect 93492 152940 93544 152992
rect 94780 152940 94832 152992
rect 201408 152940 201460 152992
rect 316592 152940 316644 152992
rect 356060 152940 356112 152992
rect 395344 152940 395396 152992
rect 529204 152940 529256 152992
rect 531412 152940 531464 152992
rect 534724 152940 534776 152992
rect 537576 152940 537628 152992
rect 575940 152940 575992 152992
rect 55128 152872 55180 152924
rect 198740 152872 198792 152924
rect 200396 152872 200448 152924
rect 354772 152872 354824 152924
rect 354864 152872 354916 152924
rect 361580 152872 361632 152924
rect 408040 152872 408092 152924
rect 555148 152872 555200 152924
rect 26792 152804 26844 152856
rect 125048 152804 125100 152856
rect 127624 152804 127676 152856
rect 289268 152804 289320 152856
rect 334992 152804 335044 152856
rect 378784 152804 378836 152856
rect 407028 152804 407080 152856
rect 554136 152804 554188 152856
rect 32496 152736 32548 152788
rect 202972 152736 203024 152788
rect 310520 152736 310572 152788
rect 357440 152736 357492 152788
rect 381544 152736 381596 152788
rect 391664 152736 391716 152788
rect 406936 152736 406988 152788
rect 563888 152736 563940 152788
rect 37924 152668 37976 152720
rect 209780 152668 209832 152720
rect 315028 152668 315080 152720
rect 393964 152668 394016 152720
rect 409604 152668 409656 152720
rect 566556 152668 566608 152720
rect 32312 152600 32364 152652
rect 208768 152600 208820 152652
rect 287980 152600 288032 152652
rect 377864 152600 377916 152652
rect 381636 152600 381688 152652
rect 545120 152600 545172 152652
rect 36636 152532 36688 152584
rect 297640 152532 297692 152584
rect 309232 152532 309284 152584
rect 357532 152532 357584 152584
rect 376116 152532 376168 152584
rect 542268 152532 542320 152584
rect 547328 152532 547380 152584
rect 555332 152532 555384 152584
rect 36452 152464 36504 152516
rect 326620 152464 326672 152516
rect 344008 152464 344060 152516
rect 351920 152464 351972 152516
rect 354772 152464 354824 152516
rect 360844 152464 360896 152516
rect 50344 152396 50396 152448
rect 82544 152396 82596 152448
rect 341800 152396 341852 152448
rect 54576 152328 54628 152380
rect 65800 152328 65852 152380
rect 68744 152328 68796 152380
rect 69664 152328 69716 152380
rect 61292 152260 61344 152312
rect 68284 152260 68336 152312
rect 355324 152328 355376 152380
rect 403256 152464 403308 152516
rect 403808 152464 403860 152516
rect 580264 152464 580316 152516
rect 367744 152396 367796 152448
rect 385776 152396 385828 152448
rect 414848 152396 414900 152448
rect 457444 152396 457496 152448
rect 499856 152396 499908 152448
rect 503076 152396 503128 152448
rect 400864 152328 400916 152380
rect 410340 152328 410392 152380
rect 499580 152328 499632 152380
rect 507676 152328 507728 152380
rect 529204 152396 529256 152448
rect 534632 152396 534684 152448
rect 537484 152396 537536 152448
rect 537852 152396 537904 152448
rect 540336 152396 540388 152448
rect 536840 152328 536892 152380
rect 541992 152328 542044 152380
rect 409144 152260 409196 152312
rect 419356 152260 419408 152312
rect 505652 152260 505704 152312
rect 508504 152260 508556 152312
rect 199108 151784 199160 151836
rect 360200 151784 360252 151836
rect 49056 151716 49108 151768
rect 76012 151716 76064 151768
rect 398656 151716 398708 151768
rect 563520 151716 563572 151768
rect 54208 151648 54260 151700
rect 96620 151648 96672 151700
rect 324320 151648 324372 151700
rect 543188 151648 543240 151700
rect 57888 151580 57940 151632
rect 58900 151580 58952 151632
rect 60004 151580 60056 151632
rect 226340 151580 226392 151632
rect 252560 151580 252612 151632
rect 548432 151580 548484 151632
rect 30840 151512 30892 151564
rect 360108 151512 360160 151564
rect 390100 151512 390152 151564
rect 567752 151512 567804 151564
rect 53472 151444 53524 151496
rect 113364 151444 113416 151496
rect 222200 151444 222252 151496
rect 551744 151444 551796 151496
rect 44732 151376 44784 151428
rect 375472 151376 375524 151428
rect 394240 151376 394292 151428
rect 572812 151376 572864 151428
rect 46388 151308 46440 151360
rect 414020 151308 414072 151360
rect 537668 151308 537720 151360
rect 548156 151308 548208 151360
rect 51816 151240 51868 151292
rect 126980 151240 127032 151292
rect 158720 151240 158772 151292
rect 547052 151240 547104 151292
rect 547880 151240 547932 151292
rect 559288 151240 559340 151292
rect 45928 151172 45980 151224
rect 460940 151172 460992 151224
rect 536104 151172 536156 151224
rect 552296 151172 552348 151224
rect 58164 151104 58216 151156
rect 111800 151104 111852 151156
rect 111892 151104 111944 151156
rect 545304 151104 545356 151156
rect 547236 151104 547288 151156
rect 574836 151104 574888 151156
rect 35072 151036 35124 151088
rect 551376 151036 551428 151088
rect 50712 150968 50764 151020
rect 70492 150968 70544 151020
rect 380440 150968 380492 151020
rect 541900 150968 541952 151020
rect 51908 150900 51960 150952
rect 65524 150900 65576 150952
rect 408960 150900 409012 150952
rect 562232 150900 562284 150952
rect 56508 150832 56560 150884
rect 60004 150832 60056 150884
rect 406752 150832 406804 150884
rect 553124 150832 553176 150884
rect 50068 150764 50120 150816
rect 60740 150764 60792 150816
rect 549076 150628 549128 150680
rect 556620 150628 556672 150680
rect 538864 150424 538916 150476
rect 540980 150424 541032 150476
rect 539048 150356 539100 150408
rect 549628 150356 549680 150408
rect 540612 150288 540664 150340
rect 495440 150220 495492 150272
rect 496636 150220 496688 150272
rect 539324 150084 539376 150136
rect 546500 150084 546552 150136
rect 474648 150016 474700 150068
rect 480076 150016 480128 150068
rect 515036 150016 515088 150068
rect 54576 149948 54628 150000
rect 59544 149948 59596 150000
rect 537944 150016 537996 150068
rect 540428 150016 540480 150068
rect 51448 149880 51500 149932
rect 349712 149880 349764 149932
rect 49608 149812 49660 149864
rect 370964 149880 371016 149932
rect 403164 149880 403216 149932
rect 53012 149744 53064 149796
rect 459560 149880 459612 149932
rect 3516 149676 3568 149728
rect 474648 149880 474700 149932
rect 474740 149880 474792 149932
rect 480076 149880 480128 149932
rect 515036 149880 515088 149932
rect 537760 149948 537812 150000
rect 538864 149880 538916 149932
rect 538956 149880 539008 149932
rect 540152 149880 540204 149932
rect 552848 149948 552900 150000
rect 551100 149880 551152 149932
rect 565360 149812 565412 149864
rect 546132 149744 546184 149796
rect 548524 149744 548576 149796
rect 560300 149744 560352 149796
rect 544384 149676 544436 149728
rect 550088 149676 550140 149728
rect 57152 149064 57204 149116
rect 59636 149064 59688 149116
rect 543648 149064 543700 149116
rect 545212 149064 545264 149116
rect 554136 149064 554188 149116
rect 555424 149064 555476 149116
rect 546040 148996 546092 149048
rect 547880 148996 547932 149048
rect 549904 148384 549956 148436
rect 559012 148384 559064 148436
rect 549996 148316 550048 148368
rect 567568 148316 567620 148368
rect 541716 147636 541768 147688
rect 543740 147636 543792 147688
rect 543556 147568 543608 147620
rect 561864 147568 561916 147620
rect 541532 147500 541584 147552
rect 543924 147500 543976 147552
rect 50252 147296 50304 147348
rect 55772 147296 55824 147348
rect 542912 147296 542964 147348
rect 54668 146956 54720 147008
rect 58624 146956 58676 147008
rect 59084 146956 59136 147008
rect 59544 146956 59596 147008
rect 542544 146956 542596 147008
rect 542820 146956 542872 147008
rect 542912 146956 542964 147008
rect 540704 146888 540756 146940
rect 549812 146820 549864 146872
rect 549904 146820 549956 146872
rect 550824 146820 550876 146872
rect 541256 146616 541308 146668
rect 544660 146616 544712 146668
rect 52920 146208 52972 146260
rect 56508 146208 56560 146260
rect 59820 146276 59872 146328
rect 541808 146276 541860 146328
rect 543556 146276 543608 146328
rect 540704 146208 540756 146260
rect 540980 146208 541032 146260
rect 542176 146208 542228 146260
rect 544108 146208 544160 146260
rect 545948 146208 546000 146260
rect 550364 146208 550416 146260
rect 59268 146140 59320 146192
rect 543096 146140 543148 146192
rect 545212 146140 545264 146192
rect 55772 146072 55824 146124
rect 59452 146072 59504 146124
rect 540520 146072 540572 146124
rect 543464 146072 543516 146124
rect 546408 146072 546460 146124
rect 547972 146072 548024 146124
rect 546040 145596 546092 145648
rect 549352 145596 549404 145648
rect 541716 145528 541768 145580
rect 545764 145528 545816 145580
rect 545856 145460 545908 145512
rect 549352 145460 549404 145512
rect 540152 144848 540204 144900
rect 543280 144848 543332 144900
rect 543648 144848 543700 144900
rect 544752 144848 544804 144900
rect 541624 144780 541676 144832
rect 544384 144780 544436 144832
rect 543188 144712 543240 144764
rect 544292 144712 544344 144764
rect 540520 144168 540572 144220
rect 541164 144168 541216 144220
rect 544476 144100 544528 144152
rect 549444 144100 549496 144152
rect 542084 143896 542136 143948
rect 544016 143896 544068 143948
rect 543004 143556 543056 143608
rect 543740 143556 543792 143608
rect 547972 143556 548024 143608
rect 549260 143556 549312 143608
rect 55864 143488 55916 143540
rect 56968 143488 57020 143540
rect 540888 143488 540940 143540
rect 542820 143488 542872 143540
rect 543188 143488 543240 143540
rect 563336 143488 563388 143540
rect 540796 143420 540848 143472
rect 543924 143420 543976 143472
rect 540612 143352 540664 143404
rect 542820 143352 542872 143404
rect 541992 143284 542044 143336
rect 545488 143284 545540 143336
rect 543096 143148 543148 143200
rect 545028 143148 545080 143200
rect 50804 142808 50856 142860
rect 58624 142808 58676 142860
rect 49700 142196 49752 142248
rect 57152 142196 57204 142248
rect 541164 142128 541216 142180
rect 544200 142128 544252 142180
rect 55036 142060 55088 142112
rect 57888 142060 57940 142112
rect 543648 142060 543700 142112
rect 583576 142060 583628 142112
rect 550180 141992 550232 142044
rect 554228 141992 554280 142044
rect 543188 141652 543240 141704
rect 546592 141652 546644 141704
rect 53840 141380 53892 141432
rect 58716 141380 58768 141432
rect 542176 141108 542228 141160
rect 543280 141108 543332 141160
rect 56508 140836 56560 140888
rect 59544 140836 59596 140888
rect 541532 140836 541584 140888
rect 543832 140836 543884 140888
rect 57060 140768 57112 140820
rect 59728 140768 59780 140820
rect 542268 140768 542320 140820
rect 543556 140768 543608 140820
rect 563704 140768 563756 140820
rect 565176 140768 565228 140820
rect 31300 140700 31352 140752
rect 57888 140700 57940 140752
rect 40316 140632 40368 140684
rect 57152 140632 57204 140684
rect 545120 140020 545172 140072
rect 548064 140020 548116 140072
rect 540796 139544 540848 139596
rect 541716 139544 541768 139596
rect 540612 139476 540664 139528
rect 540888 139476 540940 139528
rect 541256 139476 541308 139528
rect 545396 139476 545448 139528
rect 563796 139476 563848 139528
rect 565176 139476 565228 139528
rect 565268 139476 565320 139528
rect 566648 139476 566700 139528
rect 541164 139408 541216 139460
rect 541808 139408 541860 139460
rect 565360 139408 565412 139460
rect 565820 139408 565872 139460
rect 543556 139340 543608 139392
rect 559472 139340 559524 139392
rect 567936 139340 567988 139392
rect 580448 139340 580500 139392
rect 555608 138660 555660 138712
rect 563796 138660 563848 138712
rect 542176 137980 542228 138032
rect 545212 137980 545264 138032
rect 21548 137912 21600 137964
rect 57888 137912 57940 137964
rect 3148 137844 3200 137896
rect 32404 137844 32456 137896
rect 558184 137708 558236 137760
rect 559472 137708 559524 137760
rect 544752 137504 544804 137556
rect 545948 137504 546000 137556
rect 541992 137368 542044 137420
rect 544752 137368 544804 137420
rect 540428 137300 540480 137352
rect 540980 137300 541032 137352
rect 542820 137300 542872 137352
rect 544660 137300 544712 137352
rect 558368 137300 558420 137352
rect 559012 137300 559064 137352
rect 540244 137232 540296 137284
rect 549812 137232 549864 137284
rect 51448 136552 51500 136604
rect 53196 136552 53248 136604
rect 55128 136552 55180 136604
rect 55864 136552 55916 136604
rect 543556 136552 543608 136604
rect 572720 136552 572772 136604
rect 55772 136484 55824 136536
rect 59636 136484 59688 136536
rect 543648 136484 543700 136536
rect 564716 136484 564768 136536
rect 50988 136144 51040 136196
rect 53012 136144 53064 136196
rect 54116 135872 54168 135924
rect 59452 135872 59504 135924
rect 549444 135872 549496 135924
rect 558184 135872 558236 135924
rect 543648 135396 543700 135448
rect 546500 135396 546552 135448
rect 52368 135328 52420 135380
rect 52920 135328 52972 135380
rect 545028 135260 545080 135312
rect 549444 135260 549496 135312
rect 24676 135192 24728 135244
rect 57888 135192 57940 135244
rect 543556 135192 543608 135244
rect 568580 135192 568632 135244
rect 546040 135124 546092 135176
rect 549260 135124 549312 135176
rect 58900 134716 58952 134768
rect 59084 134716 59136 134768
rect 25872 133832 25924 133884
rect 57888 133832 57940 133884
rect 545120 133900 545172 133952
rect 542268 133832 542320 133884
rect 542544 133832 542596 133884
rect 543280 133832 543332 133884
rect 545580 133832 545632 133884
rect 554228 133832 554280 133884
rect 556988 133832 557040 133884
rect 542268 133696 542320 133748
rect 546408 133152 546460 133204
rect 548524 133152 548576 133204
rect 545948 133084 546000 133136
rect 552020 133084 552072 133136
rect 546408 133016 546460 133068
rect 547972 133016 548024 133068
rect 545856 132744 545908 132796
rect 552112 132744 552164 132796
rect 57060 132676 57112 132728
rect 57888 132676 57940 132728
rect 56508 132472 56560 132524
rect 57152 132472 57204 132524
rect 32588 132404 32640 132456
rect 57060 132404 57112 132456
rect 543556 132404 543608 132456
rect 578792 132404 578844 132456
rect 56508 132336 56560 132388
rect 59268 132336 59320 132388
rect 546132 132336 546184 132388
rect 548984 132336 549036 132388
rect 543648 131452 543700 131504
rect 548064 131452 548116 131504
rect 541716 131248 541768 131300
rect 548248 131248 548300 131300
rect 541992 131180 542044 131232
rect 546960 131180 547012 131232
rect 53380 131112 53432 131164
rect 54576 131112 54628 131164
rect 58532 131112 58584 131164
rect 59636 131112 59688 131164
rect 540980 131112 541032 131164
rect 542176 131112 542228 131164
rect 543740 131112 543792 131164
rect 540796 131044 540848 131096
rect 543556 131044 543608 131096
rect 578240 131044 578292 131096
rect 545948 130976 546000 131028
rect 546592 130976 546644 131028
rect 548616 130976 548668 131028
rect 551284 130976 551336 131028
rect 544752 130908 544804 130960
rect 545028 130908 545080 130960
rect 540704 130840 540756 130892
rect 546960 130840 547012 130892
rect 544660 130772 544712 130824
rect 547236 130772 547288 130824
rect 544476 130024 544528 130076
rect 545396 130024 545448 130076
rect 54576 129684 54628 129736
rect 55864 129684 55916 129736
rect 551468 129684 551520 129736
rect 552112 129684 552164 129736
rect 54852 129616 54904 129668
rect 57060 129616 57112 129668
rect 551284 129616 551336 129668
rect 552020 129616 552072 129668
rect 55128 129548 55180 129600
rect 56968 129548 57020 129600
rect 56416 128324 56468 128376
rect 56876 128324 56928 128376
rect 39488 128256 39540 128308
rect 57244 128256 57296 128308
rect 543556 128256 543608 128308
rect 563060 128256 563112 128308
rect 542084 128188 542136 128240
rect 544016 128188 544068 128240
rect 50988 127780 51040 127832
rect 54392 127780 54444 127832
rect 53748 127576 53800 127628
rect 58532 127576 58584 127628
rect 540980 127576 541032 127628
rect 545028 127576 545080 127628
rect 49608 126896 49660 126948
rect 50344 126896 50396 126948
rect 54760 126896 54812 126948
rect 57244 126896 57296 126948
rect 58992 126896 59044 126948
rect 59360 126896 59412 126948
rect 541900 126896 541952 126948
rect 543188 126896 543240 126948
rect 541624 126828 541676 126880
rect 543464 126828 543516 126880
rect 53748 126216 53800 126268
rect 57152 126216 57204 126268
rect 540336 126216 540388 126268
rect 556896 126216 556948 126268
rect 542268 125672 542320 125724
rect 544568 125672 544620 125724
rect 540796 125604 540848 125656
rect 541992 125604 542044 125656
rect 28908 125536 28960 125588
rect 57244 125536 57296 125588
rect 542084 125536 542136 125588
rect 543740 125604 543792 125656
rect 543556 125536 543608 125588
rect 562324 125536 562376 125588
rect 52368 125468 52420 125520
rect 55036 125468 55088 125520
rect 59268 124448 59320 124500
rect 59820 124448 59872 124500
rect 22836 124108 22888 124160
rect 57244 124108 57296 124160
rect 58900 124108 58952 124160
rect 59452 124108 59504 124160
rect 544384 124108 544436 124160
rect 545396 124108 545448 124160
rect 562324 124108 562376 124160
rect 565268 124108 565320 124160
rect 56508 124040 56560 124092
rect 58716 124040 58768 124092
rect 543372 123360 543424 123412
rect 552480 123360 552532 123412
rect 55128 122884 55180 122936
rect 55312 122816 55364 122868
rect 544108 122816 544160 122868
rect 546408 122816 546460 122868
rect 543556 122748 543608 122800
rect 574928 122748 574980 122800
rect 546500 122680 546552 122732
rect 549076 122680 549128 122732
rect 57152 121660 57204 121712
rect 57888 121660 57940 121712
rect 58992 121592 59044 121644
rect 59360 121592 59412 121644
rect 57336 121524 57388 121576
rect 57888 121524 57940 121576
rect 545120 121456 545172 121508
rect 548524 121456 548576 121508
rect 36176 121388 36228 121440
rect 57336 121388 57388 121440
rect 543556 121388 543608 121440
rect 560852 121388 560904 121440
rect 543188 121252 543240 121304
rect 547880 121252 547932 121304
rect 54576 120708 54628 120760
rect 55220 120708 55272 120760
rect 546040 120368 546092 120420
rect 549260 120368 549312 120420
rect 59176 120164 59228 120216
rect 59820 120164 59872 120216
rect 59268 120096 59320 120148
rect 59452 120096 59504 120148
rect 540888 120096 540940 120148
rect 543096 120096 543148 120148
rect 549996 120096 550048 120148
rect 552112 120096 552164 120148
rect 40592 119960 40644 120012
rect 57336 119960 57388 120012
rect 54760 119348 54812 119400
rect 59636 119348 59688 119400
rect 548524 119348 548576 119400
rect 565820 119348 565872 119400
rect 58716 118668 58768 118720
rect 59544 118668 59596 118720
rect 54116 118600 54168 118652
rect 56600 118600 56652 118652
rect 56508 118124 56560 118176
rect 59728 118124 59780 118176
rect 57152 117988 57204 118040
rect 59728 117988 59780 118040
rect 59176 117920 59228 117972
rect 59360 117920 59412 117972
rect 540704 117512 540756 117564
rect 546960 117512 547012 117564
rect 546132 117308 546184 117360
rect 546592 117308 546644 117360
rect 22928 117240 22980 117292
rect 57336 117240 57388 117292
rect 543556 117240 543608 117292
rect 568028 117240 568080 117292
rect 545028 117172 545080 117224
rect 546592 117172 546644 117224
rect 549076 117172 549128 117224
rect 552112 117172 552164 117224
rect 547788 116628 547840 116680
rect 548800 116628 548852 116680
rect 541808 116560 541860 116612
rect 552204 116560 552256 116612
rect 54852 116424 54904 116476
rect 56876 116424 56928 116476
rect 43168 115880 43220 115932
rect 57336 115880 57388 115932
rect 541808 115880 541860 115932
rect 542820 115880 542872 115932
rect 545764 115880 545816 115932
rect 547236 115880 547288 115932
rect 543556 115812 543608 115864
rect 558276 115880 558328 115932
rect 541992 115472 542044 115524
rect 548800 115472 548852 115524
rect 541440 115404 541492 115456
rect 542360 115404 542412 115456
rect 24308 115200 24360 115252
rect 57152 115200 57204 115252
rect 544384 114996 544436 115048
rect 545488 114996 545540 115048
rect 547788 114860 547840 114912
rect 547972 114860 548024 114912
rect 545120 114588 545172 114640
rect 547880 114588 547932 114640
rect 547328 114520 547380 114572
rect 548064 114520 548116 114572
rect 542084 114452 542136 114504
rect 542360 114452 542412 114504
rect 543556 114452 543608 114504
rect 572168 114452 572220 114504
rect 543648 114384 543700 114436
rect 559564 114384 559616 114436
rect 540520 114316 540572 114368
rect 545488 114316 545540 114368
rect 540612 113976 540664 114028
rect 546132 113976 546184 114028
rect 54668 113772 54720 113824
rect 58716 113772 58768 113824
rect 543004 113500 543056 113552
rect 547880 113500 547932 113552
rect 545120 113160 545172 113212
rect 547972 113160 548024 113212
rect 557080 113160 557132 113212
rect 558276 113160 558328 113212
rect 542268 113092 542320 113144
rect 549904 113092 549956 113144
rect 576216 113092 576268 113144
rect 580448 113092 580500 113144
rect 48872 112888 48924 112940
rect 57336 112888 57388 112940
rect 59636 112072 59688 112124
rect 59820 112072 59872 112124
rect 59268 111936 59320 111988
rect 59820 111936 59872 111988
rect 558184 111868 558236 111920
rect 565820 111868 565872 111920
rect 58900 111800 58952 111852
rect 59544 111800 59596 111852
rect 546408 111800 546460 111852
rect 549996 111800 550048 111852
rect 556988 111052 557040 111104
rect 561680 111052 561732 111104
rect 543096 110576 543148 110628
rect 543832 110576 543884 110628
rect 540888 110508 540940 110560
rect 543372 110508 543424 110560
rect 56508 110440 56560 110492
rect 59636 110440 59688 110492
rect 543004 110440 543056 110492
rect 544016 110440 544068 110492
rect 543556 110372 543608 110424
rect 551376 110372 551428 110424
rect 543188 109692 543240 109744
rect 550732 109692 550784 109744
rect 43260 108944 43312 108996
rect 57428 108944 57480 108996
rect 542268 108944 542320 108996
rect 543096 108944 543148 108996
rect 44640 108876 44692 108928
rect 57520 108876 57572 108928
rect 547880 108876 547932 108928
rect 550088 108876 550140 108928
rect 543648 108808 543700 108860
rect 544200 108808 544252 108860
rect 543740 108400 543792 108452
rect 549628 108400 549680 108452
rect 542176 108332 542228 108384
rect 542820 108332 542872 108384
rect 545028 108332 545080 108384
rect 551284 108332 551336 108384
rect 546224 108264 546276 108316
rect 550640 108264 550692 108316
rect 57888 108196 57940 108248
rect 58808 108196 58860 108248
rect 542176 108196 542228 108248
rect 544476 108196 544528 108248
rect 545948 108060 546000 108112
rect 546592 108060 546644 108112
rect 543188 107856 543240 107908
rect 548984 107856 549036 107908
rect 50252 107584 50304 107636
rect 54668 107584 54720 107636
rect 540796 107584 540848 107636
rect 541164 107584 541216 107636
rect 540796 107448 540848 107500
rect 543832 107652 543884 107704
rect 543280 107584 543332 107636
rect 562416 107584 562468 107636
rect 546040 106224 546092 106276
rect 547420 106224 547472 106276
rect 548708 105884 548760 105936
rect 552112 105884 552164 105936
rect 542360 104864 542412 104916
rect 53288 104796 53340 104848
rect 57428 104796 57480 104848
rect 543832 104796 543884 104848
rect 50436 104728 50488 104780
rect 57520 104728 57572 104780
rect 541532 104728 541584 104780
rect 544016 104728 544068 104780
rect 543464 104184 543516 104236
rect 545028 104184 545080 104236
rect 541900 104116 541952 104168
rect 558368 104184 558420 104236
rect 547236 104116 547288 104168
rect 563796 104116 563848 104168
rect 24492 103436 24544 103488
rect 57520 103436 57572 103488
rect 24400 103368 24452 103420
rect 57428 103368 57480 103420
rect 549904 103096 549956 103148
rect 552480 103096 552532 103148
rect 540888 102280 540940 102332
rect 545028 102280 545080 102332
rect 542176 102212 542228 102264
rect 543648 102212 543700 102264
rect 542268 102144 542320 102196
rect 542820 102144 542872 102196
rect 563796 102144 563848 102196
rect 565820 102144 565872 102196
rect 542176 102076 542228 102128
rect 548800 102076 548852 102128
rect 53748 101940 53800 101992
rect 55404 101940 55456 101992
rect 543096 101804 543148 101856
rect 549628 101804 549680 101856
rect 544476 100716 544528 100768
rect 545580 100716 545632 100768
rect 549996 100716 550048 100768
rect 550732 100716 550784 100768
rect 560208 100716 560260 100768
rect 560852 100716 560904 100768
rect 27344 100648 27396 100700
rect 57520 100648 57572 100700
rect 540980 99968 541032 100020
rect 570144 99968 570196 100020
rect 559564 99356 559616 99408
rect 561680 99356 561732 99408
rect 540704 98812 540756 98864
rect 542360 98812 542412 98864
rect 541440 98676 541492 98728
rect 541992 98676 542044 98728
rect 543556 98608 543608 98660
rect 551284 98608 551336 98660
rect 57980 97996 58032 98048
rect 59728 97996 59780 98048
rect 540520 97996 540572 98048
rect 542176 97996 542228 98048
rect 46112 97928 46164 97980
rect 57520 97928 57572 97980
rect 57888 97928 57940 97980
rect 58808 97928 58860 97980
rect 543556 97928 543608 97980
rect 570052 97928 570104 97980
rect 53196 97860 53248 97912
rect 55864 97860 55916 97912
rect 58532 97860 58584 97912
rect 59728 97860 59780 97912
rect 2872 97724 2924 97776
rect 4804 97724 4856 97776
rect 543096 97248 543148 97300
rect 547328 97248 547380 97300
rect 543556 96568 543608 96620
rect 575572 96568 575624 96620
rect 54760 96092 54812 96144
rect 57428 96092 57480 96144
rect 547420 95276 547472 95328
rect 547880 95276 547932 95328
rect 53288 95208 53340 95260
rect 55312 95208 55364 95260
rect 547328 95208 547380 95260
rect 547972 95208 548024 95260
rect 28172 95140 28224 95192
rect 57520 95140 57572 95192
rect 542268 95140 542320 95192
rect 543372 95140 543424 95192
rect 543556 95140 543608 95192
rect 555516 95140 555568 95192
rect 548800 94188 548852 94240
rect 554136 94188 554188 94240
rect 543280 94052 543332 94104
rect 544568 94052 544620 94104
rect 57520 93916 57572 93968
rect 57888 93916 57940 93968
rect 543556 93916 543608 93968
rect 545120 93916 545172 93968
rect 51632 93780 51684 93832
rect 57888 93780 57940 93832
rect 51632 92488 51684 92540
rect 55404 92488 55456 92540
rect 543556 91196 543608 91248
rect 549720 91196 549772 91248
rect 41236 90992 41288 91044
rect 57888 90992 57940 91044
rect 542268 90856 542320 90908
rect 549720 90856 549772 90908
rect 543464 90516 543516 90568
rect 544108 90516 544160 90568
rect 540888 89768 540940 89820
rect 543740 89768 543792 89820
rect 542636 89700 542688 89752
rect 544200 89700 544252 89752
rect 30104 89632 30156 89684
rect 57888 89632 57940 89684
rect 543556 89632 543608 89684
rect 581736 89632 581788 89684
rect 546132 89564 546184 89616
rect 547880 89564 547932 89616
rect 546408 89496 546460 89548
rect 547972 89496 548024 89548
rect 547420 89428 547472 89480
rect 549628 89428 549680 89480
rect 540612 88272 540664 88324
rect 543832 88272 543884 88324
rect 545028 88272 545080 88324
rect 545948 88272 546000 88324
rect 543464 87592 543516 87644
rect 550640 87592 550692 87644
rect 540520 85756 540572 85808
rect 543464 85756 543516 85808
rect 543832 85756 543884 85808
rect 549260 85756 549312 85808
rect 3516 85484 3568 85536
rect 21364 85484 21416 85536
rect 540796 85484 540848 85536
rect 547328 85484 547380 85536
rect 542360 84600 542412 84652
rect 544936 84600 544988 84652
rect 543556 84124 543608 84176
rect 552572 84124 552624 84176
rect 543740 83920 543792 83972
rect 547880 83920 547932 83972
rect 545028 83852 545080 83904
rect 546500 83852 546552 83904
rect 552940 83444 552992 83496
rect 565176 83444 565228 83496
rect 544568 82968 544620 83020
rect 547972 82968 548024 83020
rect 57060 82900 57112 82952
rect 57612 82900 57664 82952
rect 540520 82900 540572 82952
rect 546132 82900 546184 82952
rect 54760 82832 54812 82884
rect 55220 82832 55272 82884
rect 546040 82832 546092 82884
rect 547420 82832 547472 82884
rect 552848 82832 552900 82884
rect 556620 82832 556672 82884
rect 23388 82764 23440 82816
rect 57612 82764 57664 82816
rect 543556 82764 543608 82816
rect 552388 82764 552440 82816
rect 47584 82696 47636 82748
rect 57888 82696 57940 82748
rect 48964 82084 49016 82136
rect 55956 82084 56008 82136
rect 551376 80044 551428 80096
rect 552480 80044 552532 80096
rect 540152 79296 540204 79348
rect 540428 79296 540480 79348
rect 543648 78616 543700 78668
rect 563980 78616 564032 78668
rect 543556 78548 543608 78600
rect 561036 78548 561088 78600
rect 543556 77188 543608 77240
rect 559656 77188 559708 77240
rect 51724 75828 51776 75880
rect 57612 75828 57664 75880
rect 540612 75828 540664 75880
rect 542452 75828 542504 75880
rect 543556 75216 543608 75268
rect 550272 75216 550324 75268
rect 545948 74536 546000 74588
rect 549812 74536 549864 74588
rect 53288 73652 53340 73704
rect 56968 73652 57020 73704
rect 542176 73176 542228 73228
rect 544108 73176 544160 73228
rect 546040 73176 546092 73228
rect 549904 73176 549956 73228
rect 556896 73176 556948 73228
rect 548248 73108 548300 73160
rect 576124 73108 576176 73160
rect 580264 73108 580316 73160
rect 543556 72428 543608 72480
rect 562508 72428 562560 72480
rect 545120 72224 545172 72276
rect 549996 72224 550048 72276
rect 547328 71680 547380 71732
rect 549812 71680 549864 71732
rect 542820 71000 542872 71052
rect 566740 71000 566792 71052
rect 542084 70592 542136 70644
rect 546500 70592 546552 70644
rect 546500 70456 546552 70508
rect 549260 70456 549312 70508
rect 543556 70320 543608 70372
rect 552296 70320 552348 70372
rect 542636 69844 542688 69896
rect 544108 69844 544160 69896
rect 45100 69640 45152 69692
rect 57060 69640 57112 69692
rect 543740 69640 543792 69692
rect 546960 69640 547012 69692
rect 18972 68960 19024 69012
rect 57612 68960 57664 69012
rect 540888 68960 540940 69012
rect 542636 68960 542688 69012
rect 56968 68076 57020 68128
rect 57612 68076 57664 68128
rect 546040 67600 546092 67652
rect 546500 67600 546552 67652
rect 50528 67124 50580 67176
rect 56692 67124 56744 67176
rect 540612 66648 540664 66700
rect 545120 66648 545172 66700
rect 543556 66172 543608 66224
rect 577320 66172 577372 66224
rect 20444 64812 20496 64864
rect 56968 64812 57020 64864
rect 46204 64744 46256 64796
rect 57888 64744 57940 64796
rect 543556 63996 543608 64048
rect 549536 63996 549588 64048
rect 57796 63656 57848 63708
rect 43536 63452 43588 63504
rect 57704 63452 57756 63504
rect 57796 63452 57848 63504
rect 41788 62024 41840 62076
rect 57704 62024 57756 62076
rect 543556 62024 543608 62076
rect 560760 62024 560812 62076
rect 543648 61956 543700 62008
rect 560576 61956 560628 62008
rect 574744 60664 574796 60716
rect 580264 60664 580316 60716
rect 26056 59304 26108 59356
rect 57704 59304 57756 59356
rect 543556 57876 543608 57928
rect 574100 57876 574152 57928
rect 54944 57264 54996 57316
rect 57704 57264 57756 57316
rect 49240 53728 49292 53780
rect 57704 53728 57756 53780
rect 543556 53728 543608 53780
rect 569224 53728 569276 53780
rect 543464 50804 543516 50856
rect 547052 50804 547104 50856
rect 543556 49648 543608 49700
rect 551192 49648 551244 49700
rect 30196 48220 30248 48272
rect 57704 48220 57756 48272
rect 543556 48220 543608 48272
rect 575480 48220 575532 48272
rect 543556 45500 543608 45552
rect 579896 45500 579948 45552
rect 543648 45432 543700 45484
rect 563152 45432 563204 45484
rect 543556 44072 543608 44124
rect 560484 44072 560536 44124
rect 542360 42304 542412 42356
rect 544200 42304 544252 42356
rect 46296 41352 46348 41404
rect 57704 41352 57756 41404
rect 543556 41352 543608 41404
rect 563888 41352 563940 41404
rect 47032 39992 47084 40044
rect 57704 39992 57756 40044
rect 543556 37204 543608 37256
rect 562048 37204 562100 37256
rect 540888 36728 540940 36780
rect 542544 36728 542596 36780
rect 543556 35844 543608 35896
rect 581644 35844 581696 35896
rect 24584 34416 24636 34468
rect 57704 34416 57756 34468
rect 33692 33056 33744 33108
rect 57704 33056 57756 33108
rect 570604 33056 570656 33108
rect 579804 33056 579856 33108
rect 34060 32988 34112 33040
rect 57796 32988 57848 33040
rect 46572 31696 46624 31748
rect 57704 31696 57756 31748
rect 543556 31696 543608 31748
rect 583300 31696 583352 31748
rect 540888 31084 540940 31136
rect 567752 31084 567804 31136
rect 540704 31016 540756 31068
rect 568856 31016 568908 31068
rect 540612 30268 540664 30320
rect 544476 30268 544528 30320
rect 168380 29860 168432 29912
rect 169500 29860 169552 29912
rect 340880 29860 340932 29912
rect 342092 29860 342144 29912
rect 361580 29860 361632 29912
rect 362700 29860 362752 29912
rect 445852 29860 445904 29912
rect 447064 29860 447116 29912
rect 458180 29860 458232 29912
rect 459300 29860 459352 29912
rect 474740 29860 474792 29912
rect 476044 29860 476096 29912
rect 525800 29860 525852 29912
rect 526920 29860 526972 29912
rect 536840 29656 536892 29708
rect 545856 29656 545908 29708
rect 45284 29588 45336 29640
rect 69020 29588 69072 29640
rect 531412 29588 531464 29640
rect 534816 29588 534868 29640
rect 535460 29588 535512 29640
rect 581828 29588 581880 29640
rect 52828 29520 52880 29572
rect 63224 29520 63276 29572
rect 474648 29520 474700 29572
rect 474832 29520 474884 29572
rect 515956 29520 516008 29572
rect 548156 29520 548208 29572
rect 43076 29452 43128 29504
rect 69664 29452 69716 29504
rect 514024 29452 514076 29504
rect 548340 29452 548392 29504
rect 33968 29384 34020 29436
rect 71596 29384 71648 29436
rect 509516 29384 509568 29436
rect 546776 29384 546828 29436
rect 42524 29316 42576 29368
rect 159824 29316 159876 29368
rect 506940 29316 506992 29368
rect 565912 29316 565964 29368
rect 51816 29248 51868 29300
rect 170772 29248 170824 29300
rect 443184 29248 443236 29300
rect 561956 29248 562008 29300
rect 47216 29180 47268 29232
rect 199752 29180 199804 29232
rect 372988 29180 373040 29232
rect 535460 29180 535512 29232
rect 537852 29180 537904 29232
rect 546316 29180 546368 29232
rect 29736 29112 29788 29164
rect 187516 29112 187568 29164
rect 356888 29112 356940 29164
rect 560944 29112 560996 29164
rect 42248 29044 42300 29096
rect 205548 29044 205600 29096
rect 287336 29044 287388 29096
rect 31116 28976 31168 29028
rect 109592 28976 109644 29028
rect 158536 28976 158588 29028
rect 531228 28976 531280 29028
rect 534816 29044 534868 29096
rect 550916 29044 550968 29096
rect 539508 28976 539560 29028
rect 52092 28908 52144 28960
rect 70952 28908 71004 28960
rect 247408 28908 247460 28960
rect 511264 28908 511316 28960
rect 49424 28840 49476 28892
rect 67732 28840 67784 28892
rect 381360 28840 381412 28892
rect 553952 28840 554004 28892
rect 39856 28772 39908 28824
rect 82544 28772 82596 28824
rect 82820 28772 82872 28824
rect 249984 28772 250036 28824
rect 451556 28772 451608 28824
rect 561128 28772 561180 28824
rect 45468 28704 45520 28756
rect 204904 28704 204956 28756
rect 275744 28704 275796 28756
rect 387064 28704 387116 28756
rect 531228 28704 531280 28756
rect 583392 28704 583444 28756
rect 41696 28636 41748 28688
rect 195244 28636 195296 28688
rect 523040 28636 523092 28688
rect 579712 28636 579764 28688
rect 34796 28568 34848 28620
rect 103796 28568 103848 28620
rect 105636 28568 105688 28620
rect 211344 28568 211396 28620
rect 322112 28568 322164 28620
rect 504180 28568 504232 28620
rect 512092 28568 512144 28620
rect 583208 28568 583260 28620
rect 35440 28500 35492 28552
rect 73528 28500 73580 28552
rect 74632 28500 74684 28552
rect 190736 28500 190788 28552
rect 271236 28500 271288 28552
rect 474004 28500 474056 28552
rect 493416 28500 493468 28552
rect 573180 28500 573232 28552
rect 46756 28432 46808 28484
rect 105084 28432 105136 28484
rect 105544 28432 105596 28484
rect 272524 28432 272576 28484
rect 295708 28432 295760 28484
rect 527824 28432 527876 28484
rect 529480 28432 529532 28484
rect 577412 28432 577464 28484
rect 41328 28364 41380 28416
rect 89628 28364 89680 28416
rect 89720 28364 89772 28416
rect 259000 28364 259052 28416
rect 266084 28364 266136 28416
rect 522304 28364 522356 28416
rect 527180 28364 527232 28416
rect 72516 28296 72568 28348
rect 252560 28296 252612 28348
rect 268016 28296 268068 28348
rect 528560 28296 528612 28348
rect 537208 28364 537260 28416
rect 546868 28364 546920 28416
rect 539508 28296 539560 28348
rect 55588 28228 55640 28280
rect 87696 28228 87748 28280
rect 89076 28228 89128 28280
rect 213276 28228 213328 28280
rect 484400 28228 484452 28280
rect 485044 28228 485096 28280
rect 505652 28228 505704 28280
rect 548892 28228 548944 28280
rect 39120 28160 39172 28212
rect 124404 28160 124456 28212
rect 147680 28160 147732 28212
rect 148876 28160 148928 28212
rect 165620 28160 165672 28212
rect 166264 28160 166316 28212
rect 167000 28160 167052 28212
rect 168196 28160 168248 28212
rect 191840 28160 191892 28212
rect 192668 28160 192720 28212
rect 194692 28160 194744 28212
rect 195888 28160 195940 28212
rect 215300 28160 215352 28212
rect 216496 28160 216548 28212
rect 300860 28160 300912 28212
rect 302148 28160 302200 28212
rect 320180 28160 320232 28212
rect 321468 28160 321520 28212
rect 321560 28160 321612 28212
rect 322756 28160 322808 28212
rect 329840 28160 329892 28212
rect 331128 28160 331180 28212
rect 347780 28160 347832 28212
rect 348516 28160 348568 28212
rect 368480 28160 368532 28212
rect 369768 28160 369820 28212
rect 426440 28160 426492 28212
rect 427728 28160 427780 28212
rect 427820 28160 427872 28212
rect 429016 28160 429068 28212
rect 436100 28160 436152 28212
rect 437388 28160 437440 28212
rect 444380 28160 444432 28212
rect 445116 28160 445168 28212
rect 447140 28160 447192 28212
rect 448336 28160 448388 28212
rect 463700 28160 463752 28212
rect 464436 28160 464488 28212
rect 474832 28160 474884 28212
rect 552664 28160 552716 28212
rect 69756 28092 69808 28144
rect 120540 28092 120592 28144
rect 155960 28092 156012 28144
rect 157248 28092 157300 28144
rect 291200 28092 291252 28144
rect 291844 28092 291896 28144
rect 378140 28092 378192 28144
rect 379428 28092 379480 28144
rect 484492 28092 484544 28144
rect 485688 28092 485740 28144
rect 505100 28092 505152 28144
rect 506296 28092 506348 28144
rect 506388 28092 506440 28144
rect 569960 28092 570012 28144
rect 39396 28024 39448 28076
rect 128912 28024 128964 28076
rect 483112 28024 483164 28076
rect 536840 28024 536892 28076
rect 43996 27956 44048 28008
rect 217784 27956 217836 28008
rect 360108 27956 360160 28008
rect 527180 27956 527232 28008
rect 43812 27888 43864 27940
rect 92204 27888 92256 27940
rect 127624 27888 127676 27940
rect 579988 27888 580040 27940
rect 389088 27820 389140 27872
rect 534724 27820 534776 27872
rect 502340 27752 502392 27804
rect 506388 27752 506440 27804
rect 88984 27616 89036 27668
rect 89628 27616 89680 27668
rect 52184 27548 52236 27600
rect 70308 27548 70360 27600
rect 528192 27548 528244 27600
rect 553032 27548 553084 27600
rect 50896 27480 50948 27532
rect 62580 27480 62632 27532
rect 492772 27480 492824 27532
rect 555332 27480 555384 27532
rect 28816 27412 28868 27464
rect 123760 27412 123812 27464
rect 174636 27412 174688 27464
rect 578332 27412 578384 27464
rect 54484 27344 54536 27396
rect 441252 27344 441304 27396
rect 511448 27344 511500 27396
rect 545304 27344 545356 27396
rect 44456 27276 44508 27328
rect 389732 27276 389784 27328
rect 398748 27276 398800 27328
rect 582840 27276 582892 27328
rect 41880 27208 41932 27260
rect 116676 27208 116728 27260
rect 224224 27208 224276 27260
rect 548616 27208 548668 27260
rect 45192 27140 45244 27192
rect 363972 27140 364024 27192
rect 365904 27140 365956 27192
rect 579896 27140 579948 27192
rect 35624 27072 35676 27124
rect 244188 27072 244240 27124
rect 268660 27072 268712 27124
rect 578608 27072 578660 27124
rect 52000 27004 52052 27056
rect 293132 27004 293184 27056
rect 327264 27004 327316 27056
rect 560668 27004 560720 27056
rect 43628 26936 43680 26988
rect 100576 26936 100628 26988
rect 344008 26936 344060 26988
rect 562140 26936 562192 26988
rect 26884 26868 26936 26920
rect 71780 26868 71832 26920
rect 410340 26868 410392 26920
rect 556804 26868 556856 26920
rect 417424 26800 417476 26852
rect 560392 26800 560444 26852
rect 409696 26732 409748 26784
rect 540888 26732 540940 26784
rect 42064 26664 42116 26716
rect 473452 26664 473504 26716
rect 516600 26664 516652 26716
rect 574836 26664 574888 26716
rect 37648 26596 37700 26648
rect 520464 26596 520516 26648
rect 27436 26188 27488 26240
rect 523040 26188 523092 26240
rect 538220 26188 538272 26240
rect 555700 26188 555752 26240
rect 35716 26120 35768 26172
rect 494060 26120 494112 26172
rect 509240 26120 509292 26172
rect 574560 26120 574612 26172
rect 29828 26052 29880 26104
rect 470876 26052 470928 26104
rect 476212 26052 476264 26104
rect 553124 26052 553176 26104
rect 20260 25984 20312 26036
rect 391940 25984 391992 26036
rect 423680 25984 423732 26036
rect 567660 25984 567712 26036
rect 40868 25916 40920 25968
rect 387800 25916 387852 25968
rect 389272 25916 389324 25968
rect 580080 25916 580132 25968
rect 23112 25848 23164 25900
rect 213920 25848 213972 25900
rect 280160 25848 280212 25900
rect 575848 25848 575900 25900
rect 59728 25780 59780 25832
rect 211252 25780 211304 25832
rect 322940 25780 322992 25832
rect 578516 25780 578568 25832
rect 32128 25712 32180 25764
rect 165712 25712 165764 25764
rect 325792 25712 325844 25764
rect 578424 25712 578476 25764
rect 33600 25644 33652 25696
rect 156052 25644 156104 25696
rect 430580 25644 430632 25696
rect 540704 25644 540756 25696
rect 22560 25576 22612 25628
rect 131212 25576 131264 25628
rect 477500 25576 477552 25628
rect 572996 25576 573048 25628
rect 53564 25508 53616 25560
rect 100760 25508 100812 25560
rect 396080 25508 396132 25560
rect 547696 25508 547748 25560
rect 52276 25440 52328 25492
rect 98000 25440 98052 25492
rect 513380 25440 513432 25492
rect 569040 25440 569092 25492
rect 53656 25372 53708 25424
rect 81440 25372 81492 25424
rect 520280 25372 520332 25424
rect 571524 25372 571576 25424
rect 54300 25304 54352 25356
rect 77300 25304 77352 25356
rect 516140 25304 516192 25356
rect 568120 25304 568172 25356
rect 49056 24760 49108 24812
rect 191932 24760 191984 24812
rect 534724 24760 534776 24812
rect 544016 24760 544068 24812
rect 54208 24692 54260 24744
rect 397460 24692 397512 24744
rect 409880 24692 409932 24744
rect 555424 24692 555476 24744
rect 37004 24624 37056 24676
rect 325700 24624 325752 24676
rect 385132 24624 385184 24676
rect 580356 24624 580408 24676
rect 21916 24556 21968 24608
rect 285680 24556 285732 24608
rect 465172 24556 465224 24608
rect 561772 24556 561824 24608
rect 47676 24488 47728 24540
rect 291292 24488 291344 24540
rect 502524 24488 502576 24540
rect 582656 24488 582708 24540
rect 24216 24420 24268 24472
rect 266360 24420 266412 24472
rect 465264 24420 465316 24472
rect 541072 24420 541124 24472
rect 31208 24352 31260 24404
rect 256700 24352 256752 24404
rect 503720 24352 503772 24404
rect 555240 24352 555292 24404
rect 33784 24284 33836 24336
rect 219440 24284 219492 24336
rect 502432 24284 502484 24336
rect 548432 24284 548484 24336
rect 44824 24216 44876 24268
rect 219532 24216 219584 24268
rect 245660 24216 245712 24268
rect 564900 24216 564952 24268
rect 51908 24148 51960 24200
rect 209780 24148 209832 24200
rect 220820 24148 220872 24200
rect 568672 24148 568724 24200
rect 55496 24080 55548 24132
rect 197360 24080 197412 24132
rect 209872 24080 209924 24132
rect 566188 24080 566240 24132
rect 47768 24012 47820 24064
rect 161480 24012 161532 24064
rect 510620 24012 510672 24064
rect 551652 24012 551704 24064
rect 53472 23944 53524 23996
rect 142160 23944 142212 23996
rect 171140 23944 171192 23996
rect 578240 23944 578292 23996
rect 51540 23876 51592 23928
rect 95332 23876 95384 23928
rect 503720 23468 503772 23520
rect 504364 23468 504416 23520
rect 48044 23400 48096 23452
rect 69756 23400 69808 23452
rect 138020 23400 138072 23452
rect 581092 23400 581144 23452
rect 185032 23332 185084 23384
rect 581368 23332 581420 23384
rect 38476 23264 38528 23316
rect 426532 23264 426584 23316
rect 434812 23264 434864 23316
rect 564624 23264 564676 23316
rect 38568 23196 38620 23248
rect 382280 23196 382332 23248
rect 383660 23196 383712 23248
rect 574652 23196 574704 23248
rect 50068 23128 50120 23180
rect 368480 23128 368532 23180
rect 376760 23128 376812 23180
rect 576952 23128 577004 23180
rect 25688 23060 25740 23112
rect 306380 23060 306432 23112
rect 361580 23060 361632 23112
rect 552940 23060 552992 23112
rect 27160 22992 27212 23044
rect 307760 22992 307812 23044
rect 447140 22992 447192 23044
rect 565084 22992 565136 23044
rect 47308 22924 47360 22976
rect 324320 22924 324372 22976
rect 484492 22924 484544 22976
rect 563612 22924 563664 22976
rect 50712 22856 50764 22908
rect 296720 22856 296772 22908
rect 434720 22856 434772 22908
rect 559104 22856 559156 22908
rect 40960 22788 41012 22840
rect 183560 22788 183612 22840
rect 389180 22788 389232 22840
rect 556344 22788 556396 22840
rect 39672 22720 39724 22772
rect 182180 22720 182232 22772
rect 360200 22720 360252 22772
rect 547604 22720 547656 22772
rect 57244 22652 57296 22704
rect 116032 22652 116084 22704
rect 498200 22652 498252 22704
rect 545672 22652 545724 22704
rect 46848 22584 46900 22636
rect 102140 22584 102192 22636
rect 31392 22516 31444 22568
rect 131120 22516 131172 22568
rect 41052 22448 41104 22500
rect 193220 22448 193272 22500
rect 56048 22040 56100 22092
rect 69572 22040 69624 22092
rect 26148 21972 26200 22024
rect 448612 21972 448664 22024
rect 488540 21972 488592 22024
rect 577504 21972 577556 22024
rect 49148 21904 49200 21956
rect 411260 21904 411312 21956
rect 420920 21904 420972 21956
rect 552204 21904 552256 21956
rect 53104 21836 53156 21888
rect 400220 21836 400272 21888
rect 419540 21836 419592 21888
rect 543924 21836 543976 21888
rect 46480 21768 46532 21820
rect 270500 21768 270552 21820
rect 523040 21768 523092 21820
rect 575664 21768 575716 21820
rect 37924 21700 37976 21752
rect 229100 21700 229152 21752
rect 470600 21700 470652 21752
rect 556160 21700 556212 21752
rect 48872 21632 48924 21684
rect 205640 21632 205692 21684
rect 416780 21632 416832 21684
rect 557816 21632 557868 21684
rect 49516 21564 49568 21616
rect 179420 21564 179472 21616
rect 407120 21564 407172 21616
rect 555792 21564 555844 21616
rect 36912 21496 36964 21548
rect 147680 21496 147732 21548
rect 249800 21496 249852 21548
rect 568948 21496 569000 21548
rect 53380 21428 53432 21480
rect 155960 21428 156012 21480
rect 229100 21428 229152 21480
rect 574376 21428 574428 21480
rect 40224 21360 40276 21412
rect 139400 21360 139452 21412
rect 176660 21360 176712 21412
rect 572904 21360 572956 21412
rect 55864 21292 55916 21344
rect 140780 21292 140832 21344
rect 58716 21224 58768 21276
rect 128452 21224 128504 21276
rect 17776 21156 17828 21208
rect 505100 21156 505152 21208
rect 179420 20816 179472 20868
rect 569960 20816 570012 20868
rect 161480 20748 161532 20800
rect 560300 20748 560352 20800
rect 135260 20680 135312 20732
rect 571432 20680 571484 20732
rect 20352 20612 20404 20664
rect 458180 20612 458232 20664
rect 527180 20612 527232 20664
rect 547236 20612 547288 20664
rect 28540 20544 28592 20596
rect 462320 20544 462372 20596
rect 469220 20544 469272 20596
rect 567476 20544 567528 20596
rect 19064 20476 19116 20528
rect 364432 20476 364484 20528
rect 449900 20476 449952 20528
rect 558092 20476 558144 20528
rect 25504 20408 25556 20460
rect 356060 20408 356112 20460
rect 459560 20408 459612 20460
rect 544292 20408 544344 20460
rect 27528 20340 27580 20392
rect 354680 20340 354732 20392
rect 477592 20340 477644 20392
rect 554044 20340 554096 20392
rect 23020 20272 23072 20324
rect 342260 20272 342312 20324
rect 463700 20272 463752 20324
rect 540060 20272 540112 20324
rect 19156 20204 19208 20256
rect 333980 20204 334032 20256
rect 474740 20204 474792 20256
rect 551100 20204 551152 20256
rect 18880 20136 18932 20188
rect 311900 20136 311952 20188
rect 452660 20136 452712 20188
rect 557724 20136 557776 20188
rect 44732 20068 44784 20120
rect 202880 20068 202932 20120
rect 427912 20068 427964 20120
rect 543188 20068 543240 20120
rect 59820 20000 59872 20052
rect 216772 20000 216824 20052
rect 296720 20000 296772 20052
rect 563704 20000 563756 20052
rect 33048 19932 33100 19984
rect 167000 19932 167052 19984
rect 271880 19932 271932 19984
rect 556712 19932 556764 19984
rect 38108 19864 38160 19916
rect 149060 19864 149112 19916
rect 504180 19864 504232 19916
rect 544660 19864 544712 19916
rect 37096 19796 37148 19848
rect 125600 19796 125652 19848
rect 533344 19796 533396 19848
rect 550088 19796 550140 19848
rect 41144 19728 41196 19780
rect 95240 19728 95292 19780
rect 461032 19728 461084 19780
rect 562232 19728 562284 19780
rect 201592 19320 201644 19372
rect 445852 19320 445904 19372
rect 58992 19252 59044 19304
rect 88984 19252 89036 19304
rect 527824 19252 527876 19304
rect 549812 19252 549864 19304
rect 57428 19184 57480 19236
rect 72516 19184 72568 19236
rect 426440 19184 426492 19236
rect 570696 19184 570748 19236
rect 54668 19116 54720 19168
rect 336740 19116 336792 19168
rect 465080 19116 465132 19168
rect 571984 19116 572036 19168
rect 57520 19048 57572 19100
rect 215300 19048 215352 19100
rect 291200 19048 291252 19100
rect 569132 19048 569184 19100
rect 54760 18980 54812 19032
rect 293960 18980 294012 19032
rect 353300 18980 353352 19032
rect 540336 18980 540388 19032
rect 38200 18912 38252 18964
rect 194692 18912 194744 18964
rect 339592 18912 339644 18964
rect 574192 18912 574244 18964
rect 39212 18844 39264 18896
rect 189080 18844 189132 18896
rect 321560 18844 321612 18896
rect 567384 18844 567436 18896
rect 39764 18776 39816 18828
rect 150440 18776 150492 18828
rect 314752 18776 314804 18828
rect 569408 18776 569460 18828
rect 43720 18708 43772 18760
rect 146300 18708 146352 18760
rect 307760 18708 307812 18760
rect 570328 18708 570380 18760
rect 55128 18640 55180 18692
rect 154580 18640 154632 18692
rect 276112 18640 276164 18692
rect 571524 18640 571576 18692
rect 56508 18572 56560 18624
rect 105636 18572 105688 18624
rect 267740 18572 267792 18624
rect 573548 18572 573600 18624
rect 58900 18504 58952 18556
rect 89076 18504 89128 18556
rect 440332 18504 440384 18556
rect 544108 18504 544160 18556
rect 47952 18436 48004 18488
rect 164332 18436 164384 18488
rect 160100 18368 160152 18420
rect 564992 18368 565044 18420
rect 38016 18300 38068 18352
rect 364340 18300 364392 18352
rect 39304 17892 39356 17944
rect 444380 17892 444432 17944
rect 445760 17892 445812 17944
rect 577228 17892 577280 17944
rect 190552 17824 190604 17876
rect 577596 17824 577648 17876
rect 47860 17756 47912 17808
rect 427820 17756 427872 17808
rect 448520 17756 448572 17808
rect 566556 17756 566608 17808
rect 236000 17688 236052 17740
rect 582748 17688 582800 17740
rect 39580 17620 39632 17672
rect 375380 17620 375432 17672
rect 438860 17620 438912 17672
rect 541808 17620 541860 17672
rect 46664 17552 46716 17604
rect 245752 17552 245804 17604
rect 251272 17552 251324 17604
rect 583024 17552 583076 17604
rect 59636 17484 59688 17536
rect 251180 17484 251232 17536
rect 260932 17484 260984 17536
rect 581276 17484 581328 17536
rect 50344 17416 50396 17468
rect 234620 17416 234672 17468
rect 299480 17416 299532 17468
rect 543280 17416 543332 17468
rect 58808 17348 58860 17400
rect 227720 17348 227772 17400
rect 259460 17348 259512 17400
rect 542176 17348 542228 17400
rect 35532 17280 35584 17332
rect 191840 17280 191892 17332
rect 256700 17280 256752 17332
rect 543372 17280 543424 17332
rect 55956 17212 56008 17264
rect 165620 17212 165672 17264
rect 234620 17212 234672 17264
rect 553768 17212 553820 17264
rect 46388 17144 46440 17196
rect 147680 17144 147732 17196
rect 460940 17144 460992 17196
rect 542912 17144 542964 17196
rect 31484 17076 31536 17128
rect 117320 17076 117372 17128
rect 511264 17076 511316 17128
rect 580172 17076 580224 17128
rect 59268 17008 59320 17060
rect 105544 17008 105596 17060
rect 31576 16940 31628 16992
rect 201500 16940 201552 16992
rect 51632 16872 51684 16924
rect 237380 16872 237432 16924
rect 522304 16532 522356 16584
rect 549720 16532 549772 16584
rect 310612 16464 310664 16516
rect 566280 16464 566332 16516
rect 403072 16396 403124 16448
rect 582472 16396 582524 16448
rect 382372 16328 382424 16380
rect 548524 16328 548576 16380
rect 364616 16260 364668 16312
rect 541164 16260 541216 16312
rect 349160 16192 349212 16244
rect 543004 16192 543056 16244
rect 357532 16124 357584 16176
rect 562324 16124 562376 16176
rect 346952 16056 347004 16108
rect 559472 16056 559524 16108
rect 342904 15988 342956 16040
rect 575756 15988 575808 16040
rect 293224 15920 293276 15972
rect 554964 15920 555016 15972
rect 120632 15852 120684 15904
rect 576032 15852 576084 15904
rect 403624 15784 403676 15836
rect 541900 15784 541952 15836
rect 433340 15716 433392 15768
rect 551744 15716 551796 15768
rect 300860 15648 300912 15700
rect 582380 15648 582432 15700
rect 220912 15104 220964 15156
rect 564716 15104 564768 15156
rect 324412 15036 324464 15088
rect 542084 15036 542136 15088
rect 380900 14968 380952 15020
rect 567568 14968 567620 15020
rect 367744 14900 367796 14952
rect 581000 14900 581052 14952
rect 254216 14832 254268 14884
rect 540520 14832 540572 14884
rect 247592 14764 247644 14816
rect 551376 14764 551428 14816
rect 264980 14696 265032 14748
rect 570512 14696 570564 14748
rect 233424 14628 233476 14680
rect 544568 14628 544620 14680
rect 253480 14560 253532 14612
rect 576860 14560 576912 14612
rect 175464 14492 175516 14544
rect 568764 14492 568816 14544
rect 171968 14424 172020 14476
rect 564808 14424 564860 14476
rect 414296 14356 414348 14408
rect 579252 14356 579304 14408
rect 474004 14288 474056 14340
rect 540244 14288 540296 14340
rect 233240 13744 233292 13796
rect 563796 13744 563848 13796
rect 320180 13676 320232 13728
rect 544844 13676 544896 13728
rect 340880 13608 340932 13660
rect 559564 13608 559616 13660
rect 351920 13540 351972 13592
rect 551284 13540 551336 13592
rect 357440 13472 357492 13524
rect 544384 13472 544436 13524
rect 363052 13404 363104 13456
rect 545948 13404 546000 13456
rect 378140 13336 378192 13388
rect 549444 13336 549496 13388
rect 404360 13268 404412 13320
rect 560852 13268 560904 13320
rect 386420 13200 386472 13252
rect 542452 13200 542504 13252
rect 398932 13132 398984 13184
rect 576308 13132 576360 13184
rect 143540 13064 143592 13116
rect 553400 13064 553452 13116
rect 393320 12996 393372 13048
rect 548708 12996 548760 13048
rect 410800 12928 410852 12980
rect 559748 12928 559800 12980
rect 456892 12860 456944 12912
rect 551008 12860 551060 12912
rect 23204 12384 23256 12436
rect 544200 12384 544252 12436
rect 313280 12316 313332 12368
rect 542636 12316 542688 12368
rect 335452 12248 335504 12300
rect 541992 12248 542044 12300
rect 347780 12180 347832 12232
rect 549352 12180 549404 12232
rect 398840 12112 398892 12164
rect 581184 12112 581236 12164
rect 467472 12044 467524 12096
rect 545396 12044 545448 12096
rect 299480 11976 299532 12028
rect 583668 11976 583720 12028
rect 228272 11908 228324 11960
rect 545488 11908 545540 11960
rect 194416 11840 194468 11892
rect 551560 11840 551612 11892
rect 36820 11772 36872 11824
rect 132960 11772 133012 11824
rect 504364 11772 504416 11824
rect 56784 11704 56836 11756
rect 574468 11704 574520 11756
rect 314660 10956 314712 11008
rect 548248 10956 548300 11008
rect 328460 10888 328512 10940
rect 546960 10888 547012 10940
rect 338120 10820 338172 10872
rect 540612 10820 540664 10872
rect 339500 10752 339552 10804
rect 540152 10752 540204 10804
rect 346400 10684 346452 10736
rect 546040 10684 546092 10736
rect 387064 10616 387116 10668
rect 540428 10616 540480 10668
rect 141240 10276 141292 10328
rect 557908 10276 557960 10328
rect 371700 8984 371752 9036
rect 553676 8984 553728 9036
rect 258264 8916 258316 8968
rect 553492 8916 553544 8968
rect 421380 7556 421432 7608
rect 559840 7556 559892 7608
rect 567844 7556 567896 7608
rect 579804 7556 579856 7608
rect 506480 6808 506532 6860
rect 566464 6808 566516 6860
rect 499396 6740 499448 6792
rect 571892 6740 571944 6792
rect 460388 6672 460440 6724
rect 541624 6672 541676 6724
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 485228 6604 485280 6656
rect 567292 6604 567344 6656
rect 463976 6536 464028 6588
rect 548800 6536 548852 6588
rect 446220 6468 446272 6520
rect 543096 6468 543148 6520
rect 449808 6400 449860 6452
rect 558000 6400 558052 6452
rect 442632 6332 442684 6384
rect 559380 6332 559432 6384
rect 439136 6264 439188 6316
rect 563520 6264 563572 6316
rect 432052 6196 432104 6248
rect 573272 6196 573324 6248
rect 332692 6128 332744 6180
rect 556252 6128 556304 6180
rect 288440 5448 288492 5500
rect 550364 5448 550416 5500
rect 375288 4836 375340 4888
rect 557540 4836 557592 4888
rect 318524 4768 318576 4820
rect 547144 4768 547196 4820
rect 38292 4088 38344 4140
rect 125876 4088 125928 4140
rect 492312 4088 492364 4140
rect 553860 4088 553912 4140
rect 42340 4020 42392 4072
rect 134156 4020 134208 4072
rect 488816 4020 488868 4072
rect 566372 4020 566424 4072
rect 48780 3952 48832 4004
rect 151820 3952 151872 4004
rect 424968 3952 425020 4004
rect 555148 3952 555200 4004
rect 565820 3952 565872 4004
rect 566096 3952 566148 4004
rect 43904 3884 43956 3936
rect 158904 3884 158956 3936
rect 286600 3884 286652 3936
rect 578700 3884 578752 3936
rect 48228 3816 48280 3868
rect 173164 3816 173216 3868
rect 239312 3816 239364 3868
rect 533344 3816 533396 3868
rect 534908 3816 534960 3868
rect 573456 3816 573508 3868
rect 45008 3748 45060 3800
rect 189724 3748 189776 3800
rect 244096 3748 244148 3800
rect 545764 3748 545816 3800
rect 552664 3748 552716 3800
rect 574284 3748 574336 3800
rect 34428 3680 34480 3732
rect 193220 3680 193272 3732
rect 218152 3680 218204 3732
rect 34152 3612 34204 3664
rect 196808 3612 196860 3664
rect 237012 3680 237064 3732
rect 581552 3680 581604 3732
rect 571616 3612 571668 3664
rect 31668 3544 31720 3596
rect 212172 3544 212224 3596
rect 218060 3544 218112 3596
rect 219256 3544 219308 3596
rect 219348 3544 219400 3596
rect 573088 3544 573140 3596
rect 41972 3476 42024 3528
rect 37188 3408 37240 3460
rect 161296 3408 161348 3460
rect 168380 3408 168432 3460
rect 42432 3340 42484 3392
rect 130568 3340 130620 3392
rect 135260 3340 135312 3392
rect 136456 3340 136508 3392
rect 50252 3272 50304 3324
rect 110512 3272 110564 3324
rect 184940 3476 184992 3528
rect 186136 3476 186188 3528
rect 190828 3476 190880 3528
rect 552848 3476 552900 3528
rect 572076 3476 572128 3528
rect 573916 3476 573968 3528
rect 187332 3340 187384 3392
rect 565820 3408 565872 3460
rect 215668 3340 215720 3392
rect 219348 3340 219400 3392
rect 234620 3340 234672 3392
rect 235816 3340 235868 3392
rect 259460 3340 259512 3392
rect 260656 3340 260708 3392
rect 299480 3340 299532 3392
rect 300768 3340 300820 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 495900 3340 495952 3392
rect 556436 3340 556488 3392
rect 510068 3272 510120 3324
rect 563428 3272 563480 3324
rect 578976 3272 579028 3324
rect 582196 3272 582248 3324
rect 545488 3204 545540 3256
rect 571708 3204 571760 3256
rect 527824 3136 527876 3188
rect 546684 3136 546736 3188
rect 552756 3000 552808 3052
rect 556160 3000 556212 3052
rect 324320 2048 324372 2100
rect 325608 2048 325660 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 6932 692102 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700369 24348 703520
rect 24306 700360 24362 700369
rect 24306 700295 24362 700304
rect 6920 692096 6972 692102
rect 6920 692038 6972 692044
rect 40052 687954 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 690674 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 693462 88380 702406
rect 105464 698970 105492 703520
rect 105452 698964 105504 698970
rect 105452 698906 105504 698912
rect 137848 697610 137876 703520
rect 137836 697604 137888 697610
rect 137836 697546 137888 697552
rect 154132 696250 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 696244 154172 696250
rect 154120 696186 154172 696192
rect 88340 693456 88392 693462
rect 88340 693398 88392 693404
rect 71780 690668 71832 690674
rect 71780 690610 71832 690616
rect 40040 687948 40092 687954
rect 40040 687890 40092 687896
rect 21362 683360 21418 683369
rect 21362 683295 21418 683304
rect 3424 682576 3476 682582
rect 3424 682518 3476 682524
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3436 553897 3464 682518
rect 9680 679108 9732 679114
rect 9680 679050 9732 679056
rect 3608 679040 3660 679046
rect 3608 678982 3660 678988
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 588606 3556 671191
rect 3620 658209 3648 678982
rect 7564 677612 7616 677618
rect 7564 677554 7616 677560
rect 3606 658200 3662 658209
rect 3606 658135 3662 658144
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3516 588600 3568 588606
rect 3516 588542 3568 588548
rect 3620 574802 3648 619103
rect 3698 606112 3754 606121
rect 3698 606047 3754 606056
rect 3712 584361 3740 606047
rect 3698 584352 3754 584361
rect 3698 584287 3754 584296
rect 3608 574796 3660 574802
rect 3608 574738 3660 574744
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 2962 201920 3018 201929
rect 2962 201855 3018 201864
rect 2976 194585 3004 201855
rect 3436 197334 3464 501735
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3528 345166 3556 345335
rect 3516 345160 3568 345166
rect 3516 345102 3568 345108
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3424 197328 3476 197334
rect 3424 197270 3476 197276
rect 2962 194576 3018 194585
rect 2962 194511 3018 194520
rect 2778 192536 2834 192545
rect 2778 192471 2834 192480
rect 4804 192500 4856 192506
rect 2792 16574 2820 192471
rect 4804 192442 4856 192448
rect 3424 191276 3476 191282
rect 3424 191218 3476 191224
rect 3148 137896 3200 137902
rect 3148 137838 3200 137844
rect 3160 136785 3188 137838
rect 3146 136776 3202 136785
rect 3146 136711 3202 136720
rect 2872 97776 2924 97782
rect 2872 97718 2924 97724
rect 2884 97617 2912 97718
rect 2870 97608 2926 97617
rect 2870 97543 2926 97552
rect 3436 58585 3464 191218
rect 3516 188964 3568 188970
rect 3516 188906 3568 188912
rect 3528 188873 3556 188906
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3528 149734 3556 149767
rect 3516 149728 3568 149734
rect 3516 149670 3568 149676
rect 4816 97782 4844 192442
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 2792 16546 2912 16574
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1688 480 1716 7511
rect 2884 480 2912 16546
rect 7576 6662 7604 677554
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 679050
rect 17224 565888 17276 565894
rect 17224 565830 17276 565836
rect 17236 193662 17264 565830
rect 19248 564732 19300 564738
rect 19248 564674 19300 564680
rect 18972 529984 19024 529990
rect 18972 529926 19024 529932
rect 17868 520328 17920 520334
rect 17868 520270 17920 520276
rect 17316 448588 17368 448594
rect 17316 448530 17368 448536
rect 17328 197062 17356 448530
rect 17408 397520 17460 397526
rect 17408 397462 17460 397468
rect 17420 199442 17448 397462
rect 17776 389224 17828 389230
rect 17776 389166 17828 389172
rect 17500 292596 17552 292602
rect 17500 292538 17552 292544
rect 17408 199436 17460 199442
rect 17408 199378 17460 199384
rect 17316 197056 17368 197062
rect 17316 196998 17368 197004
rect 17224 193656 17276 193662
rect 17224 193598 17276 193604
rect 17512 191826 17540 292538
rect 17500 191820 17552 191826
rect 17500 191762 17552 191768
rect 13820 170400 13872 170406
rect 13820 170342 13872 170348
rect 13832 16574 13860 170342
rect 17788 21214 17816 389166
rect 17776 21208 17828 21214
rect 17776 21150 17828 21156
rect 17880 19825 17908 520270
rect 18880 463752 18932 463758
rect 18880 463694 18932 463700
rect 18892 20194 18920 463694
rect 18984 69018 19012 529926
rect 19156 505164 19208 505170
rect 19156 505106 19208 505112
rect 19064 483064 19116 483070
rect 19064 483006 19116 483012
rect 18972 69012 19024 69018
rect 18972 68954 19024 68960
rect 19076 20534 19104 483006
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19168 20262 19196 505106
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 18880 20188 18932 20194
rect 18880 20130 18932 20136
rect 17866 19816 17922 19825
rect 17866 19751 17922 19760
rect 19260 19009 19288 564674
rect 20628 562012 20680 562018
rect 20628 561954 20680 561960
rect 19984 462392 20036 462398
rect 19984 462334 20036 462340
rect 19996 190466 20024 462334
rect 20168 414044 20220 414050
rect 20168 413986 20220 413992
rect 20180 194546 20208 413986
rect 20444 398880 20496 398886
rect 20444 398822 20496 398828
rect 20352 345092 20404 345098
rect 20352 345034 20404 345040
rect 20260 298172 20312 298178
rect 20260 298114 20312 298120
rect 20168 194540 20220 194546
rect 20168 194482 20220 194488
rect 19984 190460 20036 190466
rect 19984 190402 20036 190408
rect 20272 26042 20300 298114
rect 20260 26036 20312 26042
rect 20260 25978 20312 25984
rect 20364 20670 20392 345034
rect 20456 64870 20484 398822
rect 20536 394732 20588 394738
rect 20536 394674 20588 394680
rect 20444 64864 20496 64870
rect 20444 64806 20496 64812
rect 20352 20664 20404 20670
rect 20352 20606 20404 20612
rect 20548 20505 20576 394674
rect 20640 152697 20668 561954
rect 21272 300892 21324 300898
rect 21272 300834 21324 300840
rect 21284 189038 21312 300834
rect 21272 189032 21324 189038
rect 21272 188974 21324 188980
rect 20626 152688 20682 152697
rect 20626 152623 20682 152632
rect 21376 85542 21404 683295
rect 26882 683224 26938 683233
rect 26882 683159 26938 683168
rect 24674 681456 24730 681465
rect 24674 681391 24730 681400
rect 21824 587852 21876 587858
rect 21824 587794 21876 587800
rect 21732 561400 21784 561406
rect 21732 561342 21784 561348
rect 21640 484424 21692 484430
rect 21640 484366 21692 484372
rect 21456 407176 21508 407182
rect 21456 407118 21508 407124
rect 21468 196858 21496 407118
rect 21548 349172 21600 349178
rect 21548 349114 21600 349120
rect 21456 196852 21508 196858
rect 21456 196794 21508 196800
rect 21560 137970 21588 349114
rect 21652 151201 21680 484366
rect 21744 193730 21772 561342
rect 21836 198694 21864 587794
rect 23386 587208 23442 587217
rect 23386 587143 23442 587152
rect 22744 587036 22796 587042
rect 22744 586978 22796 586984
rect 22650 560960 22706 560969
rect 22650 560895 22706 560904
rect 22008 541000 22060 541006
rect 22008 540942 22060 540948
rect 21916 460964 21968 460970
rect 21916 460906 21968 460912
rect 21824 198688 21876 198694
rect 21824 198630 21876 198636
rect 21732 193724 21784 193730
rect 21732 193666 21784 193672
rect 21638 151192 21694 151201
rect 21638 151127 21694 151136
rect 21548 137964 21600 137970
rect 21548 137906 21600 137912
rect 21364 85536 21416 85542
rect 21364 85478 21416 85484
rect 21928 24614 21956 460906
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 22020 23361 22048 540942
rect 22560 302252 22612 302258
rect 22560 302194 22612 302200
rect 22572 25634 22600 302194
rect 22664 194274 22692 560895
rect 22756 198286 22784 586978
rect 22928 562624 22980 562630
rect 22928 562566 22980 562572
rect 22836 561944 22888 561950
rect 22836 561886 22888 561892
rect 22744 198280 22796 198286
rect 22744 198222 22796 198228
rect 22652 194268 22704 194274
rect 22652 194210 22704 194216
rect 22848 124166 22876 561886
rect 22836 124160 22888 124166
rect 22836 124102 22888 124108
rect 22940 117298 22968 562566
rect 23296 520396 23348 520402
rect 23296 520338 23348 520344
rect 23204 492720 23256 492726
rect 23204 492662 23256 492668
rect 23112 476128 23164 476134
rect 23112 476070 23164 476076
rect 23020 467900 23072 467906
rect 23020 467842 23072 467848
rect 22928 117292 22980 117298
rect 22928 117234 22980 117240
rect 22560 25628 22612 25634
rect 22560 25570 22612 25576
rect 22006 23352 22062 23361
rect 22006 23287 22062 23296
rect 20534 20496 20590 20505
rect 20534 20431 20590 20440
rect 23032 20330 23060 467842
rect 23124 25906 23152 476070
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 19246 19000 19302 19009
rect 19246 18935 19302 18944
rect 13832 16546 14320 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 23216 12442 23244 492662
rect 23308 29073 23336 520338
rect 23400 82822 23428 587143
rect 24492 563304 24544 563310
rect 24492 563246 24544 563252
rect 24308 563236 24360 563242
rect 24308 563178 24360 563184
rect 24124 423700 24176 423706
rect 24124 423642 24176 423648
rect 24032 281580 24084 281586
rect 24032 281522 24084 281528
rect 24044 193118 24072 281522
rect 24032 193112 24084 193118
rect 24032 193054 24084 193060
rect 24136 153134 24164 423642
rect 24216 415472 24268 415478
rect 24216 415414 24268 415420
rect 24124 153128 24176 153134
rect 24124 153070 24176 153076
rect 23388 82816 23440 82822
rect 23388 82758 23440 82764
rect 23294 29064 23350 29073
rect 23294 28999 23350 29008
rect 24228 24478 24256 415414
rect 24320 115258 24348 563178
rect 24400 561876 24452 561882
rect 24400 561818 24452 561824
rect 24308 115252 24360 115258
rect 24308 115194 24360 115200
rect 24412 103426 24440 561818
rect 24504 103494 24532 563246
rect 24582 560824 24638 560833
rect 24582 560759 24638 560768
rect 24492 103488 24544 103494
rect 24492 103430 24544 103436
rect 24400 103420 24452 103426
rect 24400 103362 24452 103368
rect 24596 34474 24624 560759
rect 24688 135250 24716 681391
rect 25780 589552 25832 589558
rect 25780 589494 25832 589500
rect 24768 563372 24820 563378
rect 24768 563314 24820 563320
rect 24676 135244 24728 135250
rect 24676 135186 24728 135192
rect 24584 34468 24636 34474
rect 24584 34410 24636 34416
rect 24216 24472 24268 24478
rect 24216 24414 24268 24420
rect 24780 17105 24808 563314
rect 25596 561264 25648 561270
rect 25596 561206 25648 561212
rect 25412 336796 25464 336802
rect 25412 336738 25464 336744
rect 25320 277432 25372 277438
rect 25320 277374 25372 277380
rect 25332 193186 25360 277374
rect 25320 193180 25372 193186
rect 25320 193122 25372 193128
rect 25424 162178 25452 336738
rect 25504 314696 25556 314702
rect 25504 314638 25556 314644
rect 25412 162172 25464 162178
rect 25412 162114 25464 162120
rect 25516 20466 25544 314638
rect 25608 199102 25636 561206
rect 25688 392012 25740 392018
rect 25688 391954 25740 391960
rect 25596 199096 25648 199102
rect 25596 199038 25648 199044
rect 25700 23118 25728 391954
rect 25792 197946 25820 589494
rect 26056 567248 26108 567254
rect 26056 567190 26108 567196
rect 25962 562048 26018 562057
rect 25962 561983 26018 561992
rect 25872 531344 25924 531350
rect 25872 531286 25924 531292
rect 25780 197940 25832 197946
rect 25780 197882 25832 197888
rect 25884 133890 25912 531286
rect 25976 160818 26004 561983
rect 25964 160812 26016 160818
rect 25964 160754 26016 160760
rect 25872 133884 25924 133890
rect 25872 133826 25924 133832
rect 26068 59362 26096 567190
rect 26146 561912 26202 561921
rect 26146 561847 26202 561856
rect 26056 59356 26108 59362
rect 26056 59298 26108 59304
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 26160 22030 26188 561847
rect 26792 419552 26844 419558
rect 26792 419494 26844 419500
rect 26700 305040 26752 305046
rect 26700 304982 26752 304988
rect 26712 193050 26740 304982
rect 26700 193044 26752 193050
rect 26700 192986 26752 192992
rect 26804 152862 26832 419494
rect 26896 255270 26924 683159
rect 169772 678298 169800 702406
rect 201512 694822 201540 702986
rect 218992 700466 219020 703520
rect 218980 700460 219032 700466
rect 218980 700402 219032 700408
rect 201500 694816 201552 694822
rect 201500 694758 201552 694764
rect 234632 688022 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700330 267688 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 300136 700398 300164 703520
rect 332520 700670 332548 703520
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 348804 700466 348832 703520
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 342996 700460 343048 700466
rect 342996 700402 343048 700408
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 234620 688016 234672 688022
rect 234620 687958 234672 687964
rect 171782 681320 171838 681329
rect 171782 681255 171838 681264
rect 165528 678292 165580 678298
rect 165528 678234 165580 678240
rect 169760 678292 169812 678298
rect 169760 678234 169812 678240
rect 165540 678201 165568 678234
rect 165526 678192 165582 678201
rect 165526 678127 165582 678136
rect 153108 677680 153160 677686
rect 153106 677648 153108 677657
rect 171140 677680 171192 677686
rect 153160 677648 153162 677657
rect 171140 677622 171192 677628
rect 153106 677583 153162 677592
rect 32862 628280 32918 628289
rect 32862 628215 32918 628224
rect 31574 628008 31630 628017
rect 31574 627943 31630 627952
rect 31390 625424 31446 625433
rect 31390 625359 31446 625368
rect 28906 587344 28962 587353
rect 28906 587279 28962 587288
rect 27526 562184 27582 562193
rect 27526 562119 27582 562128
rect 27342 561368 27398 561377
rect 27342 561303 27398 561312
rect 27252 561128 27304 561134
rect 27252 561070 27304 561076
rect 26976 514820 27028 514826
rect 26976 514762 27028 514768
rect 26884 255264 26936 255270
rect 26884 255206 26936 255212
rect 26882 254008 26938 254017
rect 26882 253943 26938 253952
rect 26792 152856 26844 152862
rect 26792 152798 26844 152804
rect 26896 26926 26924 253943
rect 26988 197198 27016 514762
rect 27068 444440 27120 444446
rect 27068 444382 27120 444388
rect 26976 197192 27028 197198
rect 26976 197134 27028 197140
rect 27080 151065 27108 444382
rect 27160 362976 27212 362982
rect 27160 362918 27212 362924
rect 27066 151056 27122 151065
rect 27066 150991 27122 151000
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 27172 23050 27200 362918
rect 27264 199170 27292 561070
rect 27252 199164 27304 199170
rect 27252 199106 27304 199112
rect 27356 100706 27384 561303
rect 27436 532772 27488 532778
rect 27436 532714 27488 532720
rect 27344 100700 27396 100706
rect 27344 100642 27396 100648
rect 27448 26246 27476 532714
rect 27436 26240 27488 26246
rect 27436 26182 27488 26188
rect 27160 23044 27212 23050
rect 27160 22986 27212 22992
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 27540 20398 27568 562119
rect 28724 561196 28776 561202
rect 28724 561138 28776 561144
rect 28632 489932 28684 489938
rect 28632 489874 28684 489880
rect 28356 419620 28408 419626
rect 28356 419562 28408 419568
rect 28264 372632 28316 372638
rect 28264 372574 28316 372580
rect 28080 357468 28132 357474
rect 28080 357410 28132 357416
rect 28092 198529 28120 357410
rect 28172 285728 28224 285734
rect 28172 285670 28224 285676
rect 28078 198520 28134 198529
rect 28078 198455 28134 198464
rect 27618 184512 27674 184521
rect 27618 184447 27674 184456
rect 27528 20392 27580 20398
rect 27528 20334 27580 20340
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 27632 16574 27660 184447
rect 28184 95198 28212 285670
rect 28276 151337 28304 372574
rect 28368 197266 28396 419562
rect 28448 380928 28500 380934
rect 28448 380870 28500 380876
rect 28356 197260 28408 197266
rect 28356 197202 28408 197208
rect 28460 155281 28488 380870
rect 28540 310548 28592 310554
rect 28540 310490 28592 310496
rect 28446 155272 28502 155281
rect 28446 155207 28502 155216
rect 28262 151328 28318 151337
rect 28262 151263 28318 151272
rect 28172 95192 28224 95198
rect 28172 95134 28224 95140
rect 28552 20602 28580 310490
rect 28644 155650 28672 489874
rect 28736 198626 28764 561138
rect 28816 415540 28868 415546
rect 28816 415482 28868 415488
rect 28724 198620 28776 198626
rect 28724 198562 28776 198568
rect 28632 155644 28684 155650
rect 28632 155586 28684 155592
rect 28828 27470 28856 415482
rect 28920 125594 28948 587279
rect 31404 577522 31432 625359
rect 31482 619712 31538 619721
rect 31482 619647 31538 619656
rect 31392 577516 31444 577522
rect 31392 577458 31444 577464
rect 31496 572014 31524 619647
rect 31588 591394 31616 627943
rect 32770 622432 32826 622441
rect 32770 622367 32826 622376
rect 31666 601760 31722 601769
rect 31666 601695 31722 601704
rect 31576 591388 31628 591394
rect 31576 591330 31628 591336
rect 31576 587444 31628 587450
rect 31576 587386 31628 587392
rect 31484 572008 31536 572014
rect 31484 571950 31536 571956
rect 31208 565412 31260 565418
rect 31208 565354 31260 565360
rect 30102 561776 30158 561785
rect 30102 561711 30158 561720
rect 29920 561536 29972 561542
rect 29920 561478 29972 561484
rect 29644 445800 29696 445806
rect 29644 445742 29696 445748
rect 29552 346452 29604 346458
rect 29552 346394 29604 346400
rect 29460 345160 29512 345166
rect 29460 345102 29512 345108
rect 29472 198393 29500 345102
rect 29458 198384 29514 198393
rect 29458 198319 29514 198328
rect 29564 194478 29592 346394
rect 29552 194472 29604 194478
rect 29552 194414 29604 194420
rect 29656 153202 29684 445742
rect 29828 386436 29880 386442
rect 29828 386378 29880 386384
rect 29736 371272 29788 371278
rect 29736 371214 29788 371220
rect 29644 153196 29696 153202
rect 29644 153138 29696 153144
rect 28908 125588 28960 125594
rect 28908 125530 28960 125536
rect 29748 29170 29776 371214
rect 29736 29164 29788 29170
rect 29736 29106 29788 29112
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 29840 26110 29868 386378
rect 29932 198558 29960 561478
rect 30010 561096 30066 561105
rect 30010 561031 30066 561040
rect 29920 198552 29972 198558
rect 29920 198494 29972 198500
rect 30024 192914 30052 561031
rect 30012 192908 30064 192914
rect 30012 192850 30064 192856
rect 30116 89690 30144 561711
rect 30196 549296 30248 549302
rect 30196 549238 30248 549244
rect 30104 89684 30156 89690
rect 30104 89626 30156 89632
rect 30208 48278 30236 549238
rect 30288 547936 30340 547942
rect 30288 547878 30340 547884
rect 30196 48272 30248 48278
rect 30196 48214 30248 48220
rect 30300 28937 30328 547878
rect 31024 328500 31076 328506
rect 31024 328442 31076 328448
rect 30932 267776 30984 267782
rect 30932 267718 30984 267724
rect 30840 234660 30892 234666
rect 30840 234602 30892 234608
rect 30852 151570 30880 234602
rect 30944 152998 30972 267718
rect 31036 159390 31064 328442
rect 31220 325650 31248 565354
rect 31484 561740 31536 561746
rect 31484 561682 31536 561688
rect 31392 458244 31444 458250
rect 31392 458186 31444 458192
rect 31300 379568 31352 379574
rect 31300 379510 31352 379516
rect 31208 325644 31260 325650
rect 31208 325586 31260 325592
rect 31116 223644 31168 223650
rect 31116 223586 31168 223592
rect 31024 159384 31076 159390
rect 31024 159326 31076 159332
rect 30932 152992 30984 152998
rect 30932 152934 30984 152940
rect 30840 151564 30892 151570
rect 30840 151506 30892 151512
rect 31128 29034 31156 223586
rect 31208 220856 31260 220862
rect 31208 220798 31260 220804
rect 31116 29028 31168 29034
rect 31116 28970 31168 28976
rect 30286 28928 30342 28937
rect 30286 28863 30342 28872
rect 29828 26104 29880 26110
rect 29828 26046 29880 26052
rect 31220 24410 31248 220798
rect 31312 140758 31340 379510
rect 31404 193225 31432 458186
rect 31496 198150 31524 561682
rect 31588 198218 31616 587386
rect 31680 198762 31708 601695
rect 32678 600400 32734 600409
rect 32678 600335 32734 600344
rect 32692 592006 32720 600335
rect 32680 592000 32732 592006
rect 32680 591942 32732 591948
rect 32404 591388 32456 591394
rect 32404 591330 32456 591336
rect 32416 386374 32444 591330
rect 32784 591326 32812 622367
rect 32876 591394 32904 628215
rect 33046 624200 33102 624209
rect 33046 624135 33102 624144
rect 32954 621344 33010 621353
rect 32954 621279 33010 621288
rect 32864 591388 32916 591394
rect 32864 591330 32916 591336
rect 32772 591320 32824 591326
rect 32772 591262 32824 591268
rect 32864 590028 32916 590034
rect 32864 589970 32916 589976
rect 32496 563168 32548 563174
rect 32496 563110 32548 563116
rect 32508 411262 32536 563110
rect 32772 560516 32824 560522
rect 32772 560458 32824 560464
rect 32678 560008 32734 560017
rect 32678 559943 32734 559952
rect 32496 411256 32548 411262
rect 32496 411198 32548 411204
rect 32404 386368 32456 386374
rect 32404 386310 32456 386316
rect 32128 367124 32180 367130
rect 32128 367066 32180 367072
rect 31668 198756 31720 198762
rect 31668 198698 31720 198704
rect 31576 198212 31628 198218
rect 31576 198154 31628 198160
rect 31484 198144 31536 198150
rect 31484 198086 31536 198092
rect 31390 193216 31446 193225
rect 31390 193151 31446 193160
rect 31576 192432 31628 192438
rect 31576 192374 31628 192380
rect 31392 181824 31444 181830
rect 31392 181766 31444 181772
rect 31300 140752 31352 140758
rect 31300 140694 31352 140700
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 31404 22574 31432 181766
rect 31484 181688 31536 181694
rect 31484 181630 31536 181636
rect 31392 22568 31444 22574
rect 31392 22510 31444 22516
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 31496 17134 31524 181630
rect 31484 17128 31536 17134
rect 31484 17070 31536 17076
rect 31588 16998 31616 192374
rect 31668 189780 31720 189786
rect 31668 189722 31720 189728
rect 31576 16992 31628 16998
rect 31576 16934 31628 16940
rect 27632 16546 28488 16574
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 19430 6216 19486 6225
rect 19430 6151 19486 6160
rect 19444 480 19472 6151
rect 24214 3496 24270 3505
rect 24214 3431 24270 3440
rect 24228 480 24256 3431
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 31680 3602 31708 189722
rect 31758 187232 31814 187241
rect 31758 187167 31814 187176
rect 31772 16574 31800 187167
rect 32140 25770 32168 367066
rect 32692 331226 32720 559943
rect 32784 367062 32812 560458
rect 32772 367056 32824 367062
rect 32772 366998 32824 367004
rect 32680 331220 32732 331226
rect 32680 331162 32732 331168
rect 32404 320204 32456 320210
rect 32404 320146 32456 320152
rect 32220 240168 32272 240174
rect 32220 240110 32272 240116
rect 32232 195906 32260 240110
rect 32312 227792 32364 227798
rect 32312 227734 32364 227740
rect 32220 195900 32272 195906
rect 32220 195842 32272 195848
rect 32324 152658 32352 227734
rect 32416 195770 32444 320146
rect 32496 292596 32548 292602
rect 32496 292538 32548 292544
rect 32404 195764 32456 195770
rect 32404 195706 32456 195712
rect 32402 186960 32458 186969
rect 32402 186895 32458 186904
rect 32312 152652 32364 152658
rect 32312 152594 32364 152600
rect 32416 137902 32444 186895
rect 32508 152794 32536 292538
rect 32588 281648 32640 281654
rect 32588 281590 32640 281596
rect 32496 152788 32548 152794
rect 32496 152730 32548 152736
rect 32404 137896 32456 137902
rect 32404 137838 32456 137844
rect 32600 132462 32628 281590
rect 32680 273284 32732 273290
rect 32680 273226 32732 273232
rect 32588 132456 32640 132462
rect 32588 132398 32640 132404
rect 32128 25764 32180 25770
rect 32128 25706 32180 25712
rect 32692 20641 32720 273226
rect 32876 198422 32904 589970
rect 32968 202842 32996 621279
rect 32956 202836 33008 202842
rect 32956 202778 33008 202784
rect 33060 198801 33088 624135
rect 78864 591388 78916 591394
rect 78864 591330 78916 591336
rect 153660 591388 153712 591394
rect 153660 591330 153712 591336
rect 37004 590708 37056 590714
rect 37004 590650 37056 590656
rect 35254 589928 35310 589937
rect 35254 589863 35310 589872
rect 34888 587648 34940 587654
rect 34888 587590 34940 587596
rect 34428 565888 34480 565894
rect 34428 565830 34480 565836
rect 33968 564868 34020 564874
rect 33968 564810 34020 564816
rect 33600 469260 33652 469266
rect 33600 469202 33652 469208
rect 33046 198792 33102 198801
rect 33046 198727 33102 198736
rect 32864 198416 32916 198422
rect 32864 198358 32916 198364
rect 33048 181892 33100 181898
rect 33048 181834 33100 181840
rect 32678 20632 32734 20641
rect 32678 20567 32734 20576
rect 33060 19990 33088 181834
rect 33612 25702 33640 469202
rect 33876 433356 33928 433362
rect 33876 433298 33928 433304
rect 33784 427848 33836 427854
rect 33784 427790 33836 427796
rect 33692 309188 33744 309194
rect 33692 309130 33744 309136
rect 33704 194410 33732 309130
rect 33692 194404 33744 194410
rect 33692 194346 33744 194352
rect 33690 184784 33746 184793
rect 33690 184719 33746 184728
rect 33704 33114 33732 184719
rect 33796 184550 33824 427790
rect 33784 184544 33836 184550
rect 33784 184486 33836 184492
rect 33784 181756 33836 181762
rect 33784 181698 33836 181704
rect 33692 33108 33744 33114
rect 33692 33050 33744 33056
rect 33600 25696 33652 25702
rect 33600 25638 33652 25644
rect 33796 24342 33824 181698
rect 33888 158030 33916 433298
rect 33980 268394 34008 564810
rect 34152 563780 34204 563786
rect 34152 563722 34204 563728
rect 34060 560992 34112 560998
rect 34060 560934 34112 560940
rect 33968 268388 34020 268394
rect 33968 268330 34020 268336
rect 33968 231872 34020 231878
rect 33968 231814 34020 231820
rect 33876 158024 33928 158030
rect 33876 157966 33928 157972
rect 33980 29442 34008 231814
rect 34072 198966 34100 560934
rect 34164 199209 34192 563722
rect 34336 545148 34388 545154
rect 34336 545090 34388 545096
rect 34244 516180 34296 516186
rect 34244 516122 34296 516128
rect 34150 199200 34206 199209
rect 34150 199135 34206 199144
rect 34060 198960 34112 198966
rect 34060 198902 34112 198908
rect 34060 192840 34112 192846
rect 34060 192782 34112 192788
rect 34072 33046 34100 192782
rect 34152 188420 34204 188426
rect 34152 188362 34204 188368
rect 34060 33040 34112 33046
rect 34060 32982 34112 32988
rect 33968 29436 34020 29442
rect 33968 29378 34020 29384
rect 33784 24336 33836 24342
rect 33784 24278 33836 24284
rect 33048 19984 33100 19990
rect 33048 19926 33100 19932
rect 31772 16546 31984 16574
rect 31668 3596 31720 3602
rect 31668 3538 31720 3544
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 34164 3670 34192 188362
rect 34256 152969 34284 516122
rect 34348 177478 34376 545090
rect 34440 451246 34468 565830
rect 34428 451240 34480 451246
rect 34428 451182 34480 451188
rect 34796 222216 34848 222222
rect 34796 222158 34848 222164
rect 34428 181620 34480 181626
rect 34428 181562 34480 181568
rect 34336 177472 34388 177478
rect 34336 177414 34388 177420
rect 34242 152960 34298 152969
rect 34242 152895 34298 152904
rect 34440 3738 34468 181562
rect 34808 28626 34836 222158
rect 34900 198665 34928 587590
rect 34980 564800 35032 564806
rect 34980 564742 35032 564748
rect 34992 211857 35020 564742
rect 35164 420980 35216 420986
rect 35164 420922 35216 420928
rect 35072 256012 35124 256018
rect 35072 255954 35124 255960
rect 35084 224233 35112 255954
rect 35070 224224 35126 224233
rect 35070 224159 35126 224168
rect 34978 211848 35034 211857
rect 34978 211783 35034 211792
rect 35072 211200 35124 211206
rect 35072 211142 35124 211148
rect 34886 198656 34942 198665
rect 34886 198591 34942 198600
rect 35084 151094 35112 211142
rect 35176 172310 35204 420922
rect 35268 293962 35296 589863
rect 36728 587172 36780 587178
rect 36728 587114 36780 587120
rect 36544 568608 36596 568614
rect 36544 568550 36596 568556
rect 35624 565956 35676 565962
rect 35624 565898 35676 565904
rect 35348 564936 35400 564942
rect 35348 564878 35400 564884
rect 35256 293956 35308 293962
rect 35256 293898 35308 293904
rect 35256 230512 35308 230518
rect 35256 230454 35308 230460
rect 35268 197130 35296 230454
rect 35360 221746 35388 564878
rect 35532 561332 35584 561338
rect 35532 561274 35584 561280
rect 35348 221740 35400 221746
rect 35348 221682 35400 221688
rect 35440 218068 35492 218074
rect 35440 218010 35492 218016
rect 35256 197124 35308 197130
rect 35256 197066 35308 197072
rect 35256 181552 35308 181558
rect 35256 181494 35308 181500
rect 35164 172304 35216 172310
rect 35164 172246 35216 172252
rect 35072 151088 35124 151094
rect 35072 151030 35124 151036
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 35268 17513 35296 181494
rect 35452 28558 35480 218010
rect 35544 199238 35572 561274
rect 35636 463690 35664 565898
rect 35808 562284 35860 562290
rect 35808 562226 35860 562232
rect 35624 463684 35676 463690
rect 35624 463626 35676 463632
rect 35624 411324 35676 411330
rect 35624 411266 35676 411272
rect 35532 199232 35584 199238
rect 35532 199174 35584 199180
rect 35532 189916 35584 189922
rect 35532 189858 35584 189864
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 35254 17504 35310 17513
rect 35254 17439 35310 17448
rect 35544 17338 35572 189858
rect 35636 27130 35664 411266
rect 35716 202904 35768 202910
rect 35716 202846 35768 202852
rect 35624 27124 35676 27130
rect 35624 27066 35676 27072
rect 35728 26178 35756 202846
rect 35820 153105 35848 562226
rect 36268 562216 36320 562222
rect 36268 562158 36320 562164
rect 36176 385076 36228 385082
rect 36176 385018 36228 385024
rect 35900 191140 35952 191146
rect 35900 191082 35952 191088
rect 35806 153096 35862 153105
rect 35806 153031 35862 153040
rect 35716 26172 35768 26178
rect 35716 26114 35768 26120
rect 35532 17332 35584 17338
rect 35532 17274 35584 17280
rect 35912 16574 35940 191082
rect 36188 121446 36216 385018
rect 36280 195090 36308 562158
rect 36452 380996 36504 381002
rect 36452 380938 36504 380944
rect 36464 253706 36492 380938
rect 36556 353258 36584 568550
rect 36636 564528 36688 564534
rect 36636 564470 36688 564476
rect 36544 353252 36596 353258
rect 36544 353194 36596 353200
rect 36544 322992 36596 322998
rect 36544 322934 36596 322940
rect 36452 253700 36504 253706
rect 36452 253642 36504 253648
rect 36452 247104 36504 247110
rect 36452 247046 36504 247052
rect 36360 221740 36412 221746
rect 36360 221682 36412 221688
rect 36372 209098 36400 221682
rect 36360 209092 36412 209098
rect 36360 209034 36412 209040
rect 36268 195084 36320 195090
rect 36268 195026 36320 195032
rect 36464 152522 36492 247046
rect 36556 199753 36584 322934
rect 36648 310486 36676 564470
rect 36740 383654 36768 587114
rect 36912 565072 36964 565078
rect 36912 565014 36964 565020
rect 36820 559564 36872 559570
rect 36820 559506 36872 559512
rect 36728 383648 36780 383654
rect 36728 383590 36780 383596
rect 36636 310480 36688 310486
rect 36636 310422 36688 310428
rect 36636 298580 36688 298586
rect 36636 298522 36688 298528
rect 36648 256018 36676 298522
rect 36832 269822 36860 559506
rect 36820 269816 36872 269822
rect 36820 269758 36872 269764
rect 36820 267844 36872 267850
rect 36820 267786 36872 267792
rect 36636 256012 36688 256018
rect 36636 255954 36688 255960
rect 36636 253972 36688 253978
rect 36636 253914 36688 253920
rect 36542 199744 36598 199753
rect 36542 199679 36598 199688
rect 36648 152590 36676 253914
rect 36636 152584 36688 152590
rect 36636 152526 36688 152532
rect 36452 152516 36504 152522
rect 36452 152458 36504 152464
rect 36176 121440 36228 121446
rect 36176 121382 36228 121388
rect 35912 16546 36032 16574
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34152 3664 34204 3670
rect 34152 3606 34204 3612
rect 36004 480 36032 16546
rect 36832 11830 36860 267786
rect 36924 218754 36952 565014
rect 37016 238746 37044 590650
rect 50066 590608 50122 590617
rect 50066 590543 50122 590552
rect 55862 590608 55918 590617
rect 55862 590543 55918 590552
rect 60370 590608 60426 590617
rect 60370 590543 60426 590552
rect 69018 590608 69074 590617
rect 69018 590543 69074 590552
rect 74814 590608 74870 590617
rect 74814 590543 74870 590552
rect 77850 590608 77906 590617
rect 77850 590543 77906 590552
rect 48964 590300 49016 590306
rect 48964 590242 49016 590248
rect 42616 590232 42668 590238
rect 42616 590174 42668 590180
rect 42522 590064 42578 590073
rect 42522 589999 42578 590008
rect 41236 589960 41288 589966
rect 41236 589902 41288 589908
rect 41144 589484 41196 589490
rect 41144 589426 41196 589432
rect 38384 589416 38436 589422
rect 38384 589358 38436 589364
rect 37096 563848 37148 563854
rect 37096 563790 37148 563796
rect 37004 238740 37056 238746
rect 37004 238682 37056 238688
rect 37004 238060 37056 238066
rect 37004 238002 37056 238008
rect 37016 221474 37044 238002
rect 37004 221468 37056 221474
rect 37004 221410 37056 221416
rect 36912 218748 36964 218754
rect 36912 218690 36964 218696
rect 36912 216776 36964 216782
rect 36912 216718 36964 216724
rect 36924 197742 36952 216718
rect 37004 216708 37056 216714
rect 37004 216650 37056 216656
rect 36912 197736 36964 197742
rect 36912 197678 36964 197684
rect 36912 192636 36964 192642
rect 36912 192578 36964 192584
rect 36924 21554 36952 192578
rect 37016 24682 37044 216650
rect 37108 196790 37136 563790
rect 38108 563508 38160 563514
rect 38108 563450 38160 563456
rect 37832 560312 37884 560318
rect 37832 560254 37884 560260
rect 37844 358766 37872 560254
rect 38016 513392 38068 513398
rect 38016 513334 38068 513340
rect 37924 392080 37976 392086
rect 37924 392022 37976 392028
rect 37832 358760 37884 358766
rect 37832 358702 37884 358708
rect 37832 354748 37884 354754
rect 37832 354690 37884 354696
rect 37188 257372 37240 257378
rect 37188 257314 37240 257320
rect 37200 247722 37228 257314
rect 37188 247716 37240 247722
rect 37188 247658 37240 247664
rect 37648 220312 37700 220318
rect 37648 220254 37700 220260
rect 37660 209774 37688 220254
rect 37740 215348 37792 215354
rect 37740 215290 37792 215296
rect 37568 209746 37688 209774
rect 37188 205692 37240 205698
rect 37188 205634 37240 205640
rect 37200 199889 37228 205634
rect 37568 201113 37596 209746
rect 37646 201376 37702 201385
rect 37646 201311 37702 201320
rect 37554 201104 37610 201113
rect 37554 201039 37610 201048
rect 37186 199880 37242 199889
rect 37186 199815 37242 199824
rect 37096 196784 37148 196790
rect 37096 196726 37148 196732
rect 37096 192364 37148 192370
rect 37096 192306 37148 192312
rect 37004 24676 37056 24682
rect 37004 24618 37056 24624
rect 36912 21548 36964 21554
rect 36912 21490 36964 21496
rect 37108 19854 37136 192306
rect 37188 176248 37240 176254
rect 37188 176190 37240 176196
rect 37096 19848 37148 19854
rect 37096 19790 37148 19796
rect 36820 11824 36872 11830
rect 36820 11766 36872 11772
rect 37200 3466 37228 176190
rect 37660 26654 37688 201311
rect 37752 155582 37780 215290
rect 37844 156806 37872 354690
rect 37936 170678 37964 392022
rect 38028 173330 38056 513334
rect 38120 218686 38148 563450
rect 38292 562080 38344 562086
rect 38292 562022 38344 562028
rect 38200 561060 38252 561066
rect 38200 561002 38252 561008
rect 38108 218680 38160 218686
rect 38108 218622 38160 218628
rect 38212 195809 38240 561002
rect 38198 195800 38254 195809
rect 38198 195735 38254 195744
rect 38304 195362 38332 562022
rect 38396 197849 38424 589358
rect 40960 587784 41012 587790
rect 40960 587726 41012 587732
rect 40868 587716 40920 587722
rect 40868 587658 40920 587664
rect 39948 587308 40000 587314
rect 39948 587250 40000 587256
rect 39580 566500 39632 566506
rect 39580 566442 39632 566448
rect 39304 563576 39356 563582
rect 39304 563518 39356 563524
rect 38568 514820 38620 514826
rect 38568 514762 38620 514768
rect 38476 443012 38528 443018
rect 38476 442954 38528 442960
rect 38382 197840 38438 197849
rect 38382 197775 38438 197784
rect 38292 195356 38344 195362
rect 38292 195298 38344 195304
rect 38108 184272 38160 184278
rect 38108 184214 38160 184220
rect 38016 173324 38068 173330
rect 38016 173266 38068 173272
rect 37924 170672 37976 170678
rect 37924 170614 37976 170620
rect 37832 156800 37884 156806
rect 37832 156742 37884 156748
rect 37740 155576 37792 155582
rect 37740 155518 37792 155524
rect 38016 155236 38068 155242
rect 38016 155178 38068 155184
rect 37924 152720 37976 152726
rect 37924 152662 37976 152668
rect 37648 26648 37700 26654
rect 37648 26590 37700 26596
rect 37936 21758 37964 152662
rect 37924 21752 37976 21758
rect 37924 21694 37976 21700
rect 38028 18358 38056 155178
rect 38120 19922 38148 184214
rect 38200 184204 38252 184210
rect 38200 184146 38252 184152
rect 38108 19916 38160 19922
rect 38108 19858 38160 19864
rect 38212 18970 38240 184146
rect 38290 176080 38346 176089
rect 38290 176015 38346 176024
rect 38200 18964 38252 18970
rect 38200 18906 38252 18912
rect 38016 18352 38068 18358
rect 38016 18294 38068 18300
rect 38304 4146 38332 176015
rect 38488 23322 38516 442954
rect 38476 23316 38528 23322
rect 38476 23258 38528 23264
rect 38580 23254 38608 514762
rect 39120 495508 39172 495514
rect 39120 495450 39172 495456
rect 38660 179104 38712 179110
rect 38660 179046 38712 179052
rect 38568 23248 38620 23254
rect 38568 23190 38620 23196
rect 38672 16574 38700 179046
rect 39132 28218 39160 495450
rect 39212 281716 39264 281722
rect 39212 281658 39264 281664
rect 39224 198490 39252 281658
rect 39316 220318 39344 563518
rect 39488 560448 39540 560454
rect 39488 560390 39540 560396
rect 39396 559632 39448 559638
rect 39396 559574 39448 559580
rect 39408 298586 39436 559574
rect 39500 460902 39528 560390
rect 39488 460896 39540 460902
rect 39488 460838 39540 460844
rect 39488 418192 39540 418198
rect 39488 418134 39540 418140
rect 39396 298580 39448 298586
rect 39396 298522 39448 298528
rect 39396 296744 39448 296750
rect 39396 296686 39448 296692
rect 39304 220312 39356 220318
rect 39304 220254 39356 220260
rect 39304 218136 39356 218142
rect 39304 218078 39356 218084
rect 39212 198484 39264 198490
rect 39212 198426 39264 198432
rect 39212 155780 39264 155786
rect 39212 155722 39264 155728
rect 39120 28212 39172 28218
rect 39120 28154 39172 28160
rect 39224 18902 39252 155722
rect 39212 18896 39264 18902
rect 39212 18838 39264 18844
rect 39316 17950 39344 218078
rect 39408 28082 39436 296686
rect 39500 128314 39528 418134
rect 39592 208350 39620 566442
rect 39856 564596 39908 564602
rect 39856 564538 39908 564544
rect 39672 563916 39724 563922
rect 39672 563858 39724 563864
rect 39580 208344 39632 208350
rect 39580 208286 39632 208292
rect 39684 199306 39712 563858
rect 39764 562352 39816 562358
rect 39764 562294 39816 562300
rect 39672 199300 39724 199306
rect 39672 199242 39724 199248
rect 39776 195974 39804 562294
rect 39868 510610 39896 564538
rect 39856 510604 39908 510610
rect 39856 510546 39908 510552
rect 39960 502110 39988 587250
rect 40776 566024 40828 566030
rect 40776 565966 40828 565972
rect 40684 565004 40736 565010
rect 40684 564946 40736 564952
rect 40408 528624 40460 528630
rect 40408 528566 40460 528572
rect 39948 502104 40000 502110
rect 39948 502046 40000 502052
rect 39856 485852 39908 485858
rect 39856 485794 39908 485800
rect 39764 195968 39816 195974
rect 39764 195910 39816 195916
rect 39762 195528 39818 195537
rect 39762 195463 39818 195472
rect 39670 178936 39726 178945
rect 39670 178871 39726 178880
rect 39580 154148 39632 154154
rect 39580 154090 39632 154096
rect 39488 128308 39540 128314
rect 39488 128250 39540 128256
rect 39396 28076 39448 28082
rect 39396 28018 39448 28024
rect 39304 17944 39356 17950
rect 39304 17886 39356 17892
rect 39592 17678 39620 154090
rect 39684 22778 39712 178871
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39776 18834 39804 195463
rect 39868 28830 39896 485794
rect 39948 221740 40000 221746
rect 39948 221682 40000 221688
rect 39960 198898 39988 221682
rect 39948 198892 40000 198898
rect 39948 198834 40000 198840
rect 40224 194880 40276 194886
rect 40224 194822 40276 194828
rect 39856 28824 39908 28830
rect 39856 28766 39908 28772
rect 40236 21418 40264 194822
rect 40314 183288 40370 183297
rect 40314 183223 40370 183232
rect 40328 140690 40356 183223
rect 40420 183122 40448 528566
rect 40696 508366 40724 564946
rect 40684 508360 40736 508366
rect 40684 508302 40736 508308
rect 40788 496806 40816 565966
rect 40880 500954 40908 587658
rect 40972 521558 41000 587726
rect 41052 558952 41104 558958
rect 41052 558894 41104 558900
rect 40960 521552 41012 521558
rect 40960 521494 41012 521500
rect 40868 500948 40920 500954
rect 40868 500890 40920 500896
rect 40776 496800 40828 496806
rect 40776 496742 40828 496748
rect 40868 490000 40920 490006
rect 40868 489942 40920 489948
rect 40776 467968 40828 467974
rect 40776 467910 40828 467916
rect 40592 464160 40644 464166
rect 40592 464102 40644 464108
rect 40500 427916 40552 427922
rect 40500 427858 40552 427864
rect 40408 183116 40460 183122
rect 40408 183058 40460 183064
rect 40512 180402 40540 427858
rect 40604 196654 40632 464102
rect 40684 439000 40736 439006
rect 40684 438942 40736 438948
rect 40592 196648 40644 196654
rect 40592 196590 40644 196596
rect 40592 187332 40644 187338
rect 40592 187274 40644 187280
rect 40500 180396 40552 180402
rect 40500 180338 40552 180344
rect 40316 140684 40368 140690
rect 40316 140626 40368 140632
rect 40604 120018 40632 187274
rect 40696 164966 40724 438942
rect 40788 166462 40816 467910
rect 40880 179246 40908 489942
rect 41064 195673 41092 558894
rect 41156 198354 41184 589426
rect 41144 198348 41196 198354
rect 41144 198290 41196 198296
rect 41050 195664 41106 195673
rect 41050 195599 41106 195608
rect 41248 194342 41276 589902
rect 41972 586560 42024 586566
rect 41972 586502 42024 586508
rect 41880 562488 41932 562494
rect 41880 562430 41932 562436
rect 41328 561808 41380 561814
rect 41328 561750 41380 561756
rect 41236 194336 41288 194342
rect 41236 194278 41288 194284
rect 40868 179240 40920 179246
rect 40868 179182 40920 179188
rect 41052 178492 41104 178498
rect 41052 178434 41104 178440
rect 40960 176044 41012 176050
rect 40960 175986 41012 175992
rect 40776 166456 40828 166462
rect 40776 166398 40828 166404
rect 40684 164960 40736 164966
rect 40684 164902 40736 164908
rect 40868 155304 40920 155310
rect 40868 155246 40920 155252
rect 40592 120012 40644 120018
rect 40592 119954 40644 119960
rect 40880 25974 40908 155246
rect 40868 25968 40920 25974
rect 40868 25910 40920 25916
rect 40972 22846 41000 175986
rect 40960 22840 41012 22846
rect 40960 22782 41012 22788
rect 41064 22506 41092 178434
rect 41144 177540 41196 177546
rect 41144 177482 41196 177488
rect 41052 22500 41104 22506
rect 41052 22442 41104 22448
rect 40224 21412 40276 21418
rect 40224 21354 40276 21360
rect 41156 19786 41184 177482
rect 41236 166592 41288 166598
rect 41236 166534 41288 166540
rect 41248 91050 41276 166534
rect 41236 91044 41288 91050
rect 41236 90986 41288 90992
rect 41340 28422 41368 561750
rect 41788 551200 41840 551206
rect 41788 551142 41840 551148
rect 41696 438932 41748 438938
rect 41696 438874 41748 438880
rect 41708 28694 41736 438874
rect 41800 62082 41828 551142
rect 41892 480486 41920 562430
rect 41984 495446 42012 586502
rect 42156 565276 42208 565282
rect 42156 565218 42208 565224
rect 42064 563984 42116 563990
rect 42064 563926 42116 563932
rect 41972 495440 42024 495446
rect 41972 495382 42024 495388
rect 41880 480480 41932 480486
rect 41880 480422 41932 480428
rect 41972 403028 42024 403034
rect 41972 402970 42024 402976
rect 41984 195294 42012 402970
rect 42076 221746 42104 563926
rect 42168 402150 42196 565218
rect 42432 565140 42484 565146
rect 42432 565082 42484 565088
rect 42246 560144 42302 560153
rect 42246 560079 42302 560088
rect 42156 402144 42208 402150
rect 42156 402086 42208 402092
rect 42156 400240 42208 400246
rect 42156 400182 42208 400188
rect 42064 221740 42116 221746
rect 42064 221682 42116 221688
rect 42062 209536 42118 209545
rect 42062 209471 42118 209480
rect 41972 195288 42024 195294
rect 41972 195230 42024 195236
rect 41880 188556 41932 188562
rect 41880 188498 41932 188504
rect 41788 62076 41840 62082
rect 41788 62018 41840 62024
rect 41696 28688 41748 28694
rect 41696 28630 41748 28636
rect 41328 28416 41380 28422
rect 41328 28358 41380 28364
rect 41892 27266 41920 188498
rect 41972 176180 42024 176186
rect 41972 176122 42024 176128
rect 41880 27260 41932 27266
rect 41880 27202 41932 27208
rect 41144 19780 41196 19786
rect 41144 19722 41196 19728
rect 39764 18828 39816 18834
rect 39764 18770 39816 18776
rect 39580 17672 39632 17678
rect 39580 17614 39632 17620
rect 38672 16546 39160 16574
rect 38292 4140 38344 4146
rect 38292 4082 38344 4088
rect 37188 3460 37240 3466
rect 37188 3402 37240 3408
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41984 3534 42012 176122
rect 42076 26722 42104 209471
rect 42168 163606 42196 400182
rect 42260 321570 42288 560079
rect 42340 550860 42392 550866
rect 42340 550802 42392 550808
rect 42248 321564 42300 321570
rect 42248 321506 42300 321512
rect 42248 318980 42300 318986
rect 42248 318922 42300 318928
rect 42156 163600 42208 163606
rect 42156 163542 42208 163548
rect 42260 29102 42288 318922
rect 42352 196722 42380 550802
rect 42444 206990 42472 565082
rect 42536 498166 42564 589999
rect 42524 498160 42576 498166
rect 42524 498102 42576 498108
rect 42628 489870 42656 590174
rect 45284 590164 45336 590170
rect 45284 590106 45336 590112
rect 45100 590096 45152 590102
rect 45100 590038 45152 590044
rect 43720 589892 43772 589898
rect 43720 589834 43772 589840
rect 43444 564120 43496 564126
rect 43444 564062 43496 564068
rect 43352 562148 43404 562154
rect 43352 562090 43404 562096
rect 43364 562018 43392 562090
rect 43352 562012 43404 562018
rect 43352 561954 43404 561960
rect 43350 558920 43406 558929
rect 43350 558855 43406 558864
rect 43076 543788 43128 543794
rect 43076 543730 43128 543736
rect 42616 489864 42668 489870
rect 42616 489806 42668 489812
rect 42524 431996 42576 432002
rect 42524 431938 42576 431944
rect 42432 206984 42484 206990
rect 42432 206926 42484 206932
rect 42340 196716 42392 196722
rect 42340 196658 42392 196664
rect 42432 187264 42484 187270
rect 42432 187206 42484 187212
rect 42340 179036 42392 179042
rect 42340 178978 42392 178984
rect 42248 29096 42300 29102
rect 42248 29038 42300 29044
rect 42064 26716 42116 26722
rect 42064 26658 42116 26664
rect 42352 4078 42380 178978
rect 42340 4072 42392 4078
rect 42340 4014 42392 4020
rect 41972 3528 42024 3534
rect 41972 3470 42024 3476
rect 42444 3398 42472 187206
rect 42536 29374 42564 431938
rect 42708 236020 42760 236026
rect 42708 235962 42760 235968
rect 42616 219496 42668 219502
rect 42616 219438 42668 219444
rect 42628 199578 42656 219438
rect 42616 199572 42668 199578
rect 42616 199514 42668 199520
rect 42720 196994 42748 235962
rect 42708 196988 42760 196994
rect 42708 196930 42760 196936
rect 43088 29510 43116 543730
rect 43364 323542 43392 558855
rect 43456 538218 43484 564062
rect 43628 563712 43680 563718
rect 43628 563654 43680 563660
rect 43536 560380 43588 560386
rect 43536 560322 43588 560328
rect 43444 538212 43496 538218
rect 43444 538154 43496 538160
rect 43548 474638 43576 560322
rect 43536 474632 43588 474638
rect 43536 474574 43588 474580
rect 43536 436144 43588 436150
rect 43536 436086 43588 436092
rect 43444 425128 43496 425134
rect 43444 425070 43496 425076
rect 43352 323536 43404 323542
rect 43352 323478 43404 323484
rect 43352 321632 43404 321638
rect 43352 321574 43404 321580
rect 43260 294024 43312 294030
rect 43260 293966 43312 293972
rect 43168 253700 43220 253706
rect 43168 253642 43220 253648
rect 43180 218618 43208 253642
rect 43272 236026 43300 293966
rect 43260 236020 43312 236026
rect 43260 235962 43312 235968
rect 43168 218612 43220 218618
rect 43168 218554 43220 218560
rect 43168 188760 43220 188766
rect 43168 188702 43220 188708
rect 43180 115938 43208 188702
rect 43260 188624 43312 188630
rect 43260 188566 43312 188572
rect 43168 115932 43220 115938
rect 43168 115874 43220 115880
rect 43272 109002 43300 188566
rect 43364 166326 43392 321574
rect 43456 176390 43484 425070
rect 43548 185774 43576 436086
rect 43640 292641 43668 563654
rect 43732 302190 43760 589834
rect 44640 589824 44692 589830
rect 44640 589766 44692 589772
rect 44088 587376 44140 587382
rect 44088 587318 44140 587324
rect 43996 587240 44048 587246
rect 43996 587182 44048 587188
rect 43904 580508 43956 580514
rect 43904 580450 43956 580456
rect 43810 561232 43866 561241
rect 43810 561167 43866 561176
rect 43824 371210 43852 561167
rect 43812 371204 43864 371210
rect 43812 371146 43864 371152
rect 43812 368552 43864 368558
rect 43812 368494 43864 368500
rect 43720 302184 43772 302190
rect 43720 302126 43772 302132
rect 43626 292632 43682 292641
rect 43626 292567 43682 292576
rect 43720 291236 43772 291242
rect 43720 291178 43772 291184
rect 43628 284708 43680 284714
rect 43628 284650 43680 284656
rect 43640 253706 43668 284650
rect 43628 253700 43680 253706
rect 43628 253642 43680 253648
rect 43628 218680 43680 218686
rect 43628 218622 43680 218628
rect 43536 185768 43588 185774
rect 43536 185710 43588 185716
rect 43536 182980 43588 182986
rect 43536 182922 43588 182928
rect 43444 176384 43496 176390
rect 43444 176326 43496 176332
rect 43352 166320 43404 166326
rect 43352 166262 43404 166268
rect 43260 108996 43312 109002
rect 43260 108938 43312 108944
rect 43548 63510 43576 182922
rect 43536 63504 43588 63510
rect 43536 63446 43588 63452
rect 43076 29504 43128 29510
rect 43076 29446 43128 29452
rect 42524 29368 42576 29374
rect 42524 29310 42576 29316
rect 43640 26994 43668 218622
rect 43732 195401 43760 291178
rect 43718 195392 43774 195401
rect 43718 195327 43774 195336
rect 43720 185904 43772 185910
rect 43720 185846 43772 185852
rect 43628 26988 43680 26994
rect 43628 26930 43680 26936
rect 43732 18766 43760 185846
rect 43824 27946 43852 368494
rect 43916 234054 43944 580450
rect 44008 456754 44036 587182
rect 44100 525774 44128 587318
rect 44548 556232 44600 556238
rect 44548 556174 44600 556180
rect 44088 525768 44140 525774
rect 44088 525710 44140 525716
rect 43996 456748 44048 456754
rect 43996 456690 44048 456696
rect 43996 434784 44048 434790
rect 43996 434726 44048 434732
rect 43904 234048 43956 234054
rect 43904 233990 43956 233996
rect 43904 230580 43956 230586
rect 43904 230522 43956 230528
rect 43916 199510 43944 230522
rect 43904 199504 43956 199510
rect 43904 199446 43956 199452
rect 43904 171896 43956 171902
rect 43904 171838 43956 171844
rect 43812 27940 43864 27946
rect 43812 27882 43864 27888
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43916 3942 43944 171838
rect 44008 28014 44036 434726
rect 44180 402144 44232 402150
rect 44180 402086 44232 402092
rect 44192 294030 44220 402086
rect 44180 294024 44232 294030
rect 44180 293966 44232 293972
rect 44456 258120 44508 258126
rect 44456 258062 44508 258068
rect 44088 234864 44140 234870
rect 44088 234806 44140 234812
rect 44100 230790 44128 234806
rect 44088 230784 44140 230790
rect 44088 230726 44140 230732
rect 44088 217388 44140 217394
rect 44088 217330 44140 217336
rect 44100 196926 44128 217330
rect 44088 196920 44140 196926
rect 44088 196862 44140 196868
rect 43996 28008 44048 28014
rect 43996 27950 44048 27956
rect 44468 27334 44496 258062
rect 44560 198082 44588 556174
rect 44652 488238 44680 589766
rect 44732 589756 44784 589762
rect 44732 589698 44784 589704
rect 44640 488232 44692 488238
rect 44640 488174 44692 488180
rect 44744 478718 44772 589698
rect 44916 589348 44968 589354
rect 44916 589290 44968 589296
rect 44824 587104 44876 587110
rect 44824 587046 44876 587052
rect 44732 478712 44784 478718
rect 44732 478654 44784 478660
rect 44640 323536 44692 323542
rect 44640 323478 44692 323484
rect 44652 245478 44680 323478
rect 44730 321600 44786 321609
rect 44730 321535 44786 321544
rect 44640 245472 44692 245478
rect 44640 245414 44692 245420
rect 44640 245336 44692 245342
rect 44640 245278 44692 245284
rect 44652 210594 44680 245278
rect 44744 241505 44772 321535
rect 44836 281722 44864 587046
rect 44928 509318 44956 589290
rect 45008 563100 45060 563106
rect 45008 563042 45060 563048
rect 44916 509312 44968 509318
rect 44916 509254 44968 509260
rect 44916 508360 44968 508366
rect 44916 508302 44968 508308
rect 44928 322930 44956 508302
rect 45020 381002 45048 563042
rect 45112 474706 45140 590038
rect 45192 564052 45244 564058
rect 45192 563994 45244 564000
rect 45100 474700 45152 474706
rect 45100 474642 45152 474648
rect 45008 380996 45060 381002
rect 45008 380938 45060 380944
rect 45006 373008 45062 373017
rect 45006 372943 45062 372952
rect 44916 322924 44968 322930
rect 44916 322866 44968 322872
rect 44914 283248 44970 283257
rect 44914 283183 44970 283192
rect 44824 281716 44876 281722
rect 44824 281658 44876 281664
rect 44824 253700 44876 253706
rect 44824 253642 44876 253648
rect 44836 245546 44864 253642
rect 44824 245540 44876 245546
rect 44824 245482 44876 245488
rect 44822 242992 44878 243001
rect 44822 242927 44878 242936
rect 44730 241496 44786 241505
rect 44730 241431 44786 241440
rect 44640 210588 44692 210594
rect 44640 210530 44692 210536
rect 44732 210452 44784 210458
rect 44732 210394 44784 210400
rect 44548 198076 44600 198082
rect 44548 198018 44600 198024
rect 44640 192772 44692 192778
rect 44640 192714 44692 192720
rect 44652 108934 44680 192714
rect 44744 152833 44772 210394
rect 44836 182850 44864 242927
rect 44928 198014 44956 283183
rect 45020 199714 45048 372943
rect 45098 359408 45154 359417
rect 45098 359343 45154 359352
rect 45008 199708 45060 199714
rect 45008 199650 45060 199656
rect 44916 198008 44968 198014
rect 44916 197950 44968 197956
rect 44916 187196 44968 187202
rect 44916 187138 44968 187144
rect 44824 182844 44876 182850
rect 44824 182786 44876 182792
rect 44824 176656 44876 176662
rect 44824 176598 44876 176604
rect 44730 152824 44786 152833
rect 44730 152759 44786 152768
rect 44732 151428 44784 151434
rect 44732 151370 44784 151376
rect 44640 108928 44692 108934
rect 44640 108870 44692 108876
rect 44456 27328 44508 27334
rect 44456 27270 44508 27276
rect 44744 20126 44772 151370
rect 44836 24274 44864 176598
rect 44928 31113 44956 187138
rect 45008 178764 45060 178770
rect 45008 178706 45060 178712
rect 44914 31104 44970 31113
rect 44914 31039 44970 31048
rect 44824 24268 44876 24274
rect 44824 24210 44876 24216
rect 44732 20120 44784 20126
rect 44732 20062 44784 20068
rect 43904 3936 43956 3942
rect 43904 3878 43956 3884
rect 45020 3806 45048 178706
rect 45112 69698 45140 359343
rect 45204 264761 45232 563994
rect 45296 361554 45324 590106
rect 47584 589620 47636 589626
rect 47584 589562 47636 589568
rect 47032 587580 47084 587586
rect 47032 587522 47084 587528
rect 46664 581732 46716 581738
rect 46664 581674 46716 581680
rect 46388 578944 46440 578950
rect 46388 578886 46440 578892
rect 45376 573640 45428 573646
rect 45376 573582 45428 573588
rect 45284 361548 45336 361554
rect 45284 361490 45336 361496
rect 45282 339552 45338 339561
rect 45282 339487 45338 339496
rect 45190 264752 45246 264761
rect 45190 264687 45246 264696
rect 45190 237416 45246 237425
rect 45190 237351 45246 237360
rect 45100 69692 45152 69698
rect 45100 69634 45152 69640
rect 45204 27198 45232 237351
rect 45296 29646 45324 339487
rect 45388 251841 45416 573582
rect 46204 570852 46256 570858
rect 46204 570794 46256 570800
rect 45836 562080 45888 562086
rect 46020 562080 46072 562086
rect 45888 562040 46020 562068
rect 45836 562022 45888 562028
rect 46020 562022 46072 562028
rect 45744 559972 45796 559978
rect 45744 559914 45796 559920
rect 45756 521801 45784 559914
rect 46110 556608 46166 556617
rect 46110 556543 46166 556552
rect 46124 556238 46152 556543
rect 46112 556232 46164 556238
rect 45926 556200 45982 556209
rect 46112 556174 46164 556180
rect 45926 556135 45982 556144
rect 45742 521792 45798 521801
rect 45742 521727 45798 521736
rect 45650 520704 45706 520713
rect 45650 520639 45706 520648
rect 45558 520432 45614 520441
rect 45558 520367 45560 520376
rect 45612 520367 45614 520376
rect 45560 520338 45612 520344
rect 45664 520334 45692 520639
rect 45652 520328 45704 520334
rect 45652 520270 45704 520276
rect 45836 519580 45888 519586
rect 45836 519522 45888 519528
rect 45558 516624 45614 516633
rect 45558 516559 45614 516568
rect 45572 516186 45600 516559
rect 45560 516180 45612 516186
rect 45560 516122 45612 516128
rect 45558 515264 45614 515273
rect 45558 515199 45614 515208
rect 45572 514826 45600 515199
rect 45560 514820 45612 514826
rect 45560 514762 45612 514768
rect 45848 514078 45876 519522
rect 45836 514072 45888 514078
rect 45836 514014 45888 514020
rect 45836 502104 45888 502110
rect 45836 502046 45888 502052
rect 45848 501401 45876 502046
rect 45834 501392 45890 501401
rect 45834 501327 45890 501336
rect 45836 498160 45888 498166
rect 45836 498102 45888 498108
rect 45848 497321 45876 498102
rect 45834 497312 45890 497321
rect 45834 497247 45890 497256
rect 45836 480480 45888 480486
rect 45836 480422 45888 480428
rect 45650 463856 45706 463865
rect 45650 463791 45706 463800
rect 45664 463758 45692 463791
rect 45652 463752 45704 463758
rect 45652 463694 45704 463700
rect 45650 425232 45706 425241
rect 45650 425167 45706 425176
rect 45664 425134 45692 425167
rect 45652 425128 45704 425134
rect 45652 425070 45704 425076
rect 45650 421016 45706 421025
rect 45650 420951 45652 420960
rect 45704 420951 45706 420960
rect 45652 420922 45704 420928
rect 45650 419656 45706 419665
rect 45650 419591 45652 419600
rect 45704 419591 45706 419600
rect 45652 419562 45704 419568
rect 45650 415576 45706 415585
rect 45650 415511 45652 415520
rect 45704 415511 45706 415520
rect 45652 415482 45704 415488
rect 45652 371204 45704 371210
rect 45652 371146 45704 371152
rect 45664 284714 45692 371146
rect 45744 322924 45796 322930
rect 45744 322866 45796 322872
rect 45652 284708 45704 284714
rect 45652 284650 45704 284656
rect 45650 281616 45706 281625
rect 45650 281551 45652 281560
rect 45704 281551 45706 281560
rect 45652 281522 45704 281528
rect 45560 269816 45612 269822
rect 45560 269758 45612 269764
rect 45572 268002 45600 269758
rect 45480 267974 45600 268002
rect 45480 267730 45508 267974
rect 45480 267702 45692 267730
rect 45468 266416 45520 266422
rect 45468 266358 45520 266364
rect 45480 256766 45508 266358
rect 45664 257378 45692 267702
rect 45652 257372 45704 257378
rect 45652 257314 45704 257320
rect 45468 256760 45520 256766
rect 45468 256702 45520 256708
rect 45374 251832 45430 251841
rect 45374 251767 45430 251776
rect 45560 247716 45612 247722
rect 45560 247658 45612 247664
rect 45468 245608 45520 245614
rect 45468 245550 45520 245556
rect 45480 233442 45508 245550
rect 45572 245154 45600 247658
rect 45652 245472 45704 245478
rect 45652 245414 45704 245420
rect 45664 245274 45692 245414
rect 45756 245342 45784 322866
rect 45744 245336 45796 245342
rect 45744 245278 45796 245284
rect 45652 245268 45704 245274
rect 45652 245210 45704 245216
rect 45572 245126 45784 245154
rect 45652 245064 45704 245070
rect 45652 245006 45704 245012
rect 45468 233436 45520 233442
rect 45468 233378 45520 233384
rect 45558 232248 45614 232257
rect 45558 232183 45614 232192
rect 45572 231878 45600 232183
rect 45560 231872 45612 231878
rect 45560 231814 45612 231820
rect 45558 230616 45614 230625
rect 45558 230551 45614 230560
rect 45572 230518 45600 230551
rect 45560 230512 45612 230518
rect 45560 230454 45612 230460
rect 45558 227896 45614 227905
rect 45558 227831 45614 227840
rect 45572 227798 45600 227831
rect 45560 227792 45612 227798
rect 45560 227734 45612 227740
rect 45466 214024 45522 214033
rect 45466 213959 45522 213968
rect 45284 29640 45336 29646
rect 45284 29582 45336 29588
rect 45480 28762 45508 213959
rect 45558 211304 45614 211313
rect 45558 211239 45614 211248
rect 45572 211206 45600 211239
rect 45560 211200 45612 211206
rect 45560 211142 45612 211148
rect 45664 210458 45692 245006
rect 45756 238066 45784 245126
rect 45744 238060 45796 238066
rect 45744 238002 45796 238008
rect 45744 233436 45796 233442
rect 45744 233378 45796 233384
rect 45756 217394 45784 233378
rect 45848 219502 45876 480422
rect 45940 430001 45968 556135
rect 46110 551304 46166 551313
rect 46110 551239 46166 551248
rect 46124 551206 46152 551239
rect 46112 551200 46164 551206
rect 46112 551142 46164 551148
rect 46110 550896 46166 550905
rect 46110 550831 46112 550840
rect 46164 550831 46166 550840
rect 46112 550802 46164 550808
rect 46110 549808 46166 549817
rect 46110 549743 46166 549752
rect 46124 549302 46152 549743
rect 46112 549296 46164 549302
rect 46112 549238 46164 549244
rect 46110 548312 46166 548321
rect 46110 548247 46166 548256
rect 46124 547942 46152 548247
rect 46112 547936 46164 547942
rect 46112 547878 46164 547884
rect 46112 546032 46164 546038
rect 46112 545974 46164 545980
rect 46124 544241 46152 545974
rect 46110 544232 46166 544241
rect 46110 544167 46166 544176
rect 46110 529000 46166 529009
rect 46110 528935 46166 528944
rect 46124 528630 46152 528935
rect 46112 528624 46164 528630
rect 46112 528566 46164 528572
rect 46020 524476 46072 524482
rect 46020 524418 46072 524424
rect 46032 519586 46060 524418
rect 46020 519580 46072 519586
rect 46020 519522 46072 519528
rect 46216 514570 46244 570794
rect 46296 567860 46348 567866
rect 46296 567802 46348 567808
rect 46308 526561 46336 567802
rect 46294 526552 46350 526561
rect 46294 526487 46350 526496
rect 46296 521552 46348 521558
rect 46296 521494 46348 521500
rect 46032 514542 46244 514570
rect 46032 510921 46060 514542
rect 46112 514072 46164 514078
rect 46112 514014 46164 514020
rect 46018 510912 46074 510921
rect 46018 510847 46074 510856
rect 46020 497072 46072 497078
rect 46020 497014 46072 497020
rect 46032 494601 46060 497014
rect 46018 494592 46074 494601
rect 46018 494527 46074 494536
rect 46124 474201 46152 514014
rect 46202 513904 46258 513913
rect 46202 513839 46258 513848
rect 46216 513398 46244 513839
rect 46204 513392 46256 513398
rect 46204 513334 46256 513340
rect 46204 509312 46256 509318
rect 46204 509254 46256 509260
rect 46110 474192 46166 474201
rect 46110 474127 46166 474136
rect 46018 439648 46074 439657
rect 46018 439583 46074 439592
rect 46032 438938 46060 439583
rect 46020 438932 46072 438938
rect 46020 438874 46072 438880
rect 45926 429992 45982 430001
rect 45926 429927 45982 429936
rect 45926 420064 45982 420073
rect 45926 419999 45982 420008
rect 45940 419558 45968 419999
rect 45928 419552 45980 419558
rect 45928 419494 45980 419500
rect 45926 418704 45982 418713
rect 45926 418639 45982 418648
rect 45940 418198 45968 418639
rect 45928 418192 45980 418198
rect 45928 418134 45980 418140
rect 45926 415984 45982 415993
rect 45926 415919 45982 415928
rect 45940 415478 45968 415919
rect 45928 415472 45980 415478
rect 45928 415414 45980 415420
rect 46110 392728 46166 392737
rect 46110 392663 46166 392672
rect 46018 392184 46074 392193
rect 46018 392119 46074 392128
rect 46032 392086 46060 392119
rect 46020 392080 46072 392086
rect 46020 392022 46072 392028
rect 46124 392018 46152 392663
rect 46112 392012 46164 392018
rect 46112 391954 46164 391960
rect 46112 386368 46164 386374
rect 46112 386310 46164 386316
rect 46124 385801 46152 386310
rect 46110 385792 46166 385801
rect 46110 385727 46166 385736
rect 46020 367056 46072 367062
rect 46020 366998 46072 367004
rect 46032 366081 46060 366998
rect 46018 366072 46074 366081
rect 46018 366007 46074 366016
rect 46110 310992 46166 311001
rect 46110 310927 46166 310936
rect 46124 310554 46152 310927
rect 46112 310548 46164 310554
rect 46112 310490 46164 310496
rect 46110 309224 46166 309233
rect 46110 309159 46112 309168
rect 46164 309159 46166 309168
rect 46112 309130 46164 309136
rect 46112 293956 46164 293962
rect 46112 293898 46164 293904
rect 46124 292641 46152 293898
rect 46110 292632 46166 292641
rect 46110 292567 46166 292576
rect 46018 258360 46074 258369
rect 46018 258295 46074 258304
rect 46032 258126 46060 258295
rect 46020 258120 46072 258126
rect 46020 258062 46072 258068
rect 46020 256760 46072 256766
rect 46020 256702 46072 256708
rect 46032 245614 46060 256702
rect 46020 245608 46072 245614
rect 46020 245550 46072 245556
rect 45928 245540 45980 245546
rect 45928 245482 45980 245488
rect 45940 234870 45968 245482
rect 45928 234864 45980 234870
rect 45928 234806 45980 234812
rect 45928 234048 45980 234054
rect 45928 233990 45980 233996
rect 45940 233481 45968 233990
rect 45926 233472 45982 233481
rect 45926 233407 45982 233416
rect 46018 230888 46074 230897
rect 46018 230823 46074 230832
rect 46032 230586 46060 230823
rect 46020 230580 46072 230586
rect 46020 230522 46072 230528
rect 45928 221468 45980 221474
rect 45928 221410 45980 221416
rect 45836 219496 45888 219502
rect 45836 219438 45888 219444
rect 45744 217388 45796 217394
rect 45744 217330 45796 217336
rect 45940 215294 45968 221410
rect 46110 218648 46166 218657
rect 46020 218612 46072 218618
rect 46110 218583 46166 218592
rect 46020 218554 46072 218560
rect 45756 215266 45968 215294
rect 45652 210452 45704 210458
rect 45652 210394 45704 210400
rect 45560 208344 45612 208350
rect 45560 208286 45612 208292
rect 45572 207641 45600 208286
rect 45558 207632 45614 207641
rect 45558 207567 45614 207576
rect 45756 207482 45784 215266
rect 45834 212664 45890 212673
rect 45834 212599 45890 212608
rect 45572 207454 45784 207482
rect 45572 178498 45600 207454
rect 45652 206984 45704 206990
rect 45650 206952 45652 206961
rect 45704 206952 45706 206961
rect 45650 206887 45706 206896
rect 45650 206000 45706 206009
rect 45650 205935 45706 205944
rect 45664 205698 45692 205935
rect 45652 205692 45704 205698
rect 45652 205634 45704 205640
rect 45560 178492 45612 178498
rect 45560 178434 45612 178440
rect 45848 176662 45876 212599
rect 46032 205634 46060 218554
rect 46124 218074 46152 218583
rect 46112 218068 46164 218074
rect 46112 218010 46164 218016
rect 45940 205606 46060 205634
rect 45940 194886 45968 205606
rect 46216 198121 46244 509254
rect 46308 327078 46336 521494
rect 46400 497078 46428 578886
rect 46572 570920 46624 570926
rect 46572 570862 46624 570868
rect 46480 569356 46532 569362
rect 46480 569298 46532 569304
rect 46388 497072 46440 497078
rect 46388 497014 46440 497020
rect 46386 496088 46442 496097
rect 46386 496023 46442 496032
rect 46400 495514 46428 496023
rect 46388 495508 46440 495514
rect 46388 495450 46440 495456
rect 46386 489968 46442 489977
rect 46386 489903 46388 489912
rect 46440 489903 46442 489912
rect 46388 489874 46440 489880
rect 46388 488232 46440 488238
rect 46388 488174 46440 488180
rect 46296 327072 46348 327078
rect 46296 327014 46348 327020
rect 46296 323196 46348 323202
rect 46296 323138 46348 323144
rect 46308 318481 46336 323138
rect 46294 318472 46350 318481
rect 46294 318407 46350 318416
rect 46294 314800 46350 314809
rect 46294 314735 46350 314744
rect 46308 314702 46336 314735
rect 46296 314696 46348 314702
rect 46296 314638 46348 314644
rect 46296 310480 46348 310486
rect 46296 310422 46348 310428
rect 46308 310321 46336 310422
rect 46294 310312 46350 310321
rect 46294 310247 46350 310256
rect 46400 306374 46428 488174
rect 46492 482361 46520 569298
rect 46478 482352 46534 482361
rect 46478 482287 46534 482296
rect 46584 475561 46612 570862
rect 46676 480321 46704 581674
rect 46848 577584 46900 577590
rect 46848 577526 46900 577532
rect 46756 566636 46808 566642
rect 46756 566578 46808 566584
rect 46768 546038 46796 566578
rect 46756 546032 46808 546038
rect 46756 545974 46808 545980
rect 46754 545728 46810 545737
rect 46754 545663 46810 545672
rect 46768 545154 46796 545663
rect 46756 545148 46808 545154
rect 46756 545090 46808 545096
rect 46754 544368 46810 544377
rect 46754 544303 46810 544312
rect 46768 543794 46796 544303
rect 46756 543788 46808 543794
rect 46756 543730 46808 543736
rect 46754 541104 46810 541113
rect 46754 541039 46810 541048
rect 46768 541006 46796 541039
rect 46756 541000 46808 541006
rect 46756 540942 46808 540948
rect 46756 538212 46808 538218
rect 46756 538154 46808 538160
rect 46768 538121 46796 538154
rect 46754 538112 46810 538121
rect 46754 538047 46810 538056
rect 46754 533352 46810 533361
rect 46754 533287 46810 533296
rect 46768 532778 46796 533287
rect 46756 532772 46808 532778
rect 46756 532714 46808 532720
rect 46754 532128 46810 532137
rect 46754 532063 46810 532072
rect 46768 531350 46796 532063
rect 46756 531344 46808 531350
rect 46756 531286 46808 531292
rect 46756 529984 46808 529990
rect 46754 529952 46756 529961
rect 46808 529952 46810 529961
rect 46754 529887 46810 529896
rect 46756 525768 46808 525774
rect 46756 525710 46808 525716
rect 46768 525201 46796 525710
rect 46754 525192 46810 525201
rect 46754 525127 46810 525136
rect 46756 510604 46808 510610
rect 46756 510546 46808 510552
rect 46768 509561 46796 510546
rect 46754 509552 46810 509561
rect 46754 509487 46810 509496
rect 46754 505200 46810 505209
rect 46754 505135 46756 505144
rect 46808 505135 46810 505144
rect 46756 505106 46808 505112
rect 46756 500948 46808 500954
rect 46756 500890 46808 500896
rect 46768 500721 46796 500890
rect 46754 500712 46810 500721
rect 46754 500647 46810 500656
rect 46756 496800 46808 496806
rect 46756 496742 46808 496748
rect 46768 495961 46796 496742
rect 46754 495952 46810 495961
rect 46754 495887 46810 495896
rect 46756 495440 46808 495446
rect 46756 495382 46808 495388
rect 46768 495281 46796 495382
rect 46754 495272 46810 495281
rect 46754 495207 46810 495216
rect 46754 493232 46810 493241
rect 46754 493167 46810 493176
rect 46768 492726 46796 493167
rect 46756 492720 46808 492726
rect 46756 492662 46808 492668
rect 46754 490648 46810 490657
rect 46754 490583 46810 490592
rect 46768 490006 46796 490583
rect 46756 490000 46808 490006
rect 46756 489942 46808 489948
rect 46756 489864 46808 489870
rect 46754 489832 46756 489841
rect 46808 489832 46810 489841
rect 46754 489767 46810 489776
rect 46754 485888 46810 485897
rect 46754 485823 46756 485832
rect 46808 485823 46810 485832
rect 46756 485794 46808 485800
rect 46754 484800 46810 484809
rect 46754 484735 46810 484744
rect 46768 484430 46796 484735
rect 46756 484424 46808 484430
rect 46756 484366 46808 484372
rect 46754 483440 46810 483449
rect 46754 483375 46810 483384
rect 46768 483070 46796 483375
rect 46756 483064 46808 483070
rect 46756 483006 46808 483012
rect 46662 480312 46718 480321
rect 46662 480247 46718 480256
rect 46664 478712 46716 478718
rect 46664 478654 46716 478660
rect 46570 475552 46626 475561
rect 46570 475487 46626 475496
rect 46480 474700 46532 474706
rect 46480 474642 46532 474648
rect 46492 390561 46520 474642
rect 46572 474632 46624 474638
rect 46572 474574 46624 474580
rect 46584 473521 46612 474574
rect 46570 473512 46626 473521
rect 46570 473447 46626 473456
rect 46570 468344 46626 468353
rect 46570 468279 46626 468288
rect 46584 467906 46612 468279
rect 46572 467900 46624 467906
rect 46572 467842 46624 467848
rect 46572 460896 46624 460902
rect 46572 460838 46624 460844
rect 46584 459921 46612 460838
rect 46570 459912 46626 459921
rect 46570 459847 46626 459856
rect 46676 442921 46704 478654
rect 46754 476504 46810 476513
rect 46754 476439 46810 476448
rect 46768 476134 46796 476439
rect 46756 476128 46808 476134
rect 46756 476070 46808 476076
rect 46754 469704 46810 469713
rect 46754 469639 46810 469648
rect 46768 469266 46796 469639
rect 46756 469260 46808 469266
rect 46756 469202 46808 469208
rect 46754 468072 46810 468081
rect 46754 468007 46810 468016
rect 46768 467974 46796 468007
rect 46756 467968 46808 467974
rect 46756 467910 46808 467916
rect 46754 464264 46810 464273
rect 46754 464199 46810 464208
rect 46768 464166 46796 464199
rect 46756 464160 46808 464166
rect 46756 464102 46808 464108
rect 46756 463684 46808 463690
rect 46756 463626 46808 463632
rect 46768 463321 46796 463626
rect 46754 463312 46810 463321
rect 46754 463247 46810 463256
rect 46754 461000 46810 461009
rect 46754 460935 46756 460944
rect 46808 460935 46810 460944
rect 46756 460906 46808 460912
rect 46754 458280 46810 458289
rect 46754 458215 46756 458224
rect 46808 458215 46810 458224
rect 46756 458186 46808 458192
rect 46756 456748 46808 456754
rect 46756 456690 46808 456696
rect 46768 456521 46796 456690
rect 46754 456512 46810 456521
rect 46754 456447 46810 456456
rect 46756 451240 46808 451246
rect 46756 451182 46808 451188
rect 46768 450401 46796 451182
rect 46754 450392 46810 450401
rect 46754 450327 46810 450336
rect 46754 445904 46810 445913
rect 46754 445839 46810 445848
rect 46768 445806 46796 445839
rect 46756 445800 46808 445806
rect 46756 445742 46808 445748
rect 46754 445088 46810 445097
rect 46754 445023 46810 445032
rect 46768 444446 46796 445023
rect 46756 444440 46808 444446
rect 46756 444382 46808 444388
rect 46754 443320 46810 443329
rect 46754 443255 46810 443264
rect 46768 443018 46796 443255
rect 46756 443012 46808 443018
rect 46756 442954 46808 442960
rect 46662 442912 46718 442921
rect 46662 442847 46718 442856
rect 46754 439104 46810 439113
rect 46754 439039 46810 439048
rect 46768 439006 46796 439039
rect 46756 439000 46808 439006
rect 46756 438942 46808 438948
rect 46754 436520 46810 436529
rect 46754 436455 46810 436464
rect 46768 436150 46796 436455
rect 46756 436144 46808 436150
rect 46756 436086 46808 436092
rect 46756 434784 46808 434790
rect 46754 434752 46756 434761
rect 46808 434752 46810 434761
rect 46754 434687 46810 434696
rect 46754 433664 46810 433673
rect 46754 433599 46810 433608
rect 46768 433362 46796 433599
rect 46756 433356 46808 433362
rect 46756 433298 46808 433304
rect 46754 432032 46810 432041
rect 46754 431967 46756 431976
rect 46808 431967 46810 431976
rect 46756 431938 46808 431944
rect 46662 428360 46718 428369
rect 46662 428295 46718 428304
rect 46676 427922 46704 428295
rect 46754 427952 46810 427961
rect 46664 427916 46716 427922
rect 46754 427887 46810 427896
rect 46664 427858 46716 427864
rect 46768 427854 46796 427887
rect 46756 427848 46808 427854
rect 46756 427790 46808 427796
rect 46662 425368 46718 425377
rect 46662 425303 46718 425312
rect 46570 421288 46626 421297
rect 46570 421223 46626 421232
rect 46478 390552 46534 390561
rect 46478 390487 46534 390496
rect 46478 389328 46534 389337
rect 46478 389263 46534 389272
rect 46492 389230 46520 389263
rect 46480 389224 46532 389230
rect 46480 389166 46532 389172
rect 46478 386472 46534 386481
rect 46478 386407 46480 386416
rect 46532 386407 46534 386416
rect 46480 386378 46532 386384
rect 46478 385112 46534 385121
rect 46478 385047 46480 385056
rect 46532 385047 46534 385056
rect 46480 385018 46532 385024
rect 46480 383648 46532 383654
rect 46480 383590 46532 383596
rect 46492 383081 46520 383590
rect 46478 383072 46534 383081
rect 46478 383007 46534 383016
rect 46480 381132 46532 381138
rect 46480 381074 46532 381080
rect 46492 376281 46520 381074
rect 46478 376272 46534 376281
rect 46478 376207 46534 376216
rect 46480 361548 46532 361554
rect 46480 361490 46532 361496
rect 46492 357814 46520 361490
rect 46480 357808 46532 357814
rect 46480 357750 46532 357756
rect 46478 354784 46534 354793
rect 46478 354719 46480 354728
rect 46532 354719 46534 354728
rect 46480 354690 46532 354696
rect 46480 353252 46532 353258
rect 46480 353194 46532 353200
rect 46492 353161 46520 353194
rect 46478 353152 46534 353161
rect 46478 353087 46534 353096
rect 46478 349208 46534 349217
rect 46478 349143 46480 349152
rect 46532 349143 46534 349152
rect 46480 349114 46532 349120
rect 46478 347168 46534 347177
rect 46478 347103 46534 347112
rect 46492 346458 46520 347103
rect 46480 346452 46532 346458
rect 46480 346394 46532 346400
rect 46478 345128 46534 345137
rect 46478 345063 46480 345072
rect 46532 345063 46534 345072
rect 46480 345034 46532 345040
rect 46478 336832 46534 336841
rect 46478 336767 46480 336776
rect 46532 336767 46534 336776
rect 46480 336738 46532 336744
rect 46480 331220 46532 331226
rect 46480 331162 46532 331168
rect 46492 330721 46520 331162
rect 46478 330712 46534 330721
rect 46478 330647 46534 330656
rect 46478 328944 46534 328953
rect 46478 328879 46534 328888
rect 46492 328506 46520 328879
rect 46480 328500 46532 328506
rect 46480 328442 46532 328448
rect 46480 325644 46532 325650
rect 46480 325586 46532 325592
rect 46492 325281 46520 325586
rect 46478 325272 46534 325281
rect 46478 325207 46534 325216
rect 46480 321564 46532 321570
rect 46480 321506 46532 321512
rect 46308 306346 46428 306374
rect 46308 302297 46336 306346
rect 46386 302968 46442 302977
rect 46386 302903 46442 302912
rect 46294 302288 46350 302297
rect 46400 302258 46428 302903
rect 46294 302223 46350 302232
rect 46388 302252 46440 302258
rect 46388 302194 46440 302200
rect 46296 302184 46348 302190
rect 46296 302126 46348 302132
rect 46308 226681 46336 302126
rect 46386 300928 46442 300937
rect 46386 300863 46388 300872
rect 46440 300863 46442 300872
rect 46388 300834 46440 300840
rect 46386 298208 46442 298217
rect 46386 298143 46388 298152
rect 46440 298143 46442 298152
rect 46388 298114 46440 298120
rect 46386 297120 46442 297129
rect 46386 297055 46442 297064
rect 46400 296750 46428 297055
rect 46388 296744 46440 296750
rect 46388 296686 46440 296692
rect 46386 292904 46442 292913
rect 46386 292839 46442 292848
rect 46400 292602 46428 292839
rect 46388 292596 46440 292602
rect 46388 292538 46440 292544
rect 46386 291544 46442 291553
rect 46386 291479 46442 291488
rect 46400 291242 46428 291479
rect 46388 291236 46440 291242
rect 46388 291178 46440 291184
rect 46386 285832 46442 285841
rect 46386 285767 46442 285776
rect 46400 285734 46428 285767
rect 46388 285728 46440 285734
rect 46388 285670 46440 285676
rect 46492 276078 46520 321506
rect 46480 276072 46532 276078
rect 46480 276014 46532 276020
rect 46480 274712 46532 274718
rect 46480 274654 46532 274660
rect 46492 272610 46520 274654
rect 46480 272604 46532 272610
rect 46480 272546 46532 272552
rect 46478 268288 46534 268297
rect 46478 268223 46534 268232
rect 46386 267880 46442 267889
rect 46386 267815 46388 267824
rect 46440 267815 46442 267824
rect 46388 267786 46440 267792
rect 46492 267782 46520 268223
rect 46480 267776 46532 267782
rect 46480 267718 46532 267724
rect 46478 256728 46534 256737
rect 46478 256663 46534 256672
rect 46386 236056 46442 236065
rect 46386 235991 46442 236000
rect 46400 229770 46428 235991
rect 46388 229764 46440 229770
rect 46388 229706 46440 229712
rect 46294 226672 46350 226681
rect 46294 226607 46350 226616
rect 46386 224904 46442 224913
rect 46386 224839 46442 224848
rect 46294 217288 46350 217297
rect 46294 217223 46350 217232
rect 46308 216782 46336 217223
rect 46296 216776 46348 216782
rect 46296 216718 46348 216724
rect 46296 209092 46348 209098
rect 46296 209034 46348 209040
rect 46308 205634 46336 209034
rect 46400 208350 46428 224839
rect 46388 208344 46440 208350
rect 46388 208286 46440 208292
rect 46308 205606 46428 205634
rect 46400 205578 46428 205606
rect 46308 205550 46428 205578
rect 46202 198112 46258 198121
rect 46202 198047 46258 198056
rect 45928 194880 45980 194886
rect 45928 194822 45980 194828
rect 46308 192302 46336 205550
rect 46386 202872 46442 202881
rect 46386 202807 46388 202816
rect 46440 202807 46442 202816
rect 46388 202778 46440 202784
rect 46386 201648 46442 201657
rect 46386 201583 46442 201592
rect 46296 192296 46348 192302
rect 46296 192238 46348 192244
rect 46020 185632 46072 185638
rect 46020 185574 46072 185580
rect 45836 176656 45888 176662
rect 45836 176598 45888 176604
rect 45928 151224 45980 151230
rect 45928 151166 45980 151172
rect 45940 142154 45968 151166
rect 46032 150521 46060 185574
rect 46112 180260 46164 180266
rect 46112 180202 46164 180208
rect 46018 150512 46074 150521
rect 46018 150447 46074 150456
rect 45940 142126 46060 142154
rect 46032 100065 46060 142126
rect 46018 100056 46074 100065
rect 46018 99991 46074 100000
rect 46124 97986 46152 180202
rect 46204 177336 46256 177342
rect 46204 177278 46256 177284
rect 46112 97980 46164 97986
rect 46112 97922 46164 97928
rect 46216 64802 46244 177278
rect 46296 174616 46348 174622
rect 46296 174558 46348 174564
rect 46204 64796 46256 64802
rect 46204 64738 46256 64744
rect 46308 41410 46336 174558
rect 46400 155718 46428 201583
rect 46492 173194 46520 256663
rect 46584 244361 46612 421223
rect 46676 247081 46704 425303
rect 46754 423736 46810 423745
rect 46754 423671 46756 423680
rect 46808 423671 46810 423680
rect 46756 423642 46808 423648
rect 46754 414080 46810 414089
rect 46754 414015 46756 414024
rect 46808 414015 46810 414024
rect 46756 413986 46808 413992
rect 46754 411360 46810 411369
rect 46754 411295 46756 411304
rect 46808 411295 46810 411304
rect 46756 411266 46808 411272
rect 46754 407688 46810 407697
rect 46754 407623 46810 407632
rect 46768 407182 46796 407623
rect 46756 407176 46808 407182
rect 46756 407118 46808 407124
rect 46754 403608 46810 403617
rect 46754 403543 46810 403552
rect 46768 403034 46796 403543
rect 46756 403028 46808 403034
rect 46756 402970 46808 402976
rect 46754 400344 46810 400353
rect 46754 400279 46810 400288
rect 46768 400246 46796 400279
rect 46756 400240 46808 400246
rect 46756 400182 46808 400188
rect 46754 399528 46810 399537
rect 46754 399463 46810 399472
rect 46768 398886 46796 399463
rect 46756 398880 46808 398886
rect 46756 398822 46808 398828
rect 46754 394768 46810 394777
rect 46754 394703 46756 394712
rect 46808 394703 46810 394712
rect 46756 394674 46808 394680
rect 46754 393544 46810 393553
rect 46754 393479 46810 393488
rect 46662 247072 46718 247081
rect 46662 247007 46718 247016
rect 46570 244352 46626 244361
rect 46570 244287 46626 244296
rect 46664 238740 46716 238746
rect 46664 238682 46716 238688
rect 46676 238241 46704 238682
rect 46662 238232 46718 238241
rect 46662 238167 46718 238176
rect 46662 234696 46718 234705
rect 46662 234631 46664 234640
rect 46716 234631 46718 234640
rect 46664 234602 46716 234608
rect 46572 229764 46624 229770
rect 46572 229706 46624 229712
rect 46584 222154 46612 229706
rect 46662 224088 46718 224097
rect 46662 224023 46718 224032
rect 46676 223650 46704 224023
rect 46664 223644 46716 223650
rect 46664 223586 46716 223592
rect 46662 222456 46718 222465
rect 46662 222391 46718 222400
rect 46676 222222 46704 222391
rect 46664 222216 46716 222222
rect 46664 222158 46716 222164
rect 46572 222148 46624 222154
rect 46572 222090 46624 222096
rect 46570 221368 46626 221377
rect 46570 221303 46626 221312
rect 46584 200114 46612 221303
rect 46662 221096 46718 221105
rect 46662 221031 46718 221040
rect 46676 220862 46704 221031
rect 46664 220856 46716 220862
rect 46664 220798 46716 220804
rect 46662 218376 46718 218385
rect 46662 218311 46718 218320
rect 46676 218142 46704 218311
rect 46664 218136 46716 218142
rect 46664 218078 46716 218084
rect 46662 216744 46718 216753
rect 46662 216679 46664 216688
rect 46716 216679 46718 216688
rect 46664 216650 46716 216656
rect 46662 215384 46718 215393
rect 46662 215319 46664 215328
rect 46716 215319 46718 215328
rect 46664 215290 46716 215296
rect 46662 203688 46718 203697
rect 46662 203623 46718 203632
rect 46676 202910 46704 203623
rect 46664 202904 46716 202910
rect 46664 202846 46716 202852
rect 46768 200161 46796 393479
rect 46860 381138 46888 577526
rect 47044 438841 47072 587522
rect 47216 562556 47268 562562
rect 47216 562498 47268 562504
rect 47124 561604 47176 561610
rect 47124 561546 47176 561552
rect 47030 438832 47086 438841
rect 47030 438767 47086 438776
rect 46848 381132 46900 381138
rect 46848 381074 46900 381080
rect 46846 381032 46902 381041
rect 46846 380967 46902 380976
rect 46860 380934 46888 380967
rect 46848 380928 46900 380934
rect 46848 380870 46900 380876
rect 46846 379808 46902 379817
rect 46846 379743 46902 379752
rect 46860 379574 46888 379743
rect 46848 379568 46900 379574
rect 46848 379510 46900 379516
rect 46846 372736 46902 372745
rect 46846 372671 46902 372680
rect 46860 372638 46888 372671
rect 46848 372632 46900 372638
rect 46848 372574 46900 372580
rect 46846 371512 46902 371521
rect 46846 371447 46902 371456
rect 46860 371278 46888 371447
rect 46848 371272 46900 371278
rect 46848 371214 46900 371220
rect 46846 368928 46902 368937
rect 46846 368863 46902 368872
rect 46860 368558 46888 368863
rect 46848 368552 46900 368558
rect 46848 368494 46900 368500
rect 46846 367568 46902 367577
rect 46846 367503 46902 367512
rect 46860 367130 46888 367503
rect 46848 367124 46900 367130
rect 46848 367066 46900 367072
rect 46846 363488 46902 363497
rect 46846 363423 46902 363432
rect 46860 362982 46888 363423
rect 46848 362976 46900 362982
rect 46848 362918 46900 362924
rect 46848 358760 46900 358766
rect 46848 358702 46900 358708
rect 46860 357921 46888 358702
rect 46846 357912 46902 357921
rect 46846 357847 46902 357856
rect 46848 357808 46900 357814
rect 46848 357750 46900 357756
rect 46860 323202 46888 357750
rect 47030 335472 47086 335481
rect 47030 335407 47086 335416
rect 46940 327072 46992 327078
rect 46940 327014 46992 327020
rect 46848 323196 46900 323202
rect 46848 323138 46900 323144
rect 46846 323096 46902 323105
rect 46846 323031 46902 323040
rect 46860 322998 46888 323031
rect 46848 322992 46900 322998
rect 46848 322934 46900 322940
rect 46846 321736 46902 321745
rect 46846 321671 46902 321680
rect 46860 321638 46888 321671
rect 46848 321632 46900 321638
rect 46848 321574 46900 321580
rect 46846 320240 46902 320249
rect 46846 320175 46848 320184
rect 46900 320175 46902 320184
rect 46848 320146 46900 320152
rect 46846 319016 46902 319025
rect 46846 318951 46848 318960
rect 46900 318951 46902 318960
rect 46848 318922 46900 318928
rect 46952 316034 46980 327014
rect 46860 316006 46980 316034
rect 46860 282962 46888 316006
rect 46860 282934 46980 282962
rect 46846 281888 46902 281897
rect 46846 281823 46902 281832
rect 46860 281654 46888 281823
rect 46848 281648 46900 281654
rect 46848 281590 46900 281596
rect 46846 277808 46902 277817
rect 46846 277743 46902 277752
rect 46860 277438 46888 277743
rect 46848 277432 46900 277438
rect 46848 277374 46900 277380
rect 46846 273728 46902 273737
rect 46846 273663 46902 273672
rect 46860 273290 46888 273663
rect 46848 273284 46900 273290
rect 46848 273226 46900 273232
rect 46848 272604 46900 272610
rect 46848 272546 46900 272552
rect 46860 257242 46888 272546
rect 46952 266422 46980 282934
rect 46940 266416 46992 266422
rect 46940 266358 46992 266364
rect 46848 257236 46900 257242
rect 46848 257178 46900 257184
rect 46846 254008 46902 254017
rect 46846 253943 46848 253952
rect 46900 253943 46902 253952
rect 46848 253914 46900 253920
rect 46846 247480 46902 247489
rect 46846 247415 46902 247424
rect 46860 247110 46888 247415
rect 46848 247104 46900 247110
rect 46848 247046 46900 247052
rect 46846 245848 46902 245857
rect 46846 245783 46902 245792
rect 46754 200152 46810 200161
rect 46584 200086 46704 200114
rect 46754 200087 46810 200096
rect 46676 198830 46704 200086
rect 46664 198824 46716 198830
rect 46664 198766 46716 198772
rect 46756 195696 46808 195702
rect 46756 195638 46808 195644
rect 46572 183048 46624 183054
rect 46572 182990 46624 182996
rect 46480 173188 46532 173194
rect 46480 173130 46532 173136
rect 46478 155952 46534 155961
rect 46478 155887 46534 155896
rect 46388 155712 46440 155718
rect 46388 155654 46440 155660
rect 46388 151360 46440 151366
rect 46388 151302 46440 151308
rect 46296 41404 46348 41410
rect 46296 41346 46348 41352
rect 45468 28756 45520 28762
rect 45468 28698 45520 28704
rect 45192 27192 45244 27198
rect 45192 27134 45244 27140
rect 46400 17202 46428 151302
rect 46492 21826 46520 155887
rect 46584 31754 46612 182990
rect 46664 172032 46716 172038
rect 46664 171974 46716 171980
rect 46572 31748 46624 31754
rect 46572 31690 46624 31696
rect 46480 21820 46532 21826
rect 46480 21762 46532 21768
rect 46676 17610 46704 171974
rect 46768 28490 46796 195638
rect 46860 195265 46888 245783
rect 46940 230784 46992 230790
rect 46940 230726 46992 230732
rect 46952 210497 46980 230726
rect 46938 210488 46994 210497
rect 46938 210423 46994 210432
rect 46846 195256 46902 195265
rect 46846 195191 46902 195200
rect 46848 191480 46900 191486
rect 46848 191422 46900 191428
rect 46756 28484 46808 28490
rect 46756 28426 46808 28432
rect 46860 22642 46888 191422
rect 47044 40050 47072 335407
rect 47136 270201 47164 561546
rect 47228 298081 47256 562498
rect 47308 562420 47360 562426
rect 47308 562362 47360 562368
rect 47320 328001 47348 562362
rect 47492 561468 47544 561474
rect 47492 561410 47544 561416
rect 47398 524648 47454 524657
rect 47398 524583 47454 524592
rect 47306 327992 47362 328001
rect 47306 327927 47362 327936
rect 47306 305008 47362 305017
rect 47306 304943 47362 304952
rect 47214 298072 47270 298081
rect 47214 298007 47270 298016
rect 47320 274718 47348 304943
rect 47412 282985 47440 524583
rect 47504 504121 47532 561410
rect 47596 524482 47624 589562
rect 47676 569424 47728 569430
rect 47676 569366 47728 569372
rect 47584 524476 47636 524482
rect 47584 524418 47636 524424
rect 47490 504112 47546 504121
rect 47490 504047 47546 504056
rect 47490 329896 47546 329905
rect 47490 329831 47546 329840
rect 47398 282976 47454 282985
rect 47398 282911 47454 282920
rect 47308 274712 47360 274718
rect 47308 274654 47360 274660
rect 47214 273320 47270 273329
rect 47214 273255 47270 273264
rect 47122 270192 47178 270201
rect 47122 270127 47178 270136
rect 47124 268388 47176 268394
rect 47124 268330 47176 268336
rect 47136 209681 47164 268330
rect 47122 209672 47178 209681
rect 47122 209607 47178 209616
rect 47032 40044 47084 40050
rect 47032 39986 47084 39992
rect 47228 29238 47256 273255
rect 47400 257236 47452 257242
rect 47400 257178 47452 257184
rect 47412 220833 47440 257178
rect 47398 220824 47454 220833
rect 47398 220759 47454 220768
rect 47400 208344 47452 208350
rect 47400 208286 47452 208292
rect 47306 201240 47362 201249
rect 47306 201175 47362 201184
rect 47216 29232 47268 29238
rect 47216 29174 47268 29180
rect 47320 22982 47348 201175
rect 47412 199073 47440 208286
rect 47504 199646 47532 329831
rect 47584 276072 47636 276078
rect 47584 276014 47636 276020
rect 47596 229809 47624 276014
rect 47688 257961 47716 569366
rect 48976 567194 49004 590242
rect 50080 590238 50108 590543
rect 50068 590232 50120 590238
rect 50068 590174 50120 590180
rect 55876 589694 55904 590543
rect 60384 590306 60412 590543
rect 60372 590300 60424 590306
rect 60372 590242 60424 590248
rect 69032 590034 69060 590543
rect 69020 590028 69072 590034
rect 69020 589970 69072 589976
rect 55864 589688 55916 589694
rect 55864 589630 55916 589636
rect 67638 589656 67694 589665
rect 67638 589591 67694 589600
rect 51078 589520 51134 589529
rect 51078 589455 51134 589464
rect 53838 589520 53894 589529
rect 53838 589455 53894 589464
rect 60646 589520 60702 589529
rect 60646 589455 60702 589464
rect 62210 589520 62266 589529
rect 62210 589455 62266 589464
rect 49056 576224 49108 576230
rect 49056 576166 49108 576172
rect 48884 567166 49004 567194
rect 47860 564664 47912 564670
rect 47860 564606 47912 564612
rect 47766 562320 47822 562329
rect 47766 562255 47822 562264
rect 47780 558929 47808 562255
rect 47766 558920 47822 558929
rect 47766 558855 47822 558864
rect 47674 257952 47730 257961
rect 47674 257887 47730 257896
rect 47582 229800 47638 229809
rect 47582 229735 47638 229744
rect 47584 222148 47636 222154
rect 47584 222090 47636 222096
rect 47492 199640 47544 199646
rect 47492 199582 47544 199588
rect 47398 199064 47454 199073
rect 47398 198999 47454 199008
rect 47596 82754 47624 222090
rect 47676 218748 47728 218754
rect 47676 218690 47728 218696
rect 47688 155922 47716 218690
rect 47768 210588 47820 210594
rect 47768 210530 47820 210536
rect 47780 200977 47808 210530
rect 47766 200968 47822 200977
rect 47766 200903 47822 200912
rect 47768 171964 47820 171970
rect 47768 171906 47820 171912
rect 47676 155916 47728 155922
rect 47676 155858 47728 155864
rect 47674 151464 47730 151473
rect 47674 151399 47730 151408
rect 47584 82748 47636 82754
rect 47584 82690 47636 82696
rect 47688 24546 47716 151399
rect 47676 24540 47728 24546
rect 47676 24482 47728 24488
rect 47780 24070 47808 171906
rect 47872 158098 47900 564606
rect 48228 562012 48280 562018
rect 48228 561954 48280 561960
rect 48240 559994 48268 561954
rect 48070 559966 48268 559994
rect 48884 559978 48912 567166
rect 48962 562592 49018 562601
rect 48962 562527 49018 562536
rect 48976 559994 49004 562527
rect 49068 562018 49096 576166
rect 51092 565146 51120 589455
rect 51170 589384 51226 589393
rect 51170 589319 51226 589328
rect 53746 589384 53802 589393
rect 53746 589319 53802 589328
rect 51080 565140 51132 565146
rect 51080 565082 51132 565088
rect 50344 562488 50396 562494
rect 50344 562430 50396 562436
rect 50356 562154 50384 562430
rect 50252 562148 50304 562154
rect 50252 562090 50304 562096
rect 50344 562148 50396 562154
rect 50344 562090 50396 562096
rect 49056 562012 49108 562018
rect 49056 561954 49108 561960
rect 50264 559994 50292 562090
rect 51184 561542 51212 589319
rect 52736 573368 52788 573374
rect 52736 573310 52788 573316
rect 51540 561876 51592 561882
rect 51540 561818 51592 561824
rect 52000 561876 52052 561882
rect 52000 561818 52052 561824
rect 51172 561536 51224 561542
rect 51172 561478 51224 561484
rect 51552 559994 51580 561818
rect 48872 559972 48924 559978
rect 48976 559966 49358 559994
rect 50264 559966 50600 559994
rect 51552 559966 51934 559994
rect 52012 559978 52040 561818
rect 52748 559994 52776 573310
rect 53760 566409 53788 589319
rect 53746 566400 53802 566409
rect 53746 566335 53802 566344
rect 52828 562012 52880 562018
rect 52828 561954 52880 561960
rect 52840 560046 52868 561954
rect 53852 561406 53880 589455
rect 56690 589384 56746 589393
rect 56690 589319 56746 589328
rect 57978 589384 58034 589393
rect 57978 589319 58034 589328
rect 53840 561400 53892 561406
rect 53840 561342 53892 561348
rect 56704 560969 56732 589319
rect 57992 576854 58020 589319
rect 57992 576826 58112 576854
rect 57978 562184 58034 562193
rect 57978 562119 58034 562128
rect 57426 562048 57482 562057
rect 57426 561983 57482 561992
rect 56690 560960 56746 560969
rect 56690 560895 56746 560904
rect 52000 559972 52052 559978
rect 48872 559914 48924 559920
rect 52578 559966 52776 559994
rect 52828 560040 52880 560046
rect 52828 559982 52880 559988
rect 57440 559994 57468 561983
rect 57992 559994 58020 562119
rect 58084 561270 58112 576826
rect 60660 570722 60688 589455
rect 60738 589384 60794 589393
rect 60738 589319 60794 589328
rect 62118 589384 62174 589393
rect 62118 589319 62174 589328
rect 60752 576854 60780 589319
rect 60752 576826 60872 576854
rect 60648 570716 60700 570722
rect 60648 570658 60700 570664
rect 58992 564664 59044 564670
rect 58992 564606 59044 564612
rect 59004 562494 59032 564606
rect 59818 564496 59874 564505
rect 59818 564431 59874 564440
rect 58992 562488 59044 562494
rect 58992 562430 59044 562436
rect 58530 562048 58586 562057
rect 58530 561983 58586 561992
rect 58072 561264 58124 561270
rect 58072 561206 58124 561212
rect 58544 560153 58572 561983
rect 58530 560144 58586 560153
rect 58530 560079 58586 560088
rect 59832 559994 59860 564431
rect 59910 561912 59966 561921
rect 59910 561847 59966 561856
rect 60738 561912 60794 561921
rect 60738 561847 60794 561856
rect 57440 559966 57730 559994
rect 57992 559966 58374 559994
rect 59662 559966 59860 559994
rect 59924 559994 59952 561847
rect 60752 561241 60780 561847
rect 60738 561232 60794 561241
rect 60738 561167 60794 561176
rect 60844 561134 60872 576826
rect 62132 561202 62160 589319
rect 62224 566506 62252 589455
rect 63498 589384 63554 589393
rect 63498 589319 63554 589328
rect 64786 589384 64842 589393
rect 64786 589319 64842 589328
rect 65430 589384 65486 589393
rect 65430 589319 65486 589328
rect 66258 589384 66314 589393
rect 66258 589319 66314 589328
rect 67546 589384 67602 589393
rect 67546 589319 67602 589328
rect 62212 566500 62264 566506
rect 62212 566442 62264 566448
rect 62488 564664 62540 564670
rect 62488 564606 62540 564612
rect 62120 561196 62172 561202
rect 62120 561138 62172 561144
rect 60832 561128 60884 561134
rect 60832 561070 60884 561076
rect 62500 559994 62528 564606
rect 63512 561105 63540 589319
rect 64800 566545 64828 589319
rect 65444 585818 65472 589319
rect 65432 585812 65484 585818
rect 65432 585754 65484 585760
rect 64786 566536 64842 566545
rect 64786 566471 64842 566480
rect 64788 565140 64840 565146
rect 64788 565082 64840 565088
rect 63498 561096 63554 561105
rect 63498 561031 63554 561040
rect 63222 560416 63278 560425
rect 63222 560351 63278 560360
rect 63236 559994 63264 560351
rect 64800 560266 64828 565082
rect 65708 562624 65760 562630
rect 65708 562566 65760 562572
rect 59924 559966 60260 559994
rect 62238 559966 62528 559994
rect 62882 559966 63264 559994
rect 64754 560238 64828 560266
rect 64754 559980 64782 560238
rect 65720 559994 65748 562566
rect 66272 561610 66300 589319
rect 67560 570654 67588 589319
rect 67548 570648 67600 570654
rect 67548 570590 67600 570596
rect 66260 561604 66312 561610
rect 66260 561546 66312 561552
rect 67652 560998 67680 589591
rect 72422 589520 72478 589529
rect 72422 589455 72478 589464
rect 74538 589520 74594 589529
rect 74538 589455 74594 589464
rect 67730 589384 67786 589393
rect 67730 589319 67786 589328
rect 70306 589384 70362 589393
rect 70306 589319 70362 589328
rect 71134 589384 71190 589393
rect 71134 589319 71190 589328
rect 71778 589384 71834 589393
rect 71778 589319 71834 589328
rect 67744 561338 67772 589319
rect 70320 562698 70348 589319
rect 71148 583001 71176 589319
rect 71134 582992 71190 583001
rect 71134 582927 71190 582936
rect 70308 562692 70360 562698
rect 70308 562634 70360 562640
rect 67732 561332 67784 561338
rect 67732 561274 67784 561280
rect 71792 561066 71820 589319
rect 72436 584497 72464 589455
rect 73158 589384 73214 589393
rect 73158 589319 73214 589328
rect 72422 584488 72478 584497
rect 72422 584423 72478 584432
rect 73172 561474 73200 589319
rect 74552 562562 74580 589455
rect 74828 588674 74856 590543
rect 75182 590472 75238 590481
rect 75182 590407 75238 590416
rect 77298 590472 77354 590481
rect 77298 590407 77354 590416
rect 75196 589801 75224 590407
rect 77312 590170 77340 590407
rect 77300 590164 77352 590170
rect 77300 590106 77352 590112
rect 75182 589792 75238 589801
rect 75182 589727 75238 589736
rect 75642 589384 75698 589393
rect 75642 589319 75698 589328
rect 75918 589384 75974 589393
rect 75918 589319 75974 589328
rect 74816 588668 74868 588674
rect 74816 588610 74868 588616
rect 75656 566710 75684 589319
rect 75736 584452 75788 584458
rect 75736 584394 75788 584400
rect 75748 576854 75776 584394
rect 75748 576826 75868 576854
rect 75644 566704 75696 566710
rect 75644 566646 75696 566652
rect 74540 562556 74592 562562
rect 74540 562498 74592 562504
rect 73160 561468 73212 561474
rect 73160 561410 73212 561416
rect 71780 561060 71832 561066
rect 71780 561002 71832 561008
rect 67640 560992 67692 560998
rect 67640 560934 67692 560940
rect 75840 559994 75868 576826
rect 75932 562426 75960 589319
rect 77864 588577 77892 590543
rect 78678 590472 78734 590481
rect 78678 590407 78734 590416
rect 78692 590102 78720 590407
rect 78680 590096 78732 590102
rect 78680 590038 78732 590044
rect 78678 589520 78734 589529
rect 78678 589455 78734 589464
rect 77850 588568 77906 588577
rect 77850 588503 77906 588512
rect 78692 587450 78720 589455
rect 78680 587444 78732 587450
rect 78680 587386 78732 587392
rect 77942 564632 77998 564641
rect 77942 564567 77998 564576
rect 76656 562556 76708 562562
rect 76656 562498 76708 562504
rect 75920 562420 75972 562426
rect 75920 562362 75972 562368
rect 76668 559994 76696 562498
rect 77956 559994 77984 564567
rect 78876 560266 78904 591330
rect 99930 590608 99986 590617
rect 99930 590543 99986 590552
rect 107566 590608 107622 590617
rect 107566 590543 107622 590552
rect 127346 590608 127402 590617
rect 127346 590543 127402 590552
rect 129738 590608 129794 590617
rect 129738 590543 129794 590552
rect 92478 590472 92534 590481
rect 92478 590407 92534 590416
rect 92492 589898 92520 590407
rect 92480 589892 92532 589898
rect 92480 589834 92532 589840
rect 81346 589520 81402 589529
rect 81346 589455 81402 589464
rect 82726 589520 82782 589529
rect 82726 589455 82782 589464
rect 84198 589520 84254 589529
rect 84198 589455 84254 589464
rect 88246 589520 88302 589529
rect 88246 589455 88302 589464
rect 89626 589520 89682 589529
rect 89626 589455 89682 589464
rect 91006 589520 91062 589529
rect 99944 589490 99972 590543
rect 104898 589520 104954 589529
rect 91006 589455 91062 589464
rect 99932 589484 99984 589490
rect 81360 576162 81388 589455
rect 81438 589384 81494 589393
rect 81438 589319 81494 589328
rect 82634 589384 82690 589393
rect 82634 589319 82690 589328
rect 81348 576156 81400 576162
rect 81348 576098 81400 576104
rect 81452 563786 81480 589319
rect 82648 577658 82676 589319
rect 82636 577652 82688 577658
rect 82636 577594 82688 577600
rect 82740 573442 82768 589455
rect 84106 589384 84162 589393
rect 84106 589319 84162 589328
rect 82728 573436 82780 573442
rect 82728 573378 82780 573384
rect 84120 570994 84148 589319
rect 84108 570988 84160 570994
rect 84108 570930 84160 570936
rect 84212 563854 84240 589455
rect 85578 589384 85634 589393
rect 85578 589319 85634 589328
rect 86958 589384 87014 589393
rect 86958 589319 87014 589328
rect 85486 566808 85542 566817
rect 85486 566743 85542 566752
rect 84200 563848 84252 563854
rect 83094 563816 83150 563825
rect 81440 563780 81492 563786
rect 84200 563790 84252 563796
rect 83094 563751 83150 563760
rect 81440 563722 81492 563728
rect 81624 562352 81676 562358
rect 81624 562294 81676 562300
rect 78876 560238 78950 560266
rect 65720 559966 66102 559994
rect 75762 559966 75868 559994
rect 76406 559966 76696 559994
rect 77694 559966 77984 559994
rect 78922 559980 78950 560238
rect 81636 559994 81664 562294
rect 83108 559994 83136 563751
rect 83740 562284 83792 562290
rect 83740 562226 83792 562232
rect 81558 559966 81664 559994
rect 82846 559966 83136 559994
rect 83752 559994 83780 562226
rect 85500 559994 85528 566743
rect 85592 563922 85620 589319
rect 86040 587444 86092 587450
rect 86040 587386 86092 587392
rect 86052 576854 86080 587386
rect 86052 576826 86172 576854
rect 85580 563916 85632 563922
rect 85580 563858 85632 563864
rect 86144 559994 86172 576826
rect 86972 563990 87000 589319
rect 88260 574870 88288 589455
rect 88248 574864 88300 574870
rect 88248 574806 88300 574812
rect 89640 566574 89668 589455
rect 89718 589384 89774 589393
rect 89718 589319 89774 589328
rect 90914 589384 90970 589393
rect 90914 589319 90970 589328
rect 89628 566568 89680 566574
rect 89628 566510 89680 566516
rect 87696 565208 87748 565214
rect 87696 565150 87748 565156
rect 86960 563984 87012 563990
rect 86960 563926 87012 563932
rect 86316 563576 86368 563582
rect 86316 563518 86368 563524
rect 83752 559966 84088 559994
rect 85422 559966 85528 559994
rect 86066 559966 86172 559994
rect 86328 559994 86356 563518
rect 87708 559994 87736 565150
rect 89732 564058 89760 589319
rect 90928 572121 90956 589319
rect 90914 572112 90970 572121
rect 90914 572047 90970 572056
rect 91020 570790 91048 589455
rect 107580 589490 107608 590543
rect 127360 589830 127388 590543
rect 127348 589824 127400 589830
rect 122562 589792 122618 589801
rect 127348 589766 127400 589772
rect 129752 589762 129780 590543
rect 122562 589727 122618 589736
rect 129740 589756 129792 589762
rect 104898 589455 104954 589464
rect 107568 589484 107620 589490
rect 99932 589426 99984 589432
rect 91098 589384 91154 589393
rect 91098 589319 91154 589328
rect 93766 589384 93822 589393
rect 93766 589319 93822 589328
rect 95146 589384 95202 589393
rect 95146 589319 95202 589328
rect 103426 589384 103482 589393
rect 103426 589319 103482 589328
rect 91008 570784 91060 570790
rect 91008 570726 91060 570732
rect 89720 564052 89772 564058
rect 89720 563994 89772 564000
rect 91112 563718 91140 589319
rect 93780 581670 93808 589319
rect 93768 581664 93820 581670
rect 93768 581606 93820 581612
rect 95160 573510 95188 589319
rect 100852 587512 100904 587518
rect 100852 587454 100904 587460
rect 100864 576854 100892 587454
rect 103440 583030 103468 589319
rect 104912 587042 104940 589455
rect 107568 589426 107620 589432
rect 110326 589384 110382 589393
rect 110326 589319 110382 589328
rect 113086 589384 113142 589393
rect 113086 589319 113142 589328
rect 115846 589384 115902 589393
rect 115846 589319 115902 589328
rect 117318 589384 117374 589393
rect 117318 589319 117374 589328
rect 119986 589384 120042 589393
rect 119986 589319 120042 589328
rect 104900 587036 104952 587042
rect 104900 586978 104952 586984
rect 103428 583024 103480 583030
rect 103428 582966 103480 582972
rect 100864 576826 100984 576854
rect 95148 573504 95200 573510
rect 95148 573446 95200 573452
rect 91100 563712 91152 563718
rect 91100 563654 91152 563660
rect 91284 562692 91336 562698
rect 91284 562634 91336 562640
rect 90824 562624 90876 562630
rect 90824 562566 90876 562572
rect 89718 562456 89774 562465
rect 89718 562391 89774 562400
rect 86328 559966 86710 559994
rect 87354 559966 87736 559994
rect 89732 559994 89760 562391
rect 90836 559994 90864 562566
rect 91296 559994 91324 562634
rect 94780 562216 94832 562222
rect 94780 562158 94832 562164
rect 89732 559966 89930 559994
rect 90574 559966 90864 559994
rect 91218 559966 91324 559994
rect 94792 559994 94820 562158
rect 99380 562148 99432 562154
rect 99380 562090 99432 562096
rect 99392 559994 99420 562090
rect 100956 559994 100984 576826
rect 109960 567316 110012 567322
rect 109960 567258 110012 567264
rect 109590 566128 109646 566137
rect 109590 566063 109646 566072
rect 106186 565992 106242 566001
rect 106186 565927 106242 565936
rect 104346 562320 104402 562329
rect 104346 562255 104402 562264
rect 94792 559966 95082 559994
rect 99392 559966 99590 559994
rect 100878 559966 100984 559994
rect 104360 559994 104388 562255
rect 105084 562080 105136 562086
rect 105084 562022 105136 562028
rect 105096 559994 105124 562022
rect 106200 559994 106228 565927
rect 108304 563780 108356 563786
rect 108304 563722 108356 563728
rect 108316 559994 108344 563722
rect 109604 559994 109632 566063
rect 109972 559994 110000 567258
rect 110340 565350 110368 589319
rect 113100 574938 113128 589319
rect 113088 574932 113140 574938
rect 113088 574874 113140 574880
rect 115860 569226 115888 589319
rect 117332 580514 117360 589319
rect 117320 580508 117372 580514
rect 117320 580450 117372 580456
rect 117320 580372 117372 580378
rect 117320 580314 117372 580320
rect 115848 569220 115900 569226
rect 115848 569162 115900 569168
rect 110328 565344 110380 565350
rect 110328 565286 110380 565292
rect 111892 565072 111944 565078
rect 111892 565014 111944 565020
rect 111904 559994 111932 565014
rect 113456 561944 113508 561950
rect 113456 561886 113508 561892
rect 104360 559966 104742 559994
rect 105096 559966 105386 559994
rect 106030 559966 106228 559994
rect 107962 559966 108344 559994
rect 109250 559966 109632 559994
rect 109894 559966 110000 559994
rect 111826 559966 111932 559994
rect 113468 559994 113496 561886
rect 116584 560584 116636 560590
rect 116584 560526 116636 560532
rect 116596 559994 116624 560526
rect 113468 559966 113758 559994
rect 116334 559966 116624 559994
rect 117332 559994 117360 580314
rect 120000 569294 120028 589319
rect 122576 587858 122604 589727
rect 129740 589698 129792 589704
rect 137282 589656 137338 589665
rect 137282 589591 137338 589600
rect 125506 589384 125562 589393
rect 125506 589319 125562 589328
rect 132498 589384 132554 589393
rect 132498 589319 132554 589328
rect 133878 589384 133934 589393
rect 133878 589319 133934 589328
rect 122564 587852 122616 587858
rect 122564 587794 122616 587800
rect 119988 569288 120040 569294
rect 119988 569230 120040 569236
rect 125520 566506 125548 589319
rect 132512 584458 132540 589319
rect 132500 584452 132552 584458
rect 132500 584394 132552 584400
rect 133892 569430 133920 589319
rect 137296 587110 137324 589591
rect 140686 589384 140742 589393
rect 140686 589319 140742 589328
rect 137284 587104 137336 587110
rect 137284 587046 137336 587052
rect 135628 581800 135680 581806
rect 135628 581742 135680 581748
rect 135640 576854 135668 581742
rect 140700 577726 140728 589319
rect 150440 585880 150492 585886
rect 150440 585822 150492 585828
rect 140780 584452 140832 584458
rect 140780 584394 140832 584400
rect 140688 577720 140740 577726
rect 140688 577662 140740 577668
rect 140792 576854 140820 584394
rect 147220 583092 147272 583098
rect 147220 583034 147272 583040
rect 147232 576854 147260 583034
rect 147864 577652 147916 577658
rect 147864 577594 147916 577600
rect 147876 576854 147904 577594
rect 150452 576854 150480 585822
rect 153672 576854 153700 591330
rect 171152 589966 171180 677622
rect 171230 671256 171286 671265
rect 171230 671191 171286 671200
rect 171140 589960 171192 589966
rect 171140 589902 171192 589908
rect 157246 589384 157302 589393
rect 157246 589319 157302 589328
rect 158626 589384 158682 589393
rect 158626 589319 158682 589328
rect 154580 577652 154632 577658
rect 154580 577594 154632 577600
rect 154592 576854 154620 577594
rect 135640 576826 135760 576854
rect 140792 576826 140912 576854
rect 147232 576826 147352 576854
rect 147876 576826 147996 576854
rect 150452 576826 150572 576854
rect 153672 576826 153792 576854
rect 154592 576826 155264 576854
rect 133880 569424 133932 569430
rect 133880 569366 133932 569372
rect 130566 568848 130622 568857
rect 130566 568783 130622 568792
rect 126058 568712 126114 568721
rect 126058 568647 126114 568656
rect 125508 566500 125560 566506
rect 125508 566442 125560 566448
rect 124956 564800 125008 564806
rect 124956 564742 125008 564748
rect 121550 562728 121606 562737
rect 121550 562663 121606 562672
rect 121564 559994 121592 562663
rect 117332 559966 117576 559994
rect 121486 559966 121592 559994
rect 124968 559994 124996 564742
rect 126072 559994 126100 568647
rect 130580 559994 130608 568783
rect 131212 567384 131264 567390
rect 131212 567326 131264 567332
rect 124968 559966 125350 559994
rect 125994 559966 126100 559994
rect 130502 559966 130608 559994
rect 131224 559994 131252 567326
rect 135732 559994 135760 576826
rect 138020 562012 138072 562018
rect 138020 561954 138072 561960
rect 131224 559966 131744 559994
rect 135654 559966 135760 559994
rect 138032 559994 138060 561954
rect 138572 561740 138624 561746
rect 138572 561682 138624 561688
rect 140504 561740 140556 561746
rect 140504 561682 140556 561688
rect 138584 559994 138612 561682
rect 140516 559994 140544 561682
rect 140884 559994 140912 576826
rect 143446 566264 143502 566273
rect 143446 566199 143502 566208
rect 143460 559994 143488 566199
rect 146208 564800 146260 564806
rect 146208 564742 146260 564748
rect 146220 559994 146248 564742
rect 147324 559994 147352 576826
rect 147968 559994 147996 576826
rect 148784 562352 148836 562358
rect 148784 562294 148836 562300
rect 148796 559994 148824 562294
rect 150544 559994 150572 576826
rect 153764 559994 153792 576826
rect 138032 559966 138230 559994
rect 138584 559966 138874 559994
rect 140162 559966 140544 559994
rect 140806 559966 140912 559994
rect 143382 559966 143488 559994
rect 145958 559966 146248 559994
rect 147246 559966 147352 559994
rect 147890 559966 147996 559994
rect 148534 559966 148824 559994
rect 148980 559978 149178 559994
rect 148968 559972 149178 559978
rect 52000 559914 52052 559920
rect 149020 559966 149178 559972
rect 150466 559966 150572 559994
rect 153686 559966 153792 559994
rect 155236 559994 155264 576826
rect 157260 573578 157288 589319
rect 158640 579018 158668 589319
rect 163320 585948 163372 585954
rect 163320 585890 163372 585896
rect 160100 584520 160152 584526
rect 160100 584462 160152 584468
rect 158628 579012 158680 579018
rect 158628 578954 158680 578960
rect 160112 576854 160140 584462
rect 163332 576854 163360 585890
rect 171244 585886 171272 671191
rect 171322 605704 171378 605713
rect 171322 605639 171378 605648
rect 171336 591394 171364 605639
rect 171324 591388 171376 591394
rect 171324 591330 171376 591336
rect 171692 587852 171744 587858
rect 171692 587794 171744 587800
rect 171232 585880 171284 585886
rect 171232 585822 171284 585828
rect 163964 577720 164016 577726
rect 163964 577662 164016 577668
rect 163976 576854 164004 577662
rect 160112 576826 160232 576854
rect 163332 576826 163452 576854
rect 163976 576826 164096 576854
rect 157248 573572 157300 573578
rect 157248 573514 157300 573520
rect 157800 562420 157852 562426
rect 157800 562362 157852 562368
rect 157812 559994 157840 562362
rect 160204 559994 160232 576826
rect 162308 565004 162360 565010
rect 162308 564946 162360 564952
rect 155236 559966 155572 559994
rect 157550 559966 157840 559994
rect 160126 559966 160232 559994
rect 162320 559994 162348 564946
rect 163424 559994 163452 576826
rect 164068 559994 164096 576826
rect 168564 564936 168616 564942
rect 168564 564878 168616 564884
rect 164332 562488 164384 562494
rect 164332 562430 164384 562436
rect 162320 559966 162702 559994
rect 163346 559966 163452 559994
rect 163990 559966 164096 559994
rect 164344 559994 164372 562430
rect 168576 559994 168604 564878
rect 170770 562048 170826 562057
rect 170770 561983 170826 561992
rect 164344 559966 164634 559994
rect 168498 559966 168604 559994
rect 170784 559994 170812 561983
rect 171704 560130 171732 587794
rect 171796 562630 171824 681255
rect 174544 681216 174596 681222
rect 174544 681158 174596 681164
rect 172610 611416 172666 611425
rect 172610 611351 172666 611360
rect 172518 606928 172574 606937
rect 172518 606863 172574 606872
rect 172532 565282 172560 606863
rect 172624 581738 172652 611351
rect 173806 609784 173862 609793
rect 173806 609719 173862 609728
rect 173820 608666 173848 609719
rect 173808 608660 173860 608666
rect 173808 608602 173860 608608
rect 173806 608424 173862 608433
rect 173806 608359 173862 608368
rect 173820 607238 173848 608359
rect 173808 607232 173860 607238
rect 173808 607174 173860 607180
rect 172612 581732 172664 581738
rect 172612 581674 172664 581680
rect 172520 565276 172572 565282
rect 172520 565218 172572 565224
rect 171784 562624 171836 562630
rect 171784 562566 171836 562572
rect 174556 562562 174584 681158
rect 342904 681012 342956 681018
rect 342904 680954 342956 680960
rect 337568 678292 337620 678298
rect 337568 678234 337620 678240
rect 325056 677748 325108 677754
rect 325056 677690 325108 677696
rect 325068 677657 325096 677690
rect 325792 677680 325844 677686
rect 325054 677648 325110 677657
rect 337580 677657 337608 678234
rect 325792 677622 325844 677628
rect 337566 677648 337622 677657
rect 325054 677583 325110 677592
rect 325804 677113 325832 677622
rect 337566 677583 337622 677592
rect 325790 677104 325846 677113
rect 325790 677039 325846 677048
rect 337580 676870 337608 677583
rect 337568 676864 337620 676870
rect 337568 676806 337620 676812
rect 204166 628280 204222 628289
rect 204166 628215 204222 628224
rect 203522 628008 203578 628017
rect 203522 627943 203578 627952
rect 202144 608660 202196 608666
rect 202144 608602 202196 608608
rect 199384 607232 199436 607238
rect 199384 607174 199436 607180
rect 175924 601724 175976 601730
rect 175924 601666 175976 601672
rect 175936 566642 175964 601666
rect 198188 568744 198240 568750
rect 198188 568686 198240 568692
rect 188528 568676 188580 568682
rect 188528 568618 188580 568624
rect 175924 566636 175976 566642
rect 175924 566578 175976 566584
rect 179696 563848 179748 563854
rect 179696 563790 179748 563796
rect 179144 563440 179196 563446
rect 179144 563382 179196 563388
rect 174544 562556 174596 562562
rect 174544 562498 174596 562504
rect 173898 561912 173954 561921
rect 173898 561847 173954 561856
rect 171704 560102 171824 560130
rect 171796 559994 171824 560102
rect 170784 559966 171074 559994
rect 171718 559966 171824 559994
rect 173912 559994 173940 561847
rect 179156 559994 179184 563382
rect 179708 559994 179736 563790
rect 180706 563408 180762 563417
rect 180706 563343 180762 563352
rect 180720 560130 180748 563343
rect 181076 563100 181128 563106
rect 181076 563042 181128 563048
rect 180720 560102 180794 560130
rect 180766 559994 180794 560102
rect 173912 559966 174294 559994
rect 178802 559966 179184 559994
rect 179446 559966 179736 559994
rect 180734 559966 180794 559994
rect 181088 559994 181116 563042
rect 186872 561944 186924 561950
rect 184846 561912 184902 561921
rect 181628 561876 181680 561882
rect 186872 561886 186924 561892
rect 184846 561847 184902 561856
rect 181628 561818 181680 561824
rect 181640 559994 181668 561818
rect 183008 560652 183060 560658
rect 183008 560594 183060 560600
rect 183020 559994 183048 560594
rect 184860 559994 184888 561847
rect 186884 559994 186912 561886
rect 188540 559994 188568 568618
rect 190366 566672 190422 566681
rect 190366 566607 190422 566616
rect 189446 562184 189502 562193
rect 189446 562119 189502 562128
rect 189460 559994 189488 562119
rect 190380 560130 190408 566607
rect 195886 564768 195942 564777
rect 195886 564703 195942 564712
rect 191380 563508 191432 563514
rect 191380 563450 191432 563456
rect 190380 560102 190454 560130
rect 190426 559994 190454 560102
rect 181088 559966 181378 559994
rect 181640 559966 182022 559994
rect 182666 559966 183048 559994
rect 184598 559966 184888 559994
rect 186530 559966 186912 559994
rect 188462 559966 188568 559994
rect 189106 559966 189488 559994
rect 190394 559966 190454 559994
rect 191392 559994 191420 563450
rect 192576 561876 192628 561882
rect 192576 561818 192628 561824
rect 192588 559994 192616 561818
rect 193864 561808 193916 561814
rect 193864 561750 193916 561756
rect 191392 559966 191682 559994
rect 192326 559966 192616 559994
rect 193876 559994 193904 561750
rect 195900 559994 195928 564703
rect 198200 559994 198228 568686
rect 199396 565282 199424 607174
rect 202156 580310 202184 608602
rect 203062 601760 203118 601769
rect 203062 601695 203064 601704
rect 203116 601695 203118 601704
rect 203064 601666 203116 601672
rect 203536 587722 203564 627943
rect 203614 625424 203670 625433
rect 203614 625359 203670 625368
rect 203628 587790 203656 625359
rect 204074 624200 204130 624209
rect 204074 624135 204130 624144
rect 203982 622432 204038 622441
rect 203982 622367 204038 622376
rect 203890 619712 203946 619721
rect 203890 619647 203946 619656
rect 203798 599448 203854 599457
rect 203798 599383 203854 599392
rect 203616 587784 203668 587790
rect 203616 587726 203668 587732
rect 203524 587716 203576 587722
rect 203524 587658 203576 587664
rect 202880 581732 202932 581738
rect 202880 581674 202932 581680
rect 202144 580304 202196 580310
rect 202144 580246 202196 580252
rect 202892 576854 202920 581674
rect 202892 576826 203380 576854
rect 199384 565276 199436 565282
rect 199384 565218 199436 565224
rect 201408 562692 201460 562698
rect 201408 562634 201460 562640
rect 201038 562048 201094 562057
rect 201038 561983 201094 561992
rect 201052 559994 201080 561983
rect 201420 559994 201448 562634
rect 203156 562488 203208 562494
rect 203156 562430 203208 562436
rect 203168 560294 203196 562430
rect 203352 560294 203380 576826
rect 203812 568002 203840 599383
rect 203904 571062 203932 619647
rect 203892 571056 203944 571062
rect 203892 570998 203944 571004
rect 203800 567996 203852 568002
rect 203800 567938 203852 567944
rect 203996 567934 204024 622367
rect 203984 567928 204036 567934
rect 203984 567870 204036 567876
rect 204088 566642 204116 624135
rect 204180 568070 204208 628215
rect 205546 621986 205602 621995
rect 205546 621921 205602 621930
rect 204902 600400 204958 600409
rect 204902 600335 204958 600344
rect 204916 592006 204944 600335
rect 204904 592000 204956 592006
rect 204904 591942 204956 591948
rect 204916 580514 204944 591942
rect 204904 580508 204956 580514
rect 204904 580450 204956 580456
rect 205560 580446 205588 621921
rect 306288 591320 306340 591326
rect 306288 591262 306340 591268
rect 220818 590608 220874 590617
rect 220818 590543 220874 590552
rect 223026 590608 223082 590617
rect 223026 590543 223082 590552
rect 238390 590608 238446 590617
rect 238390 590543 238446 590552
rect 241518 590608 241574 590617
rect 241518 590543 241574 590552
rect 246670 590608 246726 590617
rect 246670 590543 246726 590552
rect 252374 590608 252430 590617
rect 252374 590543 252430 590552
rect 273258 590608 273314 590617
rect 273258 590543 273314 590552
rect 289542 590608 289598 590617
rect 289542 590543 289598 590552
rect 292118 590608 292174 590617
rect 292118 590543 292174 590552
rect 215484 587104 215536 587110
rect 215484 587046 215536 587052
rect 205548 580440 205600 580446
rect 205548 580382 205600 580388
rect 215496 576854 215524 587046
rect 215496 576826 215616 576854
rect 211712 574932 211764 574938
rect 211712 574874 211764 574880
rect 204168 568064 204220 568070
rect 204168 568006 204220 568012
rect 204076 566636 204128 566642
rect 204076 566578 204128 566584
rect 208032 563712 208084 563718
rect 208032 563654 208084 563660
rect 207478 560960 207534 560969
rect 207478 560895 207534 560904
rect 203168 560266 203288 560294
rect 203352 560266 203472 560294
rect 203260 560130 203288 560266
rect 203260 560102 203380 560130
rect 203352 559994 203380 560102
rect 193876 559966 194212 559994
rect 195546 559966 195928 559994
rect 198122 559966 198228 559994
rect 200698 559966 201080 559994
rect 201342 559966 201448 559994
rect 203274 559966 203380 559994
rect 203444 559994 203472 560266
rect 207492 559994 207520 560895
rect 208044 559994 208072 563654
rect 208766 562320 208822 562329
rect 208766 562255 208822 562264
rect 208780 559994 208808 562255
rect 211724 559994 211752 574874
rect 214472 562080 214524 562086
rect 214472 562022 214524 562028
rect 214484 559994 214512 562022
rect 215588 559994 215616 576826
rect 220832 576230 220860 590543
rect 223040 589558 223068 590543
rect 225144 590028 225196 590034
rect 225144 589970 225196 589976
rect 223028 589552 223080 589558
rect 223028 589494 223080 589500
rect 223578 589384 223634 589393
rect 223578 589319 223634 589328
rect 222200 581664 222252 581670
rect 222200 581606 222252 581612
rect 220820 576224 220872 576230
rect 220820 576166 220872 576172
rect 222016 568812 222068 568818
rect 222016 568754 222068 568760
rect 216862 567216 216918 567225
rect 216862 567151 216918 567160
rect 216876 559994 216904 567151
rect 219716 565344 219768 565350
rect 219716 565286 219768 565292
rect 217784 563644 217836 563650
rect 217784 563586 217836 563592
rect 217796 559994 217824 563586
rect 203444 559966 203872 559994
rect 207138 559966 207520 559994
rect 207782 559966 208072 559994
rect 208426 559966 208808 559994
rect 211646 559966 211752 559994
rect 214222 559966 214512 559994
rect 215510 559966 215616 559994
rect 216798 559966 216904 559994
rect 217442 559966 217824 559994
rect 219728 559994 219756 565286
rect 222028 559994 222056 568754
rect 219728 559966 220018 559994
rect 221950 559966 222056 559994
rect 222212 559994 222240 581606
rect 223592 573646 223620 589319
rect 225156 576854 225184 589970
rect 226432 589960 226484 589966
rect 226432 589902 226484 589908
rect 225326 589384 225382 589393
rect 225326 589319 225382 589328
rect 225340 587654 225368 589319
rect 225328 587648 225380 587654
rect 225328 587590 225380 587596
rect 226444 576854 226472 589902
rect 227076 589688 227128 589694
rect 227076 589630 227128 589636
rect 226614 589384 226670 589393
rect 226614 589319 226670 589328
rect 226628 585886 226656 589319
rect 226616 585880 226668 585886
rect 226616 585822 226668 585828
rect 227088 576854 227116 589630
rect 238404 589558 238432 590543
rect 240598 589792 240654 589801
rect 240598 589727 240654 589736
rect 238392 589552 238444 589558
rect 230202 589520 230258 589529
rect 230202 589455 230258 589464
rect 230478 589520 230534 589529
rect 230478 589455 230534 589464
rect 234526 589520 234582 589529
rect 234526 589455 234582 589464
rect 235998 589520 236054 589529
rect 238392 589494 238444 589500
rect 239954 589520 240010 589529
rect 235998 589455 236054 589464
rect 239954 589455 240010 589464
rect 229006 589384 229062 589393
rect 229006 589319 229062 589328
rect 225156 576826 225276 576854
rect 226444 576826 226564 576854
rect 227088 576826 227208 576854
rect 223580 573640 223632 573646
rect 223580 573582 223632 573588
rect 224224 563576 224276 563582
rect 224224 563518 224276 563524
rect 224236 559994 224264 563518
rect 224776 563508 224828 563514
rect 224776 563450 224828 563456
rect 224788 559994 224816 563450
rect 225248 559994 225276 576826
rect 225420 566704 225472 566710
rect 225420 566646 225472 566652
rect 222212 559966 222548 559994
rect 223882 559966 224264 559994
rect 224526 559966 224816 559994
rect 225170 559966 225276 559994
rect 225432 559994 225460 566646
rect 226536 559994 226564 576826
rect 227180 559994 227208 576826
rect 229020 569430 229048 589319
rect 230216 571130 230244 589455
rect 230386 589384 230442 589393
rect 230386 589319 230442 589328
rect 230296 577720 230348 577726
rect 230296 577662 230348 577668
rect 230204 571124 230256 571130
rect 230204 571066 230256 571072
rect 229008 569424 229060 569430
rect 229008 569366 229060 569372
rect 230308 567194 230336 577662
rect 230400 569498 230428 589319
rect 230388 569492 230440 569498
rect 230388 569434 230440 569440
rect 230308 567166 230428 567194
rect 230400 559994 230428 567166
rect 230492 563786 230520 589455
rect 231858 589384 231914 589393
rect 231858 589319 231914 589328
rect 233238 589384 233294 589393
rect 233238 589319 233294 589328
rect 231872 585954 231900 589319
rect 231860 585948 231912 585954
rect 231860 585890 231912 585896
rect 233252 580378 233280 589319
rect 233240 580372 233292 580378
rect 233240 580314 233292 580320
rect 234540 569566 234568 589455
rect 234618 589384 234674 589393
rect 234618 589319 234674 589328
rect 234528 569560 234580 569566
rect 234528 569502 234580 569508
rect 234632 567866 234660 589319
rect 236012 577590 236040 589455
rect 236090 589384 236146 589393
rect 236090 589319 236146 589328
rect 237286 589384 237342 589393
rect 237286 589319 237342 589328
rect 236104 587858 236132 589319
rect 236092 587852 236144 587858
rect 236092 587794 236144 587800
rect 236000 577584 236052 577590
rect 236000 577526 236052 577532
rect 237300 574938 237328 589319
rect 239312 587648 239364 587654
rect 239312 587590 239364 587596
rect 239324 576854 239352 587590
rect 239968 580378 239996 589455
rect 240046 589384 240102 589393
rect 240046 589319 240102 589328
rect 239956 580372 240008 580378
rect 239956 580314 240008 580320
rect 240060 577590 240088 589319
rect 240612 587722 240640 589727
rect 241532 589626 241560 590543
rect 246684 589626 246712 590543
rect 241520 589620 241572 589626
rect 241520 589562 241572 589568
rect 246672 589620 246724 589626
rect 246672 589562 246724 589568
rect 242806 589520 242862 589529
rect 242806 589455 242862 589464
rect 244278 589520 244334 589529
rect 244278 589455 244334 589464
rect 248418 589520 248474 589529
rect 248418 589455 248474 589464
rect 251178 589520 251234 589529
rect 251178 589455 251234 589464
rect 240600 587716 240652 587722
rect 240600 587658 240652 587664
rect 240048 577584 240100 577590
rect 240048 577526 240100 577532
rect 239324 576826 239444 576854
rect 237288 574932 237340 574938
rect 237288 574874 237340 574880
rect 236184 571396 236236 571402
rect 236184 571338 236236 571344
rect 234620 567860 234672 567866
rect 234620 567802 234672 567808
rect 233792 566160 233844 566166
rect 233792 566102 233844 566108
rect 232504 564936 232556 564942
rect 232504 564878 232556 564884
rect 230480 563780 230532 563786
rect 230480 563722 230532 563728
rect 232516 559994 232544 564878
rect 233804 559994 233832 566102
rect 235080 565072 235132 565078
rect 235080 565014 235132 565020
rect 235092 559994 235120 565014
rect 235816 560720 235868 560726
rect 235816 560662 235868 560668
rect 235828 559994 235856 560662
rect 236196 559994 236224 571338
rect 237380 570988 237432 570994
rect 237380 570930 237432 570936
rect 237392 560266 237420 570930
rect 238668 567452 238720 567458
rect 238668 567394 238720 567400
rect 225432 559966 225814 559994
rect 226458 559966 226564 559994
rect 227102 559966 227208 559994
rect 230322 559966 230428 559994
rect 232254 559966 232544 559994
rect 233542 559966 233832 559994
rect 234830 559966 235120 559994
rect 235474 559966 235856 559994
rect 236118 559966 236224 559994
rect 237346 560238 237420 560266
rect 237346 559980 237374 560238
rect 238680 560130 238708 567394
rect 238680 560102 238754 560130
rect 238726 559994 238754 560102
rect 239416 559994 239444 576826
rect 241336 567520 241388 567526
rect 241336 567462 241388 567468
rect 240046 562456 240102 562465
rect 240046 562391 240102 562400
rect 240060 559994 240088 562391
rect 240968 560788 241020 560794
rect 240968 560730 241020 560736
rect 240980 559994 241008 560730
rect 241348 559994 241376 567462
rect 242820 565350 242848 589455
rect 242898 589384 242954 589393
rect 242898 589319 242954 589328
rect 244186 589384 244242 589393
rect 244186 589319 244242 589328
rect 242912 581738 242940 589319
rect 242900 581732 242952 581738
rect 242900 581674 242952 581680
rect 244200 567866 244228 589319
rect 244188 567860 244240 567866
rect 244188 567802 244240 567808
rect 242808 565344 242860 565350
rect 242808 565286 242860 565292
rect 243636 565276 243688 565282
rect 243636 565218 243688 565224
rect 243544 562216 243596 562222
rect 243544 562158 243596 562164
rect 243556 559994 243584 562158
rect 238694 559966 238754 559994
rect 239338 559966 239444 559994
rect 239982 559966 240088 559994
rect 240626 559966 241008 559994
rect 241270 559966 241376 559994
rect 243202 559966 243584 559994
rect 243648 559994 243676 565218
rect 244292 565214 244320 589455
rect 245566 589384 245622 589393
rect 245566 589319 245622 589328
rect 247038 589384 247094 589393
rect 247038 589319 247094 589328
rect 248326 589384 248382 589393
rect 248326 589319 248382 589328
rect 245580 572082 245608 589319
rect 245844 572144 245896 572150
rect 245844 572086 245896 572092
rect 245568 572076 245620 572082
rect 245568 572018 245620 572024
rect 244280 565208 244332 565214
rect 244280 565150 244332 565156
rect 244924 564868 244976 564874
rect 244924 564810 244976 564816
rect 244832 560856 244884 560862
rect 244832 560798 244884 560804
rect 244844 559994 244872 560798
rect 243648 559966 243846 559994
rect 244490 559966 244872 559994
rect 244936 559994 244964 564810
rect 245856 559994 245884 572086
rect 247052 565146 247080 589319
rect 248340 570994 248368 589319
rect 248432 572257 248460 589455
rect 251192 589422 251220 589455
rect 252388 589422 252416 590543
rect 257344 590096 257396 590102
rect 257344 590038 257396 590044
rect 256054 589792 256110 589801
rect 256054 589727 256110 589736
rect 253938 589520 253994 589529
rect 253938 589455 253994 589464
rect 251180 589416 251232 589422
rect 248510 589384 248566 589393
rect 248510 589319 248566 589328
rect 249798 589384 249854 589393
rect 252376 589416 252428 589422
rect 251180 589358 251232 589364
rect 251270 589384 251326 589393
rect 249798 589319 249854 589328
rect 252376 589358 252428 589364
rect 253846 589384 253902 589393
rect 251270 589319 251326 589328
rect 253846 589319 253902 589328
rect 248524 581806 248552 589319
rect 248512 581800 248564 581806
rect 248512 581742 248564 581748
rect 248418 572248 248474 572257
rect 248418 572183 248474 572192
rect 248328 570988 248380 570994
rect 248328 570930 248380 570936
rect 249812 569362 249840 589319
rect 250444 580508 250496 580514
rect 250444 580450 250496 580456
rect 249800 569356 249852 569362
rect 249800 569298 249852 569304
rect 247040 565140 247092 565146
rect 247040 565082 247092 565088
rect 248328 564868 248380 564874
rect 248328 564810 248380 564816
rect 248340 560130 248368 564810
rect 250456 562018 250484 580450
rect 251284 577658 251312 589319
rect 251272 577652 251324 577658
rect 251272 577594 251324 577600
rect 253860 566710 253888 589319
rect 253952 574841 253980 589455
rect 254122 589384 254178 589393
rect 254122 589319 254178 589328
rect 254136 584526 254164 589319
rect 256068 587790 256096 589727
rect 256056 587784 256108 587790
rect 256056 587726 256108 587732
rect 254124 584520 254176 584526
rect 254124 584462 254176 584468
rect 257356 576854 257384 590038
rect 257986 589520 258042 589529
rect 257986 589455 258042 589464
rect 259458 589520 259514 589529
rect 259458 589455 259514 589464
rect 260838 589520 260894 589529
rect 260838 589455 260894 589464
rect 264886 589520 264942 589529
rect 264886 589455 264942 589464
rect 266358 589520 266414 589529
rect 266358 589455 266414 589464
rect 257894 589384 257950 589393
rect 257894 589319 257950 589328
rect 257356 576826 257476 576854
rect 253938 574832 253994 574841
rect 253938 574767 253994 574776
rect 253848 566704 253900 566710
rect 253848 566646 253900 566652
rect 253940 566568 253992 566574
rect 253940 566510 253992 566516
rect 251824 565140 251876 565146
rect 251824 565082 251876 565088
rect 250444 562012 250496 562018
rect 250444 561954 250496 561960
rect 248340 560102 248414 560130
rect 248386 559994 248414 560102
rect 250456 559994 250484 561954
rect 251836 559994 251864 565082
rect 244936 559966 245134 559994
rect 245778 559966 245884 559994
rect 248354 559966 248414 559994
rect 250286 559966 250484 559994
rect 251574 559966 251864 559994
rect 253952 559994 253980 566510
rect 255136 565004 255188 565010
rect 255136 564946 255188 564952
rect 255148 559994 255176 564946
rect 255504 563372 255556 563378
rect 255504 563314 255556 563320
rect 255516 559994 255544 563314
rect 255688 563304 255740 563310
rect 255688 563246 255740 563252
rect 253952 559966 254150 559994
rect 254794 559966 255176 559994
rect 255438 559966 255544 559994
rect 255700 559994 255728 563246
rect 257448 559994 257476 576826
rect 257908 571198 257936 589319
rect 257896 571192 257948 571198
rect 257896 571134 257948 571140
rect 258000 569362 258028 589455
rect 258078 589384 258134 589393
rect 258078 589319 258134 589328
rect 259274 589384 259330 589393
rect 259472 589354 259500 589455
rect 260746 589384 260802 589393
rect 259274 589319 259330 589328
rect 259460 589348 259512 589354
rect 257988 569356 258040 569362
rect 257988 569298 258040 569304
rect 258092 563854 258120 589319
rect 259288 568138 259316 589319
rect 260746 589319 260802 589328
rect 259460 589290 259512 589296
rect 259276 568132 259328 568138
rect 259276 568074 259328 568080
rect 258080 563848 258132 563854
rect 258080 563790 258132 563796
rect 260760 563786 260788 589319
rect 260852 570926 260880 589455
rect 262126 589384 262182 589393
rect 262126 589319 262182 589328
rect 263506 589384 263562 589393
rect 263506 589319 263562 589328
rect 264794 589384 264850 589393
rect 264794 589319 264850 589328
rect 260840 570920 260892 570926
rect 260840 570862 260892 570868
rect 262140 566574 262168 589319
rect 263520 570926 263548 589319
rect 264808 575006 264836 589319
rect 264796 575000 264848 575006
rect 264796 574942 264848 574948
rect 264900 571266 264928 589455
rect 266266 589384 266322 589393
rect 266266 589319 266322 589328
rect 265072 585948 265124 585954
rect 265072 585890 265124 585896
rect 264888 571260 264940 571266
rect 264888 571202 264940 571208
rect 263508 570920 263560 570926
rect 263508 570862 263560 570868
rect 263232 567588 263284 567594
rect 263232 567530 263284 567536
rect 262128 566568 262180 566574
rect 262128 566510 262180 566516
rect 260748 563780 260800 563786
rect 260748 563722 260800 563728
rect 260748 563304 260800 563310
rect 260748 563246 260800 563252
rect 260288 562148 260340 562154
rect 260288 562090 260340 562096
rect 260300 559994 260328 562090
rect 260760 559994 260788 563246
rect 263244 559994 263272 567530
rect 265084 567194 265112 585890
rect 265164 568880 265216 568886
rect 265164 568822 265216 568828
rect 264992 567166 265112 567194
rect 264992 560294 265020 567166
rect 265176 560294 265204 568822
rect 266280 563854 266308 589319
rect 266372 585721 266400 589455
rect 270406 589384 270462 589393
rect 270406 589319 270462 589328
rect 271878 589384 271934 589393
rect 271878 589319 271934 589328
rect 266358 585712 266414 585721
rect 266358 585647 266414 585656
rect 270224 579012 270276 579018
rect 270224 578954 270276 578960
rect 270236 576854 270264 578954
rect 270236 576826 270356 576854
rect 269856 565208 269908 565214
rect 269856 565150 269908 565156
rect 266268 563848 266320 563854
rect 266268 563790 266320 563796
rect 267922 561776 267978 561785
rect 267922 561711 267978 561720
rect 264992 560266 265112 560294
rect 265176 560266 265296 560294
rect 265084 560130 265112 560266
rect 265084 560102 265204 560130
rect 265176 559994 265204 560102
rect 255700 559966 256036 559994
rect 257370 559966 257476 559994
rect 259946 559966 260328 559994
rect 260590 559966 260788 559994
rect 263166 559966 263272 559994
rect 265098 559966 265204 559994
rect 265268 559994 265296 560266
rect 267936 559994 267964 561711
rect 269868 559994 269896 565150
rect 270328 559994 270356 576826
rect 270420 576230 270448 589319
rect 271892 583098 271920 589319
rect 271880 583092 271932 583098
rect 271880 583034 271932 583040
rect 270408 576224 270460 576230
rect 270408 576166 270460 576172
rect 273272 576065 273300 590543
rect 278962 589656 279018 589665
rect 278962 589591 279018 589600
rect 277306 589384 277362 589393
rect 277306 589319 277362 589328
rect 277320 581670 277348 589319
rect 278976 587110 279004 589591
rect 282826 589384 282882 589393
rect 282826 589319 282882 589328
rect 284298 589384 284354 589393
rect 289556 589354 289584 590543
rect 292132 589694 292160 590543
rect 292764 590164 292816 590170
rect 292764 590106 292816 590112
rect 292120 589688 292172 589694
rect 292120 589630 292172 589636
rect 284298 589319 284354 589328
rect 289544 589348 289596 589354
rect 278964 587104 279016 587110
rect 278964 587046 279016 587052
rect 277308 581664 277360 581670
rect 277308 581606 277360 581612
rect 278596 580440 278648 580446
rect 278596 580382 278648 580388
rect 278608 576854 278636 580382
rect 282840 579018 282868 589319
rect 282828 579012 282880 579018
rect 282828 578954 282880 578960
rect 278608 576826 278728 576854
rect 273258 576056 273314 576065
rect 273258 575991 273314 576000
rect 273168 566092 273220 566098
rect 273168 566034 273220 566040
rect 273180 559994 273208 566034
rect 275006 564904 275062 564913
rect 275006 564839 275062 564848
rect 274454 562728 274510 562737
rect 274454 562663 274510 562672
rect 274468 559994 274496 562663
rect 275020 559994 275048 564839
rect 277030 563680 277086 563689
rect 277030 563615 277086 563624
rect 277044 559994 277072 563615
rect 278320 562284 278372 562290
rect 278320 562226 278372 562232
rect 278332 559994 278360 562226
rect 278700 559994 278728 576826
rect 284312 567905 284340 589319
rect 289544 589290 289596 589296
rect 292776 576854 292804 590106
rect 293958 589520 294014 589529
rect 293958 589455 294014 589464
rect 296718 589520 296774 589529
rect 296718 589455 296774 589464
rect 299478 589520 299534 589529
rect 299478 589455 299534 589464
rect 300858 589520 300914 589529
rect 300858 589455 300914 589464
rect 293972 585954 294000 589455
rect 295984 588668 296036 588674
rect 295984 588610 296036 588616
rect 293960 585948 294012 585954
rect 293960 585890 294012 585896
rect 295996 576854 296024 588610
rect 292776 576826 292896 576854
rect 295996 576826 296116 576854
rect 290924 569968 290976 569974
rect 290924 569910 290976 569916
rect 284298 567896 284354 567905
rect 284298 567831 284354 567840
rect 289176 567656 289228 567662
rect 289176 567598 289228 567604
rect 281540 565344 281592 565350
rect 281540 565286 281592 565292
rect 265268 559966 265696 559994
rect 267936 559966 268318 559994
rect 269606 559966 269896 559994
rect 270250 559966 270356 559994
rect 272826 559966 273208 559994
rect 274114 559966 274496 559994
rect 274758 559966 275048 559994
rect 276690 559966 277072 559994
rect 277978 559966 278360 559994
rect 278622 559966 278728 559994
rect 281552 559994 281580 565286
rect 287888 560924 287940 560930
rect 287888 560866 287940 560872
rect 287900 559994 287928 560866
rect 281552 559966 281842 559994
rect 287638 559966 287928 559994
rect 289188 559994 289216 567598
rect 290936 559994 290964 569910
rect 292868 559994 292896 576826
rect 294326 563272 294382 563281
rect 294326 563207 294382 563216
rect 289188 559966 289524 559994
rect 290858 559966 290964 559994
rect 292790 559966 292896 559994
rect 294340 559994 294368 563207
rect 296088 559994 296116 576826
rect 296732 570858 296760 589455
rect 297916 580440 297968 580446
rect 297916 580382 297968 580388
rect 297928 576854 297956 580382
rect 299492 578950 299520 589455
rect 299480 578944 299532 578950
rect 299480 578886 299532 578892
rect 297928 576826 298048 576854
rect 296720 570852 296772 570858
rect 296720 570794 296772 570800
rect 297638 563272 297694 563281
rect 297638 563207 297694 563216
rect 297652 559994 297680 563207
rect 298020 559994 298048 576826
rect 300872 574705 300900 589455
rect 300858 574696 300914 574705
rect 300858 574631 300914 574640
rect 303988 568948 304040 568954
rect 303988 568890 304040 568896
rect 301412 564732 301464 564738
rect 301412 564674 301464 564680
rect 298926 563544 298982 563553
rect 298926 563479 298982 563488
rect 298940 559994 298968 563479
rect 299388 560992 299440 560998
rect 299388 560934 299440 560940
rect 299400 559994 299428 560934
rect 294340 559966 294676 559994
rect 296010 559966 296116 559994
rect 297298 559966 297680 559994
rect 297942 559966 298048 559994
rect 298586 559966 298968 559994
rect 299230 559966 299428 559994
rect 301424 559994 301452 564674
rect 304000 562426 304028 568890
rect 304080 562556 304132 562562
rect 304080 562498 304132 562504
rect 303988 562420 304040 562426
rect 303988 562362 304040 562368
rect 304092 559994 304120 562498
rect 305920 562420 305972 562426
rect 305920 562362 305972 562368
rect 305932 559994 305960 562362
rect 306300 560130 306328 591262
rect 312082 590608 312138 590617
rect 312082 590543 312138 590552
rect 306378 589520 306434 589529
rect 309138 589520 309194 589529
rect 306378 589455 306434 589464
rect 308404 589484 308456 589490
rect 306392 577726 306420 589455
rect 312096 589490 312124 590543
rect 317420 590232 317472 590238
rect 317420 590174 317472 590180
rect 309138 589455 309194 589464
rect 312084 589484 312136 589490
rect 308404 589426 308456 589432
rect 306380 577720 306432 577726
rect 306380 577662 306432 577668
rect 308416 576298 308444 589426
rect 308404 576292 308456 576298
rect 308404 576234 308456 576240
rect 307024 576224 307076 576230
rect 307024 576166 307076 576172
rect 307760 576224 307812 576230
rect 307760 576166 307812 576172
rect 306300 560102 306374 560130
rect 306346 559994 306374 560102
rect 307036 559994 307064 576166
rect 307772 563378 307800 576166
rect 309152 571985 309180 589455
rect 312084 589426 312136 589432
rect 317432 576854 317460 590174
rect 329746 589656 329802 589665
rect 329746 589591 329802 589600
rect 329654 589520 329710 589529
rect 329654 589455 329710 589464
rect 320456 583092 320508 583098
rect 320456 583034 320508 583040
rect 320468 576854 320496 583034
rect 317432 576826 318104 576854
rect 320468 576826 320588 576854
rect 309138 571976 309194 571985
rect 309138 571911 309194 571920
rect 308310 567352 308366 567361
rect 308310 567287 308366 567296
rect 307760 563372 307812 563378
rect 307760 563314 307812 563320
rect 307668 561196 307720 561202
rect 307668 561138 307720 561144
rect 307680 559994 307708 561138
rect 308324 559994 308352 567287
rect 315948 565276 316000 565282
rect 315948 565218 316000 565224
rect 314936 564732 314988 564738
rect 314936 564674 314988 564680
rect 308496 563372 308548 563378
rect 308496 563314 308548 563320
rect 313096 563372 313148 563378
rect 313096 563314 313148 563320
rect 301424 559966 301806 559994
rect 303738 559966 304120 559994
rect 305670 559966 305960 559994
rect 306314 559966 306374 559994
rect 306958 559966 307064 559994
rect 307602 559966 307708 559994
rect 308246 559966 308352 559994
rect 308508 559994 308536 563314
rect 311162 560824 311218 560833
rect 311162 560759 311218 560768
rect 311176 559994 311204 560759
rect 313108 559994 313136 563314
rect 314948 559994 314976 564674
rect 315672 561060 315724 561066
rect 315672 561002 315724 561008
rect 315684 559994 315712 561002
rect 315960 560130 315988 565218
rect 317972 562624 318024 562630
rect 317972 562566 318024 562572
rect 315960 560102 316080 560130
rect 316052 559994 316080 560102
rect 317984 559994 318012 562566
rect 308508 559966 308844 559994
rect 311176 559966 311466 559994
rect 312754 559966 313136 559994
rect 314686 559966 314976 559994
rect 315330 559966 315712 559994
rect 315974 559966 316080 559994
rect 317906 559966 318012 559994
rect 318076 559994 318104 576826
rect 319168 561740 319220 561746
rect 319168 561682 319220 561688
rect 319180 560046 319208 561682
rect 319168 560040 319220 560046
rect 318076 559966 318504 559994
rect 320560 559994 320588 576826
rect 329668 568206 329696 589455
rect 329656 568200 329708 568206
rect 329656 568142 329708 568148
rect 329760 566778 329788 589591
rect 330208 576292 330260 576298
rect 330208 576234 330260 576240
rect 329748 566772 329800 566778
rect 329748 566714 329800 566720
rect 322112 564460 322164 564466
rect 322112 564402 322164 564408
rect 322124 559994 322152 564402
rect 324688 563916 324740 563922
rect 324688 563858 324740 563864
rect 324700 559994 324728 563858
rect 325976 563236 326028 563242
rect 325976 563178 326028 563184
rect 325608 561740 325660 561746
rect 325608 561682 325660 561688
rect 325620 560130 325648 561682
rect 325620 560102 325694 560130
rect 325666 559994 325694 560102
rect 319168 559982 319220 559988
rect 320482 559966 320588 559994
rect 321770 559966 322152 559994
rect 324346 559966 324728 559994
rect 325634 559966 325694 559994
rect 325988 559994 326016 563178
rect 328366 560688 328422 560697
rect 328366 560623 328422 560632
rect 328380 559994 328408 560623
rect 330220 559994 330248 576234
rect 331496 573504 331548 573510
rect 331496 573446 331548 573452
rect 330482 561368 330538 561377
rect 330482 561303 330538 561312
rect 325988 559966 326278 559994
rect 327566 559978 327764 559994
rect 327566 559972 327776 559978
rect 327566 559966 327724 559972
rect 148968 559914 149020 559920
rect 328210 559966 328408 559994
rect 330142 559966 330248 559994
rect 330496 559994 330524 561303
rect 331508 559994 331536 573446
rect 336280 566228 336332 566234
rect 336280 566170 336332 566176
rect 334992 563236 335044 563242
rect 334992 563178 335044 563184
rect 335004 559994 335032 563178
rect 336186 563136 336242 563145
rect 336186 563071 336242 563080
rect 336200 562358 336228 563071
rect 336188 562352 336240 562358
rect 336188 562294 336240 562300
rect 336292 559994 336320 566170
rect 340144 563100 340196 563106
rect 340144 563042 340196 563048
rect 338028 563032 338080 563038
rect 338028 562974 338080 562980
rect 337568 561128 337620 561134
rect 337568 561070 337620 561076
rect 337580 559994 337608 561070
rect 338040 559994 338068 562974
rect 340156 562494 340184 563042
rect 342916 563038 342944 680954
rect 343008 670682 343036 700402
rect 389916 697604 389968 697610
rect 389916 697546 389968 697552
rect 383016 690668 383068 690674
rect 383016 690610 383068 690616
rect 373632 687948 373684 687954
rect 373632 687890 373684 687896
rect 367744 686112 367796 686118
rect 367744 686054 367796 686060
rect 364248 682644 364300 682650
rect 364248 682586 364300 682592
rect 360844 682168 360896 682174
rect 360844 682110 360896 682116
rect 358084 679244 358136 679250
rect 358084 679186 358136 679192
rect 343732 677748 343784 677754
rect 343732 677690 343784 677696
rect 343638 671256 343694 671265
rect 343638 671191 343694 671200
rect 342996 670676 343048 670682
rect 342996 670618 343048 670624
rect 343652 576230 343680 671191
rect 343744 590238 343772 677690
rect 353944 677680 353996 677686
rect 353944 677622 353996 677628
rect 347044 648644 347096 648650
rect 347044 648586 347096 648592
rect 344284 641776 344336 641782
rect 344284 641718 344336 641724
rect 343732 590232 343784 590238
rect 343732 590174 343784 590180
rect 343640 576224 343692 576230
rect 343640 576166 343692 576172
rect 344296 572150 344324 641718
rect 346306 611416 346362 611425
rect 346306 611351 346308 611360
rect 346360 611351 346362 611360
rect 346308 611322 346360 611328
rect 345018 609784 345074 609793
rect 345018 609719 345074 609728
rect 345032 587586 345060 609719
rect 345110 608424 345166 608433
rect 345110 608359 345166 608368
rect 345124 607238 345152 608359
rect 345112 607232 345164 607238
rect 345112 607174 345164 607180
rect 345570 606928 345626 606937
rect 345570 606863 345626 606872
rect 345584 605878 345612 606863
rect 345572 605872 345624 605878
rect 345572 605814 345624 605820
rect 345110 605704 345166 605713
rect 345110 605639 345166 605648
rect 345020 587580 345072 587586
rect 345020 587522 345072 587528
rect 345124 584458 345152 605639
rect 345112 584452 345164 584458
rect 345112 584394 345164 584400
rect 347056 580446 347084 648586
rect 348516 589688 348568 589694
rect 348516 589630 348568 589636
rect 347044 580440 347096 580446
rect 347044 580382 347096 580388
rect 348056 577516 348108 577522
rect 348056 577458 348108 577464
rect 347780 576156 347832 576162
rect 347780 576098 347832 576104
rect 344284 572144 344336 572150
rect 344284 572086 344336 572092
rect 347596 566160 347648 566166
rect 347596 566102 347648 566108
rect 346492 563848 346544 563854
rect 346492 563790 346544 563796
rect 343732 563780 343784 563786
rect 343732 563722 343784 563728
rect 342904 563032 342956 563038
rect 342904 562974 342956 562980
rect 340144 562488 340196 562494
rect 340144 562430 340196 562436
rect 340144 561944 340196 561950
rect 340144 561886 340196 561892
rect 340052 561808 340104 561814
rect 340052 561750 340104 561756
rect 340064 559994 340092 561750
rect 340156 561105 340184 561886
rect 341982 561776 342038 561785
rect 341982 561711 342038 561720
rect 340142 561096 340198 561105
rect 340142 561031 340198 561040
rect 341996 559994 342024 561711
rect 343744 559994 343772 563722
rect 330496 559966 330786 559994
rect 331430 559966 331536 559994
rect 334650 559966 335032 559994
rect 335938 559966 336320 559994
rect 336582 559978 336688 559994
rect 336582 559972 336700 559978
rect 336582 559966 336648 559972
rect 327724 559914 327776 559920
rect 337226 559966 337608 559994
rect 337870 559966 338068 559994
rect 339802 559966 340092 559994
rect 340446 559978 340736 559994
rect 340446 559972 340748 559978
rect 340446 559966 340696 559972
rect 336648 559914 336700 559920
rect 341734 559966 342024 559994
rect 343666 559966 343772 559994
rect 346504 559994 346532 563790
rect 347228 562284 347280 562290
rect 347228 562226 347280 562232
rect 346504 559966 346886 559994
rect 347240 559978 347268 562226
rect 347320 562080 347372 562086
rect 347320 562022 347372 562028
rect 347332 559978 347360 562022
rect 347608 560250 347636 566102
rect 347688 562080 347740 562086
rect 347688 562022 347740 562028
rect 347596 560244 347648 560250
rect 347596 560186 347648 560192
rect 347700 559994 347728 562022
rect 347228 559972 347280 559978
rect 340696 559914 340748 559920
rect 347228 559914 347280 559920
rect 347320 559972 347372 559978
rect 347530 559966 347728 559994
rect 347320 559914 347372 559920
rect 347792 471209 347820 576098
rect 347964 574932 348016 574938
rect 347964 574874 348016 574880
rect 347872 573572 347924 573578
rect 347872 573514 347924 573520
rect 347778 471200 347834 471209
rect 347778 471135 347834 471144
rect 347884 451489 347912 573514
rect 347870 451480 347926 451489
rect 347870 451415 347926 451424
rect 347870 445768 347926 445777
rect 347870 445703 347926 445712
rect 347686 200424 347742 200433
rect 347686 200359 347742 200368
rect 48056 197946 48084 200124
rect 48700 198694 48728 200124
rect 48688 198688 48740 198694
rect 48688 198630 48740 198636
rect 48044 197940 48096 197946
rect 48044 197882 48096 197888
rect 49240 197872 49292 197878
rect 49240 197814 49292 197820
rect 48044 192704 48096 192710
rect 48044 192646 48096 192652
rect 47952 174548 48004 174554
rect 47952 174490 48004 174496
rect 47860 158092 47912 158098
rect 47860 158034 47912 158040
rect 47860 155848 47912 155854
rect 47860 155790 47912 155796
rect 47768 24064 47820 24070
rect 47768 24006 47820 24012
rect 47308 22976 47360 22982
rect 47308 22918 47360 22924
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 47872 17814 47900 155790
rect 47964 18494 47992 174490
rect 48056 23458 48084 192646
rect 48228 191344 48280 191350
rect 48228 191286 48280 191292
rect 48044 23452 48096 23458
rect 48044 23394 48096 23400
rect 47952 18488 48004 18494
rect 47952 18430 48004 18436
rect 47860 17808 47912 17814
rect 47860 17750 47912 17756
rect 46664 17604 46716 17610
rect 46664 17546 46716 17552
rect 46388 17196 46440 17202
rect 46388 17138 46440 17144
rect 46662 14512 46718 14521
rect 46662 14447 46718 14456
rect 45008 3800 45060 3806
rect 45008 3742 45060 3748
rect 43074 3496 43130 3505
rect 43074 3431 43130 3440
rect 42432 3392 42484 3398
rect 42432 3334 42484 3340
rect 43088 480 43116 3431
rect 46676 480 46704 14447
rect 48240 3874 48268 191286
rect 48964 188352 49016 188358
rect 48778 188320 48834 188329
rect 48964 188294 49016 188300
rect 48778 188255 48834 188264
rect 48792 4010 48820 188255
rect 48872 185700 48924 185706
rect 48872 185642 48924 185648
rect 48884 112946 48912 185642
rect 48872 112940 48924 112946
rect 48872 112882 48924 112888
rect 48870 112432 48926 112441
rect 48870 112367 48926 112376
rect 48884 21690 48912 112367
rect 48976 82142 49004 188294
rect 49148 155168 49200 155174
rect 49148 155110 49200 155116
rect 49056 151768 49108 151774
rect 49056 151710 49108 151716
rect 48964 82136 49016 82142
rect 48964 82078 49016 82084
rect 49068 24818 49096 151710
rect 49056 24812 49108 24818
rect 49056 24754 49108 24760
rect 49160 21962 49188 155110
rect 49252 53786 49280 197814
rect 49344 197402 49372 200124
rect 49988 198257 50016 200124
rect 50632 198914 50660 200124
rect 50080 198886 50660 198914
rect 49974 198248 50030 198257
rect 49974 198183 50030 198192
rect 49332 197396 49384 197402
rect 49332 197338 49384 197344
rect 49516 195832 49568 195838
rect 49516 195774 49568 195780
rect 49424 195152 49476 195158
rect 49424 195094 49476 195100
rect 49330 179208 49386 179217
rect 49330 179143 49386 179152
rect 49240 53780 49292 53786
rect 49240 53722 49292 53728
rect 49344 29617 49372 179143
rect 49330 29608 49386 29617
rect 49330 29543 49386 29552
rect 49436 28898 49464 195094
rect 49424 28892 49476 28898
rect 49424 28834 49476 28840
rect 49148 21956 49200 21962
rect 49148 21898 49200 21904
rect 48872 21684 48924 21690
rect 48872 21626 48924 21632
rect 49528 21622 49556 195774
rect 50080 180794 50108 198886
rect 50344 198824 50396 198830
rect 50344 198766 50396 198772
rect 49712 180766 50108 180794
rect 49712 169046 49740 180766
rect 49700 169040 49752 169046
rect 49700 168982 49752 168988
rect 50160 164892 50212 164898
rect 50160 164834 50212 164840
rect 50068 150816 50120 150822
rect 50068 150758 50120 150764
rect 49608 149864 49660 149870
rect 49608 149806 49660 149812
rect 49620 141409 49648 149806
rect 49700 142248 49752 142254
rect 49700 142190 49752 142196
rect 49606 141400 49662 141409
rect 49606 141335 49662 141344
rect 49712 139482 49740 142190
rect 49620 139454 49740 139482
rect 49620 126954 49648 139454
rect 49608 126948 49660 126954
rect 49608 126890 49660 126896
rect 50080 23186 50108 150758
rect 50068 23180 50120 23186
rect 50068 23122 50120 23128
rect 49516 21616 49568 21622
rect 49516 21558 49568 21564
rect 50172 16574 50200 164834
rect 50356 152454 50384 198766
rect 51276 194206 51304 200124
rect 52828 197804 52880 197810
rect 52828 197746 52880 197752
rect 52276 195628 52328 195634
rect 52276 195570 52328 195576
rect 51540 195424 51592 195430
rect 51540 195366 51592 195372
rect 51264 194200 51316 194206
rect 51264 194142 51316 194148
rect 50436 193860 50488 193866
rect 50436 193802 50488 193808
rect 50344 152448 50396 152454
rect 50344 152390 50396 152396
rect 50252 147348 50304 147354
rect 50252 147290 50304 147296
rect 50264 107642 50292 147290
rect 50344 126948 50396 126954
rect 50344 126890 50396 126896
rect 50252 107636 50304 107642
rect 50252 107578 50304 107584
rect 50356 17474 50384 126890
rect 50448 104786 50476 193802
rect 50804 191412 50856 191418
rect 50804 191354 50856 191360
rect 50620 188488 50672 188494
rect 50620 188430 50672 188436
rect 50528 172100 50580 172106
rect 50528 172042 50580 172048
rect 50436 104780 50488 104786
rect 50436 104722 50488 104728
rect 50540 67182 50568 172042
rect 50632 138689 50660 188430
rect 50712 151020 50764 151026
rect 50712 150962 50764 150968
rect 50618 138680 50674 138689
rect 50618 138615 50674 138624
rect 50528 67176 50580 67182
rect 50528 67118 50580 67124
rect 50724 22914 50752 150962
rect 50816 142866 50844 191354
rect 50894 176624 50950 176633
rect 50894 176559 50950 176568
rect 50804 142860 50856 142866
rect 50804 142802 50856 142808
rect 50802 139496 50858 139505
rect 50802 139431 50858 139440
rect 50712 22908 50764 22914
rect 50712 22850 50764 22856
rect 50816 19281 50844 139431
rect 50908 27538 50936 176559
rect 50988 155372 51040 155378
rect 50988 155314 51040 155320
rect 51000 139505 51028 155314
rect 51448 149932 51500 149938
rect 51448 149874 51500 149880
rect 50986 139496 51042 139505
rect 50986 139431 51042 139440
rect 51460 136610 51488 149874
rect 51448 136604 51500 136610
rect 51448 136546 51500 136552
rect 50988 136196 51040 136202
rect 50988 136138 51040 136144
rect 51000 127838 51028 136138
rect 50988 127832 51040 127838
rect 50988 127774 51040 127780
rect 50896 27532 50948 27538
rect 50896 27474 50948 27480
rect 51552 23934 51580 195366
rect 51724 195220 51776 195226
rect 51724 195162 51776 195168
rect 51630 178800 51686 178809
rect 51630 178735 51686 178744
rect 51644 93838 51672 178735
rect 51632 93832 51684 93838
rect 51632 93774 51684 93780
rect 51632 92540 51684 92546
rect 51632 92482 51684 92488
rect 51540 23928 51592 23934
rect 51540 23870 51592 23876
rect 50802 19272 50858 19281
rect 50802 19207 50858 19216
rect 50344 17468 50396 17474
rect 50344 17410 50396 17416
rect 51644 16930 51672 92482
rect 51736 75886 51764 195162
rect 52184 192568 52236 192574
rect 52184 192510 52236 192516
rect 52092 185836 52144 185842
rect 52092 185778 52144 185784
rect 52000 155508 52052 155514
rect 52000 155450 52052 155456
rect 51816 151292 51868 151298
rect 51816 151234 51868 151240
rect 51724 75880 51776 75886
rect 51724 75822 51776 75828
rect 51828 29306 51856 151234
rect 51908 150952 51960 150958
rect 51908 150894 51960 150900
rect 51816 29300 51868 29306
rect 51816 29242 51868 29248
rect 51920 24206 51948 150894
rect 52012 27062 52040 155450
rect 52104 28966 52132 185778
rect 52092 28960 52144 28966
rect 52092 28902 52144 28908
rect 52196 27606 52224 192510
rect 52184 27600 52236 27606
rect 52184 27542 52236 27548
rect 52000 27056 52052 27062
rect 52000 26998 52052 27004
rect 52288 25498 52316 195570
rect 52458 171728 52514 171737
rect 52458 171663 52514 171672
rect 52368 135380 52420 135386
rect 52368 135322 52420 135328
rect 52380 125526 52408 135322
rect 52368 125520 52420 125526
rect 52368 125462 52420 125468
rect 52276 25492 52328 25498
rect 52276 25434 52328 25440
rect 51908 24200 51960 24206
rect 51908 24142 51960 24148
rect 51632 16924 51684 16930
rect 51632 16866 51684 16872
rect 52472 16574 52500 171663
rect 52840 29578 52868 197746
rect 53208 197441 53236 200124
rect 53852 198665 53880 200124
rect 53838 198656 53894 198665
rect 53838 198591 53894 198600
rect 55784 198286 55812 200124
rect 55772 198280 55824 198286
rect 55772 198222 55824 198228
rect 53288 197940 53340 197946
rect 53288 197882 53340 197888
rect 53194 197432 53250 197441
rect 53104 197396 53156 197402
rect 53194 197367 53250 197376
rect 53104 197338 53156 197344
rect 53012 149796 53064 149802
rect 53012 149738 53064 149744
rect 52920 146260 52972 146266
rect 52920 146202 52972 146208
rect 52932 135386 52960 146202
rect 53024 136202 53052 149738
rect 53012 136196 53064 136202
rect 53012 136138 53064 136144
rect 52920 135380 52972 135386
rect 52920 135322 52972 135328
rect 52828 29572 52880 29578
rect 52828 29514 52880 29520
rect 53116 21894 53144 197338
rect 53196 136604 53248 136610
rect 53196 136546 53248 136552
rect 53208 97918 53236 136546
rect 53300 104854 53328 197882
rect 54482 197432 54538 197441
rect 54482 197367 54538 197376
rect 53656 187128 53708 187134
rect 53656 187070 53708 187076
rect 53380 180192 53432 180198
rect 53380 180134 53432 180140
rect 53392 132569 53420 180134
rect 53564 176316 53616 176322
rect 53564 176258 53616 176264
rect 53472 151496 53524 151502
rect 53472 151438 53524 151444
rect 53378 132560 53434 132569
rect 53378 132495 53434 132504
rect 53380 131164 53432 131170
rect 53380 131106 53432 131112
rect 53288 104848 53340 104854
rect 53288 104790 53340 104796
rect 53196 97912 53248 97918
rect 53196 97854 53248 97860
rect 53288 95260 53340 95266
rect 53288 95202 53340 95208
rect 53300 73710 53328 95202
rect 53288 73704 53340 73710
rect 53288 73646 53340 73652
rect 53104 21888 53156 21894
rect 53104 21830 53156 21836
rect 53392 21486 53420 131106
rect 53484 24002 53512 151438
rect 53576 25566 53604 176258
rect 53564 25560 53616 25566
rect 53564 25502 53616 25508
rect 53668 25430 53696 187070
rect 54298 183016 54354 183025
rect 54298 182951 54354 182960
rect 54208 151700 54260 151706
rect 54208 151642 54260 151648
rect 53840 141432 53892 141438
rect 53840 141374 53892 141380
rect 53852 136626 53880 141374
rect 53760 136598 53880 136626
rect 53760 127634 53788 136598
rect 54116 135924 54168 135930
rect 54116 135866 54168 135872
rect 53748 127628 53800 127634
rect 53748 127570 53800 127576
rect 53748 126268 53800 126274
rect 53748 126210 53800 126216
rect 53760 101998 53788 126210
rect 54128 118658 54156 135866
rect 54116 118652 54168 118658
rect 54116 118594 54168 118600
rect 53748 101992 53800 101998
rect 53748 101934 53800 101940
rect 53656 25424 53708 25430
rect 53656 25366 53708 25372
rect 54220 24750 54248 151642
rect 54312 25362 54340 182951
rect 54392 127832 54444 127838
rect 54392 127774 54444 127780
rect 54404 106729 54432 127774
rect 54390 106720 54446 106729
rect 54390 106655 54446 106664
rect 54496 27402 54524 197367
rect 58360 195650 58388 200124
rect 59004 198665 59032 200124
rect 58990 198656 59046 198665
rect 58990 198591 59046 198600
rect 60292 197169 60320 200124
rect 60278 197160 60334 197169
rect 60278 197095 60334 197104
rect 57992 195622 58388 195650
rect 54852 195560 54904 195566
rect 54852 195502 54904 195508
rect 54576 194200 54628 194206
rect 54576 194142 54628 194148
rect 54588 152386 54616 194142
rect 54760 178832 54812 178838
rect 54760 178774 54812 178780
rect 54576 152380 54628 152386
rect 54576 152322 54628 152328
rect 54576 150000 54628 150006
rect 54576 149942 54628 149948
rect 54588 131170 54616 149942
rect 54668 147008 54720 147014
rect 54668 146950 54720 146956
rect 54576 131164 54628 131170
rect 54576 131106 54628 131112
rect 54576 129736 54628 129742
rect 54576 129678 54628 129684
rect 54588 120766 54616 129678
rect 54576 120760 54628 120766
rect 54576 120702 54628 120708
rect 54680 113830 54708 146950
rect 54772 126954 54800 178774
rect 54864 129674 54892 195502
rect 56048 195492 56100 195498
rect 56048 195434 56100 195440
rect 55862 181384 55918 181393
rect 55862 181319 55918 181328
rect 55588 179172 55640 179178
rect 55588 179114 55640 179120
rect 55036 167680 55088 167686
rect 55036 167622 55088 167628
rect 54944 159452 54996 159458
rect 54944 159394 54996 159400
rect 54852 129668 54904 129674
rect 54852 129610 54904 129616
rect 54760 126948 54812 126954
rect 54760 126890 54812 126896
rect 54760 119400 54812 119406
rect 54760 119342 54812 119348
rect 54668 113824 54720 113830
rect 54668 113766 54720 113772
rect 54668 107636 54720 107642
rect 54668 107578 54720 107584
rect 54484 27396 54536 27402
rect 54484 27338 54536 27344
rect 54300 25356 54352 25362
rect 54300 25298 54352 25304
rect 54208 24744 54260 24750
rect 54208 24686 54260 24692
rect 53472 23996 53524 24002
rect 53472 23938 53524 23944
rect 53380 21480 53432 21486
rect 53380 21422 53432 21428
rect 54680 19174 54708 107578
rect 54772 96150 54800 119342
rect 54852 116476 54904 116482
rect 54852 116418 54904 116424
rect 54760 96144 54812 96150
rect 54760 96086 54812 96092
rect 54760 82884 54812 82890
rect 54760 82826 54812 82832
rect 54668 19168 54720 19174
rect 54668 19110 54720 19116
rect 54772 19038 54800 82826
rect 54864 29753 54892 116418
rect 54956 57322 54984 159394
rect 55048 142118 55076 167622
rect 55128 152924 55180 152930
rect 55128 152866 55180 152872
rect 55036 142112 55088 142118
rect 55036 142054 55088 142060
rect 55140 136610 55168 152866
rect 55494 147520 55550 147529
rect 55494 147455 55550 147464
rect 55128 136604 55180 136610
rect 55128 136546 55180 136552
rect 55128 129600 55180 129606
rect 55128 129542 55180 129548
rect 55036 125520 55088 125526
rect 55036 125462 55088 125468
rect 55048 122834 55076 125462
rect 55140 122942 55168 129542
rect 55128 122936 55180 122942
rect 55128 122878 55180 122884
rect 55312 122868 55364 122874
rect 55048 122806 55168 122834
rect 55312 122810 55364 122816
rect 54944 57316 54996 57322
rect 54944 57258 54996 57264
rect 54850 29744 54906 29753
rect 54850 29679 54906 29688
rect 54760 19032 54812 19038
rect 54760 18974 54812 18980
rect 55140 18698 55168 122806
rect 55220 120760 55272 120766
rect 55220 120702 55272 120708
rect 55232 82890 55260 120702
rect 55324 95266 55352 122810
rect 55404 101992 55456 101998
rect 55404 101934 55456 101940
rect 55312 95260 55364 95266
rect 55312 95202 55364 95208
rect 55416 92546 55444 101934
rect 55404 92540 55456 92546
rect 55404 92482 55456 92488
rect 55220 82884 55272 82890
rect 55220 82826 55272 82832
rect 55508 24138 55536 147455
rect 55600 28286 55628 179114
rect 55772 155440 55824 155446
rect 55772 155382 55824 155388
rect 55784 147354 55812 155382
rect 55772 147348 55824 147354
rect 55772 147290 55824 147296
rect 55772 146124 55824 146130
rect 55772 146066 55824 146072
rect 55784 136542 55812 146066
rect 55876 143546 55904 181319
rect 55956 167816 56008 167822
rect 55956 167758 56008 167764
rect 55864 143540 55916 143546
rect 55864 143482 55916 143488
rect 55864 136604 55916 136610
rect 55864 136546 55916 136552
rect 55772 136536 55824 136542
rect 55772 136478 55824 136484
rect 55876 129742 55904 136546
rect 55864 129736 55916 129742
rect 55864 129678 55916 129684
rect 55968 98161 55996 167758
rect 56060 119241 56088 195434
rect 56324 191752 56376 191758
rect 56324 191694 56376 191700
rect 56140 177608 56192 177614
rect 56140 177550 56192 177556
rect 56046 119232 56102 119241
rect 56046 119167 56102 119176
rect 56046 107536 56102 107545
rect 56046 107471 56102 107480
rect 55954 98152 56010 98161
rect 55954 98087 56010 98096
rect 55864 97912 55916 97918
rect 55864 97854 55916 97860
rect 55588 28280 55640 28286
rect 55588 28222 55640 28228
rect 55496 24132 55548 24138
rect 55496 24074 55548 24080
rect 55876 21350 55904 97854
rect 55956 82136 56008 82142
rect 55956 82078 56008 82084
rect 55864 21344 55916 21350
rect 55864 21286 55916 21292
rect 55128 18692 55180 18698
rect 55128 18634 55180 18640
rect 55968 17270 55996 82078
rect 56060 22098 56088 107471
rect 56152 77081 56180 177550
rect 56232 158228 56284 158234
rect 56232 158170 56284 158176
rect 56138 77072 56194 77081
rect 56138 77007 56194 77016
rect 56244 55321 56272 158170
rect 56336 86601 56364 191694
rect 56782 189952 56838 189961
rect 56782 189887 56838 189896
rect 56416 187400 56468 187406
rect 56416 187342 56468 187348
rect 56428 128382 56456 187342
rect 56508 150884 56560 150890
rect 56508 150826 56560 150832
rect 56520 146266 56548 150826
rect 56508 146260 56560 146266
rect 56508 146202 56560 146208
rect 56508 140888 56560 140894
rect 56508 140830 56560 140836
rect 56520 132530 56548 140830
rect 56508 132524 56560 132530
rect 56508 132466 56560 132472
rect 56508 132388 56560 132394
rect 56508 132330 56560 132336
rect 56416 128376 56468 128382
rect 56416 128318 56468 128324
rect 56520 124098 56548 132330
rect 56508 124092 56560 124098
rect 56508 124034 56560 124040
rect 56600 118652 56652 118658
rect 56600 118594 56652 118600
rect 56508 118176 56560 118182
rect 56508 118118 56560 118124
rect 56520 110498 56548 118118
rect 56508 110492 56560 110498
rect 56508 110434 56560 110440
rect 56612 95146 56640 118594
rect 56520 95118 56640 95146
rect 56322 86592 56378 86601
rect 56322 86527 56378 86536
rect 56230 55312 56286 55321
rect 56230 55247 56286 55256
rect 56048 22092 56100 22098
rect 56048 22034 56100 22040
rect 56520 18630 56548 95118
rect 56796 70281 56824 189887
rect 57612 178900 57664 178906
rect 57612 178842 57664 178848
rect 57520 167884 57572 167890
rect 57520 167826 57572 167832
rect 57428 165028 57480 165034
rect 57428 164970 57480 164976
rect 57336 159588 57388 159594
rect 57336 159530 57388 159536
rect 57244 158160 57296 158166
rect 57244 158102 57296 158108
rect 57152 149116 57204 149122
rect 57152 149058 57204 149064
rect 56968 143540 57020 143546
rect 56968 143482 57020 143488
rect 56980 129606 57008 143482
rect 57164 142254 57192 149058
rect 57152 142248 57204 142254
rect 57152 142190 57204 142196
rect 57060 140820 57112 140826
rect 57060 140762 57112 140768
rect 57072 132734 57100 140762
rect 57152 140684 57204 140690
rect 57152 140626 57204 140632
rect 57164 139641 57192 140626
rect 57150 139632 57206 139641
rect 57150 139567 57206 139576
rect 57060 132728 57112 132734
rect 57060 132670 57112 132676
rect 57152 132524 57204 132530
rect 57152 132466 57204 132472
rect 57060 132456 57112 132462
rect 57060 132398 57112 132404
rect 57072 131481 57100 132398
rect 57058 131472 57114 131481
rect 57058 131407 57114 131416
rect 57060 129668 57112 129674
rect 57060 129610 57112 129616
rect 56968 129600 57020 129606
rect 56968 129542 57020 129548
rect 56876 128376 56928 128382
rect 56876 128318 56928 128324
rect 56888 116482 56916 128318
rect 57072 122834 57100 129610
rect 57164 126274 57192 132466
rect 57256 130801 57284 158102
rect 57242 130792 57298 130801
rect 57242 130727 57298 130736
rect 57244 128308 57296 128314
rect 57244 128250 57296 128256
rect 57256 128081 57284 128250
rect 57242 128072 57298 128081
rect 57242 128007 57298 128016
rect 57244 126948 57296 126954
rect 57244 126890 57296 126896
rect 57256 126721 57284 126890
rect 57242 126712 57298 126721
rect 57242 126647 57298 126656
rect 57152 126268 57204 126274
rect 57152 126210 57204 126216
rect 57244 125588 57296 125594
rect 57244 125530 57296 125536
rect 57256 125361 57284 125530
rect 57242 125352 57298 125361
rect 57242 125287 57298 125296
rect 57244 124160 57296 124166
rect 57244 124102 57296 124108
rect 57256 123321 57284 124102
rect 57242 123312 57298 123321
rect 57242 123247 57298 123256
rect 57072 122806 57284 122834
rect 57152 121712 57204 121718
rect 57152 121654 57204 121660
rect 57164 118046 57192 121654
rect 57152 118040 57204 118046
rect 57152 117982 57204 117988
rect 56876 116476 56928 116482
rect 56876 116418 56928 116424
rect 57152 115252 57204 115258
rect 57152 115194 57204 115200
rect 57060 82952 57112 82958
rect 57060 82894 57112 82900
rect 57072 81161 57100 82894
rect 57058 81152 57114 81161
rect 57058 81087 57114 81096
rect 56968 73704 57020 73710
rect 56968 73646 57020 73652
rect 56782 70272 56838 70281
rect 56782 70207 56838 70216
rect 56980 68134 57008 73646
rect 57060 69692 57112 69698
rect 57060 69634 57112 69640
rect 56968 68128 57020 68134
rect 56968 68070 57020 68076
rect 56690 67552 56746 67561
rect 56690 67487 56746 67496
rect 56704 67182 56732 67487
rect 56692 67176 56744 67182
rect 56692 67118 56744 67124
rect 56968 64864 57020 64870
rect 56968 64806 57020 64812
rect 56980 64161 57008 64806
rect 56966 64152 57022 64161
rect 56966 64087 57022 64096
rect 57072 46481 57100 69634
rect 57058 46472 57114 46481
rect 57058 46407 57114 46416
rect 57164 40361 57192 115194
rect 57150 40352 57206 40361
rect 57150 40287 57206 40296
rect 57256 22710 57284 122806
rect 57348 121582 57376 159530
rect 57336 121576 57388 121582
rect 57336 121518 57388 121524
rect 57336 121440 57388 121446
rect 57336 121382 57388 121388
rect 57348 120601 57376 121382
rect 57334 120592 57390 120601
rect 57334 120527 57390 120536
rect 57336 120012 57388 120018
rect 57336 119954 57388 119960
rect 57348 119921 57376 119954
rect 57334 119912 57390 119921
rect 57334 119847 57390 119856
rect 57336 117292 57388 117298
rect 57336 117234 57388 117240
rect 57348 117201 57376 117234
rect 57334 117192 57390 117201
rect 57334 117127 57390 117136
rect 57336 115932 57388 115938
rect 57336 115874 57388 115880
rect 57348 115841 57376 115874
rect 57334 115832 57390 115841
rect 57334 115767 57390 115776
rect 57440 113121 57468 164970
rect 57426 113112 57482 113121
rect 57426 113047 57482 113056
rect 57336 112940 57388 112946
rect 57336 112882 57388 112888
rect 57348 30841 57376 112882
rect 57532 110401 57560 167826
rect 57518 110392 57574 110401
rect 57518 110327 57574 110336
rect 57428 108996 57480 109002
rect 57428 108938 57480 108944
rect 57440 107681 57468 108938
rect 57520 108928 57572 108934
rect 57520 108870 57572 108876
rect 57532 108361 57560 108870
rect 57518 108352 57574 108361
rect 57518 108287 57574 108296
rect 57426 107672 57482 107681
rect 57426 107607 57482 107616
rect 57428 104848 57480 104854
rect 57428 104790 57480 104796
rect 57440 103601 57468 104790
rect 57520 104780 57572 104786
rect 57520 104722 57572 104728
rect 57532 104281 57560 104722
rect 57518 104272 57574 104281
rect 57518 104207 57574 104216
rect 57426 103592 57482 103601
rect 57426 103527 57482 103536
rect 57520 103488 57572 103494
rect 57520 103430 57572 103436
rect 57428 103420 57480 103426
rect 57428 103362 57480 103368
rect 57440 102241 57468 103362
rect 57532 102921 57560 103430
rect 57518 102912 57574 102921
rect 57518 102847 57574 102856
rect 57426 102232 57482 102241
rect 57426 102167 57482 102176
rect 57520 100700 57572 100706
rect 57520 100642 57572 100648
rect 57532 99521 57560 100642
rect 57518 99512 57574 99521
rect 57518 99447 57574 99456
rect 57520 97980 57572 97986
rect 57520 97922 57572 97928
rect 57532 96801 57560 97922
rect 57518 96792 57574 96801
rect 57518 96727 57574 96736
rect 57428 96144 57480 96150
rect 57428 96086 57480 96092
rect 57334 30832 57390 30841
rect 57334 30767 57390 30776
rect 57244 22704 57296 22710
rect 57244 22646 57296 22652
rect 57440 19242 57468 96086
rect 57520 95192 57572 95198
rect 57520 95134 57572 95140
rect 57532 94081 57560 95134
rect 57518 94072 57574 94081
rect 57518 94007 57574 94016
rect 57520 93968 57572 93974
rect 57520 93910 57572 93916
rect 57428 19236 57480 19242
rect 57428 19178 57480 19184
rect 57532 19106 57560 93910
rect 57624 82958 57652 178842
rect 57794 169008 57850 169017
rect 57794 168943 57850 168952
rect 57704 159520 57756 159526
rect 57704 159462 57756 159468
rect 57612 82952 57664 82958
rect 57612 82894 57664 82900
rect 57612 82816 57664 82822
rect 57612 82758 57664 82764
rect 57624 82521 57652 82758
rect 57610 82512 57666 82521
rect 57610 82447 57666 82456
rect 57612 75880 57664 75886
rect 57612 75822 57664 75828
rect 57624 75721 57652 75822
rect 57610 75712 57666 75721
rect 57610 75647 57666 75656
rect 57612 69012 57664 69018
rect 57612 68954 57664 68960
rect 57624 68241 57652 68954
rect 57610 68232 57666 68241
rect 57610 68167 57666 68176
rect 57612 68128 57664 68134
rect 57612 68070 57664 68076
rect 57624 19145 57652 68070
rect 57716 63594 57744 159462
rect 57808 63714 57836 168943
rect 57992 155514 58020 195622
rect 58346 195528 58402 195537
rect 58346 195463 58402 195472
rect 57980 155508 58032 155514
rect 57980 155450 58032 155456
rect 58256 153060 58308 153066
rect 58256 153002 58308 153008
rect 57888 151632 57940 151638
rect 57888 151574 57940 151580
rect 57900 145761 57928 151574
rect 58164 151156 58216 151162
rect 58164 151098 58216 151104
rect 57886 145752 57942 145761
rect 57886 145687 57942 145696
rect 57888 142112 57940 142118
rect 57888 142054 57940 142060
rect 57900 141681 57928 142054
rect 57886 141672 57942 141681
rect 57886 141607 57942 141616
rect 57888 140752 57940 140758
rect 57888 140694 57940 140700
rect 57900 140321 57928 140694
rect 57886 140312 57942 140321
rect 57886 140247 57942 140256
rect 57888 137964 57940 137970
rect 57888 137906 57940 137912
rect 57900 137601 57928 137906
rect 57886 137592 57942 137601
rect 57886 137527 57942 137536
rect 57888 135244 57940 135250
rect 57888 135186 57940 135192
rect 57900 134881 57928 135186
rect 57886 134872 57942 134881
rect 57886 134807 57942 134816
rect 57888 133884 57940 133890
rect 57888 133826 57940 133832
rect 57900 132841 57928 133826
rect 57886 132832 57942 132841
rect 57886 132767 57942 132776
rect 57888 132728 57940 132734
rect 57888 132670 57940 132676
rect 57900 132494 57928 132670
rect 57900 132466 58020 132494
rect 57992 128466 58020 132466
rect 57900 128438 58020 128466
rect 57900 121718 57928 128438
rect 57888 121712 57940 121718
rect 57888 121654 57940 121660
rect 57888 121576 57940 121582
rect 57888 121518 57940 121524
rect 57900 114345 57928 121518
rect 57886 114336 57942 114345
rect 57886 114271 57942 114280
rect 57888 108248 57940 108254
rect 57888 108190 57940 108196
rect 57900 97986 57928 108190
rect 57980 98048 58032 98054
rect 57980 97990 58032 97996
rect 57888 97980 57940 97986
rect 57888 97922 57940 97928
rect 57992 97866 58020 97990
rect 57900 97838 58020 97866
rect 57900 93974 57928 97838
rect 57888 93968 57940 93974
rect 57888 93910 57940 93916
rect 57888 93832 57940 93838
rect 57888 93774 57940 93780
rect 57900 92721 57928 93774
rect 57886 92712 57942 92721
rect 57886 92647 57942 92656
rect 57888 91044 57940 91050
rect 57888 90986 57940 90992
rect 57900 90681 57928 90986
rect 57886 90672 57942 90681
rect 57886 90607 57942 90616
rect 57888 89684 57940 89690
rect 57888 89626 57940 89632
rect 57900 89321 57928 89626
rect 57886 89312 57942 89321
rect 57886 89247 57942 89256
rect 57888 82748 57940 82754
rect 57888 82690 57940 82696
rect 57900 81841 57928 82690
rect 57886 81832 57942 81841
rect 57886 81767 57942 81776
rect 57886 64832 57942 64841
rect 57886 64767 57888 64776
rect 57940 64767 57942 64776
rect 57888 64738 57940 64744
rect 57796 63708 57848 63714
rect 57796 63650 57848 63656
rect 57716 63566 57928 63594
rect 57704 63504 57756 63510
rect 57702 63472 57704 63481
rect 57796 63504 57848 63510
rect 57756 63472 57758 63481
rect 57796 63446 57848 63452
rect 57702 63407 57758 63416
rect 57702 62112 57758 62121
rect 57702 62047 57704 62056
rect 57756 62047 57758 62056
rect 57704 62018 57756 62024
rect 57808 59401 57836 63446
rect 57794 59392 57850 59401
rect 57704 59356 57756 59362
rect 57794 59327 57850 59336
rect 57704 59298 57756 59304
rect 57716 58721 57744 59298
rect 57702 58712 57758 58721
rect 57702 58647 57758 58656
rect 57702 57352 57758 57361
rect 57702 57287 57704 57296
rect 57756 57287 57758 57296
rect 57704 57258 57756 57264
rect 57900 56001 57928 63566
rect 57886 55992 57942 56001
rect 57886 55927 57942 55936
rect 57704 53780 57756 53786
rect 57704 53722 57756 53728
rect 57716 53281 57744 53722
rect 57702 53272 57758 53281
rect 57702 53207 57758 53216
rect 57704 48272 57756 48278
rect 57704 48214 57756 48220
rect 57716 47161 57744 48214
rect 57702 47152 57758 47161
rect 57702 47087 57758 47096
rect 58176 45801 58204 151098
rect 58162 45792 58218 45801
rect 58162 45727 58218 45736
rect 58268 41721 58296 153002
rect 58360 45121 58388 195463
rect 60936 195242 60964 200124
rect 61534 200002 61562 200124
rect 60752 195214 60964 195242
rect 61212 199974 61562 200002
rect 58624 191004 58676 191010
rect 58624 190946 58676 190952
rect 58532 190052 58584 190058
rect 58532 189994 58584 190000
rect 58438 138136 58494 138145
rect 58438 138071 58494 138080
rect 58452 114481 58480 138071
rect 58544 131170 58572 189994
rect 58636 147014 58664 190946
rect 58716 190324 58768 190330
rect 58716 190266 58768 190272
rect 58624 147008 58676 147014
rect 58624 146950 58676 146956
rect 58624 142860 58676 142866
rect 58624 142802 58676 142808
rect 58532 131164 58584 131170
rect 58532 131106 58584 131112
rect 58532 127628 58584 127634
rect 58532 127570 58584 127576
rect 58438 114472 58494 114481
rect 58438 114407 58494 114416
rect 58544 97918 58572 127570
rect 58532 97912 58584 97918
rect 58532 97854 58584 97860
rect 58530 89856 58586 89865
rect 58530 89791 58586 89800
rect 58346 45112 58402 45121
rect 58346 45047 58402 45056
rect 58254 41712 58310 41721
rect 58254 41647 58310 41656
rect 57704 41404 57756 41410
rect 57704 41346 57756 41352
rect 57716 41041 57744 41346
rect 57702 41032 57758 41041
rect 57702 40967 57758 40976
rect 57704 40044 57756 40050
rect 57704 39986 57756 39992
rect 57716 39681 57744 39986
rect 57702 39672 57758 39681
rect 57702 39607 57758 39616
rect 57704 34468 57756 34474
rect 57704 34410 57756 34416
rect 57716 33561 57744 34410
rect 57702 33552 57758 33561
rect 57702 33487 57758 33496
rect 57704 33108 57756 33114
rect 57704 33050 57756 33056
rect 57716 32881 57744 33050
rect 57796 33040 57848 33046
rect 57796 32982 57848 32988
rect 57702 32872 57758 32881
rect 57702 32807 57758 32816
rect 57808 32201 57836 32982
rect 57794 32192 57850 32201
rect 57794 32127 57850 32136
rect 57704 31748 57756 31754
rect 57704 31690 57756 31696
rect 57716 31521 57744 31690
rect 57702 31512 57758 31521
rect 57702 31447 57758 31456
rect 58544 28529 58572 89791
rect 58530 28520 58586 28529
rect 58530 28455 58586 28464
rect 57610 19136 57666 19145
rect 57520 19100 57572 19106
rect 57610 19071 57666 19080
rect 57520 19042 57572 19048
rect 56508 18624 56560 18630
rect 56508 18566 56560 18572
rect 58636 17377 58664 142802
rect 58728 141438 58756 190266
rect 59636 190256 59688 190262
rect 59636 190198 59688 190204
rect 59176 190120 59228 190126
rect 59176 190062 59228 190068
rect 59084 187536 59136 187542
rect 59084 187478 59136 187484
rect 58992 187468 59044 187474
rect 58992 187410 59044 187416
rect 58808 184476 58860 184482
rect 58808 184418 58860 184424
rect 58716 141432 58768 141438
rect 58716 141374 58768 141380
rect 58716 124092 58768 124098
rect 58716 124034 58768 124040
rect 58728 118726 58756 124034
rect 58716 118720 58768 118726
rect 58716 118662 58768 118668
rect 58716 113824 58768 113830
rect 58716 113766 58768 113772
rect 58728 21282 58756 113766
rect 58820 108254 58848 184418
rect 58900 154080 58952 154086
rect 58900 154022 58952 154028
rect 58912 151638 58940 154022
rect 58900 151632 58952 151638
rect 58900 151574 58952 151580
rect 58900 134768 58952 134774
rect 58900 134710 58952 134716
rect 58912 124166 58940 134710
rect 59004 126954 59032 187410
rect 59096 147014 59124 187478
rect 59084 147008 59136 147014
rect 59084 146950 59136 146956
rect 59082 146568 59138 146577
rect 59082 146503 59138 146512
rect 59096 134774 59124 146503
rect 59188 146282 59216 190062
rect 59544 189848 59596 189854
rect 59544 189790 59596 189796
rect 59452 184408 59504 184414
rect 59452 184350 59504 184356
rect 59188 146254 59400 146282
rect 59268 146192 59320 146198
rect 59268 146134 59320 146140
rect 59084 134768 59136 134774
rect 59084 134710 59136 134716
rect 59280 132394 59308 146134
rect 59372 142154 59400 146254
rect 59464 146130 59492 184350
rect 59556 150006 59584 189790
rect 59544 150000 59596 150006
rect 59544 149942 59596 149948
rect 59648 149122 59676 190198
rect 59912 190188 59964 190194
rect 59912 190130 59964 190136
rect 59820 189984 59872 189990
rect 59820 189926 59872 189932
rect 59728 184340 59780 184346
rect 59728 184282 59780 184288
rect 59636 149116 59688 149122
rect 59636 149058 59688 149064
rect 59544 147008 59596 147014
rect 59544 146950 59596 146956
rect 59452 146124 59504 146130
rect 59452 146066 59504 146072
rect 59372 142126 59492 142154
rect 59358 140992 59414 141001
rect 59358 140927 59414 140936
rect 59268 132388 59320 132394
rect 59268 132330 59320 132336
rect 59372 131186 59400 140927
rect 59464 135930 59492 142126
rect 59556 140894 59584 146950
rect 59544 140888 59596 140894
rect 59544 140830 59596 140836
rect 59740 140826 59768 184282
rect 59832 146334 59860 189926
rect 59820 146328 59872 146334
rect 59820 146270 59872 146276
rect 59728 140820 59780 140826
rect 59728 140762 59780 140768
rect 59636 136536 59688 136542
rect 59636 136478 59688 136484
rect 59452 135924 59504 135930
rect 59452 135866 59504 135872
rect 59648 132494 59676 136478
rect 59924 132494 59952 190130
rect 60004 151632 60056 151638
rect 60004 151574 60056 151580
rect 60016 150890 60044 151574
rect 60004 150884 60056 150890
rect 60004 150826 60056 150832
rect 60752 150822 60780 195214
rect 61212 180794 61240 199974
rect 64156 198218 64184 200124
rect 67088 199708 67140 199714
rect 67088 199650 67140 199656
rect 64144 198212 64196 198218
rect 64144 198154 64196 198160
rect 65064 198212 65116 198218
rect 65064 198154 65116 198160
rect 63592 198144 63644 198150
rect 63592 198086 63644 198092
rect 60844 180766 61240 180794
rect 60844 166394 60872 180766
rect 60832 166388 60884 166394
rect 60832 166330 60884 166336
rect 61934 152552 61990 152561
rect 61934 152487 61990 152496
rect 61292 152312 61344 152318
rect 61292 152254 61344 152260
rect 60740 150816 60792 150822
rect 60740 150758 60792 150764
rect 61304 149940 61332 152254
rect 61948 149940 61976 152487
rect 63604 149954 63632 198086
rect 65076 196926 65104 198154
rect 65524 198144 65576 198150
rect 65524 198086 65576 198092
rect 65064 196920 65116 196926
rect 65064 196862 65116 196868
rect 64510 159352 64566 159361
rect 64510 159287 64566 159296
rect 63604 149926 63894 149954
rect 64524 149940 64552 159287
rect 65536 150958 65564 198086
rect 66444 179308 66496 179314
rect 66444 179250 66496 179256
rect 65800 152380 65852 152386
rect 65800 152322 65852 152328
rect 65524 150952 65576 150958
rect 65524 150894 65576 150900
rect 65812 149940 65840 152322
rect 66456 149940 66484 179250
rect 67100 149940 67128 199650
rect 67376 198422 67404 200124
rect 67364 198416 67416 198422
rect 67364 198358 67416 198364
rect 68020 180794 68048 200124
rect 68284 197396 68336 197402
rect 68284 197338 68336 197344
rect 67652 180766 68048 180794
rect 67652 180169 67680 180766
rect 67638 180160 67694 180169
rect 67638 180095 67694 180104
rect 68296 152318 68324 197338
rect 69020 195084 69072 195090
rect 69020 195026 69072 195032
rect 68744 152380 68796 152386
rect 68744 152322 68796 152328
rect 68284 152312 68336 152318
rect 68284 152254 68336 152260
rect 68756 149954 68784 152322
rect 68418 149926 68784 149954
rect 69032 149940 69060 195026
rect 70596 180794 70624 200124
rect 71194 200002 71222 200124
rect 71148 199974 71222 200002
rect 71148 197402 71176 199974
rect 72528 197810 72556 200124
rect 72516 197804 72568 197810
rect 72516 197746 72568 197752
rect 71136 197396 71188 197402
rect 71136 197338 71188 197344
rect 73172 195242 73200 200124
rect 73816 198490 73844 200124
rect 73804 198484 73856 198490
rect 73804 198426 73856 198432
rect 73528 195968 73580 195974
rect 73528 195910 73580 195916
rect 73172 195214 73476 195242
rect 73344 195084 73396 195090
rect 73344 195026 73396 195032
rect 70504 180766 70624 180794
rect 69664 178968 69716 178974
rect 69664 178910 69716 178916
rect 69676 152386 69704 178910
rect 69664 152380 69716 152386
rect 69664 152322 69716 152328
rect 70504 151026 70532 180766
rect 73356 175953 73384 195026
rect 73342 175944 73398 175953
rect 73342 175879 73398 175888
rect 73448 154290 73476 195214
rect 73436 154284 73488 154290
rect 73436 154226 73488 154232
rect 72882 152416 72938 152425
rect 72882 152351 72938 152360
rect 70492 151020 70544 151026
rect 70492 150962 70544 150968
rect 72896 149940 72924 152351
rect 73540 149940 73568 195910
rect 74460 195090 74488 200124
rect 75702 200002 75730 200124
rect 75656 199974 75730 200002
rect 75460 199572 75512 199578
rect 75460 199514 75512 199520
rect 74448 195084 74500 195090
rect 74448 195026 74500 195032
rect 74816 155508 74868 155514
rect 74816 155450 74868 155456
rect 74828 149940 74856 155450
rect 75472 149940 75500 199514
rect 75656 198354 75684 199974
rect 75920 199640 75972 199646
rect 75920 199582 75972 199588
rect 75644 198348 75696 198354
rect 75644 198290 75696 198296
rect 75932 149954 75960 199582
rect 77036 180794 77064 200124
rect 77680 195242 77708 200124
rect 76024 180766 77064 180794
rect 77312 195214 77708 195242
rect 76024 151774 76052 180766
rect 77312 166598 77340 195214
rect 78324 180794 78352 200124
rect 78968 180794 78996 200124
rect 79612 197878 79640 200124
rect 79600 197872 79652 197878
rect 79600 197814 79652 197820
rect 80060 195084 80112 195090
rect 80060 195026 80112 195032
rect 77404 180766 78352 180794
rect 78784 180766 78996 180794
rect 77404 177410 77432 180766
rect 77392 177404 77444 177410
rect 77392 177346 77444 177352
rect 78036 174684 78088 174690
rect 78036 174626 78088 174632
rect 77392 171828 77444 171834
rect 77392 171770 77444 171776
rect 77300 166592 77352 166598
rect 77300 166534 77352 166540
rect 76012 151768 76064 151774
rect 76012 151710 76064 151716
rect 75932 149926 76774 149954
rect 77404 149940 77432 171770
rect 78048 149940 78076 174626
rect 78784 157214 78812 180766
rect 79324 173256 79376 173262
rect 79324 173198 79376 173204
rect 78772 157208 78824 157214
rect 78772 157150 78824 157156
rect 79336 149940 79364 173198
rect 80072 153882 80100 195026
rect 80256 190454 80284 200124
rect 80854 200002 80882 200124
rect 80808 199974 80882 200002
rect 80808 195090 80836 199974
rect 82188 196926 82216 200124
rect 82832 197849 82860 200124
rect 82818 197840 82874 197849
rect 82818 197775 82874 197784
rect 83476 197305 83504 200124
rect 84120 198937 84148 200124
rect 85362 200002 85390 200124
rect 85316 199974 85390 200002
rect 84106 198928 84162 198937
rect 84106 198863 84162 198872
rect 85316 197946 85344 199974
rect 85304 197940 85356 197946
rect 85304 197882 85356 197888
rect 83462 197296 83518 197305
rect 83462 197231 83518 197240
rect 82176 196920 82228 196926
rect 82176 196862 82228 196868
rect 85580 195356 85632 195362
rect 85580 195298 85632 195304
rect 85592 195090 85620 195298
rect 86696 195242 86724 200124
rect 87694 195664 87750 195673
rect 87694 195599 87750 195608
rect 85684 195214 86724 195242
rect 80796 195084 80848 195090
rect 80796 195026 80848 195032
rect 85580 195084 85632 195090
rect 85580 195026 85632 195032
rect 80164 190426 80284 190454
rect 80164 157078 80192 190426
rect 85684 190369 85712 195214
rect 86408 195084 86460 195090
rect 86408 195026 86460 195032
rect 85670 190360 85726 190369
rect 85670 190295 85726 190304
rect 81254 188592 81310 188601
rect 81254 188527 81310 188536
rect 80244 182912 80296 182918
rect 80244 182854 80296 182860
rect 80152 157072 80204 157078
rect 80152 157014 80204 157020
rect 80060 153876 80112 153882
rect 80060 153818 80112 153824
rect 80256 149954 80284 182854
rect 80256 149926 80638 149954
rect 81268 149940 81296 188527
rect 85764 186992 85816 186998
rect 85764 186934 85816 186940
rect 84200 170468 84252 170474
rect 84200 170410 84252 170416
rect 81900 166524 81952 166530
rect 81900 166466 81952 166472
rect 81912 149940 81940 166466
rect 82544 152448 82596 152454
rect 82544 152390 82596 152396
rect 82556 149940 82584 152390
rect 84212 149954 84240 170410
rect 84212 149926 85146 149954
rect 85776 149940 85804 186934
rect 86420 149940 86448 195026
rect 87708 149940 87736 195599
rect 88628 180794 88656 200124
rect 89272 194342 89300 200124
rect 89870 200002 89898 200124
rect 89824 199974 89898 200002
rect 89260 194336 89312 194342
rect 89260 194278 89312 194284
rect 88352 180766 88656 180794
rect 88352 175982 88380 180766
rect 88340 175976 88392 175982
rect 88340 175918 88392 175924
rect 89824 153202 89852 199974
rect 90916 198076 90968 198082
rect 90916 198018 90968 198024
rect 88984 153196 89036 153202
rect 88984 153138 89036 153144
rect 89812 153196 89864 153202
rect 89812 153138 89864 153144
rect 88996 149940 89024 153138
rect 90928 149940 90956 198018
rect 91204 180794 91232 200124
rect 91112 180766 91232 180794
rect 91112 154018 91140 180766
rect 92492 158302 92520 200124
rect 93136 198121 93164 200124
rect 94424 198121 94452 200124
rect 93122 198112 93178 198121
rect 93122 198047 93178 198056
rect 94410 198112 94466 198121
rect 94410 198047 94466 198056
rect 96356 180794 96384 200124
rect 97000 195242 97028 200124
rect 95252 180766 96384 180794
rect 96632 195214 97028 195242
rect 95252 176118 95280 180766
rect 95240 176112 95292 176118
rect 95240 176054 95292 176060
rect 92480 158296 92532 158302
rect 92480 158238 92532 158244
rect 91100 154012 91152 154018
rect 91100 153954 91152 153960
rect 93492 152992 93544 152998
rect 93492 152934 93544 152940
rect 94780 152992 94832 152998
rect 94780 152934 94832 152940
rect 93504 149940 93532 152934
rect 94792 149940 94820 152934
rect 96632 151706 96660 195214
rect 97644 180794 97672 200124
rect 100864 198830 100892 200124
rect 100852 198824 100904 198830
rect 100852 198766 100904 198772
rect 101508 198558 101536 200124
rect 101496 198552 101548 198558
rect 101496 198494 101548 198500
rect 102152 194070 102180 200124
rect 104084 199034 104112 200124
rect 104682 200002 104710 200124
rect 104636 199974 104710 200002
rect 104636 199306 104664 199974
rect 104624 199300 104676 199306
rect 104624 199242 104676 199248
rect 104072 199028 104124 199034
rect 104072 198970 104124 198976
rect 106016 198626 106044 200124
rect 106004 198620 106056 198626
rect 106004 198562 106056 198568
rect 102140 194064 102192 194070
rect 102140 194006 102192 194012
rect 106660 180794 106688 200124
rect 108592 190454 108620 200124
rect 108948 199504 109000 199510
rect 108948 199446 109000 199452
rect 96724 180766 97672 180794
rect 106292 180766 106688 180794
rect 107764 190426 108620 190454
rect 96724 172378 96752 180766
rect 99932 180328 99984 180334
rect 99932 180270 99984 180276
rect 98644 177676 98696 177682
rect 98644 177618 98696 177624
rect 96712 172372 96764 172378
rect 96712 172314 96764 172320
rect 96712 160880 96764 160886
rect 96712 160822 96764 160828
rect 96620 151700 96672 151706
rect 96620 151642 96672 151648
rect 96724 149954 96752 160822
rect 96724 149926 97382 149954
rect 98656 149940 98684 177618
rect 99288 153196 99340 153202
rect 99288 153138 99340 153144
rect 99300 149940 99328 153138
rect 99944 149940 99972 180270
rect 103796 170604 103848 170610
rect 103796 170546 103848 170552
rect 103808 149940 103836 170546
rect 106292 154222 106320 180766
rect 107764 167958 107792 190426
rect 108304 183592 108356 183598
rect 108304 183534 108356 183540
rect 107752 167952 107804 167958
rect 107752 167894 107804 167900
rect 106372 157140 106424 157146
rect 106372 157082 106424 157088
rect 106280 154216 106332 154222
rect 106280 154158 106332 154164
rect 106384 149940 106412 157082
rect 107660 153128 107712 153134
rect 107660 153070 107712 153076
rect 107672 149940 107700 153070
rect 108316 149940 108344 183534
rect 108960 149940 108988 199446
rect 111168 198082 111196 200124
rect 111156 198076 111208 198082
rect 111156 198018 111208 198024
rect 111812 195242 111840 200124
rect 111812 195214 111932 195242
rect 111800 195084 111852 195090
rect 111800 195026 111852 195032
rect 110880 162308 110932 162314
rect 110880 162250 110932 162256
rect 110892 149940 110920 162250
rect 111812 151162 111840 195026
rect 111904 151162 111932 195214
rect 112456 180794 112484 200124
rect 113100 195090 113128 200124
rect 113744 198150 113772 200124
rect 114342 200002 114370 200124
rect 114204 199974 114370 200002
rect 113732 198144 113784 198150
rect 113732 198086 113784 198092
rect 113088 195084 113140 195090
rect 113088 195026 113140 195032
rect 114204 180794 114232 199974
rect 116320 198422 116348 200124
rect 116308 198416 116360 198422
rect 116308 198358 116360 198364
rect 116964 194206 116992 200124
rect 118252 198506 118280 200124
rect 118850 199866 118878 200124
rect 118804 199838 118878 199866
rect 118804 199238 118832 199838
rect 118792 199232 118844 199238
rect 118792 199174 118844 199180
rect 117332 198478 118280 198506
rect 116952 194200 117004 194206
rect 116952 194142 117004 194148
rect 116676 191616 116728 191622
rect 116676 191558 116728 191564
rect 116032 187060 116084 187066
rect 116032 187002 116084 187008
rect 111996 180766 112484 180794
rect 113376 180766 114232 180794
rect 111996 174758 112024 180766
rect 111984 174752 112036 174758
rect 111984 174694 112036 174700
rect 113180 169108 113232 169114
rect 113180 169050 113232 169056
rect 112168 153128 112220 153134
rect 112168 153070 112220 153076
rect 111800 151156 111852 151162
rect 111800 151098 111852 151104
rect 111892 151156 111944 151162
rect 111892 151098 111944 151104
rect 112180 149940 112208 153070
rect 113192 149954 113220 169050
rect 113376 151502 113404 180766
rect 113364 151496 113416 151502
rect 113364 151438 113416 151444
rect 113192 149926 114126 149954
rect 116044 149940 116072 187002
rect 116688 149940 116716 191558
rect 117332 151609 117360 198478
rect 117964 198416 118016 198422
rect 117964 198358 118016 198364
rect 117976 157282 118004 198358
rect 120184 195974 120212 200124
rect 120724 198144 120776 198150
rect 120724 198086 120776 198092
rect 120172 195968 120224 195974
rect 120172 195910 120224 195916
rect 119896 177744 119948 177750
rect 119896 177686 119948 177692
rect 117964 157276 118016 157282
rect 117964 157218 118016 157224
rect 117318 151600 117374 151609
rect 117318 151535 117374 151544
rect 119908 149940 119936 177686
rect 120736 153134 120764 198086
rect 121472 196790 121500 200124
rect 122760 197985 122788 200124
rect 123358 199866 123386 200124
rect 123358 199838 123432 199866
rect 122746 197976 122802 197985
rect 122746 197911 122802 197920
rect 123404 197810 123432 199838
rect 123392 197804 123444 197810
rect 123392 197746 123444 197752
rect 121460 196784 121512 196790
rect 121460 196726 121512 196732
rect 121460 191208 121512 191214
rect 121460 191150 121512 191156
rect 120724 153128 120776 153134
rect 120724 153070 120776 153076
rect 121472 149954 121500 191150
rect 124692 180794 124720 200124
rect 127268 199102 127296 200124
rect 127256 199096 127308 199102
rect 127256 199038 127308 199044
rect 127912 195242 127940 200124
rect 128510 199866 128538 200124
rect 128464 199838 128538 199866
rect 127992 195356 128044 195362
rect 127992 195298 128044 195304
rect 124232 180766 124720 180794
rect 126992 195214 127940 195242
rect 124232 153950 124260 180766
rect 124404 170536 124456 170542
rect 124404 170478 124456 170484
rect 124220 153944 124272 153950
rect 124220 153886 124272 153892
rect 121472 149926 122498 149954
rect 124416 149940 124444 170478
rect 125048 152856 125100 152862
rect 125048 152798 125100 152804
rect 125060 149940 125088 152798
rect 126992 151298 127020 195214
rect 128004 194614 128032 195298
rect 128464 195158 128492 199838
rect 129844 198150 129872 200124
rect 133018 199866 133046 200124
rect 133018 199838 133092 199866
rect 133064 199102 133092 199838
rect 133052 199096 133104 199102
rect 133052 199038 133104 199044
rect 134352 198286 134380 200124
rect 134340 198280 134392 198286
rect 134340 198222 134392 198228
rect 129832 198144 129884 198150
rect 129832 198086 129884 198092
rect 128452 195152 128504 195158
rect 128452 195094 128504 195100
rect 127072 194608 127124 194614
rect 127072 194550 127124 194556
rect 127992 194608 128044 194614
rect 127992 194550 128044 194556
rect 126980 151292 127032 151298
rect 126980 151234 127032 151240
rect 127084 149954 127112 194550
rect 137572 190454 137600 200124
rect 138170 199866 138198 200124
rect 138170 199838 138244 199866
rect 138216 198558 138244 199838
rect 138204 198552 138256 198558
rect 138204 198494 138256 198500
rect 141792 196716 141844 196722
rect 141792 196658 141844 196664
rect 139398 192944 139454 192953
rect 139398 192879 139454 192888
rect 136652 190426 137600 190454
rect 135260 184544 135312 184550
rect 135260 184486 135312 184492
rect 130200 174752 130252 174758
rect 130200 174694 130252 174700
rect 129554 153096 129610 153105
rect 129554 153031 129610 153040
rect 127624 152856 127676 152862
rect 127624 152798 127676 152804
rect 127022 149926 127112 149954
rect 127636 149940 127664 152798
rect 129568 149940 129596 153031
rect 130212 149940 130240 174694
rect 135272 149954 135300 184486
rect 136652 155174 136680 190426
rect 137284 184544 137336 184550
rect 137284 184486 137336 184492
rect 136640 155168 136692 155174
rect 136640 155110 136692 155116
rect 135996 153128 136048 153134
rect 135996 153070 136048 153076
rect 135272 149926 135378 149954
rect 136008 149940 136036 153070
rect 137296 149940 137324 184486
rect 139412 149954 139440 192879
rect 141148 155916 141200 155922
rect 141148 155858 141200 155864
rect 139412 149926 139886 149954
rect 141160 149940 141188 155858
rect 141804 149940 141832 196658
rect 142080 192982 142108 200124
rect 147830 199866 147858 200124
rect 147830 199838 147904 199866
rect 147876 198354 147904 199838
rect 147864 198348 147916 198354
rect 147864 198290 147916 198296
rect 142068 192976 142120 192982
rect 142068 192918 142120 192924
rect 146300 191684 146352 191690
rect 146300 191626 146352 191632
rect 145012 167748 145064 167754
rect 145012 167690 145064 167696
rect 142436 165164 142488 165170
rect 142436 165106 142488 165112
rect 142448 149940 142476 165106
rect 145024 149940 145052 167690
rect 145654 152960 145710 152969
rect 145654 152895 145710 152904
rect 145668 149940 145696 152895
rect 146312 149940 146340 191626
rect 147678 184104 147734 184113
rect 147678 184039 147734 184048
rect 146944 172168 146996 172174
rect 146944 172110 146996 172116
rect 146956 149940 146984 172110
rect 147692 149954 147720 184039
rect 150452 160750 150480 200124
rect 151740 195158 151768 200124
rect 153672 198801 153700 200124
rect 153658 198792 153714 198801
rect 153658 198727 153714 198736
rect 150532 195152 150584 195158
rect 150532 195094 150584 195100
rect 151728 195152 151780 195158
rect 151728 195094 151780 195100
rect 150544 180130 150572 195094
rect 151820 192296 151872 192302
rect 151820 192238 151872 192244
rect 150532 180124 150584 180130
rect 150532 180066 150584 180072
rect 150440 160744 150492 160750
rect 150440 160686 150492 160692
rect 150164 158364 150216 158370
rect 150164 158306 150216 158312
rect 147692 149926 148258 149954
rect 150176 149940 150204 158306
rect 151832 149954 151860 192238
rect 154316 185910 154344 200124
rect 154304 185904 154356 185910
rect 154304 185846 154356 185852
rect 155604 180794 155632 200124
rect 156846 199866 156874 200124
rect 156846 199838 156920 199866
rect 156892 198150 156920 199838
rect 156880 198144 156932 198150
rect 156880 198086 156932 198092
rect 158180 195945 158208 200124
rect 158536 198008 158588 198014
rect 158536 197950 158588 197956
rect 158166 195936 158222 195945
rect 158166 195871 158222 195880
rect 157890 189680 157946 189689
rect 157890 189615 157946 189624
rect 154592 180766 155632 180794
rect 154592 153066 154620 180766
rect 155316 159792 155368 159798
rect 155316 159734 155368 159740
rect 154580 153060 154632 153066
rect 154580 153002 154632 153008
rect 153382 152688 153438 152697
rect 153382 152623 153438 152632
rect 151832 149926 152122 149954
rect 153396 149940 153424 152623
rect 155328 149940 155356 159734
rect 157904 149940 157932 189615
rect 158548 149940 158576 197950
rect 158824 180794 158852 200124
rect 160112 199170 160140 200124
rect 160100 199164 160152 199170
rect 160100 199106 160152 199112
rect 160756 195242 160784 200124
rect 160112 195214 160784 195242
rect 159178 181928 159234 181937
rect 159178 181863 159234 181872
rect 158732 180766 158852 180794
rect 158732 151298 158760 180766
rect 158720 151292 158772 151298
rect 158720 151234 158772 151240
rect 159192 149940 159220 181863
rect 160112 153066 160140 195214
rect 161400 195158 161428 200124
rect 160192 195152 160244 195158
rect 160192 195094 160244 195100
rect 161388 195152 161440 195158
rect 161388 195094 161440 195100
rect 160204 155786 160232 195094
rect 163332 180794 163360 200124
rect 165264 195226 165292 200124
rect 167840 198966 167868 200124
rect 167828 198960 167880 198966
rect 167828 198902 167880 198908
rect 168484 198218 168512 200124
rect 168472 198212 168524 198218
rect 168472 198154 168524 198160
rect 169128 195702 169156 200124
rect 169116 195696 169168 195702
rect 169116 195638 169168 195644
rect 165252 195220 165304 195226
rect 165252 195162 165304 195168
rect 169772 193798 169800 200124
rect 170416 198966 170444 200124
rect 170404 198960 170456 198966
rect 170404 198902 170456 198908
rect 169760 193792 169812 193798
rect 169760 193734 169812 193740
rect 172992 192370 173020 200124
rect 172980 192364 173032 192370
rect 172980 192306 173032 192312
rect 173636 190398 173664 200124
rect 174280 199374 174308 200124
rect 174268 199368 174320 199374
rect 174268 199310 174320 199316
rect 174924 198762 174952 200124
rect 175096 199368 175148 199374
rect 175096 199310 175148 199316
rect 175108 198762 175136 199310
rect 174912 198756 174964 198762
rect 174912 198698 174964 198704
rect 175096 198756 175148 198762
rect 175096 198698 175148 198704
rect 173624 190392 173676 190398
rect 173624 190334 173676 190340
rect 172058 188864 172114 188873
rect 172058 188799 172114 188808
rect 170772 181960 170824 181966
rect 170772 181902 170824 181908
rect 162872 180766 163360 180794
rect 161756 167952 161808 167958
rect 161756 167894 161808 167900
rect 160192 155780 160244 155786
rect 160192 155722 160244 155728
rect 160100 153060 160152 153066
rect 160100 153002 160152 153008
rect 161768 149940 161796 167894
rect 162872 155854 162900 180766
rect 166264 178696 166316 178702
rect 166264 178638 166316 178644
rect 163044 172236 163096 172242
rect 163044 172178 163096 172184
rect 162860 155848 162912 155854
rect 162860 155790 162912 155796
rect 163056 149940 163084 172178
rect 166276 153134 166304 178638
rect 166908 154012 166960 154018
rect 166908 153954 166960 153960
rect 166264 153128 166316 153134
rect 166264 153070 166316 153076
rect 166920 149940 166948 153954
rect 170126 152824 170182 152833
rect 170126 152759 170182 152768
rect 170140 149940 170168 152759
rect 170784 149940 170812 181902
rect 172072 149940 172100 188799
rect 176660 184680 176712 184686
rect 176660 184622 176712 184628
rect 174636 181484 174688 181490
rect 174636 181426 174688 181432
rect 174648 149940 174676 181426
rect 175924 173324 175976 173330
rect 175924 173266 175976 173272
rect 175280 155916 175332 155922
rect 175280 155858 175332 155864
rect 175292 149940 175320 155858
rect 175936 149940 175964 173266
rect 176672 149954 176700 184622
rect 178788 180794 178816 200124
rect 180076 198098 180104 200124
rect 178052 180766 178816 180794
rect 179432 198070 180104 198098
rect 178052 154018 178080 180766
rect 179432 155786 179460 198070
rect 180064 198008 180116 198014
rect 180064 197950 180116 197956
rect 180076 180794 180104 197950
rect 180720 191758 180748 200124
rect 181318 199866 181346 200124
rect 181318 199838 181392 199866
rect 181364 194138 181392 199838
rect 182652 195702 182680 200124
rect 183008 196648 183060 196654
rect 183008 196590 183060 196596
rect 182640 195696 182692 195702
rect 182640 195638 182692 195644
rect 181352 194132 181404 194138
rect 181352 194074 181404 194080
rect 180708 191752 180760 191758
rect 180708 191694 180760 191700
rect 179800 180766 180104 180794
rect 179420 155780 179472 155786
rect 179420 155722 179472 155728
rect 178040 154012 178092 154018
rect 178040 153954 178092 153960
rect 179142 152688 179198 152697
rect 179142 152623 179198 152632
rect 176672 149926 177238 149954
rect 179156 149940 179184 152623
rect 179800 149940 179828 180766
rect 180800 174888 180852 174894
rect 180800 174830 180852 174836
rect 180812 149954 180840 174830
rect 180812 149926 181746 149954
rect 183020 149940 183048 196590
rect 183940 191758 183968 200124
rect 183928 191752 183980 191758
rect 183928 191694 183980 191700
rect 184584 189718 184612 200124
rect 185826 199866 185854 200124
rect 185320 199838 185854 199866
rect 184572 189712 184624 189718
rect 184572 189654 184624 189660
rect 185320 180794 185348 199838
rect 187804 199238 187832 200124
rect 187792 199232 187844 199238
rect 187792 199174 187844 199180
rect 189092 195838 189120 200124
rect 190334 199866 190362 200124
rect 190334 199838 190408 199866
rect 190380 198218 190408 199838
rect 190368 198212 190420 198218
rect 190368 198154 190420 198160
rect 189080 195832 189132 195838
rect 189080 195774 189132 195780
rect 192956 195242 192984 200124
rect 194244 195838 194272 200124
rect 194232 195832 194284 195838
rect 194232 195774 194284 195780
rect 194888 195634 194916 200124
rect 195486 199866 195514 200124
rect 195164 199838 195514 199866
rect 194876 195628 194928 195634
rect 194876 195570 194928 195576
rect 191852 195214 192984 195242
rect 187516 187604 187568 187610
rect 187516 187546 187568 187552
rect 184952 180766 185348 180794
rect 184952 156670 184980 180766
rect 184940 156664 184992 156670
rect 184940 156606 184992 156612
rect 187528 149940 187556 187546
rect 188160 176452 188212 176458
rect 188160 176394 188212 176400
rect 188172 149940 188200 176394
rect 191852 169182 191880 195214
rect 192024 192364 192076 192370
rect 192024 192306 192076 192312
rect 191840 169176 191892 169182
rect 191840 169118 191892 169124
rect 188804 153060 188856 153066
rect 188804 153002 188856 153008
rect 188816 149940 188844 153002
rect 192036 149940 192064 192306
rect 195164 188902 195192 199838
rect 196820 196994 196848 200124
rect 196808 196988 196860 196994
rect 196808 196930 196860 196936
rect 197464 195242 197492 200124
rect 197372 195214 197492 195242
rect 195152 188896 195204 188902
rect 195152 188838 195204 188844
rect 197372 178974 197400 195214
rect 198108 189650 198136 200124
rect 198096 189644 198148 189650
rect 198096 189586 198148 189592
rect 197360 178968 197412 178974
rect 197360 178910 197412 178916
rect 193220 172304 193272 172310
rect 193220 172246 193272 172252
rect 193232 149954 193260 172246
rect 195244 170740 195296 170746
rect 195244 170682 195296 170688
rect 193232 149926 193982 149954
rect 195256 149940 195284 170682
rect 198752 152930 198780 200124
rect 199994 199866 200022 200124
rect 199994 199838 200068 199866
rect 200040 195673 200068 199838
rect 200764 198348 200816 198354
rect 200764 198290 200816 198296
rect 200026 195664 200082 195673
rect 200026 195599 200082 195608
rect 200120 195220 200172 195226
rect 200120 195162 200172 195168
rect 199752 183184 199804 183190
rect 199752 183126 199804 183132
rect 198740 152924 198792 152930
rect 198740 152866 198792 152872
rect 197174 152824 197230 152833
rect 197174 152759 197230 152768
rect 197188 149940 197216 152759
rect 199108 151836 199160 151842
rect 199108 151778 199160 151784
rect 199120 149940 199148 151778
rect 199764 149940 199792 183126
rect 200132 156942 200160 195162
rect 200776 163742 200804 198290
rect 201328 195226 201356 200124
rect 201972 198422 202000 200124
rect 201960 198416 202012 198422
rect 201960 198358 202012 198364
rect 201316 195220 201368 195226
rect 201316 195162 201368 195168
rect 204548 192302 204576 200124
rect 205146 199866 205174 200124
rect 205146 199838 205220 199866
rect 205192 194342 205220 199838
rect 208412 199170 208440 200124
rect 209654 200002 209682 200124
rect 209608 199974 209682 200002
rect 208400 199164 208452 199170
rect 208400 199106 208452 199112
rect 208124 196648 208176 196654
rect 208124 196590 208176 196596
rect 205180 194336 205232 194342
rect 205180 194278 205232 194284
rect 204536 192296 204588 192302
rect 204536 192238 204588 192244
rect 201500 188896 201552 188902
rect 201500 188838 201552 188844
rect 200764 163736 200816 163742
rect 200764 163678 200816 163684
rect 201408 159656 201460 159662
rect 201408 159598 201460 159604
rect 200120 156936 200172 156942
rect 200120 156878 200172 156884
rect 201420 152998 201448 159598
rect 201408 152992 201460 152998
rect 201408 152934 201460 152940
rect 200396 152924 200448 152930
rect 200396 152866 200448 152872
rect 200408 149940 200436 152866
rect 201512 149954 201540 188838
rect 205640 174820 205692 174826
rect 205640 174762 205692 174768
rect 204260 158092 204312 158098
rect 204260 158034 204312 158040
rect 202972 152788 203024 152794
rect 202972 152730 203024 152736
rect 201512 149926 202354 149954
rect 202984 149940 203012 152730
rect 204272 149940 204300 158034
rect 204904 155712 204956 155718
rect 204904 155654 204956 155660
rect 204916 149940 204944 155654
rect 205652 149954 205680 174762
rect 207480 173392 207532 173398
rect 207480 173334 207532 173340
rect 205652 149926 206862 149954
rect 207492 149940 207520 173334
rect 208136 149940 208164 196590
rect 209608 195226 209636 199974
rect 210988 195226 211016 200124
rect 208400 195220 208452 195226
rect 208400 195162 208452 195168
rect 209596 195220 209648 195226
rect 209596 195162 209648 195168
rect 209780 195220 209832 195226
rect 209780 195162 209832 195168
rect 210976 195220 211028 195226
rect 210976 195162 211028 195168
rect 208412 155242 208440 195162
rect 209412 191072 209464 191078
rect 209412 191014 209464 191020
rect 208400 155236 208452 155242
rect 208400 155178 208452 155184
rect 208768 152652 208820 152658
rect 208768 152594 208820 152600
rect 208780 149940 208808 152594
rect 209424 149940 209452 191014
rect 209792 152726 209820 195162
rect 209872 185904 209924 185910
rect 209872 185846 209924 185852
rect 209780 152720 209832 152726
rect 209780 152662 209832 152668
rect 209884 149954 209912 185846
rect 213564 180794 213592 200124
rect 214806 200002 214834 200124
rect 214300 199974 214834 200002
rect 214300 195242 214328 199974
rect 212552 180766 213592 180794
rect 214024 195214 214328 195242
rect 211988 177812 212040 177818
rect 211988 177754 212040 177760
rect 209884 149926 210726 149954
rect 212000 149940 212028 177754
rect 212552 156738 212580 180766
rect 214024 168094 214052 195214
rect 214104 195152 214156 195158
rect 214104 195094 214156 195100
rect 214012 168088 214064 168094
rect 214012 168030 214064 168036
rect 213276 166592 213328 166598
rect 213276 166534 213328 166540
rect 212540 156732 212592 156738
rect 212540 156674 212592 156680
rect 213288 149940 213316 166534
rect 213918 152960 213974 152969
rect 213918 152895 213974 152904
rect 213932 149940 213960 152895
rect 214116 149954 214144 195094
rect 216140 192438 216168 200124
rect 216128 192432 216180 192438
rect 216128 192374 216180 192380
rect 216784 180794 216812 200124
rect 220360 183116 220412 183122
rect 220360 183058 220412 183064
rect 216692 180766 216812 180794
rect 216496 162376 216548 162382
rect 216496 162318 216548 162324
rect 214116 149926 215234 149954
rect 216508 149940 216536 162318
rect 216692 155242 216720 180766
rect 217784 180464 217836 180470
rect 217784 180406 217836 180412
rect 216680 155236 216732 155242
rect 216680 155178 216732 155184
rect 217796 149940 217824 180406
rect 219716 158092 219768 158098
rect 219716 158034 219768 158040
rect 219728 149940 219756 158034
rect 220372 149940 220400 183058
rect 221292 180794 221320 200124
rect 221936 198898 221964 200124
rect 221924 198892 221976 198898
rect 221924 198834 221976 198840
rect 221648 196716 221700 196722
rect 221648 196658 221700 196664
rect 220832 180766 221320 180794
rect 220832 155718 220860 180766
rect 220820 155712 220872 155718
rect 220820 155654 220872 155660
rect 221660 149940 221688 196658
rect 222580 195242 222608 200124
rect 223868 198490 223896 200124
rect 223856 198484 223908 198490
rect 223856 198426 223908 198432
rect 222212 195214 222608 195242
rect 222212 151502 222240 195214
rect 222292 195152 222344 195158
rect 222292 195094 222344 195100
rect 222200 151496 222252 151502
rect 222200 151438 222252 151444
rect 222304 149940 222332 195094
rect 226156 188828 226208 188834
rect 226156 188770 226208 188776
rect 225512 180532 225564 180538
rect 225512 180474 225564 180480
rect 224868 163532 224920 163538
rect 224868 163474 224920 163480
rect 224224 154284 224276 154290
rect 224224 154226 224276 154232
rect 224236 149940 224264 154226
rect 224880 149940 224908 163474
rect 225524 149940 225552 180474
rect 226168 149940 226196 188770
rect 226444 180794 226472 200124
rect 227732 196897 227760 200124
rect 227718 196888 227774 196897
rect 227718 196823 227774 196832
rect 228376 195809 228404 200124
rect 228456 197532 228508 197538
rect 228456 197474 228508 197480
rect 228362 195800 228418 195809
rect 228362 195735 228418 195744
rect 228468 180794 228496 197474
rect 230952 192846 230980 200124
rect 230940 192840 230992 192846
rect 230940 192782 230992 192788
rect 232240 180794 232268 200124
rect 232884 197538 232912 200124
rect 233482 199866 233510 200124
rect 233482 199838 233556 199866
rect 233528 198898 233556 199838
rect 233516 198892 233568 198898
rect 233516 198834 233568 198840
rect 232872 197532 232924 197538
rect 232872 197474 232924 197480
rect 236748 190330 236776 200124
rect 238634 200002 238662 200124
rect 238588 199974 238662 200002
rect 238588 195226 238616 199974
rect 239968 195226 239996 200124
rect 237380 195220 237432 195226
rect 237380 195162 237432 195168
rect 238576 195220 238628 195226
rect 238576 195162 238628 195168
rect 238760 195220 238812 195226
rect 238760 195162 238812 195168
rect 239956 195220 240008 195226
rect 239956 195162 240008 195168
rect 236736 190324 236788 190330
rect 236736 190266 236788 190272
rect 226352 180766 226472 180794
rect 228376 180766 228496 180794
rect 231964 180766 232268 180794
rect 226352 151638 226380 180766
rect 228376 166530 228404 180766
rect 228732 168020 228784 168026
rect 228732 167962 228784 167968
rect 228364 166524 228416 166530
rect 228364 166466 228416 166472
rect 227720 163668 227772 163674
rect 227720 163610 227772 163616
rect 226800 159860 226852 159866
rect 226800 159802 226852 159808
rect 226340 151632 226392 151638
rect 226340 151574 226392 151580
rect 226812 149940 226840 159802
rect 227732 149954 227760 163610
rect 227732 149926 228114 149954
rect 228744 149940 228772 167962
rect 231964 156874 231992 180766
rect 235172 180396 235224 180402
rect 235172 180338 235224 180344
rect 234528 178968 234580 178974
rect 234528 178910 234580 178916
rect 233884 166524 233936 166530
rect 233884 166466 233936 166472
rect 231952 156868 232004 156874
rect 231952 156810 232004 156816
rect 232596 155848 232648 155854
rect 232596 155790 232648 155796
rect 229376 155780 229428 155786
rect 229376 155722 229428 155728
rect 230020 155780 230072 155786
rect 230020 155722 230072 155728
rect 229388 149940 229416 155722
rect 230032 149940 230060 155722
rect 232608 149940 232636 155790
rect 233896 149940 233924 166466
rect 234540 149940 234568 178910
rect 235184 149940 235212 180338
rect 237392 173330 237420 195162
rect 237746 182064 237802 182073
rect 237746 181999 237802 182008
rect 237380 173324 237432 173330
rect 237380 173266 237432 173272
rect 237760 149940 237788 181999
rect 238772 154154 238800 195162
rect 241256 193934 241284 200124
rect 243142 200002 243170 200124
rect 243096 199974 243170 200002
rect 243096 195566 243124 199974
rect 244476 196994 244504 200124
rect 244464 196988 244516 196994
rect 244464 196930 244516 196936
rect 243084 195560 243136 195566
rect 243084 195502 243136 195508
rect 241244 193928 241296 193934
rect 241244 193870 241296 193876
rect 246408 193730 246436 200124
rect 247052 198801 247080 200124
rect 247038 198792 247094 198801
rect 247038 198727 247094 198736
rect 247696 195498 247724 200124
rect 249628 195634 249656 200124
rect 252802 200002 252830 200124
rect 252572 199974 252830 200002
rect 249616 195628 249668 195634
rect 249616 195570 249668 195576
rect 247684 195492 247736 195498
rect 247684 195434 247736 195440
rect 246396 193724 246448 193730
rect 246396 193666 246448 193672
rect 248420 193724 248472 193730
rect 248420 193666 248472 193672
rect 242900 190324 242952 190330
rect 242900 190266 242952 190272
rect 239036 186924 239088 186930
rect 239036 186866 239088 186872
rect 238760 154148 238812 154154
rect 238760 154090 238812 154096
rect 239048 149940 239076 186866
rect 241612 173460 241664 173466
rect 241612 173402 241664 173408
rect 240140 166456 240192 166462
rect 240140 166398 240192 166404
rect 240152 149954 240180 166398
rect 240968 155644 241020 155650
rect 240968 155586 241020 155592
rect 240152 149926 240350 149954
rect 240980 149940 241008 155586
rect 241624 149940 241652 173402
rect 242256 172372 242308 172378
rect 242256 172314 242308 172320
rect 242268 149940 242296 172314
rect 242912 149940 242940 190266
rect 246120 185972 246172 185978
rect 246120 185914 246172 185920
rect 245476 170672 245528 170678
rect 245476 170614 245528 170620
rect 245488 149940 245516 170614
rect 246132 149940 246160 185914
rect 248432 149954 248460 193666
rect 249984 189576 250036 189582
rect 249984 189518 250036 189524
rect 249340 187672 249392 187678
rect 249340 187614 249392 187620
rect 248432 149926 248722 149954
rect 249352 149940 249380 187614
rect 249996 149940 250024 189518
rect 250628 167952 250680 167958
rect 250628 167894 250680 167900
rect 250640 149940 250668 167894
rect 251272 165232 251324 165238
rect 251272 165174 251324 165180
rect 251284 149940 251312 165174
rect 251916 154828 251968 154834
rect 251916 154770 251968 154776
rect 251928 149940 251956 154770
rect 252572 151638 252600 199974
rect 254780 180794 254808 200124
rect 256068 190262 256096 200124
rect 257954 199866 257982 200124
rect 257908 199838 257982 199866
rect 257908 199209 257936 199838
rect 257986 199608 258042 199617
rect 257986 199543 258042 199552
rect 258000 199238 258028 199543
rect 257988 199232 258040 199238
rect 257894 199200 257950 199209
rect 257988 199174 258040 199180
rect 257894 199135 257950 199144
rect 259000 196580 259052 196586
rect 259000 196522 259052 196528
rect 256056 190256 256108 190262
rect 256056 190198 256108 190204
rect 255780 188692 255832 188698
rect 255780 188634 255832 188640
rect 253952 180766 254808 180794
rect 253952 157010 253980 180766
rect 254492 174956 254544 174962
rect 254492 174898 254544 174904
rect 253940 157004 253992 157010
rect 253940 156946 253992 156952
rect 252652 155712 252704 155718
rect 252652 155654 252704 155660
rect 252560 151632 252612 151638
rect 252560 151574 252612 151580
rect 252664 149954 252692 155654
rect 252664 149926 253230 149954
rect 254504 149940 254532 174898
rect 255792 149940 255820 188634
rect 259012 149940 259040 196522
rect 259460 195220 259512 195226
rect 259460 195162 259512 195168
rect 259472 154834 259500 195162
rect 259932 180794 259960 200124
rect 260576 195226 260604 200124
rect 262462 199866 262490 200124
rect 262462 199838 262536 199866
rect 262508 197946 262536 199838
rect 262496 197940 262548 197946
rect 262496 197882 262548 197888
rect 260564 195220 260616 195226
rect 260564 195162 260616 195168
rect 263796 192778 263824 200124
rect 265624 197940 265676 197946
rect 265624 197882 265676 197888
rect 263784 192772 263836 192778
rect 263784 192714 263836 192720
rect 264152 186856 264204 186862
rect 264152 186798 264204 186804
rect 260840 185768 260892 185774
rect 260840 185710 260892 185716
rect 259564 180766 259960 180794
rect 259564 162246 259592 180766
rect 259644 170808 259696 170814
rect 259644 170750 259696 170756
rect 259552 162240 259604 162246
rect 259552 162182 259604 162188
rect 259460 154828 259512 154834
rect 259460 154770 259512 154776
rect 259656 149940 259684 170750
rect 260288 154148 260340 154154
rect 260288 154090 260340 154096
rect 260300 149940 260328 154090
rect 260852 149954 260880 185710
rect 260852 149926 261602 149954
rect 264164 149940 264192 186798
rect 265636 158506 265664 197882
rect 266084 186040 266136 186046
rect 266084 185982 266136 185988
rect 265624 158500 265676 158506
rect 265624 158442 265676 158448
rect 266096 149940 266124 185982
rect 266372 162450 266400 200124
rect 266970 200002 266998 200124
rect 266924 199974 266998 200002
rect 266924 195430 266952 199974
rect 266912 195424 266964 195430
rect 266912 195366 266964 195372
rect 268660 185768 268712 185774
rect 268660 185710 268712 185716
rect 266360 162444 266412 162450
rect 266360 162386 266412 162392
rect 268016 155168 268068 155174
rect 268016 155110 268068 155116
rect 268028 149940 268056 155110
rect 268672 149940 268700 185710
rect 270236 180794 270264 200124
rect 271524 199238 271552 200124
rect 272122 200002 272150 200124
rect 271984 199974 272150 200002
rect 271512 199232 271564 199238
rect 271512 199174 271564 199180
rect 270590 190088 270646 190097
rect 270590 190023 270646 190032
rect 269132 180766 270264 180794
rect 269132 155650 269160 180766
rect 269120 155644 269172 155650
rect 269120 155586 269172 155592
rect 270604 149940 270632 190023
rect 271880 184612 271932 184618
rect 271880 184554 271932 184560
rect 271236 166456 271288 166462
rect 271236 166398 271288 166404
rect 271248 149940 271276 166398
rect 271892 149940 271920 184554
rect 271984 168162 272012 199974
rect 272524 188896 272576 188902
rect 272524 188838 272576 188844
rect 271972 168156 272024 168162
rect 271972 168098 272024 168104
rect 272536 149940 272564 188838
rect 273456 180794 273484 200124
rect 275388 196790 275416 200124
rect 275376 196784 275428 196790
rect 275376 196726 275428 196732
rect 276032 196450 276060 200124
rect 276630 199866 276658 200124
rect 276630 199838 276704 199866
rect 276020 196444 276072 196450
rect 276020 196386 276072 196392
rect 276676 195566 276704 199838
rect 276664 195560 276716 195566
rect 276664 195502 276716 195508
rect 278608 192846 278636 200124
rect 278596 192840 278648 192846
rect 278596 192782 278648 192788
rect 275742 188728 275798 188737
rect 275742 188663 275798 188672
rect 273272 180766 273484 180794
rect 273272 166598 273300 180766
rect 274456 169176 274508 169182
rect 274456 169118 274508 169124
rect 273260 166592 273312 166598
rect 273260 166534 273312 166540
rect 274468 149940 274496 169118
rect 275756 149940 275784 188663
rect 279252 180794 279280 200124
rect 280540 192778 280568 200124
rect 281184 194002 281212 200124
rect 281782 199866 281810 200124
rect 281736 199838 281810 199866
rect 281172 193996 281224 194002
rect 281172 193938 281224 193944
rect 281736 193662 281764 199838
rect 281724 193656 281776 193662
rect 281724 193598 281776 193604
rect 280528 192772 280580 192778
rect 280528 192714 280580 192720
rect 283116 180794 283144 200124
rect 287624 198354 287652 200124
rect 287612 198348 287664 198354
rect 287612 198290 287664 198296
rect 283564 198144 283616 198150
rect 283564 198086 283616 198092
rect 278792 180766 279280 180794
rect 282932 180766 283144 180794
rect 277400 163804 277452 163810
rect 277400 163746 277452 163752
rect 277412 149954 277440 163746
rect 278792 162314 278820 180766
rect 279608 170672 279660 170678
rect 279608 170614 279660 170620
rect 278964 166592 279016 166598
rect 278964 166534 279016 166540
rect 278780 162308 278832 162314
rect 278780 162250 278832 162256
rect 277412 149926 278346 149954
rect 278976 149940 279004 166534
rect 279620 149940 279648 170614
rect 282932 162314 282960 180766
rect 283472 172304 283524 172310
rect 283472 172246 283524 172252
rect 282920 162308 282972 162314
rect 282920 162250 282972 162256
rect 282828 159248 282880 159254
rect 282828 159190 282880 159196
rect 281540 157072 281592 157078
rect 281540 157014 281592 157020
rect 281552 149954 281580 157014
rect 281552 149926 282210 149954
rect 282840 149940 282868 159190
rect 283484 149940 283512 172246
rect 283576 156602 283604 198086
rect 285404 195424 285456 195430
rect 285404 195366 285456 195372
rect 284760 182028 284812 182034
rect 284760 181970 284812 181976
rect 283564 156596 283616 156602
rect 283564 156538 283616 156544
rect 284116 155576 284168 155582
rect 284116 155518 284168 155524
rect 284128 149940 284156 155518
rect 284772 149940 284800 181970
rect 285416 149940 285444 195366
rect 287704 190256 287756 190262
rect 287704 190198 287756 190204
rect 285680 177880 285732 177886
rect 285680 177822 285732 177828
rect 285692 149954 285720 177822
rect 287716 152561 287744 190198
rect 290844 180794 290872 200124
rect 291442 200002 291470 200124
rect 289832 180766 290872 180794
rect 291212 199974 291470 200002
rect 289268 158432 289320 158438
rect 289268 158374 289320 158380
rect 289280 152862 289308 158374
rect 289832 155922 289860 180766
rect 289820 155916 289872 155922
rect 289820 155858 289872 155864
rect 291212 155718 291240 199974
rect 292776 180794 292804 200124
rect 294064 195242 294092 200124
rect 293972 195214 294092 195242
rect 293972 184686 294000 195214
rect 294708 190194 294736 200124
rect 295352 199073 295380 200124
rect 296074 199472 296130 199481
rect 296074 199407 296130 199416
rect 295338 199064 295394 199073
rect 295338 198999 295394 199008
rect 296088 198966 296116 199407
rect 296076 198960 296128 198966
rect 296076 198902 296128 198908
rect 295708 193656 295760 193662
rect 295708 193598 295760 193604
rect 294696 190188 294748 190194
rect 294696 190130 294748 190136
rect 293960 184680 294012 184686
rect 293960 184622 294012 184628
rect 293132 183116 293184 183122
rect 293132 183058 293184 183064
rect 292592 180766 292804 180794
rect 292592 169182 292620 180766
rect 292580 169176 292632 169182
rect 292580 169118 292632 169124
rect 291200 155712 291252 155718
rect 291200 155654 291252 155660
rect 292486 153096 292542 153105
rect 292486 153031 292542 153040
rect 289268 152856 289320 152862
rect 289268 152798 289320 152804
rect 287980 152652 288032 152658
rect 287980 152594 288032 152600
rect 287702 152552 287758 152561
rect 287702 152487 287758 152496
rect 285692 149926 286718 149954
rect 287992 149940 288020 152594
rect 291198 152552 291254 152561
rect 291198 152487 291254 152496
rect 291212 149940 291240 152487
rect 292500 149940 292528 153031
rect 293144 149940 293172 183058
rect 295720 149940 295748 193598
rect 297928 191554 297956 200124
rect 297916 191548 297968 191554
rect 297916 191490 297968 191496
rect 299860 180794 299888 200124
rect 300458 199866 300486 200124
rect 300458 199838 300532 199866
rect 300504 198966 300532 199838
rect 300492 198960 300544 198966
rect 300492 198902 300544 198908
rect 300860 186788 300912 186794
rect 300860 186730 300912 186736
rect 299492 180766 299888 180794
rect 296352 154352 296404 154358
rect 296352 154294 296404 154300
rect 296364 149940 296392 154294
rect 299492 154154 299520 180766
rect 299480 154148 299532 154154
rect 299480 154090 299532 154096
rect 297640 152584 297692 152590
rect 297640 152526 297692 152532
rect 297652 149940 297680 152526
rect 300872 149940 300900 186730
rect 301792 180794 301820 200124
rect 302148 189644 302200 189650
rect 302148 189586 302200 189592
rect 301056 180766 301820 180794
rect 301056 179382 301084 180766
rect 301044 179376 301096 179382
rect 301044 179318 301096 179324
rect 302160 149940 302188 189586
rect 303080 180794 303108 200124
rect 303724 188766 303752 200124
rect 304368 195498 304396 200124
rect 304356 195492 304408 195498
rect 304356 195434 304408 195440
rect 305012 195242 305040 200124
rect 305610 200002 305638 200124
rect 305564 199974 305638 200002
rect 305012 195214 305132 195242
rect 305000 195152 305052 195158
rect 305000 195094 305052 195100
rect 303712 188760 303764 188766
rect 303712 188702 303764 188708
rect 302252 180766 303108 180794
rect 302252 155582 302280 180766
rect 302240 155576 302292 155582
rect 302240 155518 302292 155524
rect 305012 154154 305040 195094
rect 305104 159730 305132 195214
rect 305564 195158 305592 199974
rect 305552 195152 305604 195158
rect 305552 195094 305604 195100
rect 306944 180794 306972 200124
rect 310118 200002 310146 200124
rect 309612 199974 310146 200002
rect 309612 180794 309640 199974
rect 310704 197396 310756 197402
rect 310704 197338 310756 197344
rect 310716 196858 310744 197338
rect 312740 196858 312768 200124
rect 310704 196852 310756 196858
rect 310704 196794 310756 196800
rect 312728 196852 312780 196858
rect 312728 196794 312780 196800
rect 314028 191010 314056 200124
rect 315270 199866 315298 200124
rect 315270 199838 315344 199866
rect 315316 195226 315344 199838
rect 317248 199374 317276 200124
rect 317236 199368 317288 199374
rect 317236 199310 317288 199316
rect 317892 197878 317920 200124
rect 319778 199866 319806 200124
rect 319778 199838 319852 199866
rect 319824 197946 319852 199838
rect 319812 197940 319864 197946
rect 319812 197882 319864 197888
rect 317880 197872 317932 197878
rect 317880 197814 317932 197820
rect 315304 195220 315356 195226
rect 315304 195162 315356 195168
rect 314016 191004 314068 191010
rect 314016 190946 314068 190952
rect 318248 184680 318300 184686
rect 318248 184622 318300 184628
rect 306392 180766 306972 180794
rect 309152 180766 309640 180794
rect 305092 159724 305144 159730
rect 305092 159666 305144 159672
rect 306392 157078 306420 180766
rect 306472 173528 306524 173534
rect 306472 173470 306524 173476
rect 306380 157072 306432 157078
rect 306380 157014 306432 157020
rect 305000 154148 305052 154154
rect 305000 154090 305052 154096
rect 306484 149954 306512 173470
rect 309152 170814 309180 180766
rect 312452 176520 312504 176526
rect 312452 176462 312504 176468
rect 309140 170808 309192 170814
rect 309140 170750 309192 170756
rect 309876 168156 309928 168162
rect 309876 168098 309928 168104
rect 307944 166388 307996 166394
rect 307944 166330 307996 166336
rect 306484 149926 307326 149954
rect 307956 149940 307984 166330
rect 308588 154216 308640 154222
rect 308588 154158 308640 154164
rect 308600 149940 308628 154158
rect 309232 152584 309284 152590
rect 309232 152526 309284 152532
rect 309244 149940 309272 152526
rect 309888 149940 309916 168098
rect 310520 152788 310572 152794
rect 310520 152730 310572 152736
rect 310532 149940 310560 152730
rect 312464 149940 312492 176462
rect 314384 176384 314436 176390
rect 314384 176326 314436 176332
rect 313094 175808 313150 175817
rect 313094 175743 313150 175752
rect 313108 149940 313136 175743
rect 313740 170808 313792 170814
rect 313740 170750 313792 170756
rect 313752 149940 313780 170750
rect 314396 149940 314424 176326
rect 316592 152992 316644 152998
rect 316592 152934 316644 152940
rect 315028 152720 315080 152726
rect 315028 152662 315080 152668
rect 315040 149940 315068 152662
rect 316604 149954 316632 152934
rect 317602 152280 317658 152289
rect 317602 152215 317658 152224
rect 316358 149926 316632 149954
rect 317616 149940 317644 152215
rect 318260 149940 318288 184622
rect 321112 180794 321140 200124
rect 322112 190188 322164 190194
rect 322112 190130 322164 190136
rect 320192 180766 321140 180794
rect 318892 174752 318944 174758
rect 318892 174694 318944 174700
rect 318904 149940 318932 174694
rect 320192 160954 320220 180766
rect 321468 169312 321520 169318
rect 321468 169254 321520 169260
rect 320180 160948 320232 160954
rect 320180 160890 320232 160896
rect 320824 158296 320876 158302
rect 320824 158238 320876 158244
rect 320836 149940 320864 158238
rect 321480 149940 321508 169254
rect 322124 149940 322152 190130
rect 323400 157208 323452 157214
rect 323400 157150 323452 157156
rect 322756 155644 322808 155650
rect 322756 155586 322808 155592
rect 322768 149940 322796 155586
rect 323412 149940 323440 157150
rect 324332 151706 324360 200124
rect 324930 200002 324958 200124
rect 324424 199974 324958 200002
rect 324424 188834 324452 199974
rect 326908 192642 326936 200124
rect 326988 199436 327040 199442
rect 326988 199378 327040 199384
rect 327000 198694 327028 199378
rect 326988 198688 327040 198694
rect 326988 198630 327040 198636
rect 326896 192636 326948 192642
rect 326896 192578 326948 192584
rect 324412 188828 324464 188834
rect 324412 188770 324464 188776
rect 327552 180794 327580 200124
rect 328196 199306 328224 200124
rect 328184 199300 328236 199306
rect 328184 199242 328236 199248
rect 328460 195152 328512 195158
rect 328460 195094 328512 195100
rect 327092 180766 327580 180794
rect 327092 174894 327120 180766
rect 327080 174888 327132 174894
rect 327080 174830 327132 174836
rect 328472 165102 328500 195094
rect 328840 184686 328868 200124
rect 329438 200002 329466 200124
rect 329392 199974 329466 200002
rect 329392 195158 329420 199974
rect 330484 198076 330536 198082
rect 330484 198018 330536 198024
rect 329380 195152 329432 195158
rect 329380 195094 329432 195100
rect 328828 184680 328880 184686
rect 328828 184622 328880 184628
rect 329196 179240 329248 179246
rect 329196 179182 329248 179188
rect 328460 165096 328512 165102
rect 328460 165038 328512 165044
rect 328460 161016 328512 161022
rect 328460 160958 328512 160964
rect 327264 153128 327316 153134
rect 327264 153070 327316 153076
rect 325056 153060 325108 153066
rect 325056 153002 325108 153008
rect 324320 151700 324372 151706
rect 324320 151642 324372 151648
rect 325068 149954 325096 153002
rect 326620 152516 326672 152522
rect 326620 152458 326672 152464
rect 324730 149926 325096 149954
rect 326632 149940 326660 152458
rect 327276 149940 327304 153070
rect 328472 149954 328500 160958
rect 328472 149926 328578 149954
rect 329208 149940 329236 179182
rect 330496 157214 330524 198018
rect 330772 194274 330800 200124
rect 332060 198150 332088 200124
rect 332048 198144 332100 198150
rect 332048 198086 332100 198092
rect 330760 194268 330812 194274
rect 330760 194210 330812 194216
rect 333348 192710 333376 200124
rect 333946 199866 333974 200124
rect 333946 199838 334112 199866
rect 333980 195152 334032 195158
rect 333980 195094 334032 195100
rect 333336 192704 333388 192710
rect 333336 192646 333388 192652
rect 333992 157350 334020 195094
rect 334084 158302 334112 199838
rect 335280 195158 335308 200124
rect 335268 195152 335320 195158
rect 335268 195094 335320 195100
rect 337856 192914 337884 200124
rect 339098 199866 339126 200124
rect 338960 199838 339126 199866
rect 338120 197396 338172 197402
rect 338120 197338 338172 197344
rect 338132 196450 338160 197338
rect 338120 196444 338172 196450
rect 338120 196386 338172 196392
rect 337844 192908 337896 192914
rect 337844 192850 337896 192856
rect 338960 180794 338988 199838
rect 340432 198626 340460 200124
rect 340420 198620 340472 198626
rect 340420 198562 340472 198568
rect 339500 192636 339552 192642
rect 339500 192578 339552 192584
rect 338132 180766 338988 180794
rect 335636 160812 335688 160818
rect 335636 160754 335688 160760
rect 334072 158296 334124 158302
rect 334072 158238 334124 158244
rect 333980 157344 334032 157350
rect 333980 157286 334032 157292
rect 330484 157208 330536 157214
rect 330484 157150 330536 157156
rect 334992 152856 335044 152862
rect 334992 152798 335044 152804
rect 335004 149940 335032 152798
rect 335648 149940 335676 160754
rect 338132 155650 338160 180766
rect 338120 155644 338172 155650
rect 338120 155586 338172 155592
rect 339512 149940 339540 192578
rect 341076 180794 341104 200124
rect 342364 197033 342392 200124
rect 343008 199442 343036 200124
rect 346228 199918 346256 200124
rect 346216 199912 346268 199918
rect 346216 199854 346268 199860
rect 347516 199594 347544 200124
rect 346412 199566 347544 199594
rect 347596 199572 347648 199578
rect 342996 199436 343048 199442
rect 342996 199378 343048 199384
rect 342350 197024 342406 197033
rect 342350 196959 342406 196968
rect 342720 194268 342772 194274
rect 342720 194210 342772 194216
rect 340892 180766 341104 180794
rect 340892 180266 340920 180766
rect 340880 180260 340932 180266
rect 340880 180202 340932 180208
rect 342076 166388 342128 166394
rect 342076 166330 342128 166336
rect 340144 155712 340196 155718
rect 340144 155654 340196 155660
rect 340156 149940 340184 155654
rect 341800 152448 341852 152454
rect 341800 152390 341852 152396
rect 341812 149954 341840 152390
rect 341474 149926 341840 149954
rect 342088 149940 342116 166330
rect 342732 149940 342760 194210
rect 345020 163600 345072 163606
rect 345020 163542 345072 163548
rect 343364 157276 343416 157282
rect 343364 157218 343416 157224
rect 343376 149940 343404 157218
rect 344008 152516 344060 152522
rect 344008 152458 344060 152464
rect 344020 149940 344048 152458
rect 345032 149954 345060 163542
rect 346412 155718 346440 199566
rect 347596 199514 347648 199520
rect 347504 199504 347556 199510
rect 347504 199446 347556 199452
rect 347516 180794 347544 199446
rect 347608 198694 347636 199514
rect 347700 199345 347728 200359
rect 347778 200288 347834 200297
rect 347778 200223 347780 200232
rect 347832 200223 347834 200232
rect 347780 200194 347832 200200
rect 347780 200116 347832 200122
rect 347780 200058 347832 200064
rect 347686 199336 347742 199345
rect 347686 199271 347742 199280
rect 347792 199209 347820 200058
rect 347778 199200 347834 199209
rect 347778 199135 347834 199144
rect 347596 198688 347648 198694
rect 347596 198630 347648 198636
rect 347056 180766 347544 180794
rect 347056 179178 347084 180766
rect 347044 179172 347096 179178
rect 347044 179114 347096 179120
rect 347884 173466 347912 445703
rect 347976 336569 348004 574874
rect 348068 561649 348096 577458
rect 348148 570784 348200 570790
rect 348148 570726 348200 570732
rect 348054 561640 348110 561649
rect 348054 561575 348110 561584
rect 348054 512000 348110 512009
rect 348054 511935 348110 511944
rect 347962 336560 348018 336569
rect 347962 336495 348018 336504
rect 347962 331120 348018 331129
rect 347962 331055 348018 331064
rect 347872 173460 347924 173466
rect 347872 173402 347924 173408
rect 346584 168088 346636 168094
rect 346584 168030 346636 168036
rect 346400 155712 346452 155718
rect 346400 155654 346452 155660
rect 345032 149926 345322 149954
rect 346596 149940 346624 168030
rect 347976 166394 348004 331055
rect 348068 296449 348096 511935
rect 348160 410961 348188 570726
rect 348240 569560 348292 569566
rect 348240 569502 348292 569508
rect 348252 456521 348280 569502
rect 348332 566568 348384 566574
rect 348332 566510 348384 566516
rect 348344 477601 348372 566510
rect 348422 523016 348478 523025
rect 348422 522951 348478 522960
rect 348330 477592 348386 477601
rect 348330 477527 348386 477536
rect 348238 456512 348294 456521
rect 348238 456447 348294 456456
rect 348146 410952 348202 410961
rect 348146 410887 348202 410896
rect 348238 395924 348294 395933
rect 348238 395859 348294 395868
rect 348146 391164 348202 391173
rect 348146 391099 348202 391108
rect 348054 296440 348110 296449
rect 348054 296375 348110 296384
rect 348054 262848 348110 262857
rect 348054 262783 348110 262792
rect 348068 186046 348096 262783
rect 348160 186794 348188 391099
rect 348252 191622 348280 395859
rect 348330 368724 348386 368733
rect 348330 368659 348386 368668
rect 348240 191616 348292 191622
rect 348240 191558 348292 191564
rect 348148 186788 348200 186794
rect 348148 186730 348200 186736
rect 348056 186040 348108 186046
rect 348056 185982 348108 185988
rect 348344 179314 348372 368659
rect 348436 195702 348464 522951
rect 348528 476270 348556 589630
rect 351184 589620 351236 589626
rect 351184 589562 351236 589568
rect 350816 589348 350868 589354
rect 350816 589290 350868 589296
rect 349620 583024 349672 583030
rect 349620 582966 349672 582972
rect 349252 577584 349304 577590
rect 349252 577526 349304 577532
rect 349160 572008 349212 572014
rect 349160 571950 349212 571956
rect 348608 568132 348660 568138
rect 348608 568074 348660 568080
rect 348620 511601 348648 568074
rect 349172 541521 349200 571950
rect 349158 541512 349214 541521
rect 349158 541447 349214 541456
rect 349066 540968 349122 540977
rect 349066 540903 349122 540912
rect 349080 523002 349108 540903
rect 349080 522974 349200 523002
rect 349172 513346 349200 522974
rect 349080 513318 349200 513346
rect 348606 511592 348662 511601
rect 348606 511527 348662 511536
rect 349080 485058 349108 513318
rect 349080 485030 349200 485058
rect 349172 477510 349200 485030
rect 348896 477482 349200 477510
rect 348516 476264 348568 476270
rect 348516 476206 348568 476212
rect 348698 475008 348754 475017
rect 348698 474943 348754 474952
rect 348516 281988 348568 281994
rect 348516 281930 348568 281936
rect 348528 199374 348556 281930
rect 348608 213920 348660 213926
rect 348608 213862 348660 213868
rect 348516 199368 348568 199374
rect 348516 199310 348568 199316
rect 348424 195696 348476 195702
rect 348424 195638 348476 195644
rect 348332 179308 348384 179314
rect 348332 179250 348384 179256
rect 347964 166388 348016 166394
rect 347964 166330 348016 166336
rect 348620 155854 348648 213862
rect 348712 162382 348740 474943
rect 348896 447166 348924 477482
rect 349066 469296 349122 469305
rect 349066 469231 349122 469240
rect 348976 455388 349028 455394
rect 348976 455330 349028 455336
rect 348884 447160 348936 447166
rect 348884 447102 348936 447108
rect 348884 436348 348936 436354
rect 348884 436290 348936 436296
rect 348896 392018 348924 436290
rect 348988 407794 349016 455330
rect 348976 407788 349028 407794
rect 348976 407730 349028 407736
rect 348884 392012 348936 392018
rect 348884 391954 348936 391960
rect 349080 385014 349108 469231
rect 349160 447160 349212 447166
rect 349160 447102 349212 447108
rect 349172 436354 349200 447102
rect 349160 436348 349212 436354
rect 349160 436290 349212 436296
rect 349068 385008 349120 385014
rect 349068 384950 349120 384956
rect 349068 368484 349120 368490
rect 349068 368426 349120 368432
rect 349080 313290 349108 368426
rect 349264 347041 349292 577526
rect 349436 574864 349488 574870
rect 349436 574806 349488 574812
rect 349344 571192 349396 571198
rect 349344 571134 349396 571140
rect 349356 396681 349384 571134
rect 349448 493921 349476 574806
rect 349528 566704 349580 566710
rect 349528 566646 349580 566652
rect 349434 493912 349490 493921
rect 349434 493847 349490 493856
rect 349434 465216 349490 465225
rect 349434 465151 349490 465160
rect 349342 396672 349398 396681
rect 349342 396607 349398 396616
rect 349344 392012 349396 392018
rect 349344 391954 349396 391960
rect 349356 368490 349384 391954
rect 349344 368484 349396 368490
rect 349344 368426 349396 368432
rect 349250 347032 349306 347041
rect 349250 346967 349306 346976
rect 349080 313262 349200 313290
rect 349172 306374 349200 313262
rect 349172 306346 349384 306374
rect 349158 302288 349214 302297
rect 349158 302223 349214 302232
rect 349068 279064 349120 279070
rect 349068 279006 349120 279012
rect 349080 262206 349108 279006
rect 349068 262200 349120 262206
rect 349068 262142 349120 262148
rect 349068 239760 349120 239766
rect 349068 239702 349120 239708
rect 349080 233238 349108 239702
rect 349068 233232 349120 233238
rect 349068 233174 349120 233180
rect 349172 190126 349200 302223
rect 349252 295792 349304 295798
rect 349252 295734 349304 295740
rect 349264 288561 349292 295734
rect 349250 288552 349306 288561
rect 349250 288487 349306 288496
rect 349250 280528 349306 280537
rect 349250 280463 349306 280472
rect 349160 190120 349212 190126
rect 349160 190062 349212 190068
rect 349264 177614 349292 280463
rect 349356 213926 349384 306346
rect 349448 295497 349476 465151
rect 349540 409601 349568 566646
rect 349632 455841 349660 582966
rect 350724 581664 350776 581670
rect 350724 581606 350776 581612
rect 350356 580372 350408 580378
rect 350356 580314 350408 580320
rect 349896 580304 349948 580310
rect 349896 580246 349948 580252
rect 349804 573436 349856 573442
rect 349804 573378 349856 573384
rect 349712 570988 349764 570994
rect 349712 570930 349764 570936
rect 349618 455832 349674 455841
rect 349618 455767 349674 455776
rect 349724 451081 349752 570930
rect 349816 500041 349844 573378
rect 349908 521801 349936 580246
rect 349988 559496 350040 559502
rect 349988 559438 350040 559444
rect 350000 558958 350028 559438
rect 349988 558952 350040 558958
rect 349988 558894 350040 558900
rect 350172 549228 350224 549234
rect 350172 549170 350224 549176
rect 350184 549001 350212 549170
rect 350170 548992 350226 549001
rect 350170 548927 350226 548936
rect 350262 547088 350318 547097
rect 350262 547023 350318 547032
rect 350276 546514 350304 547023
rect 350264 546508 350316 546514
rect 350264 546450 350316 546456
rect 350262 533488 350318 533497
rect 350262 533423 350318 533432
rect 350276 532846 350304 533423
rect 350264 532840 350316 532846
rect 350264 532782 350316 532788
rect 350264 524408 350316 524414
rect 350264 524350 350316 524356
rect 350276 523161 350304 524350
rect 350262 523152 350318 523161
rect 350262 523087 350318 523096
rect 349894 521792 349950 521801
rect 349894 521727 349950 521736
rect 350170 520432 350226 520441
rect 350170 520367 350226 520376
rect 350184 520334 350212 520367
rect 350172 520328 350224 520334
rect 350172 520270 350224 520276
rect 350262 516624 350318 516633
rect 350262 516559 350318 516568
rect 350276 516254 350304 516559
rect 350264 516248 350316 516254
rect 350264 516190 350316 516196
rect 350262 513496 350318 513505
rect 350262 513431 350264 513440
rect 350316 513431 350318 513440
rect 350264 513402 350316 513408
rect 350264 506456 350316 506462
rect 350264 506398 350316 506404
rect 350276 505481 350304 506398
rect 350262 505472 350318 505481
rect 350262 505407 350318 505416
rect 349802 500032 349858 500041
rect 349802 499967 349858 499976
rect 350262 492008 350318 492017
rect 350262 491943 350318 491952
rect 350276 491434 350304 491943
rect 350264 491428 350316 491434
rect 350264 491370 350316 491376
rect 350262 490240 350318 490249
rect 350262 490175 350318 490184
rect 350276 489938 350304 490175
rect 350264 489932 350316 489938
rect 350264 489874 350316 489880
rect 350172 489864 350224 489870
rect 350170 489832 350172 489841
rect 350224 489832 350226 489841
rect 350170 489767 350226 489776
rect 350264 488504 350316 488510
rect 350264 488446 350316 488452
rect 350276 487801 350304 488446
rect 350262 487792 350318 487801
rect 350262 487727 350318 487736
rect 349986 485208 350042 485217
rect 349986 485143 350042 485152
rect 350000 484430 350028 485143
rect 349988 484424 350040 484430
rect 349988 484366 350040 484372
rect 350262 483440 350318 483449
rect 350262 483375 350318 483384
rect 350276 483070 350304 483375
rect 350264 483064 350316 483070
rect 350264 483006 350316 483012
rect 350262 480720 350318 480729
rect 350262 480655 350318 480664
rect 350276 480350 350304 480655
rect 350264 480344 350316 480350
rect 350264 480286 350316 480292
rect 350170 476640 350226 476649
rect 350170 476575 350226 476584
rect 349804 476264 349856 476270
rect 349804 476206 349856 476212
rect 349710 451072 349766 451081
rect 349710 451007 349766 451016
rect 349816 433401 349844 476206
rect 350184 476202 350212 476575
rect 350262 476232 350318 476241
rect 350172 476196 350224 476202
rect 350262 476167 350318 476176
rect 350172 476138 350224 476144
rect 350276 476134 350304 476167
rect 350264 476128 350316 476134
rect 350264 476070 350316 476076
rect 350262 473512 350318 473521
rect 350262 473447 350318 473456
rect 350276 473414 350304 473447
rect 350264 473408 350316 473414
rect 350264 473350 350316 473356
rect 350264 466404 350316 466410
rect 350264 466346 350316 466352
rect 350276 466041 350304 466346
rect 350262 466032 350318 466041
rect 350262 465967 350318 465976
rect 350262 462904 350318 462913
rect 350262 462839 350318 462848
rect 350276 462466 350304 462839
rect 350264 462460 350316 462466
rect 350264 462402 350316 462408
rect 350262 461544 350318 461553
rect 350262 461479 350318 461488
rect 350276 461038 350304 461479
rect 350264 461032 350316 461038
rect 350264 460974 350316 460980
rect 350262 457328 350318 457337
rect 350262 457263 350318 457272
rect 350276 456822 350304 457263
rect 350264 456816 350316 456822
rect 350264 456758 350316 456764
rect 350262 446448 350318 446457
rect 350262 446383 350318 446392
rect 350276 445806 350304 446383
rect 350264 445800 350316 445806
rect 350264 445742 350316 445748
rect 350262 437880 350318 437889
rect 350262 437815 350318 437824
rect 350276 437510 350304 437815
rect 350264 437504 350316 437510
rect 350264 437446 350316 437452
rect 349802 433392 349858 433401
rect 349802 433327 349858 433336
rect 350262 430944 350318 430953
rect 350262 430879 350318 430888
rect 350276 430642 350304 430879
rect 350264 430636 350316 430642
rect 350264 430578 350316 430584
rect 349986 421288 350042 421297
rect 349986 421223 350042 421232
rect 350000 421054 350028 421223
rect 349988 421048 350040 421054
rect 349988 420990 350040 420996
rect 350262 414488 350318 414497
rect 350262 414423 350318 414432
rect 350276 414050 350304 414423
rect 350264 414044 350316 414050
rect 350264 413986 350316 413992
rect 349526 409592 349582 409601
rect 349526 409527 349582 409536
rect 350172 407788 350224 407794
rect 350172 407730 350224 407736
rect 349804 396840 349856 396846
rect 349804 396782 349856 396788
rect 349618 391368 349674 391377
rect 349618 391303 349674 391312
rect 349632 390590 349660 391303
rect 349620 390584 349672 390590
rect 349620 390526 349672 390532
rect 349434 295488 349490 295497
rect 349434 295423 349490 295432
rect 349434 284336 349490 284345
rect 349434 284271 349490 284280
rect 349344 213920 349396 213926
rect 349344 213862 349396 213868
rect 349342 202328 349398 202337
rect 349342 202263 349398 202272
rect 349356 199510 349384 202263
rect 349344 199504 349396 199510
rect 349344 199446 349396 199452
rect 349448 196586 349476 284271
rect 349528 248192 349580 248198
rect 349528 248134 349580 248140
rect 349540 247761 349568 248134
rect 349526 247752 349582 247761
rect 349526 247687 349582 247696
rect 349618 245712 349674 245721
rect 349618 245647 349674 245656
rect 349526 225040 349582 225049
rect 349526 224975 349582 224984
rect 349436 196580 349488 196586
rect 349436 196522 349488 196528
rect 349252 177608 349304 177614
rect 349252 177550 349304 177556
rect 348700 162376 348752 162382
rect 348700 162318 348752 162324
rect 349540 158234 349568 224975
rect 349632 184482 349660 245647
rect 349712 233232 349764 233238
rect 349712 233174 349764 233180
rect 349620 184476 349672 184482
rect 349620 184418 349672 184424
rect 349724 172242 349752 233174
rect 349816 195566 349844 396782
rect 349896 396024 349948 396030
rect 349896 395966 349948 395972
rect 349908 257961 349936 395966
rect 350078 381304 350134 381313
rect 350078 381239 350134 381248
rect 350092 381002 350120 381239
rect 350080 380996 350132 381002
rect 350080 380938 350132 380944
rect 349986 379536 350042 379545
rect 349986 379471 350042 379480
rect 350000 268841 350028 379471
rect 350080 378140 350132 378146
rect 350080 378082 350132 378088
rect 350092 376961 350120 378082
rect 350078 376952 350134 376961
rect 350078 376887 350134 376896
rect 350078 375864 350134 375873
rect 350078 375799 350134 375808
rect 350092 375426 350120 375799
rect 350080 375420 350132 375426
rect 350080 375362 350132 375368
rect 350080 371204 350132 371210
rect 350080 371146 350132 371152
rect 350092 370161 350120 371146
rect 350078 370152 350134 370161
rect 350078 370087 350134 370096
rect 350078 363352 350134 363361
rect 350078 363287 350134 363296
rect 350092 362982 350120 363287
rect 350080 362976 350132 362982
rect 350080 362918 350132 362924
rect 350078 349888 350134 349897
rect 350078 349823 350134 349832
rect 350092 349246 350120 349823
rect 350080 349240 350132 349246
rect 350080 349182 350132 349188
rect 350078 344448 350134 344457
rect 350078 344383 350134 344392
rect 350092 343670 350120 344383
rect 350080 343664 350132 343670
rect 350080 343606 350132 343612
rect 350078 311128 350134 311137
rect 350078 311063 350134 311072
rect 349986 268832 350042 268841
rect 349986 268767 350042 268776
rect 349988 262200 350040 262206
rect 349988 262142 350040 262148
rect 349894 257952 349950 257961
rect 349894 257887 349950 257896
rect 349896 255468 349948 255474
rect 349896 255410 349948 255416
rect 349908 239766 349936 255410
rect 350000 244934 350028 262142
rect 349988 244928 350040 244934
rect 349988 244870 350040 244876
rect 349986 242992 350042 243001
rect 349986 242927 350042 242936
rect 349896 239760 349948 239766
rect 349896 239702 349948 239708
rect 350000 233986 350028 242927
rect 349988 233980 350040 233986
rect 349988 233922 350040 233928
rect 349986 220008 350042 220017
rect 349986 219943 350042 219952
rect 349896 200796 349948 200802
rect 349896 200738 349948 200744
rect 349804 195560 349856 195566
rect 349804 195502 349856 195508
rect 349712 172236 349764 172242
rect 349712 172178 349764 172184
rect 349528 158228 349580 158234
rect 349528 158170 349580 158176
rect 348608 155848 348660 155854
rect 348608 155790 348660 155796
rect 347872 153196 347924 153202
rect 347872 153138 347924 153144
rect 347884 149940 347912 153138
rect 349908 151814 349936 200738
rect 350000 195537 350028 219943
rect 350092 203590 350120 311063
rect 350184 310486 350212 407730
rect 350262 404968 350318 404977
rect 350262 404903 350318 404912
rect 350276 404462 350304 404903
rect 350264 404456 350316 404462
rect 350264 404398 350316 404404
rect 350262 394768 350318 394777
rect 350262 394703 350264 394712
rect 350316 394703 350318 394712
rect 350264 394674 350316 394680
rect 350262 390008 350318 390017
rect 350262 389943 350318 389952
rect 350276 389230 350304 389943
rect 350264 389224 350316 389230
rect 350264 389166 350316 389172
rect 350264 387796 350316 387802
rect 350264 387738 350316 387744
rect 350276 387161 350304 387738
rect 350262 387152 350318 387161
rect 350262 387087 350318 387096
rect 350262 382392 350318 382401
rect 350262 382327 350318 382336
rect 350276 382294 350304 382327
rect 350264 382288 350316 382294
rect 350264 382230 350316 382236
rect 350262 381032 350318 381041
rect 350262 380967 350318 380976
rect 350276 380934 350304 380967
rect 350264 380928 350316 380934
rect 350264 380870 350316 380876
rect 350262 377224 350318 377233
rect 350262 377159 350318 377168
rect 350276 376786 350304 377159
rect 350264 376780 350316 376786
rect 350264 376722 350316 376728
rect 350264 375352 350316 375358
rect 350264 375294 350316 375300
rect 350276 374921 350304 375294
rect 350262 374912 350318 374921
rect 350262 374847 350318 374856
rect 350262 372872 350318 372881
rect 350262 372807 350318 372816
rect 350276 372638 350304 372807
rect 350264 372632 350316 372638
rect 350264 372574 350316 372580
rect 350262 371376 350318 371385
rect 350262 371311 350318 371320
rect 350276 371278 350304 371311
rect 350264 371272 350316 371278
rect 350264 371214 350316 371220
rect 350262 358864 350318 358873
rect 350262 358799 350264 358808
rect 350316 358799 350318 358808
rect 350264 358770 350316 358776
rect 350262 358320 350318 358329
rect 350262 358255 350318 358264
rect 350276 358018 350304 358255
rect 350264 358012 350316 358018
rect 350264 357954 350316 357960
rect 350262 356688 350318 356697
rect 350262 356623 350318 356632
rect 350276 356182 350304 356623
rect 350264 356176 350316 356182
rect 350264 356118 350316 356124
rect 350264 356040 350316 356046
rect 350264 355982 350316 355988
rect 350276 355881 350304 355982
rect 350262 355872 350318 355881
rect 350262 355807 350318 355816
rect 350262 354784 350318 354793
rect 350262 354719 350264 354728
rect 350316 354719 350318 354728
rect 350264 354690 350316 354696
rect 350262 350704 350318 350713
rect 350262 350639 350318 350648
rect 350276 350606 350304 350639
rect 350264 350600 350316 350606
rect 350264 350542 350316 350548
rect 350262 349480 350318 349489
rect 350262 349415 350318 349424
rect 350276 349178 350304 349415
rect 350264 349172 350316 349178
rect 350264 349114 350316 349120
rect 350262 345808 350318 345817
rect 350262 345743 350318 345752
rect 350276 345098 350304 345743
rect 350264 345092 350316 345098
rect 350264 345034 350316 345040
rect 350262 344040 350318 344049
rect 350262 343975 350318 343984
rect 350276 343738 350304 343975
rect 350264 343732 350316 343738
rect 350264 343674 350316 343680
rect 350368 335354 350396 580314
rect 350632 579012 350684 579018
rect 350632 578954 350684 578960
rect 350448 554736 350500 554742
rect 350448 554678 350500 554684
rect 350460 554441 350488 554678
rect 350446 554432 350502 554441
rect 350446 554367 350502 554376
rect 350446 551440 350502 551449
rect 350446 551375 350502 551384
rect 350460 551138 350488 551375
rect 350448 551132 350500 551138
rect 350448 551074 350500 551080
rect 350446 546680 350502 546689
rect 350446 546615 350448 546624
rect 350500 546615 350502 546624
rect 350448 546586 350500 546592
rect 350446 543008 350502 543017
rect 350446 542943 350502 542952
rect 350460 542434 350488 542943
rect 350448 542428 350500 542434
rect 350448 542370 350500 542376
rect 350446 538384 350502 538393
rect 350446 538319 350502 538328
rect 350460 538286 350488 538319
rect 350448 538280 350500 538286
rect 350448 538222 350500 538228
rect 350446 537160 350502 537169
rect 350446 537095 350502 537104
rect 350460 536858 350488 537095
rect 350448 536852 350500 536858
rect 350448 536794 350500 536800
rect 350446 534712 350502 534721
rect 350446 534647 350502 534656
rect 350460 534138 350488 534647
rect 350448 534132 350500 534138
rect 350448 534074 350500 534080
rect 350446 533080 350502 533089
rect 350446 533015 350502 533024
rect 350460 532778 350488 533015
rect 350448 532772 350500 532778
rect 350448 532714 350500 532720
rect 350446 532128 350502 532137
rect 350446 532063 350502 532072
rect 350460 531350 350488 532063
rect 350448 531344 350500 531350
rect 350448 531286 350500 531292
rect 350446 530768 350502 530777
rect 350446 530703 350502 530712
rect 350460 529990 350488 530703
rect 350448 529984 350500 529990
rect 350448 529926 350500 529932
rect 350446 527232 350502 527241
rect 350446 527167 350448 527176
rect 350500 527167 350502 527176
rect 350448 527138 350500 527144
rect 350446 526280 350502 526289
rect 350446 526215 350502 526224
rect 350460 525978 350488 526215
rect 350448 525972 350500 525978
rect 350448 525914 350500 525920
rect 350446 523288 350502 523297
rect 350446 523223 350502 523232
rect 350460 523054 350488 523223
rect 350448 523048 350500 523054
rect 350448 522990 350500 522996
rect 350446 517712 350502 517721
rect 350446 517647 350502 517656
rect 350460 517614 350488 517647
rect 350448 517608 350500 517614
rect 350448 517550 350500 517556
rect 350446 516216 350502 516225
rect 350446 516151 350448 516160
rect 350500 516151 350502 516160
rect 350448 516122 350500 516128
rect 350446 513768 350502 513777
rect 350446 513703 350502 513712
rect 350460 513398 350488 513703
rect 350448 513392 350500 513398
rect 350448 513334 350500 513340
rect 350448 509244 350500 509250
rect 350448 509186 350500 509192
rect 350460 508881 350488 509186
rect 350446 508872 350502 508881
rect 350446 508807 350502 508816
rect 350446 506968 350502 506977
rect 350446 506903 350502 506912
rect 350460 506530 350488 506903
rect 350448 506524 350500 506530
rect 350448 506466 350500 506472
rect 350446 505608 350502 505617
rect 350446 505543 350502 505552
rect 350460 505170 350488 505543
rect 350448 505164 350500 505170
rect 350448 505106 350500 505112
rect 350446 503840 350502 503849
rect 350446 503775 350502 503784
rect 350460 503742 350488 503775
rect 350448 503736 350500 503742
rect 350448 503678 350500 503684
rect 350446 500168 350502 500177
rect 350446 500103 350502 500112
rect 350460 499594 350488 500103
rect 350448 499588 350500 499594
rect 350448 499530 350500 499536
rect 350446 498264 350502 498273
rect 350446 498199 350448 498208
rect 350500 498199 350502 498208
rect 350448 498170 350500 498176
rect 350446 495544 350502 495553
rect 350446 495479 350448 495488
rect 350500 495479 350502 495488
rect 350448 495450 350500 495456
rect 350448 493468 350500 493474
rect 350448 493410 350500 493416
rect 350460 491586 350488 493410
rect 350460 491558 350580 491586
rect 350446 491464 350502 491473
rect 350446 491399 350502 491408
rect 350460 491366 350488 491399
rect 350448 491360 350500 491366
rect 350448 491302 350500 491308
rect 350446 490648 350502 490657
rect 350446 490583 350502 490592
rect 350460 490006 350488 490583
rect 350448 490000 350500 490006
rect 350448 489942 350500 489948
rect 350552 489914 350580 491558
rect 350460 489886 350580 489914
rect 350460 481794 350488 489886
rect 350460 481766 350580 481794
rect 350448 481704 350500 481710
rect 350446 481672 350448 481681
rect 350500 481672 350502 481681
rect 350446 481607 350502 481616
rect 350552 481522 350580 481766
rect 350460 481494 350580 481522
rect 350460 480434 350488 481494
rect 350460 480406 350580 480434
rect 350446 480312 350502 480321
rect 350446 480247 350448 480256
rect 350500 480247 350502 480256
rect 350448 480218 350500 480224
rect 350552 480162 350580 480406
rect 350460 480134 350580 480162
rect 350460 475402 350488 480134
rect 350460 475374 350580 475402
rect 350446 472288 350502 472297
rect 350446 472223 350502 472232
rect 350460 472054 350488 472223
rect 350448 472048 350500 472054
rect 350448 471990 350500 471996
rect 350446 466576 350502 466585
rect 350446 466511 350502 466520
rect 350460 466478 350488 466511
rect 350448 466472 350500 466478
rect 350448 466414 350500 466420
rect 350446 462632 350502 462641
rect 350446 462567 350502 462576
rect 350460 462534 350488 462567
rect 350448 462528 350500 462534
rect 350448 462470 350500 462476
rect 350446 461136 350502 461145
rect 350446 461071 350448 461080
rect 350500 461071 350502 461080
rect 350448 461042 350500 461048
rect 350446 459640 350502 459649
rect 350446 459575 350448 459584
rect 350500 459575 350502 459584
rect 350448 459546 350500 459552
rect 350446 456920 350502 456929
rect 350446 456855 350448 456864
rect 350500 456855 350502 456864
rect 350448 456826 350500 456832
rect 350552 455394 350580 475374
rect 350540 455388 350592 455394
rect 350540 455330 350592 455336
rect 350446 454200 350502 454209
rect 350446 454135 350502 454144
rect 350460 454102 350488 454135
rect 350448 454096 350500 454102
rect 350448 454038 350500 454044
rect 350446 451888 350502 451897
rect 350446 451823 350502 451832
rect 350460 451314 350488 451823
rect 350448 451308 350500 451314
rect 350448 451250 350500 451256
rect 350446 449984 350502 449993
rect 350446 449919 350448 449928
rect 350500 449919 350502 449928
rect 350448 449890 350500 449896
rect 350446 447808 350502 447817
rect 350446 447743 350502 447752
rect 350460 447166 350488 447743
rect 350448 447160 350500 447166
rect 350448 447102 350500 447108
rect 350448 445732 350500 445738
rect 350448 445674 350500 445680
rect 350460 445641 350488 445674
rect 350446 445632 350502 445641
rect 350446 445567 350502 445576
rect 350446 440600 350502 440609
rect 350446 440535 350502 440544
rect 350460 440298 350488 440535
rect 350448 440292 350500 440298
rect 350448 440234 350500 440240
rect 350448 437436 350500 437442
rect 350448 437378 350500 437384
rect 350460 436801 350488 437378
rect 350446 436792 350502 436801
rect 350446 436727 350502 436736
rect 350448 434852 350500 434858
rect 350448 434794 350500 434800
rect 350460 434761 350488 434794
rect 350446 434752 350502 434761
rect 350446 434687 350502 434696
rect 350448 430704 350500 430710
rect 350446 430672 350448 430681
rect 350500 430672 350502 430681
rect 350446 430607 350502 430616
rect 350446 427952 350502 427961
rect 350446 427887 350502 427896
rect 350460 427854 350488 427887
rect 350448 427848 350500 427854
rect 350448 427790 350500 427796
rect 350446 426592 350502 426601
rect 350446 426527 350502 426536
rect 350460 426494 350488 426527
rect 350448 426488 350500 426494
rect 350448 426430 350500 426436
rect 350446 425368 350502 425377
rect 350446 425303 350502 425312
rect 350460 425134 350488 425303
rect 350448 425128 350500 425134
rect 350448 425070 350500 425076
rect 350446 422376 350502 422385
rect 350446 422311 350448 422320
rect 350500 422311 350502 422320
rect 350448 422282 350500 422288
rect 350446 421016 350502 421025
rect 350446 420951 350448 420960
rect 350500 420951 350502 420960
rect 350448 420922 350500 420928
rect 350446 419656 350502 419665
rect 350446 419591 350448 419600
rect 350500 419591 350502 419600
rect 350448 419562 350500 419568
rect 350446 418432 350502 418441
rect 350446 418367 350502 418376
rect 350460 418266 350488 418367
rect 350448 418260 350500 418266
rect 350448 418202 350500 418208
rect 350446 416936 350502 416945
rect 350446 416871 350502 416880
rect 350460 416838 350488 416871
rect 350448 416832 350500 416838
rect 350448 416774 350500 416780
rect 350446 414216 350502 414225
rect 350446 414151 350502 414160
rect 350460 414118 350488 414151
rect 350448 414112 350500 414118
rect 350448 414054 350500 414060
rect 350446 411360 350502 411369
rect 350446 411295 350448 411304
rect 350500 411295 350502 411304
rect 350448 411266 350500 411272
rect 350446 404424 350502 404433
rect 350446 404359 350448 404368
rect 350500 404359 350502 404368
rect 350448 404330 350500 404336
rect 350446 400344 350502 400353
rect 350446 400279 350502 400288
rect 350460 400246 350488 400279
rect 350448 400240 350500 400246
rect 350448 400182 350500 400188
rect 350446 399528 350502 399537
rect 350446 399463 350502 399472
rect 350460 398886 350488 399463
rect 350448 398880 350500 398886
rect 350448 398822 350500 398828
rect 350446 397624 350502 397633
rect 350446 397559 350502 397568
rect 350460 397526 350488 397559
rect 350448 397520 350500 397526
rect 350448 397462 350500 397468
rect 350446 396808 350502 396817
rect 350446 396743 350502 396752
rect 350460 396098 350488 396743
rect 350448 396092 350500 396098
rect 350448 396034 350500 396040
rect 350448 394664 350500 394670
rect 350446 394632 350448 394641
rect 350500 394632 350502 394641
rect 350446 394567 350502 394576
rect 350446 392320 350502 392329
rect 350446 392255 350502 392264
rect 350460 392018 350488 392255
rect 350448 392012 350500 392018
rect 350448 391954 350500 391960
rect 350448 390516 350500 390522
rect 350448 390458 350500 390464
rect 350460 389881 350488 390458
rect 350446 389872 350502 389881
rect 350446 389807 350502 389816
rect 350448 387864 350500 387870
rect 350446 387832 350448 387841
rect 350500 387832 350502 387841
rect 350446 387767 350502 387776
rect 350448 386368 350500 386374
rect 350448 386310 350500 386316
rect 350460 385121 350488 386310
rect 350446 385112 350502 385121
rect 350446 385047 350502 385056
rect 350448 384328 350500 384334
rect 350448 384270 350500 384276
rect 350276 335326 350396 335354
rect 350276 324601 350304 335326
rect 350354 334112 350410 334121
rect 350354 334047 350356 334056
rect 350408 334047 350410 334056
rect 350356 334018 350408 334024
rect 350354 332752 350410 332761
rect 350354 332687 350410 332696
rect 350368 332654 350396 332687
rect 350356 332648 350408 332654
rect 350356 332590 350408 332596
rect 350354 329896 350410 329905
rect 350354 329831 350356 329840
rect 350408 329831 350410 329840
rect 350356 329802 350408 329808
rect 350354 328944 350410 328953
rect 350354 328879 350410 328888
rect 350368 328506 350396 328879
rect 350356 328500 350408 328506
rect 350356 328442 350408 328448
rect 350354 325816 350410 325825
rect 350354 325751 350410 325760
rect 350368 325718 350396 325751
rect 350356 325712 350408 325718
rect 350356 325654 350408 325660
rect 350262 324592 350318 324601
rect 350262 324527 350318 324536
rect 350354 321736 350410 321745
rect 350354 321671 350410 321680
rect 350368 321638 350396 321671
rect 350356 321632 350408 321638
rect 350356 321574 350408 321580
rect 350354 320648 350410 320657
rect 350354 320583 350410 320592
rect 350368 320210 350396 320583
rect 350356 320204 350408 320210
rect 350356 320146 350408 320152
rect 350264 320136 350316 320142
rect 350264 320078 350316 320084
rect 350276 319161 350304 320078
rect 350354 319288 350410 319297
rect 350354 319223 350410 319232
rect 350262 319152 350318 319161
rect 350262 319087 350318 319096
rect 350368 318850 350396 319223
rect 350356 318844 350408 318850
rect 350356 318786 350408 318792
rect 350354 317792 350410 317801
rect 350354 317727 350410 317736
rect 350368 317490 350396 317727
rect 350356 317484 350408 317490
rect 350356 317426 350408 317432
rect 350356 315988 350408 315994
rect 350356 315930 350408 315936
rect 350262 315208 350318 315217
rect 350262 315143 350318 315152
rect 350172 310480 350224 310486
rect 350172 310422 350224 310428
rect 350172 302320 350224 302326
rect 350172 302262 350224 302268
rect 350184 281994 350212 302262
rect 350172 281988 350224 281994
rect 350172 281930 350224 281936
rect 350276 239426 350304 315143
rect 350368 315081 350396 315930
rect 350354 315072 350410 315081
rect 350354 315007 350410 315016
rect 350354 312352 350410 312361
rect 350354 312287 350410 312296
rect 350368 311914 350396 312287
rect 350356 311908 350408 311914
rect 350356 311850 350408 311856
rect 350354 308408 350410 308417
rect 350354 308343 350410 308352
rect 350368 307834 350396 308343
rect 350356 307828 350408 307834
rect 350356 307770 350408 307776
rect 350460 306374 350488 384270
rect 350540 310480 350592 310486
rect 350540 310422 350592 310428
rect 350368 306346 350488 306374
rect 350368 294098 350396 306346
rect 350446 304328 350502 304337
rect 350446 304263 350502 304272
rect 350460 303754 350488 304263
rect 350448 303748 350500 303754
rect 350448 303690 350500 303696
rect 350446 302968 350502 302977
rect 350446 302903 350502 302912
rect 350460 302258 350488 302903
rect 350448 302252 350500 302258
rect 350448 302194 350500 302200
rect 350446 301064 350502 301073
rect 350446 300999 350502 301008
rect 350460 300966 350488 300999
rect 350448 300960 350500 300966
rect 350448 300902 350500 300908
rect 350446 300248 350502 300257
rect 350446 300183 350502 300192
rect 350460 299606 350488 300183
rect 350448 299600 350500 299606
rect 350448 299542 350500 299548
rect 350446 298888 350502 298897
rect 350446 298823 350502 298832
rect 350460 298178 350488 298823
rect 350448 298172 350500 298178
rect 350448 298114 350500 298120
rect 350446 296712 350502 296721
rect 350446 296647 350448 296656
rect 350500 296647 350502 296656
rect 350448 296618 350500 296624
rect 350448 295384 350500 295390
rect 350446 295352 350448 295361
rect 350500 295352 350502 295361
rect 350446 295287 350502 295296
rect 350356 294092 350408 294098
rect 350356 294034 350408 294040
rect 350448 294024 350500 294030
rect 350446 293992 350448 294001
rect 350500 293992 350502 294001
rect 350446 293927 350502 293936
rect 350446 288824 350502 288833
rect 350446 288759 350502 288768
rect 350460 288454 350488 288759
rect 350448 288448 350500 288454
rect 350448 288390 350500 288396
rect 350446 287192 350502 287201
rect 350446 287127 350448 287136
rect 350500 287127 350502 287136
rect 350448 287098 350500 287104
rect 350446 285832 350502 285841
rect 350446 285767 350502 285776
rect 350460 285734 350488 285767
rect 350448 285728 350500 285734
rect 350448 285670 350500 285676
rect 350356 285660 350408 285666
rect 350356 285602 350408 285608
rect 350368 285161 350396 285602
rect 350354 285152 350410 285161
rect 350354 285087 350410 285096
rect 350446 277536 350502 277545
rect 350446 277471 350502 277480
rect 350460 277438 350488 277471
rect 350448 277432 350500 277438
rect 350448 277374 350500 277380
rect 350448 276004 350500 276010
rect 350448 275946 350500 275952
rect 350460 275641 350488 275946
rect 350446 275632 350502 275641
rect 350446 275567 350502 275576
rect 350354 273864 350410 273873
rect 350354 273799 350410 273808
rect 350368 273290 350396 273799
rect 350446 273456 350502 273465
rect 350446 273391 350502 273400
rect 350460 273358 350488 273391
rect 350448 273352 350500 273358
rect 350448 273294 350500 273300
rect 350356 273284 350408 273290
rect 350356 273226 350408 273232
rect 350448 270496 350500 270502
rect 350448 270438 350500 270444
rect 350460 270201 350488 270438
rect 350446 270192 350502 270201
rect 350446 270127 350502 270136
rect 350448 269068 350500 269074
rect 350448 269010 350500 269016
rect 350460 268161 350488 269010
rect 350446 268152 350502 268161
rect 350446 268087 350502 268096
rect 350446 266792 350502 266801
rect 350446 266727 350502 266736
rect 350460 266422 350488 266727
rect 350448 266416 350500 266422
rect 350448 266358 350500 266364
rect 350446 263936 350502 263945
rect 350446 263871 350502 263880
rect 350460 263702 350488 263871
rect 350448 263696 350500 263702
rect 350448 263638 350500 263644
rect 350448 262200 350500 262206
rect 350448 262142 350500 262148
rect 350460 261361 350488 262142
rect 350446 261352 350502 261361
rect 350446 261287 350502 261296
rect 350446 258768 350502 258777
rect 350446 258703 350502 258712
rect 350460 258126 350488 258703
rect 350448 258120 350500 258126
rect 350448 258062 350500 258068
rect 350354 256048 350410 256057
rect 350354 255983 350410 255992
rect 350368 255406 350396 255983
rect 350552 255474 350580 310422
rect 350644 262721 350672 578954
rect 350736 279721 350764 581606
rect 350828 295798 350856 589290
rect 351092 585812 351144 585818
rect 351092 585754 351144 585760
rect 350908 571260 350960 571266
rect 350908 571202 350960 571208
rect 350920 302326 350948 571202
rect 351000 568064 351052 568070
rect 351000 568006 351052 568012
rect 351012 342281 351040 568006
rect 351104 365401 351132 585754
rect 351196 396030 351224 589562
rect 351460 585880 351512 585886
rect 351460 585822 351512 585828
rect 351366 560552 351422 560561
rect 351366 560487 351422 560496
rect 351276 560244 351328 560250
rect 351276 560186 351328 560192
rect 351288 493474 351316 560186
rect 351380 552022 351408 560487
rect 351368 552016 351420 552022
rect 351368 551958 351420 551964
rect 351276 493468 351328 493474
rect 351276 493410 351328 493416
rect 351184 396024 351236 396030
rect 351184 395966 351236 395972
rect 351276 390584 351328 390590
rect 351276 390526 351328 390532
rect 351182 379808 351238 379817
rect 351182 379743 351238 379752
rect 351090 365392 351146 365401
rect 351090 365327 351146 365336
rect 351090 364576 351146 364585
rect 351090 364511 351146 364520
rect 350998 342272 351054 342281
rect 350998 342207 351054 342216
rect 350998 338192 351054 338201
rect 350998 338127 351054 338136
rect 350908 302320 350960 302326
rect 350908 302262 350960 302268
rect 350816 295792 350868 295798
rect 350816 295734 350868 295740
rect 350816 294092 350868 294098
rect 350816 294034 350868 294040
rect 350722 279712 350778 279721
rect 350722 279647 350778 279656
rect 350828 279070 350856 294034
rect 350816 279064 350868 279070
rect 350816 279006 350868 279012
rect 350722 276040 350778 276049
rect 350722 275975 350778 275984
rect 350630 262712 350686 262721
rect 350630 262647 350686 262656
rect 350540 255468 350592 255474
rect 350540 255410 350592 255416
rect 350356 255400 350408 255406
rect 350356 255342 350408 255348
rect 350446 255368 350502 255377
rect 350446 255303 350448 255312
rect 350500 255303 350502 255312
rect 350448 255274 350500 255280
rect 350446 254008 350502 254017
rect 350446 253943 350448 253952
rect 350500 253943 350502 253952
rect 350448 253914 350500 253920
rect 350446 250200 350502 250209
rect 350446 250135 350502 250144
rect 350460 249830 350488 250135
rect 350448 249824 350500 249830
rect 350448 249766 350500 249772
rect 350446 248840 350502 248849
rect 350446 248775 350502 248784
rect 350460 248470 350488 248775
rect 350448 248464 350500 248470
rect 350448 248406 350500 248412
rect 350446 245984 350502 245993
rect 350446 245919 350502 245928
rect 350460 245682 350488 245919
rect 350448 245676 350500 245682
rect 350448 245618 350500 245624
rect 350538 244488 350594 244497
rect 350538 244423 350594 244432
rect 350446 244352 350502 244361
rect 350446 244287 350448 244296
rect 350500 244287 350502 244296
rect 350448 244258 350500 244264
rect 350446 243264 350502 243273
rect 350446 243199 350502 243208
rect 350460 242962 350488 243199
rect 350448 242956 350500 242962
rect 350448 242898 350500 242904
rect 350264 239420 350316 239426
rect 350264 239362 350316 239368
rect 350446 239320 350502 239329
rect 350446 239255 350502 239264
rect 350460 239018 350488 239255
rect 350448 239012 350500 239018
rect 350448 238954 350500 238960
rect 350446 238912 350502 238921
rect 350356 238876 350408 238882
rect 350446 238847 350502 238856
rect 350356 238818 350408 238824
rect 350368 224942 350396 238818
rect 350460 238814 350488 238847
rect 350448 238808 350500 238814
rect 350448 238750 350500 238756
rect 350448 237380 350500 237386
rect 350448 237322 350500 237328
rect 350460 236201 350488 237322
rect 350446 236192 350502 236201
rect 350446 236127 350502 236136
rect 350446 235104 350502 235113
rect 350446 235039 350502 235048
rect 350460 234666 350488 235039
rect 350448 234660 350500 234666
rect 350448 234602 350500 234608
rect 350446 232248 350502 232257
rect 350446 232183 350502 232192
rect 350460 231878 350488 232183
rect 350448 231872 350500 231878
rect 350448 231814 350500 231820
rect 350446 230616 350502 230625
rect 350446 230551 350502 230560
rect 350460 230518 350488 230551
rect 350448 230512 350500 230518
rect 350448 230454 350500 230460
rect 350446 229256 350502 229265
rect 350446 229191 350502 229200
rect 350460 229158 350488 229191
rect 350448 229152 350500 229158
rect 350448 229094 350500 229100
rect 350356 224936 350408 224942
rect 350356 224878 350408 224884
rect 350448 223576 350500 223582
rect 350448 223518 350500 223524
rect 350460 222601 350488 223518
rect 350446 222592 350502 222601
rect 350446 222527 350502 222536
rect 350446 221232 350502 221241
rect 350446 221167 350448 221176
rect 350500 221167 350502 221176
rect 350448 221138 350500 221144
rect 350446 218104 350502 218113
rect 350446 218039 350448 218048
rect 350500 218039 350502 218048
rect 350448 218010 350500 218016
rect 350356 218000 350408 218006
rect 350356 217942 350408 217948
rect 350368 217161 350396 217942
rect 350446 217560 350502 217569
rect 350446 217495 350502 217504
rect 350460 217258 350488 217495
rect 350448 217252 350500 217258
rect 350448 217194 350500 217200
rect 350354 217152 350410 217161
rect 350354 217087 350410 217096
rect 350446 215384 350502 215393
rect 350446 215319 350448 215328
rect 350500 215319 350502 215328
rect 350448 215290 350500 215296
rect 350446 213208 350502 213217
rect 350446 213143 350502 213152
rect 350460 212566 350488 213143
rect 350448 212560 350500 212566
rect 350448 212502 350500 212508
rect 350446 209944 350502 209953
rect 350446 209879 350448 209888
rect 350500 209879 350502 209888
rect 350448 209850 350500 209856
rect 350446 209128 350502 209137
rect 350446 209063 350502 209072
rect 350460 208418 350488 209063
rect 350448 208412 350500 208418
rect 350448 208354 350500 208360
rect 350446 207768 350502 207777
rect 350446 207703 350502 207712
rect 350354 207360 350410 207369
rect 350354 207295 350410 207304
rect 350368 207058 350396 207295
rect 350460 207126 350488 207703
rect 350448 207120 350500 207126
rect 350448 207062 350500 207068
rect 350356 207052 350408 207058
rect 350356 206994 350408 207000
rect 350448 206984 350500 206990
rect 350446 206952 350448 206961
rect 350500 206952 350502 206961
rect 350446 206887 350502 206896
rect 350354 205048 350410 205057
rect 350354 204983 350410 204992
rect 350368 204338 350396 204983
rect 350356 204332 350408 204338
rect 350356 204274 350408 204280
rect 350448 204264 350500 204270
rect 350446 204232 350448 204241
rect 350500 204232 350502 204241
rect 350446 204167 350502 204176
rect 350080 203584 350132 203590
rect 350080 203526 350132 203532
rect 350446 203280 350502 203289
rect 350446 203215 350502 203224
rect 350460 202910 350488 203215
rect 350448 202904 350500 202910
rect 350448 202846 350500 202852
rect 350446 201920 350502 201929
rect 350446 201855 350502 201864
rect 350460 201550 350488 201855
rect 350448 201544 350500 201550
rect 350448 201486 350500 201492
rect 349986 195528 350042 195537
rect 349986 195463 350042 195472
rect 350552 193662 350580 244423
rect 350540 193656 350592 193662
rect 350540 193598 350592 193604
rect 350736 170610 350764 275975
rect 350814 272232 350870 272241
rect 350814 272167 350870 272176
rect 350828 186862 350856 272167
rect 350816 186856 350868 186862
rect 350816 186798 350868 186804
rect 351012 177682 351040 338127
rect 351104 188902 351132 364511
rect 351092 188896 351144 188902
rect 351092 188838 351144 188844
rect 351092 186856 351144 186862
rect 351092 186798 351144 186804
rect 351000 177676 351052 177682
rect 351000 177618 351052 177624
rect 350724 170604 350776 170610
rect 350724 170546 350776 170552
rect 350448 166320 350500 166326
rect 350448 166262 350500 166268
rect 349724 151786 349936 151814
rect 349724 149938 349752 151786
rect 350460 149940 350488 166262
rect 351104 149940 351132 186798
rect 351196 172174 351224 379743
rect 351288 183122 351316 390526
rect 351368 274712 351420 274718
rect 351368 274654 351420 274660
rect 351380 200433 351408 274654
rect 351472 248198 351500 585822
rect 353300 572076 353352 572082
rect 353300 572018 353352 572024
rect 352564 571056 352616 571062
rect 352564 570998 352616 571004
rect 352196 570716 352248 570722
rect 352196 570658 352248 570664
rect 352012 569492 352064 569498
rect 352012 569434 352064 569440
rect 351920 567588 351972 567594
rect 351920 567530 351972 567536
rect 351828 261452 351880 261458
rect 351828 261394 351880 261400
rect 351460 248192 351512 248198
rect 351460 248134 351512 248140
rect 351460 247104 351512 247110
rect 351460 247046 351512 247052
rect 351366 200424 351422 200433
rect 351366 200359 351422 200368
rect 351472 192846 351500 247046
rect 351840 244254 351868 261394
rect 351828 244248 351880 244254
rect 351828 244190 351880 244196
rect 351460 192840 351512 192846
rect 351460 192782 351512 192788
rect 351276 183116 351328 183122
rect 351276 183058 351328 183064
rect 351184 172168 351236 172174
rect 351184 172110 351236 172116
rect 351932 152522 351960 567530
rect 352024 196518 352052 569434
rect 352104 567248 352156 567254
rect 352104 567190 352156 567196
rect 352116 549234 352144 567190
rect 352104 549228 352156 549234
rect 352104 549170 352156 549176
rect 352104 520328 352156 520334
rect 352104 520270 352156 520276
rect 352012 196512 352064 196518
rect 352012 196454 352064 196460
rect 352116 177818 352144 520270
rect 352208 386374 352236 570658
rect 352288 567860 352340 567866
rect 352288 567802 352340 567808
rect 352300 489870 352328 567802
rect 352288 489864 352340 489870
rect 352288 489806 352340 489812
rect 352288 484424 352340 484430
rect 352288 484366 352340 484372
rect 352196 386368 352248 386374
rect 352196 386310 352248 386316
rect 352300 189582 352328 484366
rect 352380 473408 352432 473414
rect 352380 473350 352432 473356
rect 352392 196722 352420 473350
rect 352472 421048 352524 421054
rect 352472 420990 352524 420996
rect 352380 196716 352432 196722
rect 352380 196658 352432 196664
rect 352288 189576 352340 189582
rect 352288 189518 352340 189524
rect 352484 186930 352512 420990
rect 352576 378146 352604 570998
rect 352656 569288 352708 569294
rect 352656 569230 352708 569236
rect 352668 396846 352696 569230
rect 353312 554742 353340 572018
rect 353392 569356 353444 569362
rect 353392 569298 353444 569304
rect 353300 554736 353352 554742
rect 353300 554678 353352 554684
rect 352656 396840 352708 396846
rect 352656 396782 352708 396788
rect 352840 394732 352892 394738
rect 352840 394674 352892 394680
rect 352656 385008 352708 385014
rect 352656 384950 352708 384956
rect 352564 378140 352616 378146
rect 352564 378082 352616 378088
rect 352564 362976 352616 362982
rect 352564 362918 352616 362924
rect 352576 192642 352604 362918
rect 352668 214577 352696 384950
rect 352748 215348 352800 215354
rect 352748 215290 352800 215296
rect 352654 214568 352710 214577
rect 352654 214503 352710 214512
rect 352656 213920 352708 213926
rect 352656 213862 352708 213868
rect 352668 193798 352696 213862
rect 352656 193792 352708 193798
rect 352656 193734 352708 193740
rect 352564 192636 352616 192642
rect 352564 192578 352616 192584
rect 352472 186924 352524 186930
rect 352472 186866 352524 186872
rect 352104 177812 352156 177818
rect 352104 177754 352156 177760
rect 352760 170746 352788 215290
rect 352748 170740 352800 170746
rect 352748 170682 352800 170688
rect 351920 152516 351972 152522
rect 351920 152458 351972 152464
rect 352852 151814 352880 394674
rect 353404 192778 353432 569298
rect 353852 569220 353904 569226
rect 353852 569162 353904 569168
rect 353760 566772 353812 566778
rect 353760 566714 353812 566720
rect 353576 566636 353628 566642
rect 353576 566578 353628 566584
rect 353484 566500 353536 566506
rect 353484 566442 353536 566448
rect 353496 195226 353524 566442
rect 353588 199918 353616 566578
rect 353668 531344 353720 531350
rect 353668 531286 353720 531292
rect 353576 199912 353628 199918
rect 353576 199854 353628 199860
rect 353484 195220 353536 195226
rect 353484 195162 353536 195168
rect 353392 192772 353444 192778
rect 353392 192714 353444 192720
rect 353680 185978 353708 531286
rect 353772 524414 353800 566714
rect 353760 524408 353812 524414
rect 353760 524350 353812 524356
rect 353760 513460 353812 513466
rect 353760 513402 353812 513408
rect 353772 187610 353800 513402
rect 353864 247110 353892 569162
rect 353956 487257 353984 677622
rect 355048 589552 355100 589558
rect 355048 589494 355100 589500
rect 354772 589484 354824 589490
rect 354772 589426 354824 589432
rect 354680 587716 354732 587722
rect 354680 587658 354732 587664
rect 354036 567384 354088 567390
rect 354036 567326 354088 567332
rect 354048 542366 354076 567326
rect 354128 563712 354180 563718
rect 354128 563654 354180 563660
rect 354036 542360 354088 542366
rect 354036 542302 354088 542308
rect 354036 498228 354088 498234
rect 354036 498170 354088 498176
rect 353942 487248 353998 487257
rect 353942 487183 353998 487192
rect 353944 472048 353996 472054
rect 353944 471990 353996 471996
rect 353852 247104 353904 247110
rect 353852 247046 353904 247052
rect 353852 231872 353904 231878
rect 353852 231814 353904 231820
rect 353760 187604 353812 187610
rect 353760 187546 353812 187552
rect 353668 185972 353720 185978
rect 353668 185914 353720 185920
rect 353864 181898 353892 231814
rect 353852 181892 353904 181898
rect 353852 181834 353904 181840
rect 353956 158166 353984 471990
rect 354048 194274 354076 498170
rect 354140 274718 354168 563654
rect 354220 563100 354272 563106
rect 354220 563042 354272 563048
rect 354128 274712 354180 274718
rect 354128 274654 354180 274660
rect 354128 253496 354180 253502
rect 354128 253438 354180 253444
rect 354036 194268 354088 194274
rect 354036 194210 354088 194216
rect 354140 189718 354168 253438
rect 354128 189712 354180 189718
rect 354128 189654 354180 189660
rect 353944 158160 353996 158166
rect 353944 158102 353996 158108
rect 354232 155786 354260 563042
rect 354692 192302 354720 587658
rect 354784 198286 354812 589426
rect 354956 575000 355008 575006
rect 354956 574942 355008 574948
rect 354864 563916 354916 563922
rect 354864 563858 354916 563864
rect 354772 198280 354824 198286
rect 354772 198222 354824 198228
rect 354680 192296 354732 192302
rect 354680 192238 354732 192244
rect 354876 191078 354904 563858
rect 354968 218006 354996 574942
rect 355060 253502 355088 589494
rect 355140 589416 355192 589422
rect 355140 589358 355192 589364
rect 355152 261458 355180 589358
rect 356152 569424 356204 569430
rect 356152 569366 356204 569372
rect 356060 567452 356112 567458
rect 356060 567394 356112 567400
rect 355416 565072 355468 565078
rect 355416 565014 355468 565020
rect 355232 561740 355284 561746
rect 355232 561682 355284 561688
rect 355140 261452 355192 261458
rect 355140 261394 355192 261400
rect 355048 253496 355100 253502
rect 355048 253438 355100 253444
rect 355140 244248 355192 244254
rect 355140 244190 355192 244196
rect 355048 218068 355100 218074
rect 355048 218010 355100 218016
rect 354956 218000 355008 218006
rect 354956 217942 355008 217948
rect 354864 191072 354916 191078
rect 354864 191014 354916 191020
rect 355060 173262 355088 218010
rect 355152 213926 355180 244190
rect 355244 238882 355272 561682
rect 355324 561196 355376 561202
rect 355324 561138 355376 561144
rect 355232 238876 355284 238882
rect 355232 238818 355284 238824
rect 355232 217252 355284 217258
rect 355232 217194 355284 217200
rect 355140 213920 355192 213926
rect 355140 213862 355192 213868
rect 355244 190058 355272 217194
rect 355232 190052 355284 190058
rect 355232 189994 355284 190000
rect 355048 173256 355100 173262
rect 355048 173198 355100 173204
rect 354312 169244 354364 169250
rect 354312 169186 354364 169192
rect 354220 155780 354272 155786
rect 354220 155722 354272 155728
rect 352760 151786 352880 151814
rect 352760 149954 352788 151786
rect 349712 149932 349764 149938
rect 352406 149926 352788 149954
rect 354324 149940 354352 169186
rect 354864 153128 354916 153134
rect 354864 153070 354916 153076
rect 354956 153128 355008 153134
rect 354956 153070 355008 153076
rect 354876 152930 354904 153070
rect 354772 152924 354824 152930
rect 354772 152866 354824 152872
rect 354864 152924 354916 152930
rect 354864 152866 354916 152872
rect 354784 152522 354812 152866
rect 354772 152516 354824 152522
rect 354772 152458 354824 152464
rect 354968 149940 354996 153070
rect 355336 152386 355364 561138
rect 355428 220794 355456 565014
rect 355508 358012 355560 358018
rect 355508 357954 355560 357960
rect 355416 220788 355468 220794
rect 355416 220730 355468 220736
rect 355520 181966 355548 357954
rect 355692 253972 355744 253978
rect 355692 253914 355744 253920
rect 355600 233912 355652 233918
rect 355600 233854 355652 233860
rect 355508 181960 355560 181966
rect 355508 181902 355560 181908
rect 355324 152380 355376 152386
rect 355324 152322 355376 152328
rect 355612 149940 355640 233854
rect 355704 191486 355732 253914
rect 355692 191480 355744 191486
rect 355692 191422 355744 191428
rect 356072 152998 356100 567394
rect 356164 194002 356192 569366
rect 357440 568880 357492 568886
rect 357440 568822 357492 568828
rect 356428 567996 356480 568002
rect 356428 567938 356480 567944
rect 356336 564460 356388 564466
rect 356336 564402 356388 564408
rect 356244 559020 356296 559026
rect 356244 558962 356296 558968
rect 356152 193996 356204 194002
rect 356152 193938 356204 193944
rect 356256 185910 356284 558962
rect 356348 191690 356376 564402
rect 356440 371210 356468 567938
rect 356702 562456 356758 562465
rect 356702 562391 356758 562400
rect 356428 371204 356480 371210
rect 356428 371146 356480 371152
rect 356428 224936 356480 224942
rect 356428 224878 356480 224884
rect 356336 191684 356388 191690
rect 356336 191626 356388 191632
rect 356244 185904 356296 185910
rect 356244 185846 356296 185852
rect 356440 170678 356468 224878
rect 356520 221196 356572 221202
rect 356520 221138 356572 221144
rect 356532 193866 356560 221138
rect 356612 209908 356664 209914
rect 356612 209850 356664 209856
rect 356520 193860 356572 193866
rect 356520 193802 356572 193808
rect 356624 185842 356652 209850
rect 356716 204921 356744 562391
rect 356796 551132 356848 551138
rect 356796 551074 356848 551080
rect 356808 210526 356836 551074
rect 356888 525972 356940 525978
rect 356888 525914 356940 525920
rect 356900 222902 356928 525914
rect 356980 419552 357032 419558
rect 356980 419494 357032 419500
rect 356888 222896 356940 222902
rect 356888 222838 356940 222844
rect 356796 210520 356848 210526
rect 356796 210462 356848 210468
rect 356702 204912 356758 204921
rect 356702 204847 356758 204856
rect 356992 199889 357020 419494
rect 357072 334076 357124 334082
rect 357072 334018 357124 334024
rect 357084 224398 357112 334018
rect 357164 287156 357216 287162
rect 357164 287098 357216 287104
rect 357176 225690 357204 287098
rect 357164 225684 357216 225690
rect 357164 225626 357216 225632
rect 357072 224392 357124 224398
rect 357072 224334 357124 224340
rect 356978 199880 357034 199889
rect 356978 199815 357034 199824
rect 356612 185836 356664 185842
rect 356612 185778 356664 185784
rect 356428 170672 356480 170678
rect 356428 170614 356480 170620
rect 356244 162444 356296 162450
rect 356244 162386 356296 162392
rect 356060 152992 356112 152998
rect 356060 152934 356112 152940
rect 356256 149940 356284 162386
rect 357452 152794 357480 568822
rect 357532 568744 357584 568750
rect 357532 568686 357584 568692
rect 357440 152788 357492 152794
rect 357440 152730 357492 152736
rect 357544 152590 357572 568686
rect 357624 220788 357676 220794
rect 357624 220730 357676 220736
rect 357636 155174 357664 220730
rect 357624 155168 357676 155174
rect 357624 155110 357676 155116
rect 358096 153134 358124 679186
rect 358176 640348 358228 640354
rect 358176 640290 358228 640296
rect 358188 159866 358216 640290
rect 359280 587784 359332 587790
rect 359280 587726 359332 587732
rect 359004 567928 359056 567934
rect 359004 567870 359056 567876
rect 358544 567520 358596 567526
rect 358544 567462 358596 567468
rect 358266 564768 358322 564777
rect 358266 564703 358322 564712
rect 358176 159860 358228 159866
rect 358176 159802 358228 159808
rect 358280 158409 358308 564703
rect 358360 561808 358412 561814
rect 358360 561750 358412 561756
rect 358372 162518 358400 561750
rect 358452 549296 358504 549302
rect 358452 549238 358504 549244
rect 358464 199238 358492 549238
rect 358556 237969 358584 567462
rect 358820 564800 358872 564806
rect 358820 564742 358872 564748
rect 358636 560584 358688 560590
rect 358636 560526 358688 560532
rect 358648 322930 358676 560526
rect 358636 322924 358688 322930
rect 358636 322866 358688 322872
rect 358636 269136 358688 269142
rect 358636 269078 358688 269084
rect 358542 237960 358598 237969
rect 358542 237895 358598 237904
rect 358544 231804 358596 231810
rect 358544 231746 358596 231752
rect 358452 199232 358504 199238
rect 358452 199174 358504 199180
rect 358556 191554 358584 231746
rect 358648 193730 358676 269078
rect 358728 244928 358780 244934
rect 358728 244870 358780 244876
rect 358740 223514 358768 244870
rect 358728 223508 358780 223514
rect 358728 223450 358780 223456
rect 358636 193724 358688 193730
rect 358636 193666 358688 193672
rect 358544 191548 358596 191554
rect 358544 191490 358596 191496
rect 358360 162512 358412 162518
rect 358360 162454 358412 162460
rect 358266 158400 358322 158409
rect 358266 158335 358322 158344
rect 358084 153128 358136 153134
rect 358084 153070 358136 153076
rect 358832 153066 358860 564742
rect 358912 532840 358964 532846
rect 358912 532782 358964 532788
rect 358924 158370 358952 532782
rect 359016 231810 359044 567870
rect 359096 491428 359148 491434
rect 359096 491370 359148 491376
rect 359004 231804 359056 231810
rect 359004 231746 359056 231752
rect 359004 229152 359056 229158
rect 359004 229094 359056 229100
rect 359016 177750 359044 229094
rect 359108 195430 359136 491370
rect 359188 425128 359240 425134
rect 359188 425070 359240 425076
rect 359096 195424 359148 195430
rect 359096 195366 359148 195372
rect 359200 192370 359228 425070
rect 359292 384334 359320 587726
rect 360200 570920 360252 570926
rect 360200 570862 360252 570868
rect 359462 562184 359518 562193
rect 359462 562119 359518 562128
rect 359280 384328 359332 384334
rect 359280 384270 359332 384276
rect 359280 332648 359332 332654
rect 359280 332590 359332 332596
rect 359188 192364 359240 192370
rect 359188 192306 359240 192312
rect 359292 187542 359320 332590
rect 359372 245676 359424 245682
rect 359372 245618 359424 245624
rect 359280 187536 359332 187542
rect 359280 187478 359332 187484
rect 359004 177744 359056 177750
rect 359004 177686 359056 177692
rect 359384 172038 359412 245618
rect 359372 172032 359424 172038
rect 359372 171974 359424 171980
rect 358912 158364 358964 158370
rect 358912 158306 358964 158312
rect 359476 156913 359504 562119
rect 359556 409896 359608 409902
rect 359556 409838 359608 409844
rect 359462 156904 359518 156913
rect 359462 156839 359518 156848
rect 359568 154086 359596 409838
rect 359648 354748 359700 354754
rect 359648 354690 359700 354696
rect 359660 224262 359688 354690
rect 359648 224256 359700 224262
rect 359648 224198 359700 224204
rect 359648 223508 359700 223514
rect 359648 223450 359700 223456
rect 359660 190398 359688 223450
rect 360212 198626 360240 570862
rect 360382 563136 360438 563145
rect 360382 563071 360438 563080
rect 360292 503736 360344 503742
rect 360292 503678 360344 503684
rect 360200 198620 360252 198626
rect 360200 198562 360252 198568
rect 359648 190392 359700 190398
rect 359648 190334 359700 190340
rect 360304 184550 360332 503678
rect 360396 265033 360424 563071
rect 360476 398880 360528 398886
rect 360476 398822 360528 398828
rect 360382 265024 360438 265033
rect 360382 264959 360438 264968
rect 360384 263628 360436 263634
rect 360384 263570 360436 263576
rect 360396 262206 360424 263570
rect 360384 262200 360436 262206
rect 360384 262142 360436 262148
rect 360384 234660 360436 234666
rect 360384 234602 360436 234608
rect 360396 192574 360424 234602
rect 360384 192568 360436 192574
rect 360384 192510 360436 192516
rect 360292 184544 360344 184550
rect 360292 184486 360344 184492
rect 360488 172106 360516 398822
rect 360476 172100 360528 172106
rect 360476 172042 360528 172048
rect 359556 154080 359608 154086
rect 359556 154022 359608 154028
rect 358820 153060 358872 153066
rect 358820 153002 358872 153008
rect 357532 152584 357584 152590
rect 357532 152526 357584 152532
rect 360856 152522 360884 682110
rect 360936 576904 360988 576910
rect 360936 576846 360988 576852
rect 360948 159798 360976 576846
rect 363604 571396 363656 571402
rect 363604 571338 363656 571344
rect 363696 571396 363748 571402
rect 363696 571338 363748 571344
rect 361672 571124 361724 571130
rect 361672 571066 361724 571072
rect 361580 563372 361632 563378
rect 361580 563314 361632 563320
rect 361028 469260 361080 469266
rect 361028 469202 361080 469208
rect 361040 199442 361068 469202
rect 361120 426556 361172 426562
rect 361120 426498 361172 426504
rect 361028 199436 361080 199442
rect 361028 199378 361080 199384
rect 361132 199034 361160 426498
rect 361304 343732 361356 343738
rect 361304 343674 361356 343680
rect 361212 299532 361264 299538
rect 361212 299474 361264 299480
rect 361120 199028 361172 199034
rect 361120 198970 361172 198976
rect 361224 179110 361252 299474
rect 361316 251870 361344 343674
rect 361304 251864 361356 251870
rect 361304 251806 361356 251812
rect 361304 249892 361356 249898
rect 361304 249834 361356 249840
rect 361212 179104 361264 179110
rect 361212 179046 361264 179052
rect 361316 165170 361344 249834
rect 361304 165164 361356 165170
rect 361304 165106 361356 165112
rect 360936 159792 360988 159798
rect 360936 159734 360988 159740
rect 361592 152930 361620 563314
rect 361684 199306 361712 571066
rect 363052 568200 363104 568206
rect 363052 568142 363104 568148
rect 361762 560688 361818 560697
rect 361762 560623 361818 560632
rect 361776 200802 361804 560623
rect 362224 534132 362276 534138
rect 362224 534074 362276 534080
rect 361856 516180 361908 516186
rect 361856 516122 361908 516128
rect 361764 200796 361816 200802
rect 361764 200738 361816 200744
rect 361672 199300 361724 199306
rect 361672 199242 361724 199248
rect 361868 191418 361896 516122
rect 361948 476196 362000 476202
rect 361948 476138 362000 476144
rect 361856 191412 361908 191418
rect 361856 191354 361908 191360
rect 361960 187406 361988 476138
rect 362040 350600 362092 350606
rect 362040 350542 362092 350548
rect 362052 187474 362080 350542
rect 362236 227254 362264 534074
rect 362960 461100 363012 461106
rect 362960 461042 363012 461048
rect 362316 460964 362368 460970
rect 362316 460906 362368 460912
rect 362224 227248 362276 227254
rect 362224 227190 362276 227196
rect 362040 187468 362092 187474
rect 362040 187410 362092 187416
rect 361948 187400 362000 187406
rect 361948 187342 362000 187348
rect 362328 165034 362356 460906
rect 362500 449948 362552 449954
rect 362500 449890 362552 449896
rect 362408 441652 362460 441658
rect 362408 441594 362460 441600
rect 362420 193934 362448 441594
rect 362512 371210 362540 449890
rect 362500 371204 362552 371210
rect 362500 371146 362552 371152
rect 362500 327140 362552 327146
rect 362500 327082 362552 327088
rect 362408 193928 362460 193934
rect 362408 193870 362460 193876
rect 362316 165028 362368 165034
rect 362316 164970 362368 164976
rect 362512 159594 362540 327082
rect 362972 184414 363000 461042
rect 363064 296682 363092 568142
rect 363144 358828 363196 358834
rect 363144 358770 363196 358776
rect 363052 296676 363104 296682
rect 363052 296618 363104 296624
rect 363052 294024 363104 294030
rect 363052 293966 363104 293972
rect 363064 188562 363092 293966
rect 363156 188630 363184 358770
rect 363328 200796 363380 200802
rect 363328 200738 363380 200744
rect 363144 188624 363196 188630
rect 363144 188566 363196 188572
rect 363052 188556 363104 188562
rect 363052 188498 363104 188504
rect 362960 184408 363012 184414
rect 362960 184350 363012 184356
rect 362500 159588 362552 159594
rect 362500 159530 362552 159536
rect 361580 152924 361632 152930
rect 361580 152866 361632 152872
rect 360844 152516 360896 152522
rect 360844 152458 360896 152464
rect 360198 152280 360254 152289
rect 360198 152215 360254 152224
rect 360212 151842 360240 152215
rect 360200 151836 360252 151842
rect 360200 151778 360252 151784
rect 360108 151564 360160 151570
rect 360108 151506 360160 151512
rect 360120 149940 360148 151506
rect 363340 149940 363368 200738
rect 363616 159633 363644 571338
rect 363708 199170 363736 571338
rect 363788 562556 363840 562562
rect 363788 562498 363840 562504
rect 363800 224330 363828 562498
rect 363880 562216 363932 562222
rect 363880 562158 363932 562164
rect 363892 240145 363920 562158
rect 363972 434784 364024 434790
rect 363972 434726 364024 434732
rect 363878 240136 363934 240145
rect 363878 240071 363934 240080
rect 363788 224324 363840 224330
rect 363788 224266 363840 224272
rect 363696 199164 363748 199170
rect 363696 199106 363748 199112
rect 363984 174690 364012 434726
rect 364064 349240 364116 349246
rect 364064 349182 364116 349188
rect 364076 307766 364104 349182
rect 364064 307760 364116 307766
rect 364064 307702 364116 307708
rect 364064 292596 364116 292602
rect 364064 292538 364116 292544
rect 364076 180538 364104 292538
rect 364260 262993 364288 682586
rect 364984 665236 365036 665242
rect 364984 665178 365036 665184
rect 364340 607232 364392 607238
rect 364340 607174 364392 607180
rect 364246 262984 364302 262993
rect 364246 262919 364302 262928
rect 364156 262268 364208 262274
rect 364156 262210 364208 262216
rect 364064 180532 364116 180538
rect 364064 180474 364116 180480
rect 364168 177886 364196 262210
rect 364352 195498 364380 607174
rect 364432 559088 364484 559094
rect 364432 559030 364484 559036
rect 364340 195492 364392 195498
rect 364340 195434 364392 195440
rect 364444 182034 364472 559030
rect 364524 461032 364576 461038
rect 364524 460974 364576 460980
rect 364536 184278 364564 460974
rect 364616 404456 364668 404462
rect 364616 404398 364668 404404
rect 364524 184272 364576 184278
rect 364524 184214 364576 184220
rect 364432 182028 364484 182034
rect 364432 181970 364484 181976
rect 364156 177880 364208 177886
rect 364156 177822 364208 177828
rect 363972 174684 364024 174690
rect 363972 174626 364024 174632
rect 364628 174622 364656 404398
rect 364708 325712 364760 325718
rect 364708 325654 364760 325660
rect 364720 322862 364748 325654
rect 364708 322856 364760 322862
rect 364708 322798 364760 322804
rect 364708 273352 364760 273358
rect 364708 273294 364760 273300
rect 364720 184929 364748 273294
rect 364996 197878 365024 665178
rect 365812 605872 365864 605878
rect 365812 605814 365864 605820
rect 365260 562624 365312 562630
rect 365260 562566 365312 562572
rect 365076 562420 365128 562426
rect 365076 562362 365128 562368
rect 365088 231130 365116 562362
rect 365168 538280 365220 538286
rect 365168 538222 365220 538228
rect 365076 231124 365128 231130
rect 365076 231066 365128 231072
rect 365180 218754 365208 538222
rect 365272 297430 365300 562566
rect 365720 561876 365772 561882
rect 365720 561818 365772 561824
rect 365444 349172 365496 349178
rect 365444 349114 365496 349120
rect 365352 303680 365404 303686
rect 365352 303622 365404 303628
rect 365260 297424 365312 297430
rect 365260 297366 365312 297372
rect 365260 295384 365312 295390
rect 365260 295326 365312 295332
rect 365272 227050 365300 295326
rect 365260 227044 365312 227050
rect 365260 226986 365312 226992
rect 365168 218748 365220 218754
rect 365168 218690 365220 218696
rect 364984 197872 365036 197878
rect 364984 197814 365036 197820
rect 365364 191282 365392 303622
rect 365456 284306 365484 349114
rect 365444 284300 365496 284306
rect 365444 284242 365496 284248
rect 365352 191276 365404 191282
rect 365352 191218 365404 191224
rect 364706 184920 364762 184929
rect 364706 184855 364762 184864
rect 364616 174616 364668 174622
rect 364616 174558 364668 174564
rect 363602 159624 363658 159633
rect 363602 159559 363658 159568
rect 365732 151473 365760 561818
rect 365824 196790 365852 605814
rect 366364 568948 366416 568954
rect 366364 568890 366416 568896
rect 365994 562320 366050 562329
rect 365994 562255 366050 562264
rect 365902 561912 365958 561921
rect 365902 561847 365958 561856
rect 365812 196784 365864 196790
rect 365812 196726 365864 196732
rect 365916 155310 365944 561847
rect 366008 155446 366036 562255
rect 366088 480344 366140 480350
rect 366088 480286 366140 480292
rect 366100 180577 366128 480286
rect 366086 180568 366142 180577
rect 366086 180503 366142 180512
rect 366376 156777 366404 568890
rect 367100 563236 367152 563242
rect 367100 563178 367152 563184
rect 366456 527196 366508 527202
rect 366456 527138 366508 527144
rect 366362 156768 366418 156777
rect 366362 156703 366418 156712
rect 366468 155961 366496 527138
rect 366548 452668 366600 452674
rect 366548 452610 366600 452616
rect 366560 191049 366588 452610
rect 366640 360256 366692 360262
rect 366640 360198 366692 360204
rect 366652 194070 366680 360198
rect 366732 300892 366784 300898
rect 366732 300834 366784 300840
rect 366640 194064 366692 194070
rect 366640 194006 366692 194012
rect 366546 191040 366602 191049
rect 366546 190975 366602 190984
rect 366744 166598 366772 300834
rect 367112 190330 367140 563178
rect 367192 456884 367244 456890
rect 367192 456826 367244 456832
rect 367100 190324 367152 190330
rect 367100 190266 367152 190272
rect 367204 181830 367232 456826
rect 367284 447160 367336 447166
rect 367284 447102 367336 447108
rect 367296 184210 367324 447102
rect 367284 184204 367336 184210
rect 367284 184146 367336 184152
rect 367192 181824 367244 181830
rect 367192 181766 367244 181772
rect 366732 166592 366784 166598
rect 366732 166534 366784 166540
rect 366454 155952 366510 155961
rect 366454 155887 366510 155896
rect 365996 155440 366048 155446
rect 365996 155382 366048 155388
rect 365904 155304 365956 155310
rect 365904 155246 365956 155252
rect 367756 152454 367784 686054
rect 373264 682304 373316 682310
rect 373264 682246 373316 682252
rect 367836 667956 367888 667962
rect 367836 667898 367888 667904
rect 367848 198218 367876 667898
rect 369124 632120 369176 632126
rect 369124 632062 369176 632068
rect 368480 569968 368532 569974
rect 368480 569910 368532 569916
rect 368204 567316 368256 567322
rect 368204 567258 368256 567264
rect 367928 491360 367980 491366
rect 367928 491302 367980 491308
rect 367940 230042 367968 491302
rect 368020 405748 368072 405754
rect 368020 405690 368072 405696
rect 367928 230036 367980 230042
rect 367928 229978 367980 229984
rect 367836 198212 367888 198218
rect 367836 198154 367888 198160
rect 368032 179042 368060 405690
rect 368112 390584 368164 390590
rect 368112 390526 368164 390532
rect 368124 195634 368152 390526
rect 368216 386374 368244 567258
rect 368296 404388 368348 404394
rect 368296 404330 368348 404336
rect 368204 386368 368256 386374
rect 368204 386310 368256 386316
rect 368308 230110 368336 404330
rect 368296 230104 368348 230110
rect 368296 230046 368348 230052
rect 368112 195628 368164 195634
rect 368112 195570 368164 195576
rect 368020 179036 368072 179042
rect 368020 178978 368072 178984
rect 368492 172310 368520 569910
rect 368572 419620 368624 419626
rect 368572 419562 368624 419568
rect 368584 185881 368612 419562
rect 369136 197946 369164 632062
rect 372068 618316 372120 618322
rect 372068 618258 372120 618264
rect 369308 615528 369360 615534
rect 369308 615470 369360 615476
rect 369216 607232 369268 607238
rect 369216 607174 369268 607180
rect 369124 197940 369176 197946
rect 369124 197882 369176 197888
rect 368570 185872 368626 185881
rect 368570 185807 368626 185816
rect 369228 180198 369256 607174
rect 369320 198937 369348 615470
rect 371332 611380 371384 611386
rect 371332 611322 371384 611328
rect 371240 568812 371292 568818
rect 371240 568754 371292 568760
rect 370688 565956 370740 565962
rect 370688 565898 370740 565904
rect 369492 565140 369544 565146
rect 369492 565082 369544 565088
rect 369400 523048 369452 523054
rect 369400 522990 369452 522996
rect 369306 198928 369362 198937
rect 369306 198863 369362 198872
rect 369216 180192 369268 180198
rect 369216 180134 369268 180140
rect 368480 172304 368532 172310
rect 368480 172246 368532 172252
rect 369412 170610 369440 522990
rect 369504 455394 369532 565082
rect 369952 564936 370004 564942
rect 369952 564878 370004 564884
rect 369492 455388 369544 455394
rect 369492 455330 369544 455336
rect 369492 426624 369544 426630
rect 369492 426566 369544 426572
rect 369504 181665 369532 426566
rect 369584 419620 369636 419626
rect 369584 419562 369636 419568
rect 369596 183054 369624 419562
rect 369676 356244 369728 356250
rect 369676 356186 369728 356192
rect 369688 195770 369716 356186
rect 369768 303748 369820 303754
rect 369768 303690 369820 303696
rect 369780 229838 369808 303690
rect 369768 229832 369820 229838
rect 369768 229774 369820 229780
rect 369676 195764 369728 195770
rect 369676 195706 369728 195712
rect 369964 189990 369992 564878
rect 370504 516180 370556 516186
rect 370504 516122 370556 516128
rect 370044 481704 370096 481710
rect 370044 481646 370096 481652
rect 369952 189984 370004 189990
rect 369952 189926 370004 189932
rect 369584 183048 369636 183054
rect 369584 182990 369636 182996
rect 370056 181762 370084 481646
rect 370136 480276 370188 480282
rect 370136 480218 370188 480224
rect 370148 184346 370176 480218
rect 370228 434852 370280 434858
rect 370228 434794 370280 434800
rect 370240 189922 370268 434794
rect 370228 189916 370280 189922
rect 370228 189858 370280 189864
rect 370136 184340 370188 184346
rect 370136 184282 370188 184288
rect 370044 181756 370096 181762
rect 370044 181698 370096 181704
rect 369490 181656 369546 181665
rect 369490 181591 369546 181600
rect 369400 170604 369452 170610
rect 369400 170546 369452 170552
rect 369124 163736 369176 163742
rect 369124 163678 369176 163684
rect 367744 152448 367796 152454
rect 367744 152390 367796 152396
rect 365718 151464 365774 151473
rect 365718 151399 365774 151408
rect 369136 149940 369164 163678
rect 370516 157146 370544 516122
rect 370596 476128 370648 476134
rect 370596 476070 370648 476076
rect 370608 207670 370636 476070
rect 370700 325650 370728 565898
rect 370964 563644 371016 563650
rect 370964 563586 371016 563592
rect 370780 445800 370832 445806
rect 370780 445742 370832 445748
rect 370792 361554 370820 445742
rect 370780 361548 370832 361554
rect 370780 361490 370832 361496
rect 370780 339516 370832 339522
rect 370780 339458 370832 339464
rect 370688 325644 370740 325650
rect 370688 325586 370740 325592
rect 370688 317484 370740 317490
rect 370688 317426 370740 317432
rect 370700 235618 370728 317426
rect 370792 237386 370820 339458
rect 370872 328500 370924 328506
rect 370872 328442 370924 328448
rect 370780 237380 370832 237386
rect 370780 237322 370832 237328
rect 370688 235612 370740 235618
rect 370688 235554 370740 235560
rect 370884 230178 370912 328442
rect 370872 230172 370924 230178
rect 370872 230114 370924 230120
rect 370596 207664 370648 207670
rect 370596 207606 370648 207612
rect 370504 157140 370556 157146
rect 370504 157082 370556 157088
rect 370594 153096 370650 153105
rect 370594 153031 370650 153040
rect 370608 149954 370636 153031
rect 370454 149926 370636 149954
rect 370976 149938 371004 563586
rect 371252 155378 371280 568754
rect 371344 199102 371372 611322
rect 371976 588600 372028 588606
rect 371976 588542 372028 588548
rect 371884 546576 371936 546582
rect 371884 546518 371936 546524
rect 371424 263696 371476 263702
rect 371424 263638 371476 263644
rect 371332 199096 371384 199102
rect 371332 199038 371384 199044
rect 371436 170474 371464 263638
rect 371896 188426 371924 546518
rect 371988 292534 372016 588542
rect 372080 488510 372108 618258
rect 372252 566024 372304 566030
rect 372252 565966 372304 565972
rect 372068 488504 372120 488510
rect 372068 488446 372120 488452
rect 372068 473408 372120 473414
rect 372068 473350 372120 473356
rect 371976 292528 372028 292534
rect 371976 292470 372028 292476
rect 371976 256760 372028 256766
rect 371976 256702 372028 256708
rect 371884 188420 371936 188426
rect 371884 188362 371936 188368
rect 371424 170468 371476 170474
rect 371424 170410 371476 170416
rect 371988 163810 372016 256702
rect 372080 183190 372108 473350
rect 372160 400240 372212 400246
rect 372160 400182 372212 400188
rect 372068 183184 372120 183190
rect 372068 183126 372120 183132
rect 371976 163804 372028 163810
rect 371976 163746 372028 163752
rect 372172 159594 372200 400182
rect 372264 336734 372292 565966
rect 372620 563304 372672 563310
rect 372620 563246 372672 563252
rect 372344 418192 372396 418198
rect 372344 418134 372396 418140
rect 372252 336728 372304 336734
rect 372252 336670 372304 336676
rect 372252 300960 372304 300966
rect 372252 300902 372304 300908
rect 372264 229974 372292 300902
rect 372252 229968 372304 229974
rect 372252 229910 372304 229916
rect 372356 223582 372384 418134
rect 372436 349172 372488 349178
rect 372436 349114 372488 349120
rect 372344 223576 372396 223582
rect 372344 223518 372396 223524
rect 372448 169114 372476 349114
rect 372632 180470 372660 563246
rect 373172 321632 373224 321638
rect 373172 321574 373224 321580
rect 373184 230246 373212 321574
rect 373172 230240 373224 230246
rect 373172 230182 373224 230188
rect 372620 180464 372672 180470
rect 372620 180406 372672 180412
rect 373276 173398 373304 682246
rect 373356 608660 373408 608666
rect 373356 608602 373408 608608
rect 373368 176225 373396 608602
rect 373448 517540 373500 517546
rect 373448 517482 373500 517488
rect 373460 189786 373488 517482
rect 373540 484424 373592 484430
rect 373540 484366 373592 484372
rect 373448 189780 373500 189786
rect 373448 189722 373500 189728
rect 373552 180334 373580 484366
rect 373644 445670 373672 687890
rect 378784 685976 378836 685982
rect 378784 685918 378836 685924
rect 377404 683664 377456 683670
rect 377404 683606 377456 683612
rect 376024 601724 376076 601730
rect 376024 601666 376076 601672
rect 374000 567656 374052 567662
rect 374000 567598 374052 567604
rect 373632 445664 373684 445670
rect 373632 445606 373684 445612
rect 373816 430704 373868 430710
rect 373816 430646 373868 430652
rect 373724 389224 373776 389230
rect 373724 389166 373776 389172
rect 373632 290488 373684 290494
rect 373632 290430 373684 290436
rect 373540 180328 373592 180334
rect 373540 180270 373592 180276
rect 373354 176216 373410 176225
rect 373354 176151 373410 176160
rect 373264 173392 373316 173398
rect 373264 173334 373316 173340
rect 372436 169108 372488 169114
rect 372436 169050 372488 169056
rect 372342 167784 372398 167793
rect 372342 167719 372398 167728
rect 372160 159588 372212 159594
rect 372160 159530 372212 159536
rect 371240 155372 371292 155378
rect 371240 155314 371292 155320
rect 372356 149940 372384 167719
rect 373644 149940 373672 290430
rect 373736 159798 373764 389166
rect 373828 231198 373856 430646
rect 373908 322992 373960 322998
rect 373908 322934 373960 322940
rect 373816 231192 373868 231198
rect 373816 231134 373868 231140
rect 373920 170814 373948 322934
rect 374012 188494 374040 567598
rect 374920 567248 374972 567254
rect 374920 567190 374972 567196
rect 374644 560924 374696 560930
rect 374644 560866 374696 560872
rect 374092 329860 374144 329866
rect 374092 329802 374144 329808
rect 374000 188488 374052 188494
rect 374000 188430 374052 188436
rect 373908 170808 373960 170814
rect 373908 170750 373960 170756
rect 374104 170542 374132 329802
rect 374092 170536 374144 170542
rect 374092 170478 374144 170484
rect 373724 159792 373776 159798
rect 373724 159734 373776 159740
rect 374656 153202 374684 560866
rect 374828 423700 374880 423706
rect 374828 423642 374880 423648
rect 374736 414112 374788 414118
rect 374736 414054 374788 414060
rect 374748 159866 374776 414054
rect 374840 176254 374868 423642
rect 374932 375358 374960 567190
rect 375380 506524 375432 506530
rect 375380 506466 375432 506472
rect 375012 427848 375064 427854
rect 375012 427790 375064 427796
rect 374920 375352 374972 375358
rect 374920 375294 374972 375300
rect 374920 372632 374972 372638
rect 374920 372574 374972 372580
rect 374828 176248 374880 176254
rect 374828 176190 374880 176196
rect 374736 159860 374788 159866
rect 374736 159802 374788 159808
rect 374932 155378 374960 372574
rect 375024 256018 375052 427790
rect 375104 411324 375156 411330
rect 375104 411266 375156 411272
rect 375012 256012 375064 256018
rect 375012 255954 375064 255960
rect 375012 245676 375064 245682
rect 375012 245618 375064 245624
rect 375024 181694 375052 245618
rect 375116 242894 375144 411266
rect 375196 307896 375248 307902
rect 375196 307838 375248 307844
rect 375104 242888 375156 242894
rect 375104 242830 375156 242836
rect 375012 181688 375064 181694
rect 375012 181630 375064 181636
rect 375208 159526 375236 307838
rect 375288 297424 375340 297430
rect 375288 297366 375340 297372
rect 375300 240009 375328 297366
rect 375286 240000 375342 240009
rect 375286 239935 375342 239944
rect 375392 176526 375420 506466
rect 375472 456816 375524 456822
rect 375472 456758 375524 456764
rect 375380 176520 375432 176526
rect 375380 176462 375432 176468
rect 375196 159520 375248 159526
rect 375196 159462 375248 159468
rect 374920 155372 374972 155378
rect 374920 155314 374972 155320
rect 374644 153196 374696 153202
rect 374644 153138 374696 153144
rect 375484 151434 375512 456758
rect 376036 160886 376064 601666
rect 376116 565276 376168 565282
rect 376116 565218 376168 565224
rect 376024 160880 376076 160886
rect 376024 160822 376076 160828
rect 376128 152590 376156 565218
rect 376206 563816 376262 563825
rect 376206 563751 376262 563760
rect 376220 240553 376248 563751
rect 376852 560856 376904 560862
rect 376852 560798 376904 560804
rect 376760 560788 376812 560794
rect 376760 560730 376812 560736
rect 376300 462460 376352 462466
rect 376300 462402 376352 462408
rect 376206 240544 376262 240553
rect 376206 240479 376262 240488
rect 376312 230450 376340 462402
rect 376576 422340 376628 422346
rect 376576 422282 376628 422288
rect 376484 414044 376536 414050
rect 376484 413986 376536 413992
rect 376392 353320 376444 353326
rect 376392 353262 376444 353268
rect 376300 230444 376352 230450
rect 376300 230386 376352 230392
rect 376404 155514 376432 353262
rect 376496 227390 376524 413986
rect 376588 345030 376616 422282
rect 376576 345024 376628 345030
rect 376576 344966 376628 344972
rect 376576 325712 376628 325718
rect 376576 325654 376628 325660
rect 376484 227384 376536 227390
rect 376484 227326 376536 227332
rect 376588 167890 376616 325654
rect 376668 274712 376720 274718
rect 376668 274654 376720 274660
rect 376680 187338 376708 274654
rect 376668 187332 376720 187338
rect 376668 187274 376720 187280
rect 376576 167884 376628 167890
rect 376576 167826 376628 167832
rect 376392 155508 376444 155514
rect 376392 155450 376444 155456
rect 376772 153134 376800 560730
rect 376864 158273 376892 560798
rect 376944 235340 376996 235346
rect 376944 235282 376996 235288
rect 376850 158264 376906 158273
rect 376850 158199 376906 158208
rect 376956 153338 376984 235282
rect 377416 190369 377444 683606
rect 378140 570648 378192 570654
rect 378140 570590 378192 570596
rect 377496 568676 377548 568682
rect 377496 568618 377548 568624
rect 377402 190360 377458 190369
rect 377402 190295 377458 190304
rect 377034 181520 377090 181529
rect 377034 181455 377090 181464
rect 376944 153332 376996 153338
rect 376944 153274 376996 153280
rect 376760 153128 376812 153134
rect 376760 153070 376812 153076
rect 376116 152584 376168 152590
rect 376116 152526 376168 152532
rect 375472 151428 375524 151434
rect 375472 151370 375524 151376
rect 377048 149954 377076 181455
rect 377508 158273 377536 568618
rect 377588 564732 377640 564738
rect 377588 564674 377640 564680
rect 377494 158264 377550 158273
rect 377494 158199 377550 158208
rect 377600 155825 377628 564674
rect 377680 512032 377732 512038
rect 377680 511974 377732 511980
rect 377692 174962 377720 511974
rect 377772 483064 377824 483070
rect 377772 483006 377824 483012
rect 377680 174956 377732 174962
rect 377680 174898 377732 174904
rect 377784 165034 377812 483006
rect 377864 390652 377916 390658
rect 377864 390594 377916 390600
rect 377772 165028 377824 165034
rect 377772 164970 377824 164976
rect 377586 155816 377642 155825
rect 377586 155751 377642 155760
rect 377220 153332 377272 153338
rect 377220 153274 377272 153280
rect 370964 149932 371016 149938
rect 349712 149874 349764 149880
rect 376878 149926 377076 149954
rect 377232 149954 377260 153274
rect 377876 152658 377904 390594
rect 377956 387864 378008 387870
rect 377956 387806 378008 387812
rect 377968 162382 377996 387806
rect 378152 269074 378180 570590
rect 378232 356176 378284 356182
rect 378232 356118 378284 356124
rect 378140 269068 378192 269074
rect 378140 269010 378192 269016
rect 378140 235272 378192 235278
rect 378140 235214 378192 235220
rect 377956 162376 378008 162382
rect 377956 162318 378008 162324
rect 377864 152652 377916 152658
rect 377864 152594 377916 152600
rect 378152 149954 378180 235214
rect 378244 187678 378272 356118
rect 378692 251864 378744 251870
rect 378692 251806 378744 251812
rect 378704 241330 378732 251806
rect 378692 241324 378744 241330
rect 378692 241266 378744 241272
rect 378692 201544 378744 201550
rect 378692 201486 378744 201492
rect 378704 200870 378732 201486
rect 378692 200864 378744 200870
rect 378692 200806 378744 200812
rect 378232 187672 378284 187678
rect 378232 187614 378284 187620
rect 378796 152862 378824 685918
rect 381544 661088 381596 661094
rect 381544 661030 381596 661036
rect 380164 652792 380216 652798
rect 380164 652734 380216 652740
rect 378968 627972 379020 627978
rect 378968 627914 379020 627920
rect 378876 599004 378928 599010
rect 378876 598946 378928 598952
rect 378888 168026 378916 598946
rect 378980 270502 379008 627914
rect 379060 562692 379112 562698
rect 379060 562634 379112 562640
rect 378968 270496 379020 270502
rect 378968 270438 379020 270444
rect 378968 266416 379020 266422
rect 378968 266358 379020 266364
rect 378876 168020 378928 168026
rect 378876 167962 378928 167968
rect 378980 160886 379008 266358
rect 379072 237289 379100 562634
rect 379520 490000 379572 490006
rect 379520 489942 379572 489948
rect 379152 416832 379204 416838
rect 379152 416774 379204 416780
rect 379058 237280 379114 237289
rect 379058 237215 379114 237224
rect 379164 225758 379192 416774
rect 379244 328500 379296 328506
rect 379244 328442 379296 328448
rect 379152 225752 379204 225758
rect 379152 225694 379204 225700
rect 379256 171902 379284 328442
rect 379336 320204 379388 320210
rect 379336 320146 379388 320152
rect 379348 230382 379376 320146
rect 379428 299600 379480 299606
rect 379428 299542 379480 299548
rect 379336 230376 379388 230382
rect 379336 230318 379388 230324
rect 379440 228410 379468 299542
rect 379532 274718 379560 489942
rect 379612 345092 379664 345098
rect 379612 345034 379664 345040
rect 379520 274712 379572 274718
rect 379520 274654 379572 274660
rect 379428 228404 379480 228410
rect 379428 228346 379480 228352
rect 379624 171970 379652 345034
rect 380176 176361 380204 652734
rect 381556 583098 381584 661030
rect 381544 583092 381596 583098
rect 381544 583034 381596 583040
rect 382924 566228 382976 566234
rect 382924 566170 382976 566176
rect 380716 565888 380768 565894
rect 380716 565830 380768 565836
rect 380346 563544 380402 563553
rect 380346 563479 380402 563488
rect 380256 560992 380308 560998
rect 380256 560934 380308 560940
rect 380162 176352 380218 176361
rect 380162 176287 380218 176296
rect 379612 171964 379664 171970
rect 379612 171906 379664 171912
rect 379244 171896 379296 171902
rect 379244 171838 379296 171844
rect 378968 160880 379020 160886
rect 378968 160822 379020 160828
rect 380268 153134 380296 560934
rect 380360 160818 380388 563479
rect 380532 558952 380584 558958
rect 380532 558894 380584 558900
rect 380440 529984 380492 529990
rect 380440 529926 380492 529932
rect 380348 160812 380400 160818
rect 380348 160754 380400 160760
rect 380256 153128 380308 153134
rect 380256 153070 380308 153076
rect 378784 152856 378836 152862
rect 378784 152798 378836 152804
rect 380452 151026 380480 529926
rect 380544 277370 380572 558894
rect 380624 454096 380676 454102
rect 380624 454038 380676 454044
rect 380532 277364 380584 277370
rect 380532 277306 380584 277312
rect 380532 260908 380584 260914
rect 380532 260850 380584 260856
rect 380544 181626 380572 260850
rect 380636 214606 380664 454038
rect 380728 416770 380756 565830
rect 381728 564596 381780 564602
rect 381728 564538 381780 564544
rect 381544 563440 381596 563446
rect 381544 563382 381596 563388
rect 380716 416764 380768 416770
rect 380716 416706 380768 416712
rect 380900 380996 380952 381002
rect 380900 380938 380952 380944
rect 380716 371272 380768 371278
rect 380716 371214 380768 371220
rect 380728 230314 380756 371214
rect 380808 287088 380860 287094
rect 380808 287030 380860 287036
rect 380716 230308 380768 230314
rect 380716 230250 380768 230256
rect 380624 214600 380676 214606
rect 380624 214542 380676 214548
rect 380820 199578 380848 287030
rect 380808 199572 380860 199578
rect 380808 199514 380860 199520
rect 380532 181620 380584 181626
rect 380532 181562 380584 181568
rect 380912 174554 380940 380938
rect 381452 277432 381504 277438
rect 381452 277374 381504 277380
rect 381464 238950 381492 277374
rect 381452 238944 381504 238950
rect 381452 238886 381504 238892
rect 380900 174548 380952 174554
rect 380900 174490 380952 174496
rect 380716 156800 380768 156806
rect 380716 156742 380768 156748
rect 380440 151020 380492 151026
rect 380440 150962 380492 150968
rect 377232 149926 377522 149954
rect 378152 149926 378810 149954
rect 380728 149940 380756 156742
rect 381556 152794 381584 563382
rect 381636 517608 381688 517614
rect 381636 517550 381688 517556
rect 381544 152788 381596 152794
rect 381544 152730 381596 152736
rect 381648 152658 381676 517550
rect 381740 241262 381768 564538
rect 381820 560516 381872 560522
rect 381820 560458 381872 560464
rect 381728 241256 381780 241262
rect 381728 241198 381780 241204
rect 381832 237153 381860 560458
rect 381912 490000 381964 490006
rect 381912 489942 381964 489948
rect 381818 237144 381874 237153
rect 381818 237079 381874 237088
rect 381924 176458 381952 489942
rect 382004 418260 382056 418266
rect 382004 418202 382056 418208
rect 381912 176452 381964 176458
rect 381912 176394 381964 176400
rect 382016 156806 382044 418202
rect 382740 396092 382792 396098
rect 382740 396034 382792 396040
rect 382188 394732 382240 394738
rect 382188 394674 382240 394680
rect 382096 302252 382148 302258
rect 382096 302194 382148 302200
rect 382108 158166 382136 302194
rect 382096 158160 382148 158166
rect 382096 158102 382148 158108
rect 382004 156800 382056 156806
rect 382004 156742 382056 156748
rect 382200 155310 382228 394674
rect 382648 318844 382700 318850
rect 382648 318786 382700 318792
rect 382660 213314 382688 318786
rect 382752 239494 382780 396034
rect 382832 343664 382884 343670
rect 382832 343606 382884 343612
rect 382740 239488 382792 239494
rect 382740 239430 382792 239436
rect 382648 213308 382700 213314
rect 382648 213250 382700 213256
rect 382278 183696 382334 183705
rect 382278 183631 382334 183640
rect 382292 183598 382320 183631
rect 382280 183592 382332 183598
rect 382280 183534 382332 183540
rect 382188 155304 382240 155310
rect 382188 155246 382240 155252
rect 382844 154290 382872 343606
rect 382936 245614 382964 566170
rect 383028 522986 383056 690610
rect 385684 682236 385736 682242
rect 385684 682178 385736 682184
rect 383568 654152 383620 654158
rect 383568 654094 383620 654100
rect 383292 579692 383344 579698
rect 383292 579634 383344 579640
rect 383016 522980 383068 522986
rect 383016 522922 383068 522928
rect 383108 505164 383160 505170
rect 383108 505106 383160 505112
rect 383016 478916 383068 478922
rect 383016 478858 383068 478864
rect 382924 245608 382976 245614
rect 382924 245550 382976 245556
rect 382924 242956 382976 242962
rect 382924 242898 382976 242904
rect 382832 154284 382884 154290
rect 382832 154226 382884 154232
rect 382936 154086 382964 242898
rect 383028 174729 383056 478858
rect 383120 229945 383148 505106
rect 383200 463752 383252 463758
rect 383200 463694 383252 463700
rect 383106 229936 383162 229945
rect 383106 229871 383162 229880
rect 383212 195362 383240 463694
rect 383304 320142 383332 579634
rect 383476 448588 383528 448594
rect 383476 448530 383528 448536
rect 383384 420980 383436 420986
rect 383384 420922 383436 420928
rect 383292 320136 383344 320142
rect 383292 320078 383344 320084
rect 383396 225622 383424 420922
rect 383488 232558 383516 448530
rect 383580 232694 383608 654094
rect 384948 644496 385000 644502
rect 384948 644438 385000 644444
rect 384672 574796 384724 574802
rect 384672 574738 384724 574744
rect 384304 546644 384356 546650
rect 384304 546586 384356 546592
rect 384120 298172 384172 298178
rect 384120 298114 384172 298120
rect 383568 232688 383620 232694
rect 383568 232630 383620 232636
rect 383476 232552 383528 232558
rect 383476 232494 383528 232500
rect 383384 225616 383436 225622
rect 383384 225558 383436 225564
rect 384132 220114 384160 298114
rect 384212 284368 384264 284374
rect 384212 284310 384264 284316
rect 384120 220108 384172 220114
rect 384120 220050 384172 220056
rect 384224 197062 384252 284310
rect 384316 213246 384344 546586
rect 384488 496868 384540 496874
rect 384488 496810 384540 496816
rect 384396 492720 384448 492726
rect 384396 492662 384448 492668
rect 384304 213240 384356 213246
rect 384304 213182 384356 213188
rect 384304 204332 384356 204338
rect 384304 204274 384356 204280
rect 384212 197056 384264 197062
rect 384212 196998 384264 197004
rect 383200 195356 383252 195362
rect 383200 195298 383252 195304
rect 384316 188222 384344 204274
rect 384304 188216 384356 188222
rect 384304 188158 384356 188164
rect 384408 174826 384436 492662
rect 384500 191350 384528 496810
rect 384580 488572 384632 488578
rect 384580 488514 384632 488520
rect 384488 191344 384540 191350
rect 384488 191286 384540 191292
rect 384592 185706 384620 488514
rect 384684 275942 384712 574738
rect 384764 499588 384816 499594
rect 384764 499530 384816 499536
rect 384672 275936 384724 275942
rect 384672 275878 384724 275884
rect 384672 256012 384724 256018
rect 384672 255954 384724 255960
rect 384684 237114 384712 255954
rect 384672 237108 384724 237114
rect 384672 237050 384724 237056
rect 384776 227186 384804 499530
rect 384856 350600 384908 350606
rect 384856 350542 384908 350548
rect 384764 227180 384816 227186
rect 384764 227122 384816 227128
rect 384580 185700 384632 185706
rect 384580 185642 384632 185648
rect 384868 182986 384896 350542
rect 384960 232665 384988 644438
rect 385592 380928 385644 380934
rect 385592 380870 385644 380876
rect 385500 245608 385552 245614
rect 385500 245550 385552 245556
rect 385040 235408 385092 235414
rect 385040 235350 385092 235356
rect 384946 232656 385002 232665
rect 384946 232591 385002 232600
rect 384856 182980 384908 182986
rect 384856 182922 384908 182928
rect 384396 174820 384448 174826
rect 384396 174762 384448 174768
rect 383014 174720 383070 174729
rect 383014 174655 383070 174664
rect 385052 171134 385080 235350
rect 385052 171106 385448 171134
rect 383936 164960 383988 164966
rect 383936 164902 383988 164908
rect 382924 154080 382976 154086
rect 382924 154022 382976 154028
rect 383292 153196 383344 153202
rect 383292 153138 383344 153144
rect 381636 152652 381688 152658
rect 381636 152594 381688 152600
rect 383304 149940 383332 153138
rect 383948 149940 383976 164902
rect 384578 156632 384634 156641
rect 384578 156567 384634 156576
rect 384592 149940 384620 156567
rect 385420 149954 385448 171106
rect 385512 158545 385540 245550
rect 385604 237318 385632 380870
rect 385592 237312 385644 237318
rect 385592 237254 385644 237260
rect 385696 166530 385724 682178
rect 387708 681964 387760 681970
rect 387708 681906 387760 681912
rect 387064 633480 387116 633486
rect 387064 633422 387116 633428
rect 386328 587920 386380 587926
rect 386328 587862 386380 587868
rect 385774 563408 385830 563417
rect 385774 563343 385830 563352
rect 385684 166524 385736 166530
rect 385684 166466 385736 166472
rect 385498 158536 385554 158545
rect 385498 158471 385554 158480
rect 385788 152454 385816 563343
rect 385960 546508 386012 546514
rect 385960 546450 386012 546456
rect 385868 523048 385920 523054
rect 385868 522990 385920 522996
rect 385880 176186 385908 522990
rect 385972 230081 386000 546450
rect 386144 532772 386196 532778
rect 386144 532714 386196 532720
rect 386052 495508 386104 495514
rect 386052 495450 386104 495456
rect 386064 456754 386092 495450
rect 386052 456748 386104 456754
rect 386052 456690 386104 456696
rect 386052 451308 386104 451314
rect 386052 451250 386104 451256
rect 385958 230072 386014 230081
rect 385958 230007 386014 230016
rect 385868 176180 385920 176186
rect 385868 176122 385920 176128
rect 386064 159934 386092 451250
rect 386156 230217 386184 532714
rect 386236 438932 386288 438938
rect 386236 438874 386288 438880
rect 386142 230208 386198 230217
rect 386142 230143 386198 230152
rect 386248 176322 386276 438874
rect 386340 236609 386368 587862
rect 386420 536852 386472 536858
rect 386420 536794 386472 536800
rect 386326 236600 386382 236609
rect 386326 236535 386382 236544
rect 386432 177721 386460 536794
rect 386972 258120 387024 258126
rect 386972 258062 387024 258068
rect 386880 238808 386932 238814
rect 386880 238750 386932 238756
rect 386892 229634 386920 238750
rect 386880 229628 386932 229634
rect 386880 229570 386932 229576
rect 386512 200864 386564 200870
rect 386512 200806 386564 200812
rect 386418 177712 386474 177721
rect 386418 177647 386474 177656
rect 386236 176316 386288 176322
rect 386236 176258 386288 176264
rect 386052 159928 386104 159934
rect 386052 159870 386104 159876
rect 385776 152448 385828 152454
rect 385776 152390 385828 152396
rect 386524 149954 386552 200806
rect 386984 163606 387012 258062
rect 387076 173534 387104 633422
rect 387248 565208 387300 565214
rect 387248 565150 387300 565156
rect 387156 516248 387208 516254
rect 387156 516190 387208 516196
rect 387064 173528 387116 173534
rect 387064 173470 387116 173476
rect 387168 167793 387196 516190
rect 387260 238649 387288 565150
rect 387340 562148 387392 562154
rect 387340 562090 387392 562096
rect 387352 256018 387380 562090
rect 387616 552084 387668 552090
rect 387616 552026 387668 552032
rect 387432 483132 387484 483138
rect 387432 483074 387484 483080
rect 387340 256012 387392 256018
rect 387340 255954 387392 255960
rect 387340 253972 387392 253978
rect 387340 253914 387392 253920
rect 387246 238640 387302 238649
rect 387246 238575 387302 238584
rect 387352 187270 387380 253914
rect 387444 196926 387472 483074
rect 387524 281512 387576 281518
rect 387524 281454 387576 281460
rect 387432 196920 387484 196926
rect 387432 196862 387484 196868
rect 387340 187264 387392 187270
rect 387340 187206 387392 187212
rect 387154 167784 387210 167793
rect 387154 167719 387210 167728
rect 386972 163600 387024 163606
rect 386972 163542 387024 163548
rect 387536 162110 387564 281454
rect 387628 232966 387656 552026
rect 387720 239873 387748 681906
rect 388536 661156 388588 661162
rect 388536 661098 388588 661104
rect 387800 566092 387852 566098
rect 387800 566034 387852 566040
rect 387812 281518 387840 566034
rect 388444 565004 388496 565010
rect 388444 564946 388496 564952
rect 388260 517608 388312 517614
rect 388260 517550 388312 517556
rect 387800 281512 387852 281518
rect 387800 281454 387852 281460
rect 388168 278792 388220 278798
rect 388168 278734 388220 278740
rect 387706 239864 387762 239873
rect 387706 239799 387762 239808
rect 388180 234122 388208 278734
rect 388272 235249 388300 517550
rect 388352 300960 388404 300966
rect 388352 300902 388404 300908
rect 388258 235240 388314 235249
rect 388258 235175 388314 235184
rect 388168 234116 388220 234122
rect 388168 234058 388220 234064
rect 387616 232960 387668 232966
rect 387616 232902 387668 232908
rect 388364 198150 388392 300902
rect 388352 198144 388404 198150
rect 388352 198086 388404 198092
rect 388456 162217 388484 564946
rect 388548 276010 388576 661098
rect 388626 562728 388682 562737
rect 388626 562663 388682 562672
rect 388536 276004 388588 276010
rect 388536 275946 388588 275952
rect 388640 162353 388668 562663
rect 389180 559700 389232 559706
rect 389180 559642 389232 559648
rect 388904 467900 388956 467906
rect 388904 467842 388956 467848
rect 388720 397520 388772 397526
rect 388720 397462 388772 397468
rect 388626 162344 388682 162353
rect 388626 162279 388682 162288
rect 388442 162208 388498 162217
rect 388442 162143 388498 162152
rect 387524 162104 387576 162110
rect 387524 162046 387576 162052
rect 388732 156534 388760 397462
rect 388812 351960 388864 351966
rect 388812 351902 388864 351908
rect 388720 156528 388772 156534
rect 388720 156470 388772 156476
rect 388824 154358 388852 351902
rect 388916 238105 388944 467842
rect 388996 414044 389048 414050
rect 388996 413986 389048 413992
rect 388902 238096 388958 238105
rect 388902 238031 388958 238040
rect 388812 154352 388864 154358
rect 388812 154294 388864 154300
rect 389008 150113 389036 413986
rect 389088 262676 389140 262682
rect 389088 262618 389140 262624
rect 389100 237046 389128 262618
rect 389088 237040 389140 237046
rect 389088 236982 389140 236988
rect 389088 188216 389140 188222
rect 389088 188158 389140 188164
rect 388994 150104 389050 150113
rect 388994 150039 389050 150048
rect 385420 149926 385894 149954
rect 386524 149926 387182 149954
rect 389100 149940 389128 188158
rect 389192 171134 389220 559642
rect 389824 543788 389876 543794
rect 389824 543730 389876 543736
rect 389732 244384 389784 244390
rect 389732 244326 389784 244332
rect 389744 176050 389772 244326
rect 389732 176044 389784 176050
rect 389732 175986 389784 175992
rect 389836 174865 389864 543730
rect 389928 513330 389956 697546
rect 396816 684684 396868 684690
rect 396816 684626 396868 684632
rect 393964 684140 394016 684146
rect 393964 684082 394016 684088
rect 393228 683800 393280 683806
rect 393228 683742 393280 683748
rect 393136 643136 393188 643142
rect 393136 643078 393188 643084
rect 390468 641844 390520 641850
rect 390468 641786 390520 641792
rect 390376 630692 390428 630698
rect 390376 630634 390428 630640
rect 390008 563576 390060 563582
rect 390008 563518 390060 563524
rect 389916 513324 389968 513330
rect 389916 513266 389968 513272
rect 389916 509312 389968 509318
rect 389916 509254 389968 509260
rect 389928 178770 389956 509254
rect 390020 238678 390048 563518
rect 390100 393372 390152 393378
rect 390100 393314 390152 393320
rect 390112 315994 390140 393314
rect 390100 315988 390152 315994
rect 390100 315930 390152 315936
rect 390284 311908 390336 311914
rect 390284 311850 390336 311856
rect 390100 307828 390152 307834
rect 390100 307770 390152 307776
rect 390008 238672 390060 238678
rect 390008 238614 390060 238620
rect 389916 178764 389968 178770
rect 389916 178706 389968 178712
rect 389822 174856 389878 174865
rect 389822 174791 389878 174800
rect 389192 171106 390048 171134
rect 390020 149954 390048 171106
rect 390112 151570 390140 307770
rect 390192 285796 390244 285802
rect 390192 285738 390244 285744
rect 390204 196450 390232 285738
rect 390296 227322 390324 311850
rect 390388 233238 390416 630634
rect 390376 233232 390428 233238
rect 390376 233174 390428 233180
rect 390480 232937 390508 641786
rect 391848 636268 391900 636274
rect 391848 636210 391900 636216
rect 391388 564868 391440 564874
rect 391388 564810 391440 564816
rect 391204 562080 391256 562086
rect 391204 562022 391256 562028
rect 391112 256012 391164 256018
rect 391112 255954 391164 255960
rect 391020 255400 391072 255406
rect 391020 255342 391072 255348
rect 390466 232928 390522 232937
rect 390466 232863 390522 232872
rect 390284 227316 390336 227322
rect 390284 227258 390336 227264
rect 390192 196444 390244 196450
rect 390192 196386 390244 196392
rect 391032 157146 391060 255342
rect 391124 237386 391152 255954
rect 391112 237380 391164 237386
rect 391112 237322 391164 237328
rect 391020 157140 391072 157146
rect 391020 157082 391072 157088
rect 391216 154358 391244 562022
rect 391296 534132 391348 534138
rect 391296 534074 391348 534080
rect 391308 161022 391336 534074
rect 391400 237862 391428 564810
rect 391480 456816 391532 456822
rect 391480 456758 391532 456764
rect 391388 237856 391440 237862
rect 391388 237798 391440 237804
rect 391492 178906 391520 456758
rect 391756 389224 391808 389230
rect 391756 389166 391808 389172
rect 391664 338156 391716 338162
rect 391664 338098 391716 338104
rect 391572 304292 391624 304298
rect 391572 304234 391624 304240
rect 391584 240106 391612 304234
rect 391572 240100 391624 240106
rect 391572 240042 391624 240048
rect 391480 178900 391532 178906
rect 391480 178842 391532 178848
rect 391676 164966 391704 338098
rect 391664 164960 391716 164966
rect 391664 164902 391716 164908
rect 391296 161016 391348 161022
rect 391296 160958 391348 160964
rect 391768 158234 391796 389166
rect 391756 158228 391808 158234
rect 391756 158170 391808 158176
rect 391204 154352 391256 154358
rect 391204 154294 391256 154300
rect 391664 152788 391716 152794
rect 391664 152730 391716 152736
rect 390100 151564 390152 151570
rect 390100 151506 390152 151512
rect 390020 149926 390402 149954
rect 391676 149940 391704 152730
rect 391860 151473 391888 636210
rect 392860 612808 392912 612814
rect 392860 612750 392912 612756
rect 392768 489932 392820 489938
rect 392768 489874 392820 489880
rect 392584 466472 392636 466478
rect 392584 466414 392636 466420
rect 392400 346452 392452 346458
rect 392400 346394 392452 346400
rect 392412 262682 392440 346394
rect 392492 310548 392544 310554
rect 392492 310490 392544 310496
rect 392400 262676 392452 262682
rect 392400 262618 392452 262624
rect 392400 244316 392452 244322
rect 392400 244258 392452 244264
rect 392412 162450 392440 244258
rect 392504 178838 392532 310490
rect 392492 178832 392544 178838
rect 392492 178774 392544 178780
rect 392596 162790 392624 466414
rect 392676 462460 392728 462466
rect 392676 462402 392728 462408
rect 392688 188970 392716 462402
rect 392780 238406 392808 489874
rect 392872 394670 392900 612750
rect 393044 488640 393096 488646
rect 393044 488582 393096 488588
rect 392952 397520 393004 397526
rect 392952 397462 393004 397468
rect 392860 394664 392912 394670
rect 392860 394606 392912 394612
rect 392860 378208 392912 378214
rect 392860 378150 392912 378156
rect 392768 238400 392820 238406
rect 392768 238342 392820 238348
rect 392676 188964 392728 188970
rect 392676 188906 392728 188912
rect 392872 186862 392900 378150
rect 392860 186856 392912 186862
rect 392860 186798 392912 186804
rect 392964 181558 392992 397462
rect 393056 284986 393084 488582
rect 393044 284980 393096 284986
rect 393044 284922 393096 284928
rect 393044 282940 393096 282946
rect 393044 282882 393096 282888
rect 393056 184618 393084 282882
rect 393148 242321 393176 643078
rect 393134 242312 393190 242321
rect 393134 242247 393190 242256
rect 393240 238241 393268 683742
rect 393872 422340 393924 422346
rect 393872 422282 393924 422288
rect 393780 273284 393832 273290
rect 393780 273226 393832 273232
rect 393226 238232 393282 238241
rect 393226 238167 393282 238176
rect 393792 235686 393820 273226
rect 393780 235680 393832 235686
rect 393780 235622 393832 235628
rect 393884 234258 393912 422282
rect 393872 234252 393924 234258
rect 393872 234194 393924 234200
rect 393044 184612 393096 184618
rect 393044 184554 393096 184560
rect 392952 181552 393004 181558
rect 392952 181494 393004 181500
rect 392584 162784 392636 162790
rect 392584 162726 392636 162732
rect 392400 162444 392452 162450
rect 392400 162386 392452 162392
rect 393976 152726 394004 684082
rect 396724 679380 396776 679386
rect 396724 679322 396776 679328
rect 395528 679176 395580 679182
rect 395528 679118 395580 679124
rect 394608 651432 394660 651438
rect 394608 651374 394660 651380
rect 394056 560652 394108 560658
rect 394056 560594 394108 560600
rect 394068 153066 394096 560594
rect 394516 556232 394568 556238
rect 394516 556174 394568 556180
rect 394148 513392 394200 513398
rect 394148 513334 394200 513340
rect 394160 310486 394188 513334
rect 394332 485852 394384 485858
rect 394332 485794 394384 485800
rect 394240 462392 394292 462398
rect 394240 462334 394292 462340
rect 394148 310480 394200 310486
rect 394148 310422 394200 310428
rect 394148 284980 394200 284986
rect 394148 284922 394200 284928
rect 394160 262954 394188 284922
rect 394148 262948 394200 262954
rect 394148 262890 394200 262896
rect 394148 261588 394200 261594
rect 394148 261530 394200 261536
rect 394160 178673 394188 261530
rect 394252 234190 394280 462334
rect 394240 234184 394292 234190
rect 394240 234126 394292 234132
rect 394344 232762 394372 485794
rect 394424 473476 394476 473482
rect 394424 473418 394476 473424
rect 394332 232756 394384 232762
rect 394332 232698 394384 232704
rect 394146 178664 394202 178673
rect 394146 178599 394202 178608
rect 394436 155446 394464 473418
rect 394528 237250 394556 556174
rect 394516 237244 394568 237250
rect 394516 237186 394568 237192
rect 394620 232830 394648 651374
rect 395436 563508 395488 563514
rect 395436 563450 395488 563456
rect 395344 561060 395396 561066
rect 395344 561002 395396 561008
rect 395160 262948 395212 262954
rect 395160 262890 395212 262896
rect 395172 237182 395200 262890
rect 395252 245744 395304 245750
rect 395252 245686 395304 245692
rect 395160 237176 395212 237182
rect 395160 237118 395212 237124
rect 394608 232824 394660 232830
rect 394608 232766 394660 232772
rect 395264 177546 395292 245686
rect 395252 177540 395304 177546
rect 395252 177482 395304 177488
rect 394424 155440 394476 155446
rect 394424 155382 394476 155388
rect 394056 153060 394108 153066
rect 394056 153002 394108 153008
rect 395356 152998 395384 561002
rect 395448 238542 395476 563450
rect 395540 390522 395568 679118
rect 396736 587450 396764 679322
rect 396724 587444 396776 587450
rect 396724 587386 396776 587392
rect 395620 563168 395672 563174
rect 395620 563110 395672 563116
rect 395632 447098 395660 563110
rect 396724 560720 396776 560726
rect 396724 560662 396776 560668
rect 395896 560448 395948 560454
rect 395896 560390 395948 560396
rect 395712 532772 395764 532778
rect 395712 532714 395764 532720
rect 395620 447092 395672 447098
rect 395620 447034 395672 447040
rect 395620 440292 395672 440298
rect 395620 440234 395672 440240
rect 395528 390516 395580 390522
rect 395528 390458 395580 390464
rect 395528 380928 395580 380934
rect 395528 380870 395580 380876
rect 395540 240038 395568 380870
rect 395528 240032 395580 240038
rect 395528 239974 395580 239980
rect 395436 238536 395488 238542
rect 395436 238478 395488 238484
rect 395632 154222 395660 440234
rect 395724 261594 395752 532714
rect 395804 462528 395856 462534
rect 395804 462470 395856 462476
rect 395712 261588 395764 261594
rect 395712 261530 395764 261536
rect 395712 259480 395764 259486
rect 395712 259422 395764 259428
rect 395724 190466 395752 259422
rect 395816 236774 395844 462470
rect 395908 441590 395936 560390
rect 395988 524476 396040 524482
rect 395988 524418 396040 524424
rect 395896 441584 395948 441590
rect 395896 441526 395948 441532
rect 395896 411324 395948 411330
rect 395896 411266 395948 411272
rect 395908 243574 395936 411266
rect 395896 243568 395948 243574
rect 395896 243510 395948 243516
rect 395804 236768 395856 236774
rect 395804 236710 395856 236716
rect 396000 235482 396028 524418
rect 396632 427916 396684 427922
rect 396632 427858 396684 427864
rect 396540 307080 396592 307086
rect 396540 307022 396592 307028
rect 396080 240032 396132 240038
rect 396080 239974 396132 239980
rect 395988 235476 396040 235482
rect 395988 235418 396040 235424
rect 395712 190460 395764 190466
rect 395712 190402 395764 190408
rect 396092 189854 396120 239974
rect 396552 235958 396580 307022
rect 396540 235952 396592 235958
rect 396540 235894 396592 235900
rect 396644 234025 396672 427858
rect 396630 234016 396686 234025
rect 396630 233951 396686 233960
rect 396080 189848 396132 189854
rect 396080 189790 396132 189796
rect 396170 177440 396226 177449
rect 396170 177375 396226 177384
rect 395620 154216 395672 154222
rect 395620 154158 395672 154164
rect 395344 152992 395396 152998
rect 395344 152934 395396 152940
rect 393964 152720 394016 152726
rect 393964 152662 394016 152668
rect 391846 151464 391902 151473
rect 391846 151399 391902 151408
rect 394240 151428 394292 151434
rect 394240 151370 394292 151376
rect 394252 149940 394280 151370
rect 396184 149940 396212 177375
rect 396736 153202 396764 560662
rect 396828 356046 396856 684626
rect 397472 663746 397500 703520
rect 398196 700664 398248 700670
rect 398196 700606 398248 700612
rect 402888 700664 402940 700670
rect 402888 700606 402940 700612
rect 398104 682100 398156 682106
rect 398104 682042 398156 682048
rect 397460 663740 397512 663746
rect 397460 663682 397512 663688
rect 397368 516248 397420 516254
rect 397368 516190 397420 516196
rect 397276 465112 397328 465118
rect 397276 465054 397328 465060
rect 396908 459604 396960 459610
rect 396908 459546 396960 459552
rect 396816 356040 396868 356046
rect 396816 355982 396868 355988
rect 396816 305040 396868 305046
rect 396816 304982 396868 304988
rect 396828 232626 396856 304982
rect 396920 239902 396948 459546
rect 397184 436144 397236 436150
rect 397184 436086 397236 436092
rect 397000 430636 397052 430642
rect 397000 430578 397052 430584
rect 396908 239896 396960 239902
rect 396908 239838 396960 239844
rect 396816 232620 396868 232626
rect 396816 232562 396868 232568
rect 397012 229702 397040 430578
rect 397092 372632 397144 372638
rect 397092 372574 397144 372580
rect 397000 229696 397052 229702
rect 397000 229638 397052 229644
rect 397104 174593 397132 372574
rect 397196 233889 397224 436086
rect 397182 233880 397238 233889
rect 397182 233815 397238 233824
rect 397288 229770 397316 465054
rect 397380 239970 397408 516190
rect 398012 342304 398064 342310
rect 398012 342246 398064 342252
rect 397920 255332 397972 255338
rect 397920 255274 397972 255280
rect 397368 239964 397420 239970
rect 397368 239906 397420 239912
rect 397276 229764 397328 229770
rect 397276 229706 397328 229712
rect 397090 174584 397146 174593
rect 397090 174519 397146 174528
rect 397932 169114 397960 255274
rect 398024 234054 398052 342246
rect 398012 234048 398064 234054
rect 398012 233990 398064 233996
rect 398116 169318 398144 682042
rect 398208 238814 398236 700606
rect 399484 700596 399536 700602
rect 399484 700538 399536 700544
rect 399392 698964 399444 698970
rect 399392 698906 399444 698912
rect 398748 684820 398800 684826
rect 398748 684762 398800 684768
rect 398656 596216 398708 596222
rect 398656 596158 398708 596164
rect 398564 592068 398616 592074
rect 398564 592010 398616 592016
rect 398286 564632 398342 564641
rect 398286 564567 398342 564576
rect 398196 238808 398248 238814
rect 398196 238750 398248 238756
rect 398104 169312 398156 169318
rect 398104 169254 398156 169260
rect 397920 169108 397972 169114
rect 397920 169050 397972 169056
rect 396724 153196 396776 153202
rect 396724 153138 396776 153144
rect 398300 152969 398328 564567
rect 398380 542428 398432 542434
rect 398380 542370 398432 542376
rect 398392 236842 398420 542370
rect 398472 437504 398524 437510
rect 398472 437446 398524 437452
rect 398380 236836 398432 236842
rect 398380 236778 398432 236784
rect 398484 221474 398512 437446
rect 398472 221468 398524 221474
rect 398472 221410 398524 221416
rect 398576 162722 398604 592010
rect 398564 162716 398616 162722
rect 398564 162658 398616 162664
rect 398286 152960 398342 152969
rect 398286 152895 398342 152904
rect 398668 151774 398696 596158
rect 398760 238474 398788 684762
rect 399404 655518 399432 698906
rect 399392 655512 399444 655518
rect 399392 655454 399444 655460
rect 398840 352028 398892 352034
rect 398840 351970 398892 351976
rect 398748 238468 398800 238474
rect 398748 238410 398800 238416
rect 398656 151768 398708 151774
rect 398656 151710 398708 151716
rect 398852 149954 398880 351970
rect 399392 256828 399444 256834
rect 399392 256770 399444 256776
rect 399404 206990 399432 256770
rect 399496 238785 399524 700538
rect 399760 687268 399812 687274
rect 399760 687210 399812 687216
rect 399576 680604 399628 680610
rect 399576 680546 399628 680552
rect 399588 506462 399616 680546
rect 399668 680400 399720 680406
rect 399668 680342 399720 680348
rect 399576 506456 399628 506462
rect 399576 506398 399628 506404
rect 399576 474768 399628 474774
rect 399576 474710 399628 474716
rect 399482 238776 399538 238785
rect 399482 238711 399538 238720
rect 399392 206984 399444 206990
rect 399392 206926 399444 206932
rect 399588 194206 399616 474710
rect 399680 445738 399708 680342
rect 399772 587382 399800 687210
rect 402428 685092 402480 685098
rect 402428 685034 402480 685040
rect 399852 684004 399904 684010
rect 399852 683946 399904 683952
rect 399864 587654 399892 683946
rect 401508 683936 401560 683942
rect 401508 683878 401560 683884
rect 400036 681352 400088 681358
rect 400036 681294 400088 681300
rect 399944 679312 399996 679318
rect 399944 679254 399996 679260
rect 399852 587648 399904 587654
rect 399852 587590 399904 587596
rect 399760 587376 399812 587382
rect 399760 587318 399812 587324
rect 399956 587314 399984 679254
rect 399944 587308 399996 587314
rect 399944 587250 399996 587256
rect 399668 445732 399720 445738
rect 399668 445674 399720 445680
rect 399668 426488 399720 426494
rect 399668 426430 399720 426436
rect 399680 238610 399708 426430
rect 399944 408536 399996 408542
rect 399944 408478 399996 408484
rect 399852 323060 399904 323066
rect 399852 323002 399904 323008
rect 399760 295384 399812 295390
rect 399760 295326 399812 295332
rect 399668 238604 399720 238610
rect 399668 238546 399720 238552
rect 399772 229906 399800 295326
rect 399864 232898 399892 323002
rect 399852 232892 399904 232898
rect 399852 232834 399904 232840
rect 399760 229900 399812 229906
rect 399760 229842 399812 229848
rect 399576 194200 399628 194206
rect 399576 194142 399628 194148
rect 399956 150113 399984 408478
rect 400048 405686 400076 681294
rect 400128 680536 400180 680542
rect 400128 680478 400180 680484
rect 400140 590034 400168 680478
rect 400864 676864 400916 676870
rect 400864 676806 400916 676812
rect 400876 651370 400904 676806
rect 400864 651364 400916 651370
rect 400864 651306 400916 651312
rect 401416 594856 401468 594862
rect 401416 594798 401468 594804
rect 400128 590028 400180 590034
rect 400128 589970 400180 589976
rect 400864 564664 400916 564670
rect 400864 564606 400916 564612
rect 400128 525836 400180 525842
rect 400128 525778 400180 525784
rect 400036 405680 400088 405686
rect 400036 405622 400088 405628
rect 400036 394800 400088 394806
rect 400036 394742 400088 394748
rect 400048 233034 400076 394742
rect 400140 245614 400168 525778
rect 400772 329860 400824 329866
rect 400772 329802 400824 329808
rect 400784 285666 400812 329802
rect 400772 285660 400824 285666
rect 400772 285602 400824 285608
rect 400772 278860 400824 278866
rect 400772 278802 400824 278808
rect 400680 249824 400732 249830
rect 400680 249766 400732 249772
rect 400128 245608 400180 245614
rect 400128 245550 400180 245556
rect 400036 233028 400088 233034
rect 400036 232970 400088 232976
rect 400220 224392 400272 224398
rect 400220 224334 400272 224340
rect 400232 151814 400260 224334
rect 400692 222970 400720 249766
rect 400784 234326 400812 278802
rect 400772 234320 400824 234326
rect 400772 234262 400824 234268
rect 400680 222964 400732 222970
rect 400680 222906 400732 222912
rect 400772 170604 400824 170610
rect 400772 170546 400824 170552
rect 400784 151814 400812 170546
rect 400876 152386 400904 564606
rect 401324 531344 401376 531350
rect 401324 531286 401376 531292
rect 401140 495508 401192 495514
rect 401140 495450 401192 495456
rect 400956 451308 401008 451314
rect 400956 451250 401008 451256
rect 400968 387802 400996 451250
rect 400956 387796 401008 387802
rect 400956 387738 401008 387744
rect 400956 382288 401008 382294
rect 400956 382230 401008 382236
rect 400968 240038 400996 382230
rect 401152 288386 401180 495450
rect 401232 487212 401284 487218
rect 401232 487154 401284 487160
rect 401140 288380 401192 288386
rect 401140 288322 401192 288328
rect 401140 287156 401192 287162
rect 401140 287098 401192 287104
rect 401048 285728 401100 285734
rect 401048 285670 401100 285676
rect 400956 240032 401008 240038
rect 400956 239974 401008 239980
rect 401060 238270 401088 285670
rect 401048 238264 401100 238270
rect 401048 238206 401100 238212
rect 401152 234394 401180 287098
rect 401140 234388 401192 234394
rect 401140 234330 401192 234336
rect 401244 155514 401272 487154
rect 401232 155508 401284 155514
rect 401232 155450 401284 155456
rect 401336 154562 401364 531286
rect 401428 155786 401456 594798
rect 401520 233170 401548 683878
rect 402336 682508 402388 682514
rect 402336 682450 402388 682456
rect 402244 682440 402296 682446
rect 402244 682382 402296 682388
rect 402152 288516 402204 288522
rect 402152 288458 402204 288464
rect 401968 267776 402020 267782
rect 401968 267718 402020 267724
rect 401980 240786 402008 267718
rect 402060 256012 402112 256018
rect 402060 255954 402112 255960
rect 401968 240780 402020 240786
rect 401968 240722 402020 240728
rect 402072 236910 402100 255954
rect 402164 253230 402192 288458
rect 402152 253224 402204 253230
rect 402152 253166 402204 253172
rect 402152 248464 402204 248470
rect 402152 248406 402204 248412
rect 402164 239834 402192 248406
rect 402152 239828 402204 239834
rect 402152 239770 402204 239776
rect 402060 236904 402112 236910
rect 402060 236846 402112 236852
rect 401508 233164 401560 233170
rect 401508 233106 401560 233112
rect 401968 177472 402020 177478
rect 401968 177414 402020 177420
rect 401416 155780 401468 155786
rect 401416 155722 401468 155728
rect 401324 154556 401376 154562
rect 401324 154498 401376 154504
rect 400864 152380 400916 152386
rect 400864 152322 400916 152328
rect 400232 151786 400352 151814
rect 400784 151786 400904 151814
rect 399942 150104 399998 150113
rect 399942 150039 399998 150048
rect 400324 149954 400352 151786
rect 400876 149954 400904 151786
rect 398852 149926 400062 149954
rect 400324 149926 400706 149954
rect 400876 149926 401350 149954
rect 401980 149940 402008 177414
rect 402256 165238 402284 682382
rect 402348 166462 402376 682450
rect 402440 590345 402468 685034
rect 402520 648712 402572 648718
rect 402520 648654 402572 648660
rect 402426 590336 402482 590345
rect 402426 590271 402482 590280
rect 402532 587178 402560 648654
rect 402612 622464 402664 622470
rect 402612 622406 402664 622412
rect 402624 587353 402652 622406
rect 402610 587344 402666 587353
rect 402610 587279 402666 587288
rect 402520 587172 402572 587178
rect 402520 587114 402572 587120
rect 402426 560008 402482 560017
rect 402426 559943 402482 559952
rect 402440 500954 402468 559943
rect 402704 521688 402756 521694
rect 402704 521630 402756 521636
rect 402428 500948 402480 500954
rect 402428 500890 402480 500896
rect 402612 429276 402664 429282
rect 402612 429218 402664 429224
rect 402428 392012 402480 392018
rect 402428 391954 402480 391960
rect 402440 215966 402468 391954
rect 402520 382288 402572 382294
rect 402520 382230 402572 382236
rect 402532 257378 402560 382230
rect 402520 257372 402572 257378
rect 402520 257314 402572 257320
rect 402520 251252 402572 251258
rect 402520 251194 402572 251200
rect 402428 215960 402480 215966
rect 402428 215902 402480 215908
rect 402336 166456 402388 166462
rect 402336 166398 402388 166404
rect 402244 165232 402296 165238
rect 402244 165174 402296 165180
rect 402532 158370 402560 251194
rect 402624 207738 402652 429218
rect 402716 292466 402744 521630
rect 402796 481704 402848 481710
rect 402796 481646 402848 481652
rect 402704 292460 402756 292466
rect 402704 292402 402756 292408
rect 402704 288380 402756 288386
rect 402704 288322 402756 288328
rect 402612 207732 402664 207738
rect 402612 207674 402664 207680
rect 402716 165238 402744 288322
rect 402808 234297 402836 481646
rect 402900 251190 402928 700606
rect 405004 700596 405056 700602
rect 405004 700538 405056 700544
rect 403808 683324 403860 683330
rect 403808 683266 403860 683272
rect 403716 682372 403768 682378
rect 403716 682314 403768 682320
rect 403440 644632 403492 644638
rect 403440 644574 403492 644580
rect 403348 474836 403400 474842
rect 403348 474778 403400 474784
rect 403164 383988 403216 383994
rect 403164 383930 403216 383936
rect 402888 251184 402940 251190
rect 402888 251126 402940 251132
rect 402794 234288 402850 234297
rect 402794 234223 402850 234232
rect 402704 165232 402756 165238
rect 402704 165174 402756 165180
rect 402520 158364 402572 158370
rect 402520 158306 402572 158312
rect 403176 149938 403204 383930
rect 403360 162858 403388 474778
rect 403452 232490 403480 644574
rect 403624 562012 403676 562018
rect 403624 561954 403676 561960
rect 403532 447160 403584 447166
rect 403532 447102 403584 447108
rect 403544 290494 403572 447102
rect 403532 290488 403584 290494
rect 403532 290430 403584 290436
rect 403532 288448 403584 288454
rect 403532 288390 403584 288396
rect 403544 238746 403572 288390
rect 403532 238740 403584 238746
rect 403532 238682 403584 238688
rect 403636 238202 403664 561954
rect 403728 437442 403756 682314
rect 403820 466410 403848 683266
rect 404084 683188 404136 683194
rect 404084 683130 404136 683136
rect 403992 681896 404044 681902
rect 403992 681838 404044 681844
rect 403808 466404 403860 466410
rect 403808 466346 403860 466352
rect 403900 458244 403952 458250
rect 403900 458186 403952 458192
rect 403716 437436 403768 437442
rect 403716 437378 403768 437384
rect 403716 375420 403768 375426
rect 403716 375362 403768 375368
rect 403624 238196 403676 238202
rect 403624 238138 403676 238144
rect 403440 232484 403492 232490
rect 403440 232426 403492 232432
rect 403348 162852 403400 162858
rect 403348 162794 403400 162800
rect 403728 162586 403756 375362
rect 403808 310616 403860 310622
rect 403808 310558 403860 310564
rect 403716 162580 403768 162586
rect 403716 162522 403768 162528
rect 403820 152522 403848 310558
rect 403912 227118 403940 458186
rect 404004 400178 404032 681838
rect 404096 469198 404124 683130
rect 404912 666596 404964 666602
rect 404912 666538 404964 666544
rect 404728 625388 404780 625394
rect 404728 625330 404780 625336
rect 404636 564460 404688 564466
rect 404636 564402 404688 564408
rect 404176 550656 404228 550662
rect 404176 550598 404228 550604
rect 404084 469192 404136 469198
rect 404084 469134 404136 469140
rect 403992 400172 404044 400178
rect 403992 400114 404044 400120
rect 403900 227112 403952 227118
rect 403900 227054 403952 227060
rect 404188 165209 404216 550598
rect 404268 247104 404320 247110
rect 404268 247046 404320 247052
rect 404280 235890 404308 247046
rect 404648 236638 404676 564402
rect 404636 236632 404688 236638
rect 404636 236574 404688 236580
rect 404268 235884 404320 235890
rect 404268 235826 404320 235832
rect 404740 224398 404768 625330
rect 404924 589937 404952 666538
rect 404910 589928 404966 589937
rect 404910 589863 404966 589872
rect 405016 573374 405044 700538
rect 413664 697610 413692 703520
rect 429856 698970 429884 703520
rect 429844 698964 429896 698970
rect 429844 698906 429896 698912
rect 413652 697604 413704 697610
rect 413652 697546 413704 697552
rect 462332 687954 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 687948 462372 687954
rect 462320 687890 462372 687896
rect 405096 687336 405148 687342
rect 405096 687278 405148 687284
rect 457352 687336 457404 687342
rect 457352 687278 457404 687284
rect 405108 589966 405136 687278
rect 407764 686044 407816 686050
rect 407764 685986 407816 685992
rect 405188 685908 405240 685914
rect 405188 685850 405240 685856
rect 405200 590209 405228 685850
rect 405372 683732 405424 683738
rect 405372 683674 405424 683680
rect 405280 679448 405332 679454
rect 405280 679390 405332 679396
rect 405186 590200 405242 590209
rect 405186 590135 405242 590144
rect 405096 589960 405148 589966
rect 405096 589902 405148 589908
rect 405292 587518 405320 679390
rect 405384 590073 405412 683674
rect 406476 683528 406528 683534
rect 406476 683470 406528 683476
rect 406384 680672 406436 680678
rect 406384 680614 406436 680620
rect 405648 637628 405700 637634
rect 405648 637570 405700 637576
rect 405370 590064 405426 590073
rect 405370 589999 405426 590008
rect 405280 587512 405332 587518
rect 405280 587454 405332 587460
rect 405004 573368 405056 573374
rect 405004 573310 405056 573316
rect 405372 572756 405424 572762
rect 405372 572698 405424 572704
rect 405004 565412 405056 565418
rect 405004 565354 405056 565360
rect 405016 438870 405044 565354
rect 405188 564528 405240 564534
rect 405188 564470 405240 564476
rect 405096 560380 405148 560386
rect 405096 560322 405148 560328
rect 405108 516118 405136 560322
rect 405200 549234 405228 564470
rect 405280 561128 405332 561134
rect 405280 561070 405332 561076
rect 405292 557258 405320 561070
rect 405280 557252 405332 557258
rect 405280 557194 405332 557200
rect 405188 549228 405240 549234
rect 405188 549170 405240 549176
rect 405188 543856 405240 543862
rect 405188 543798 405240 543804
rect 405096 516112 405148 516118
rect 405096 516054 405148 516060
rect 405004 438864 405056 438870
rect 405004 438806 405056 438812
rect 405004 400240 405056 400246
rect 405004 400182 405056 400188
rect 404912 288448 404964 288454
rect 404912 288390 404964 288396
rect 404820 261180 404872 261186
rect 404820 261122 404872 261128
rect 404832 247110 404860 261122
rect 404820 247104 404872 247110
rect 404820 247046 404872 247052
rect 404924 244730 404952 288390
rect 405016 247110 405044 400182
rect 405096 320204 405148 320210
rect 405096 320146 405148 320152
rect 405004 247104 405056 247110
rect 405004 247046 405056 247052
rect 405004 245880 405056 245886
rect 405004 245822 405056 245828
rect 404912 244724 404964 244730
rect 404912 244666 404964 244672
rect 404728 224392 404780 224398
rect 404728 224334 404780 224340
rect 404174 165200 404230 165209
rect 404174 165135 404230 165144
rect 405016 154426 405044 245822
rect 405108 159186 405136 320146
rect 405200 255270 405228 543798
rect 405280 454096 405332 454102
rect 405280 454038 405332 454044
rect 405188 255264 405240 255270
rect 405188 255206 405240 255212
rect 405188 245812 405240 245818
rect 405188 245754 405240 245760
rect 405200 160002 405228 245754
rect 405188 159996 405240 160002
rect 405188 159938 405240 159944
rect 405096 159180 405148 159186
rect 405096 159122 405148 159128
rect 405292 154494 405320 454038
rect 405384 271862 405412 572698
rect 405372 271856 405424 271862
rect 405372 271798 405424 271804
rect 405372 266416 405424 266422
rect 405372 266358 405424 266364
rect 405384 241194 405412 266358
rect 405556 248804 405608 248810
rect 405556 248746 405608 248752
rect 405464 244316 405516 244322
rect 405464 244258 405516 244264
rect 405372 241188 405424 241194
rect 405372 241130 405424 241136
rect 405476 236978 405504 244258
rect 405568 238882 405596 248746
rect 405556 238876 405608 238882
rect 405556 238818 405608 238824
rect 405464 236972 405516 236978
rect 405464 236914 405516 236920
rect 405660 231266 405688 637570
rect 406396 509250 406424 680614
rect 406488 590170 406516 683470
rect 406568 683392 406620 683398
rect 406568 683334 406620 683340
rect 406476 590164 406528 590170
rect 406476 590106 406528 590112
rect 406580 590102 406608 683334
rect 407580 681148 407632 681154
rect 407580 681090 407632 681096
rect 406660 680808 406712 680814
rect 406660 680750 406712 680756
rect 406568 590096 406620 590102
rect 406568 590038 406620 590044
rect 406384 509244 406436 509250
rect 406384 509186 406436 509192
rect 406672 461145 406700 680750
rect 406844 680740 406896 680746
rect 406844 680682 406896 680688
rect 406752 679516 406804 679522
rect 406752 679458 406804 679464
rect 406658 461136 406714 461145
rect 406658 461071 406714 461080
rect 406382 438016 406438 438025
rect 406382 437951 406438 437960
rect 406200 314696 406252 314702
rect 406200 314638 406252 314644
rect 406108 295452 406160 295458
rect 406108 295394 406160 295400
rect 406120 242457 406148 295394
rect 406106 242448 406162 242457
rect 406106 242383 406162 242392
rect 406212 233714 406240 314638
rect 406292 247104 406344 247110
rect 406292 247046 406344 247052
rect 406200 233708 406252 233714
rect 406200 233650 406252 233656
rect 405648 231260 405700 231266
rect 405648 231202 405700 231208
rect 406304 163810 406332 247046
rect 406396 245886 406424 437951
rect 406658 433256 406714 433265
rect 406658 433191 406714 433200
rect 406474 383072 406530 383081
rect 406474 383007 406530 383016
rect 406384 245880 406436 245886
rect 406384 245822 406436 245828
rect 406488 245818 406516 383007
rect 406568 257372 406620 257378
rect 406568 257314 406620 257320
rect 406476 245812 406528 245818
rect 406476 245754 406528 245760
rect 406384 244724 406436 244730
rect 406384 244666 406436 244672
rect 406292 163804 406344 163810
rect 406292 163746 406344 163752
rect 406396 161022 406424 244666
rect 406580 165170 406608 257314
rect 406672 217326 406700 433191
rect 406764 377505 406792 679458
rect 406750 377496 406806 377505
rect 406750 377431 406806 377440
rect 406856 372065 406884 680682
rect 406934 679688 406990 679697
rect 406934 679623 406990 679632
rect 406948 587246 406976 679623
rect 407118 678056 407174 678065
rect 407118 677991 407174 678000
rect 407026 677648 407082 677657
rect 407132 677618 407160 677991
rect 407026 677583 407082 677592
rect 407120 677612 407172 677618
rect 406936 587240 406988 587246
rect 406936 587182 406988 587188
rect 407040 485625 407068 677583
rect 407120 677554 407172 677560
rect 407120 670676 407172 670682
rect 407120 670618 407172 670624
rect 407132 670585 407160 670618
rect 407118 670576 407174 670585
rect 407118 670511 407174 670520
rect 407118 669216 407174 669225
rect 407118 669151 407174 669160
rect 407132 667962 407160 669151
rect 407120 667956 407172 667962
rect 407120 667898 407172 667904
rect 407118 667856 407174 667865
rect 407118 667791 407174 667800
rect 407132 666602 407160 667791
rect 407120 666596 407172 666602
rect 407120 666538 407172 666544
rect 407118 666496 407174 666505
rect 407118 666431 407174 666440
rect 407132 665242 407160 666431
rect 407120 665236 407172 665242
rect 407120 665178 407172 665184
rect 407118 663776 407174 663785
rect 407118 663711 407120 663720
rect 407172 663711 407174 663720
rect 407120 663682 407172 663688
rect 407210 662416 407266 662425
rect 407210 662351 407266 662360
rect 407118 661736 407174 661745
rect 407118 661671 407174 661680
rect 407132 661162 407160 661671
rect 407120 661156 407172 661162
rect 407120 661098 407172 661104
rect 407224 661094 407252 662351
rect 407212 661088 407264 661094
rect 407212 661030 407264 661036
rect 407120 655512 407172 655518
rect 407120 655454 407172 655460
rect 407132 654945 407160 655454
rect 407118 654936 407174 654945
rect 407118 654871 407174 654880
rect 407118 654256 407174 654265
rect 407118 654191 407174 654200
rect 407132 654158 407160 654191
rect 407120 654152 407172 654158
rect 407120 654094 407172 654100
rect 407118 652896 407174 652905
rect 407118 652831 407174 652840
rect 407132 652798 407160 652831
rect 407120 652792 407172 652798
rect 407120 652734 407172 652740
rect 407118 652216 407174 652225
rect 407118 652151 407174 652160
rect 407132 651438 407160 652151
rect 407120 651432 407172 651438
rect 407120 651374 407172 651380
rect 407592 651370 407620 681090
rect 407776 678570 407804 685986
rect 409144 685364 409196 685370
rect 409144 685306 409196 685312
rect 409052 685296 409104 685302
rect 409052 685238 409104 685244
rect 408408 685228 408460 685234
rect 408408 685170 408460 685176
rect 407948 685024 408000 685030
rect 407948 684966 408000 684972
rect 407856 683460 407908 683466
rect 407856 683402 407908 683408
rect 407764 678564 407816 678570
rect 407764 678506 407816 678512
rect 407868 678450 407896 683402
rect 407684 678422 407896 678450
rect 407580 651364 407632 651370
rect 407580 651306 407632 651312
rect 407592 650185 407620 651306
rect 407302 650176 407358 650185
rect 407302 650111 407358 650120
rect 407578 650176 407634 650185
rect 407578 650111 407634 650120
rect 407210 649496 407266 649505
rect 407210 649431 407266 649440
rect 407118 648816 407174 648825
rect 407118 648751 407174 648760
rect 407132 648718 407160 648751
rect 407120 648712 407172 648718
rect 407120 648654 407172 648660
rect 407224 648650 407252 649431
rect 407212 648644 407264 648650
rect 407212 648586 407264 648592
rect 407118 644736 407174 644745
rect 407118 644671 407174 644680
rect 407132 644638 407160 644671
rect 407120 644632 407172 644638
rect 407120 644574 407172 644580
rect 407316 644474 407344 650111
rect 407394 645416 407450 645425
rect 407394 645351 407450 645360
rect 407408 644502 407436 645351
rect 407132 644446 407344 644474
rect 407396 644496 407448 644502
rect 407132 526522 407160 644446
rect 407396 644438 407448 644444
rect 407210 644056 407266 644065
rect 407210 643991 407266 644000
rect 407224 643142 407252 643991
rect 407212 643136 407264 643142
rect 407212 643078 407264 643084
rect 407302 642152 407358 642161
rect 407302 642087 407358 642096
rect 407210 642016 407266 642025
rect 407210 641951 407266 641960
rect 407224 641782 407252 641951
rect 407316 641850 407344 642087
rect 407304 641844 407356 641850
rect 407304 641786 407356 641792
rect 407212 641776 407264 641782
rect 407212 641718 407264 641724
rect 407210 641336 407266 641345
rect 407210 641271 407266 641280
rect 407224 640354 407252 641271
rect 407212 640348 407264 640354
rect 407212 640290 407264 640296
rect 407486 638072 407542 638081
rect 407486 638007 407542 638016
rect 407500 637634 407528 638007
rect 407488 637628 407540 637634
rect 407488 637570 407540 637576
rect 407210 637256 407266 637265
rect 407210 637191 407266 637200
rect 407224 636274 407252 637191
rect 407212 636268 407264 636274
rect 407212 636210 407264 636216
rect 407210 633856 407266 633865
rect 407210 633791 407266 633800
rect 407224 633486 407252 633791
rect 407212 633480 407264 633486
rect 407212 633422 407264 633428
rect 407210 632496 407266 632505
rect 407210 632431 407266 632440
rect 407224 632126 407252 632431
rect 407212 632120 407264 632126
rect 407212 632062 407264 632068
rect 407210 631816 407266 631825
rect 407210 631751 407266 631760
rect 407224 630698 407252 631751
rect 407212 630692 407264 630698
rect 407212 630634 407264 630640
rect 407210 629096 407266 629105
rect 407210 629031 407266 629040
rect 407224 627978 407252 629031
rect 407212 627972 407264 627978
rect 407212 627914 407264 627920
rect 407394 625696 407450 625705
rect 407394 625631 407450 625640
rect 407408 625394 407436 625631
rect 407396 625388 407448 625394
rect 407396 625330 407448 625336
rect 407210 622976 407266 622985
rect 407210 622911 407266 622920
rect 407224 622470 407252 622911
rect 407212 622464 407264 622470
rect 407212 622406 407264 622412
rect 407210 618896 407266 618905
rect 407210 618831 407266 618840
rect 407224 618322 407252 618831
rect 407212 618316 407264 618322
rect 407212 618258 407264 618264
rect 407302 616856 407358 616865
rect 407302 616791 407358 616800
rect 407316 615534 407344 616791
rect 407304 615528 407356 615534
rect 407304 615470 407356 615476
rect 407302 614952 407358 614961
rect 407302 614887 407358 614896
rect 407212 612808 407264 612814
rect 407210 612776 407212 612785
rect 407264 612776 407266 612785
rect 407210 612711 407266 612720
rect 407210 608696 407266 608705
rect 407210 608631 407212 608640
rect 407264 608631 407266 608640
rect 407212 608602 407264 608608
rect 407210 607336 407266 607345
rect 407210 607271 407266 607280
rect 407224 607238 407252 607271
rect 407212 607232 407264 607238
rect 407212 607174 407264 607180
rect 407316 605834 407344 614887
rect 407684 614825 407712 678422
rect 407764 678360 407816 678366
rect 407960 678314 407988 684966
rect 408040 684548 408092 684554
rect 408040 684490 408092 684496
rect 407764 678302 407816 678308
rect 407670 614816 407726 614825
rect 407670 614751 407726 614760
rect 407776 605834 407804 678302
rect 407224 605806 407344 605834
rect 407684 605806 407804 605834
rect 407868 678286 407988 678314
rect 407120 526516 407172 526522
rect 407120 526458 407172 526464
rect 407118 525736 407174 525745
rect 407118 525671 407174 525680
rect 407132 524482 407160 525671
rect 407120 524476 407172 524482
rect 407120 524418 407172 524424
rect 407120 522980 407172 522986
rect 407120 522922 407172 522928
rect 407132 522345 407160 522922
rect 407118 522336 407174 522345
rect 407118 522271 407174 522280
rect 407120 517608 407172 517614
rect 407118 517576 407120 517585
rect 407172 517576 407174 517585
rect 407118 517511 407174 517520
rect 407120 516248 407172 516254
rect 407118 516216 407120 516225
rect 407172 516216 407174 516225
rect 407118 516151 407174 516160
rect 407120 513324 407172 513330
rect 407120 513266 407172 513272
rect 407132 512825 407160 513266
rect 407118 512816 407174 512825
rect 407118 512751 407174 512760
rect 407118 512136 407174 512145
rect 407118 512071 407174 512080
rect 407132 512038 407160 512071
rect 407120 512032 407172 512038
rect 407120 511974 407172 511980
rect 407118 509416 407174 509425
rect 407118 509351 407174 509360
rect 407132 509318 407160 509351
rect 407120 509312 407172 509318
rect 407120 509254 407172 509260
rect 407120 500948 407172 500954
rect 407120 500890 407172 500896
rect 407132 500585 407160 500890
rect 407118 500576 407174 500585
rect 407118 500511 407174 500520
rect 407118 497176 407174 497185
rect 407118 497111 407174 497120
rect 407132 496874 407160 497111
rect 407120 496868 407172 496874
rect 407120 496810 407172 496816
rect 407118 495816 407174 495825
rect 407118 495751 407174 495760
rect 407132 495514 407160 495751
rect 407120 495508 407172 495514
rect 407120 495450 407172 495456
rect 407118 493096 407174 493105
rect 407118 493031 407174 493040
rect 407132 492726 407160 493031
rect 407120 492720 407172 492726
rect 407120 492662 407172 492668
rect 407118 491056 407174 491065
rect 407118 490991 407174 491000
rect 407132 490006 407160 490991
rect 407120 490000 407172 490006
rect 407120 489942 407172 489948
rect 407118 489016 407174 489025
rect 407118 488951 407174 488960
rect 407132 488578 407160 488951
rect 407120 488572 407172 488578
rect 407120 488514 407172 488520
rect 407118 487656 407174 487665
rect 407118 487591 407174 487600
rect 407132 487218 407160 487591
rect 407120 487212 407172 487218
rect 407120 487154 407172 487160
rect 407118 486976 407174 486985
rect 407118 486911 407174 486920
rect 407132 485858 407160 486911
rect 407120 485852 407172 485858
rect 407120 485794 407172 485800
rect 407026 485616 407082 485625
rect 407026 485551 407082 485560
rect 407118 484936 407174 484945
rect 407118 484871 407174 484880
rect 407132 484430 407160 484871
rect 407120 484424 407172 484430
rect 407120 484366 407172 484372
rect 407118 484256 407174 484265
rect 407118 484191 407174 484200
rect 407026 483576 407082 483585
rect 407026 483511 407082 483520
rect 406934 478136 406990 478145
rect 406934 478071 406990 478080
rect 406842 372056 406898 372065
rect 406842 371991 406898 372000
rect 406842 356416 406898 356425
rect 406842 356351 406898 356360
rect 406750 345264 406806 345273
rect 406750 345199 406806 345208
rect 406764 254046 406792 345199
rect 406752 254040 406804 254046
rect 406752 253982 406804 253988
rect 406752 245812 406804 245818
rect 406752 245754 406804 245760
rect 406660 217320 406712 217326
rect 406660 217262 406712 217268
rect 406568 165164 406620 165170
rect 406568 165106 406620 165112
rect 406384 161016 406436 161022
rect 406384 160958 406436 160964
rect 406476 158500 406528 158506
rect 406476 158442 406528 158448
rect 405280 154488 405332 154494
rect 405280 154430 405332 154436
rect 405004 154420 405056 154426
rect 405004 154362 405056 154368
rect 403256 152516 403308 152522
rect 403256 152458 403308 152464
rect 403808 152516 403860 152522
rect 403808 152458 403860 152464
rect 403268 149940 403296 152458
rect 406488 149940 406516 158442
rect 406764 150890 406792 245754
rect 406856 162654 406884 356351
rect 406844 162648 406896 162654
rect 406844 162590 406896 162596
rect 406948 152794 406976 478071
rect 407040 152862 407068 483511
rect 407132 483138 407160 484191
rect 407120 483132 407172 483138
rect 407120 483074 407172 483080
rect 407118 482216 407174 482225
rect 407118 482151 407174 482160
rect 407132 481710 407160 482151
rect 407120 481704 407172 481710
rect 407120 481646 407172 481652
rect 407118 480176 407174 480185
rect 407118 480111 407174 480120
rect 407132 478922 407160 480111
rect 407120 478916 407172 478922
rect 407120 478858 407172 478864
rect 407118 475416 407174 475425
rect 407118 475351 407174 475360
rect 407132 474774 407160 475351
rect 407120 474768 407172 474774
rect 407120 474710 407172 474716
rect 407118 474056 407174 474065
rect 407118 473991 407174 474000
rect 407132 473482 407160 473991
rect 407120 473476 407172 473482
rect 407120 473418 407172 473424
rect 407118 469976 407174 469985
rect 407118 469911 407174 469920
rect 407132 469266 407160 469911
rect 407120 469260 407172 469266
rect 407120 469202 407172 469208
rect 407118 468208 407174 468217
rect 407118 468143 407174 468152
rect 407132 467906 407160 468143
rect 407120 467900 407172 467906
rect 407120 467842 407172 467848
rect 407118 465896 407174 465905
rect 407118 465831 407174 465840
rect 407132 465118 407160 465831
rect 407120 465112 407172 465118
rect 407120 465054 407172 465060
rect 407118 463856 407174 463865
rect 407118 463791 407174 463800
rect 407132 463758 407160 463791
rect 407120 463752 407172 463758
rect 407120 463694 407172 463700
rect 407118 462496 407174 462505
rect 407118 462431 407120 462440
rect 407172 462431 407174 462440
rect 407120 462402 407172 462408
rect 407118 461816 407174 461825
rect 407118 461751 407174 461760
rect 407132 460970 407160 461751
rect 407120 460964 407172 460970
rect 407120 460906 407172 460912
rect 407118 459096 407174 459105
rect 407118 459031 407174 459040
rect 407132 458250 407160 459031
rect 407120 458244 407172 458250
rect 407120 458186 407172 458192
rect 407118 457056 407174 457065
rect 407118 456991 407174 457000
rect 407132 456822 407160 456991
rect 407120 456816 407172 456822
rect 407120 456758 407172 456764
rect 407120 455388 407172 455394
rect 407120 455330 407172 455336
rect 407132 454345 407160 455330
rect 407118 454336 407174 454345
rect 407118 454271 407174 454280
rect 407118 453656 407174 453665
rect 407118 453591 407174 453600
rect 407132 452674 407160 453591
rect 407120 452668 407172 452674
rect 407120 452610 407172 452616
rect 407118 451344 407174 451353
rect 407118 451279 407120 451288
rect 407172 451279 407174 451288
rect 407120 451250 407172 451256
rect 407118 449576 407174 449585
rect 407118 449511 407174 449520
rect 407132 448594 407160 449511
rect 407120 448588 407172 448594
rect 407120 448530 407172 448536
rect 407120 447092 407172 447098
rect 407120 447034 407172 447040
rect 407132 446185 407160 447034
rect 407118 446176 407174 446185
rect 407118 446111 407174 446120
rect 407120 445664 407172 445670
rect 407120 445606 407172 445612
rect 407132 444825 407160 445606
rect 407118 444816 407174 444825
rect 407118 444751 407174 444760
rect 407118 442096 407174 442105
rect 407118 442031 407174 442040
rect 407132 441658 407160 442031
rect 407120 441652 407172 441658
rect 407120 441594 407172 441600
rect 407118 440056 407174 440065
rect 407118 439991 407174 440000
rect 407132 438938 407160 439991
rect 407120 438932 407172 438938
rect 407120 438874 407172 438880
rect 407118 437336 407174 437345
rect 407118 437271 407174 437280
rect 407132 436150 407160 437271
rect 407120 436144 407172 436150
rect 407120 436086 407172 436092
rect 407118 435976 407174 435985
rect 407118 435911 407174 435920
rect 407132 434790 407160 435911
rect 407120 434784 407172 434790
rect 407120 434726 407172 434732
rect 407224 434625 407252 605806
rect 407684 602585 407712 605806
rect 407670 602576 407726 602585
rect 407670 602511 407726 602520
rect 407302 601896 407358 601905
rect 407302 601831 407358 601840
rect 407316 601730 407344 601831
rect 407304 601724 407356 601730
rect 407304 601666 407356 601672
rect 407762 601216 407818 601225
rect 407762 601151 407818 601160
rect 407302 599176 407358 599185
rect 407302 599111 407358 599120
rect 407316 599010 407344 599111
rect 407304 599004 407356 599010
rect 407304 598946 407356 598952
rect 407302 597136 407358 597145
rect 407302 597071 407358 597080
rect 407316 596222 407344 597071
rect 407304 596216 407356 596222
rect 407304 596158 407356 596164
rect 407302 595096 407358 595105
rect 407302 595031 407358 595040
rect 407316 594862 407344 595031
rect 407304 594856 407356 594862
rect 407304 594798 407356 594804
rect 407302 593056 407358 593065
rect 407302 592991 407358 593000
rect 407316 592074 407344 592991
rect 407304 592068 407356 592074
rect 407304 592010 407356 592016
rect 407302 591152 407358 591161
rect 407302 591087 407358 591096
rect 407316 590714 407344 591087
rect 407304 590708 407356 590714
rect 407304 590650 407356 590656
rect 407302 588976 407358 588985
rect 407302 588911 407358 588920
rect 407316 587926 407344 588911
rect 407304 587920 407356 587926
rect 407304 587862 407356 587868
rect 407776 587217 407804 601151
rect 407762 587208 407818 587217
rect 407762 587143 407818 587152
rect 407302 586936 407358 586945
rect 407302 586871 407358 586880
rect 407316 586566 407344 586871
rect 407304 586560 407356 586566
rect 407868 586514 407896 678286
rect 407948 678224 408000 678230
rect 407948 678166 408000 678172
rect 407960 605985 407988 678166
rect 407946 605976 408002 605985
rect 407946 605911 408002 605920
rect 407946 594416 408002 594425
rect 407946 594351 408002 594360
rect 407304 586502 407356 586508
rect 407684 586486 407896 586514
rect 407684 585585 407712 586486
rect 407960 586265 407988 594351
rect 407946 586256 408002 586265
rect 407946 586191 408002 586200
rect 407670 585576 407726 585585
rect 407670 585511 407726 585520
rect 407302 580136 407358 580145
rect 407302 580071 407358 580080
rect 407316 579698 407344 580071
rect 407304 579692 407356 579698
rect 407304 579634 407356 579640
rect 407302 577416 407358 577425
rect 407302 577351 407358 577360
rect 407316 576910 407344 577351
rect 407304 576904 407356 576910
rect 407304 576846 407356 576852
rect 407394 576736 407450 576745
rect 407394 576671 407450 576680
rect 407302 572656 407358 572665
rect 407302 572591 407358 572600
rect 407316 571402 407344 572591
rect 407304 571396 407356 571402
rect 407304 571338 407356 571344
rect 407302 569936 407358 569945
rect 407302 569871 407358 569880
rect 407316 568614 407344 569871
rect 407304 568608 407356 568614
rect 407304 568550 407356 568556
rect 407408 568426 407436 576671
rect 408052 574025 408080 684490
rect 408132 682712 408184 682718
rect 408132 682654 408184 682660
rect 408038 574016 408094 574025
rect 408038 573951 408094 573960
rect 407670 573336 407726 573345
rect 407670 573271 407726 573280
rect 407684 572762 407712 573271
rect 407672 572756 407724 572762
rect 407672 572698 407724 572704
rect 407316 568398 407436 568426
rect 407316 538214 407344 568398
rect 407394 567896 407450 567905
rect 407394 567831 407450 567840
rect 407408 567254 407436 567831
rect 407396 567248 407448 567254
rect 407396 567190 407448 567196
rect 407394 564496 407450 564505
rect 407394 564431 407396 564440
rect 407448 564431 407450 564440
rect 407396 564402 407448 564408
rect 407856 564120 407908 564126
rect 407856 564062 407908 564068
rect 407394 561096 407450 561105
rect 407394 561031 407450 561040
rect 407408 560318 407436 561031
rect 407396 560312 407448 560318
rect 407396 560254 407448 560260
rect 407672 559564 407724 559570
rect 407672 559506 407724 559512
rect 407684 557534 407712 559506
rect 407684 557506 407804 557534
rect 407672 557252 407724 557258
rect 407672 557194 407724 557200
rect 407684 557025 407712 557194
rect 407670 557016 407726 557025
rect 407670 556951 407726 556960
rect 407394 556336 407450 556345
rect 407394 556271 407450 556280
rect 407408 556238 407436 556271
rect 407396 556232 407448 556238
rect 407396 556174 407448 556180
rect 407486 552936 407542 552945
rect 407486 552871 407542 552880
rect 407500 552090 407528 552871
rect 407488 552084 407540 552090
rect 407488 552026 407540 552032
rect 407396 552016 407448 552022
rect 407396 551958 407448 551964
rect 407408 551585 407436 551958
rect 407394 551576 407450 551585
rect 407394 551511 407450 551520
rect 407394 550896 407450 550905
rect 407394 550831 407450 550840
rect 407408 550662 407436 550831
rect 407396 550656 407448 550662
rect 407396 550598 407448 550604
rect 407394 550216 407450 550225
rect 407394 550151 407450 550160
rect 407408 549302 407436 550151
rect 407396 549296 407448 549302
rect 407396 549238 407448 549244
rect 407488 549228 407540 549234
rect 407488 549170 407540 549176
rect 407500 548865 407528 549170
rect 407486 548856 407542 548865
rect 407486 548791 407542 548800
rect 407394 547496 407450 547505
rect 407394 547431 407450 547440
rect 407408 546582 407436 547431
rect 407396 546576 407448 546582
rect 407396 546518 407448 546524
rect 407394 544776 407450 544785
rect 407394 544711 407450 544720
rect 407408 543794 407436 544711
rect 407486 544096 407542 544105
rect 407486 544031 407542 544040
rect 407500 543862 407528 544031
rect 407488 543856 407540 543862
rect 407488 543798 407540 543804
rect 407396 543788 407448 543794
rect 407396 543730 407448 543736
rect 407396 542360 407448 542366
rect 407396 542302 407448 542308
rect 407408 542065 407436 542302
rect 407394 542056 407450 542065
rect 407394 541991 407450 542000
rect 407316 538186 407528 538214
rect 407302 535256 407358 535265
rect 407302 535191 407358 535200
rect 407316 534138 407344 535191
rect 407304 534132 407356 534138
rect 407304 534074 407356 534080
rect 407302 533896 407358 533905
rect 407302 533831 407358 533840
rect 407316 532778 407344 533831
rect 407304 532772 407356 532778
rect 407304 532714 407356 532720
rect 407302 531856 407358 531865
rect 407302 531791 407358 531800
rect 407316 531350 407344 531791
rect 407304 531344 407356 531350
rect 407304 531286 407356 531292
rect 407304 526516 407356 526522
rect 407304 526458 407356 526464
rect 407316 525842 407344 526458
rect 407304 525836 407356 525842
rect 407304 525778 407356 525784
rect 407316 525065 407344 525778
rect 407302 525056 407358 525065
rect 407302 524991 407358 525000
rect 407302 523696 407358 523705
rect 407302 523631 407358 523640
rect 407316 523054 407344 523631
rect 407304 523048 407356 523054
rect 407304 522990 407356 522996
rect 407394 523016 407450 523025
rect 407500 522986 407528 538186
rect 407394 522951 407450 522960
rect 407488 522980 407540 522986
rect 407408 521694 407436 522951
rect 407488 522922 407540 522928
rect 407396 521688 407448 521694
rect 407396 521630 407448 521636
rect 407302 518256 407358 518265
rect 407302 518191 407358 518200
rect 407316 517546 407344 518191
rect 407304 517540 407356 517546
rect 407304 517482 407356 517488
rect 407302 516896 407358 516905
rect 407302 516831 407358 516840
rect 407316 516186 407344 516831
rect 407304 516180 407356 516186
rect 407304 516122 407356 516128
rect 407580 516112 407632 516118
rect 407580 516054 407632 516060
rect 407592 514865 407620 516054
rect 407578 514856 407634 514865
rect 407578 514791 407634 514800
rect 407776 508065 407804 557506
rect 407868 552702 407896 564062
rect 407948 559632 408000 559638
rect 407948 559574 408000 559580
rect 407960 555665 407988 559574
rect 408038 559056 408094 559065
rect 408038 558991 408094 559000
rect 407946 555656 408002 555665
rect 407946 555591 408002 555600
rect 407856 552696 407908 552702
rect 407856 552638 407908 552644
rect 407762 508056 407818 508065
rect 407762 507991 407818 508000
rect 407302 489696 407358 489705
rect 407302 489631 407358 489640
rect 407316 488646 407344 489631
rect 407304 488640 407356 488646
rect 407304 488582 407356 488588
rect 407302 476096 407358 476105
rect 407302 476031 407358 476040
rect 407316 474842 407344 476031
rect 407304 474836 407356 474842
rect 407304 474778 407356 474784
rect 407302 474736 407358 474745
rect 407302 474671 407358 474680
rect 407316 473414 407344 474671
rect 407304 473408 407356 473414
rect 407304 473350 407356 473356
rect 407304 469192 407356 469198
rect 407304 469134 407356 469140
rect 407316 467945 407344 469134
rect 407302 467936 407358 467945
rect 407302 467871 407358 467880
rect 407302 463176 407358 463185
rect 407302 463111 407358 463120
rect 407316 462398 407344 463111
rect 407304 462392 407356 462398
rect 407304 462334 407356 462340
rect 407304 456748 407356 456754
rect 407304 456690 407356 456696
rect 407316 455705 407344 456690
rect 407302 455696 407358 455705
rect 407302 455631 407358 455640
rect 407670 455016 407726 455025
rect 407670 454951 407726 454960
rect 407684 454102 407712 454951
rect 407672 454096 407724 454102
rect 407672 454038 407724 454044
rect 407302 447264 407358 447273
rect 407302 447199 407358 447208
rect 407316 447166 407344 447199
rect 407304 447160 407356 447166
rect 407304 447102 407356 447108
rect 407304 441584 407356 441590
rect 407304 441526 407356 441532
rect 407316 441425 407344 441526
rect 407302 441416 407358 441425
rect 407302 441351 407358 441360
rect 407488 438864 407540 438870
rect 407488 438806 407540 438812
rect 407500 438705 407528 438806
rect 407486 438696 407542 438705
rect 407486 438631 407542 438640
rect 407210 434616 407266 434625
rect 407210 434551 407266 434560
rect 407118 429856 407174 429865
rect 407118 429791 407174 429800
rect 407132 429282 407160 429791
rect 407120 429276 407172 429282
rect 407120 429218 407172 429224
rect 407118 429176 407174 429185
rect 407118 429111 407174 429120
rect 407132 427922 407160 429111
rect 407120 427916 407172 427922
rect 407120 427858 407172 427864
rect 407210 427816 407266 427825
rect 407210 427751 407266 427760
rect 407118 427136 407174 427145
rect 407118 427071 407174 427080
rect 407132 426562 407160 427071
rect 407224 426630 407252 427751
rect 407212 426624 407264 426630
rect 407212 426566 407264 426572
rect 407120 426556 407172 426562
rect 407120 426498 407172 426504
rect 407946 425776 408002 425785
rect 407946 425711 408002 425720
rect 407118 423736 407174 423745
rect 407118 423671 407120 423680
rect 407172 423671 407174 423680
rect 407120 423642 407172 423648
rect 407118 423056 407174 423065
rect 407118 422991 407174 423000
rect 407132 422346 407160 422991
rect 407120 422340 407172 422346
rect 407120 422282 407172 422288
rect 407854 421696 407910 421705
rect 407854 421631 407910 421640
rect 407210 420336 407266 420345
rect 407210 420271 407266 420280
rect 407118 419656 407174 419665
rect 407224 419626 407252 420271
rect 407118 419591 407174 419600
rect 407212 419620 407264 419626
rect 407132 419558 407160 419591
rect 407212 419562 407264 419568
rect 407120 419552 407172 419558
rect 407120 419494 407172 419500
rect 407118 418976 407174 418985
rect 407118 418911 407174 418920
rect 407132 418198 407160 418911
rect 407120 418192 407172 418198
rect 407120 418134 407172 418140
rect 407120 416764 407172 416770
rect 407120 416706 407172 416712
rect 407132 416265 407160 416706
rect 407118 416256 407174 416265
rect 407118 416191 407174 416200
rect 407118 414896 407174 414905
rect 407118 414831 407174 414840
rect 407132 414050 407160 414831
rect 407120 414044 407172 414050
rect 407120 413986 407172 413992
rect 407118 411496 407174 411505
rect 407118 411431 407174 411440
rect 407132 411330 407160 411431
rect 407120 411324 407172 411330
rect 407120 411266 407172 411272
rect 407118 410816 407174 410825
rect 407118 410751 407174 410760
rect 407132 409902 407160 410751
rect 407120 409896 407172 409902
rect 407120 409838 407172 409844
rect 407118 408776 407174 408785
rect 407118 408711 407174 408720
rect 407132 408542 407160 408711
rect 407120 408536 407172 408542
rect 407120 408478 407172 408484
rect 407118 406056 407174 406065
rect 407118 405991 407174 406000
rect 407132 405754 407160 405991
rect 407120 405748 407172 405754
rect 407120 405690 407172 405696
rect 407212 405680 407264 405686
rect 407212 405622 407264 405628
rect 407224 404705 407252 405622
rect 407210 404696 407266 404705
rect 407210 404631 407266 404640
rect 407762 401976 407818 401985
rect 407762 401911 407818 401920
rect 407486 400344 407542 400353
rect 407486 400279 407542 400288
rect 407500 400246 407528 400279
rect 407488 400240 407540 400246
rect 407488 400182 407540 400188
rect 407120 400172 407172 400178
rect 407120 400114 407172 400120
rect 407132 399265 407160 400114
rect 407118 399256 407174 399265
rect 407118 399191 407174 399200
rect 407118 397896 407174 397905
rect 407118 397831 407174 397840
rect 407132 397526 407160 397831
rect 407120 397520 407172 397526
rect 407120 397462 407172 397468
rect 407210 395856 407266 395865
rect 407210 395791 407266 395800
rect 407118 395176 407174 395185
rect 407118 395111 407174 395120
rect 407132 394738 407160 395111
rect 407224 394806 407252 395791
rect 407212 394800 407264 394806
rect 407212 394742 407264 394748
rect 407120 394732 407172 394738
rect 407120 394674 407172 394680
rect 407118 393816 407174 393825
rect 407118 393751 407174 393760
rect 407132 393378 407160 393751
rect 407120 393372 407172 393378
rect 407120 393314 407172 393320
rect 407578 393136 407634 393145
rect 407578 393071 407634 393080
rect 407210 391776 407266 391785
rect 407210 391711 407266 391720
rect 407118 391096 407174 391105
rect 407118 391031 407174 391040
rect 407132 390590 407160 391031
rect 407224 390658 407252 391711
rect 407212 390652 407264 390658
rect 407212 390594 407264 390600
rect 407120 390584 407172 390590
rect 407120 390526 407172 390532
rect 407118 389736 407174 389745
rect 407118 389671 407174 389680
rect 407132 389230 407160 389671
rect 407120 389224 407172 389230
rect 407120 389166 407172 389172
rect 407120 386368 407172 386374
rect 407120 386310 407172 386316
rect 407132 385665 407160 386310
rect 407118 385656 407174 385665
rect 407118 385591 407174 385600
rect 407118 384976 407174 384985
rect 407118 384911 407174 384920
rect 407132 383994 407160 384911
rect 407120 383988 407172 383994
rect 407120 383930 407172 383936
rect 407118 382936 407174 382945
rect 407118 382871 407174 382880
rect 407132 382294 407160 382871
rect 407120 382288 407172 382294
rect 407120 382230 407172 382236
rect 407118 381576 407174 381585
rect 407118 381511 407174 381520
rect 407132 380934 407160 381511
rect 407120 380928 407172 380934
rect 407120 380870 407172 380876
rect 407118 378856 407174 378865
rect 407118 378791 407174 378800
rect 407132 378214 407160 378791
rect 407120 378208 407172 378214
rect 407120 378150 407172 378156
rect 407118 373416 407174 373425
rect 407118 373351 407174 373360
rect 407132 372638 407160 373351
rect 407120 372632 407172 372638
rect 407120 372574 407172 372580
rect 407120 371204 407172 371210
rect 407120 371146 407172 371152
rect 407132 370705 407160 371146
rect 407118 370696 407174 370705
rect 407118 370631 407174 370640
rect 407120 361548 407172 361554
rect 407120 361490 407172 361496
rect 407132 361185 407160 361490
rect 407118 361176 407174 361185
rect 407118 361111 407174 361120
rect 407118 360496 407174 360505
rect 407118 360431 407174 360440
rect 407132 360262 407160 360431
rect 407120 360256 407172 360262
rect 407120 360198 407172 360204
rect 407118 357096 407174 357105
rect 407118 357031 407174 357040
rect 407132 356250 407160 357031
rect 407120 356244 407172 356250
rect 407120 356186 407172 356192
rect 407118 353696 407174 353705
rect 407118 353631 407174 353640
rect 407132 353326 407160 353631
rect 407120 353320 407172 353326
rect 407120 353262 407172 353268
rect 407210 353016 407266 353025
rect 407210 352951 407266 352960
rect 407118 352336 407174 352345
rect 407118 352271 407174 352280
rect 407132 352034 407160 352271
rect 407120 352028 407172 352034
rect 407120 351970 407172 351976
rect 407224 351966 407252 352951
rect 407212 351960 407264 351966
rect 407212 351902 407264 351908
rect 407118 351656 407174 351665
rect 407118 351591 407174 351600
rect 407132 350606 407160 351591
rect 407120 350600 407172 350606
rect 407120 350542 407172 350548
rect 407118 349208 407174 349217
rect 407118 349143 407120 349152
rect 407172 349143 407174 349152
rect 407120 349114 407172 349120
rect 407118 346896 407174 346905
rect 407118 346831 407174 346840
rect 407132 346458 407160 346831
rect 407120 346452 407172 346458
rect 407120 346394 407172 346400
rect 407120 345024 407172 345030
rect 407120 344966 407172 344972
rect 407132 344865 407160 344966
rect 407118 344856 407174 344865
rect 407118 344791 407174 344800
rect 407118 343496 407174 343505
rect 407118 343431 407174 343440
rect 407132 342310 407160 343431
rect 407120 342304 407172 342310
rect 407120 342246 407172 342252
rect 407118 340776 407174 340785
rect 407118 340711 407174 340720
rect 407132 339522 407160 340711
rect 407120 339516 407172 339522
rect 407120 339458 407172 339464
rect 407118 339416 407174 339425
rect 407118 339351 407174 339360
rect 407132 338162 407160 339351
rect 407120 338156 407172 338162
rect 407120 338098 407172 338104
rect 407120 336728 407172 336734
rect 407118 336696 407120 336705
rect 407172 336696 407174 336705
rect 407118 336631 407174 336640
rect 407394 332616 407450 332625
rect 407394 332551 407450 332560
rect 407118 330576 407174 330585
rect 407118 330511 407174 330520
rect 407132 329866 407160 330511
rect 407120 329860 407172 329866
rect 407120 329802 407172 329808
rect 407118 328536 407174 328545
rect 407118 328471 407120 328480
rect 407172 328471 407174 328480
rect 407120 328442 407172 328448
rect 407118 327856 407174 327865
rect 407118 327791 407174 327800
rect 407132 327146 407160 327791
rect 407120 327140 407172 327146
rect 407120 327082 407172 327088
rect 407118 325816 407174 325825
rect 407118 325751 407174 325760
rect 407132 325718 407160 325751
rect 407120 325712 407172 325718
rect 407120 325654 407172 325660
rect 407212 325644 407264 325650
rect 407212 325586 407264 325592
rect 407224 325145 407252 325586
rect 407210 325136 407266 325145
rect 407210 325071 407266 325080
rect 407210 323776 407266 323785
rect 407210 323711 407266 323720
rect 407118 323096 407174 323105
rect 407224 323066 407252 323711
rect 407118 323031 407174 323040
rect 407212 323060 407264 323066
rect 407132 322998 407160 323031
rect 407212 323002 407264 323008
rect 407120 322992 407172 322998
rect 407120 322934 407172 322940
rect 407212 322924 407264 322930
rect 407212 322866 407264 322872
rect 407120 322856 407172 322862
rect 407120 322798 407172 322804
rect 407132 321745 407160 322798
rect 407224 322425 407252 322866
rect 407210 322416 407266 322425
rect 407210 322351 407266 322360
rect 407118 321736 407174 321745
rect 407118 321671 407174 321680
rect 407302 321056 407358 321065
rect 407302 320991 407358 321000
rect 407316 320210 407344 320991
rect 407304 320204 407356 320210
rect 407304 320146 407356 320152
rect 407118 315616 407174 315625
rect 407118 315551 407174 315560
rect 407132 314702 407160 315551
rect 407120 314696 407172 314702
rect 407120 314638 407172 314644
rect 407210 311128 407266 311137
rect 407210 311063 407266 311072
rect 407118 310856 407174 310865
rect 407118 310791 407174 310800
rect 407132 310622 407160 310791
rect 407120 310616 407172 310622
rect 407120 310558 407172 310564
rect 407224 310554 407252 311063
rect 407212 310548 407264 310554
rect 407212 310490 407264 310496
rect 407120 310480 407172 310486
rect 407120 310422 407172 310428
rect 407132 310185 407160 310422
rect 407118 310176 407174 310185
rect 407118 310111 407174 310120
rect 407118 308136 407174 308145
rect 407118 308071 407174 308080
rect 407132 307902 407160 308071
rect 407120 307896 407172 307902
rect 407120 307838 407172 307844
rect 407120 307760 407172 307766
rect 407120 307702 407172 307708
rect 407132 306785 407160 307702
rect 407118 306776 407174 306785
rect 407118 306711 407174 306720
rect 407118 305416 407174 305425
rect 407118 305351 407174 305360
rect 407132 305046 407160 305351
rect 407120 305040 407172 305046
rect 407120 304982 407172 304988
rect 407118 304056 407174 304065
rect 407118 303991 407174 304000
rect 407132 303686 407160 303991
rect 407120 303680 407172 303686
rect 407120 303622 407172 303628
rect 407210 302016 407266 302025
rect 407210 301951 407266 301960
rect 407118 301336 407174 301345
rect 407118 301271 407174 301280
rect 407132 300966 407160 301271
rect 407120 300960 407172 300966
rect 407120 300902 407172 300908
rect 407224 300898 407252 301951
rect 407212 300892 407264 300898
rect 407212 300834 407264 300840
rect 407118 299976 407174 299985
rect 407118 299911 407174 299920
rect 407132 299538 407160 299911
rect 407120 299532 407172 299538
rect 407120 299474 407172 299480
rect 407118 295896 407174 295905
rect 407118 295831 407174 295840
rect 407132 295390 407160 295831
rect 407120 295384 407172 295390
rect 407120 295326 407172 295332
rect 407210 293856 407266 293865
rect 407210 293791 407266 293800
rect 407224 292602 407252 293791
rect 407212 292596 407264 292602
rect 407212 292538 407264 292544
rect 407120 292528 407172 292534
rect 407118 292496 407120 292505
rect 407172 292496 407174 292505
rect 407118 292431 407174 292440
rect 407212 292460 407264 292466
rect 407212 292402 407264 292408
rect 407224 291825 407252 292402
rect 407210 291816 407266 291825
rect 407210 291751 407266 291760
rect 407118 289776 407174 289785
rect 407118 289711 407174 289720
rect 407132 288522 407160 289711
rect 407302 289096 407358 289105
rect 407302 289031 407358 289040
rect 407120 288516 407172 288522
rect 407120 288458 407172 288464
rect 407316 288454 407344 289031
rect 407304 288448 407356 288454
rect 407210 288416 407266 288425
rect 407304 288390 407356 288396
rect 407210 288351 407266 288360
rect 407118 287736 407174 287745
rect 407118 287671 407174 287680
rect 407132 287162 407160 287671
rect 407120 287156 407172 287162
rect 407120 287098 407172 287104
rect 407224 287094 407252 288351
rect 407212 287088 407264 287094
rect 407118 287056 407174 287065
rect 407212 287030 407264 287036
rect 407118 286991 407174 287000
rect 407132 285802 407160 286991
rect 407120 285796 407172 285802
rect 407120 285738 407172 285744
rect 407120 284368 407172 284374
rect 407118 284336 407120 284345
rect 407172 284336 407174 284345
rect 407118 284271 407174 284280
rect 407212 284300 407264 284306
rect 407212 284242 407264 284248
rect 407224 283665 407252 284242
rect 407210 283656 407266 283665
rect 407210 283591 407266 283600
rect 407118 282976 407174 282985
rect 407118 282911 407120 282920
rect 407172 282911 407174 282920
rect 407120 282882 407172 282888
rect 407210 279576 407266 279585
rect 407210 279511 407266 279520
rect 407118 278896 407174 278905
rect 407118 278831 407120 278840
rect 407172 278831 407174 278840
rect 407120 278802 407172 278808
rect 407224 278798 407252 279511
rect 407212 278792 407264 278798
rect 407212 278734 407264 278740
rect 407120 277364 407172 277370
rect 407120 277306 407172 277312
rect 407132 276185 407160 277306
rect 407118 276176 407174 276185
rect 407118 276111 407174 276120
rect 407120 275936 407172 275942
rect 407120 275878 407172 275884
rect 407132 275505 407160 275878
rect 407118 275496 407174 275505
rect 407118 275431 407174 275440
rect 407120 271856 407172 271862
rect 407120 271798 407172 271804
rect 407132 271425 407160 271798
rect 407118 271416 407174 271425
rect 407118 271351 407174 271360
rect 407118 270056 407174 270065
rect 407118 269991 407174 270000
rect 407132 269142 407160 269991
rect 407120 269136 407172 269142
rect 407120 269078 407172 269084
rect 407118 268016 407174 268025
rect 407118 267951 407174 267960
rect 407132 267782 407160 267951
rect 407120 267776 407172 267782
rect 407120 267718 407172 267724
rect 407118 263936 407174 263945
rect 407118 263871 407174 263880
rect 407132 263634 407160 263871
rect 407120 263628 407172 263634
rect 407120 263570 407172 263576
rect 407118 262576 407174 262585
rect 407118 262511 407174 262520
rect 407132 262274 407160 262511
rect 407120 262268 407172 262274
rect 407120 262210 407172 262216
rect 407118 261896 407174 261905
rect 407118 261831 407174 261840
rect 407132 260914 407160 261831
rect 407120 260908 407172 260914
rect 407120 260850 407172 260856
rect 407118 259856 407174 259865
rect 407118 259791 407174 259800
rect 407132 259486 407160 259791
rect 407120 259480 407172 259486
rect 407120 259422 407172 259428
rect 407210 257816 407266 257825
rect 407210 257751 407266 257760
rect 407118 257136 407174 257145
rect 407118 257071 407174 257080
rect 407132 256834 407160 257071
rect 407120 256828 407172 256834
rect 407120 256770 407172 256776
rect 407224 256766 407252 257751
rect 407212 256760 407264 256766
rect 407212 256702 407264 256708
rect 407118 255096 407174 255105
rect 407118 255031 407174 255040
rect 407132 253978 407160 255031
rect 407304 254040 407356 254046
rect 407304 253982 407356 253988
rect 407120 253972 407172 253978
rect 407120 253914 407172 253920
rect 407118 251696 407174 251705
rect 407118 251631 407174 251640
rect 407132 251258 407160 251631
rect 407120 251252 407172 251258
rect 407120 251194 407172 251200
rect 407212 251184 407264 251190
rect 407212 251126 407264 251132
rect 407118 251016 407174 251025
rect 407118 250951 407174 250960
rect 407132 249898 407160 250951
rect 407224 250345 407252 251126
rect 407210 250336 407266 250345
rect 407210 250271 407266 250280
rect 407120 249892 407172 249898
rect 407120 249834 407172 249840
rect 407210 246936 407266 246945
rect 407210 246871 407266 246880
rect 407118 246256 407174 246265
rect 407118 246191 407174 246200
rect 407132 245750 407160 246191
rect 407120 245744 407172 245750
rect 407120 245686 407172 245692
rect 407224 245682 407252 246871
rect 407212 245676 407264 245682
rect 407212 245618 407264 245624
rect 407118 244896 407174 244905
rect 407118 244831 407174 244840
rect 407132 244390 407160 244831
rect 407120 244384 407172 244390
rect 407120 244326 407172 244332
rect 407316 244322 407344 253982
rect 407304 244316 407356 244322
rect 407304 244258 407356 244264
rect 407120 242888 407172 242894
rect 407120 242830 407172 242836
rect 407132 242185 407160 242830
rect 407118 242176 407174 242185
rect 407118 242111 407174 242120
rect 407304 169108 407356 169114
rect 407304 169050 407356 169056
rect 407120 167884 407172 167890
rect 407120 167826 407172 167832
rect 407028 152856 407080 152862
rect 407028 152798 407080 152804
rect 406936 152788 406988 152794
rect 406936 152730 406988 152736
rect 406752 150884 406804 150890
rect 406752 150826 406804 150832
rect 407132 149940 407160 167826
rect 407316 149954 407344 169050
rect 407408 155854 407436 332551
rect 407592 316034 407620 393071
rect 407672 369164 407724 369170
rect 407672 369106 407724 369112
rect 407500 316006 407620 316034
rect 407500 300665 407528 316006
rect 407580 307488 407632 307494
rect 407580 307430 407632 307436
rect 407592 304298 407620 307430
rect 407580 304292 407632 304298
rect 407580 304234 407632 304240
rect 407486 300656 407542 300665
rect 407486 300591 407542 300600
rect 407578 298616 407634 298625
rect 407578 298551 407634 298560
rect 407488 272604 407540 272610
rect 407488 272546 407540 272552
rect 407500 261186 407528 272546
rect 407592 261186 407620 298551
rect 407488 261180 407540 261186
rect 407488 261122 407540 261128
rect 407580 261180 407632 261186
rect 407580 261122 407632 261128
rect 407684 261066 407712 369106
rect 407776 272610 407804 401911
rect 407868 295458 407896 421631
rect 407960 307494 407988 425711
rect 408052 362545 408080 558991
rect 408144 457745 408172 682654
rect 408316 681080 408368 681086
rect 408316 681022 408368 681028
rect 408222 678328 408278 678337
rect 408222 678263 408278 678272
rect 408236 466585 408264 678263
rect 408328 565185 408356 681022
rect 408420 678230 408448 685170
rect 408960 680876 409012 680882
rect 408960 680818 409012 680824
rect 408866 680096 408922 680105
rect 408866 680031 408922 680040
rect 408880 679114 408908 680031
rect 408868 679108 408920 679114
rect 408868 679050 408920 679056
rect 408408 678224 408460 678230
rect 408408 678166 408460 678172
rect 408406 667176 408462 667185
rect 408406 667111 408462 667120
rect 408314 565176 408370 565185
rect 408314 565111 408370 565120
rect 408316 552696 408368 552702
rect 408316 552638 408368 552644
rect 408328 546145 408356 552638
rect 408314 546136 408370 546145
rect 408314 546071 408370 546080
rect 408314 501256 408370 501265
rect 408314 501191 408370 501200
rect 408222 466576 408278 466585
rect 408222 466511 408278 466520
rect 408222 466440 408278 466449
rect 408222 466375 408278 466384
rect 408130 457736 408186 457745
rect 408130 457671 408186 457680
rect 408130 433936 408186 433945
rect 408130 433871 408186 433880
rect 408144 378826 408172 433871
rect 408132 378820 408184 378826
rect 408132 378762 408184 378768
rect 408130 374096 408186 374105
rect 408130 374031 408186 374040
rect 408144 369170 408172 374031
rect 408132 369164 408184 369170
rect 408132 369106 408184 369112
rect 408038 362536 408094 362545
rect 408038 362471 408094 362480
rect 408130 335336 408186 335345
rect 408130 335271 408186 335280
rect 408038 312896 408094 312905
rect 408038 312831 408094 312840
rect 407948 307488 408000 307494
rect 407948 307430 408000 307436
rect 407946 302696 408002 302705
rect 407946 302631 408002 302640
rect 407856 295452 407908 295458
rect 407856 295394 407908 295400
rect 407854 276856 407910 276865
rect 407854 276791 407910 276800
rect 407764 272604 407816 272610
rect 407764 272546 407816 272552
rect 407762 267336 407818 267345
rect 407762 267271 407818 267280
rect 407776 266422 407804 267271
rect 407764 266416 407816 266422
rect 407764 266358 407816 266364
rect 407500 261038 407712 261066
rect 407500 256018 407528 261038
rect 407580 260976 407632 260982
rect 407580 260918 407632 260924
rect 407488 256012 407540 256018
rect 407488 255954 407540 255960
rect 407488 255264 407540 255270
rect 407488 255206 407540 255212
rect 407500 254425 407528 255206
rect 407486 254416 407542 254425
rect 407486 254351 407542 254360
rect 407592 245818 407620 260918
rect 407762 249656 407818 249665
rect 407762 249591 407818 249600
rect 407776 248810 407804 249591
rect 407764 248804 407816 248810
rect 407764 248746 407816 248752
rect 407580 245812 407632 245818
rect 407580 245754 407632 245760
rect 407764 244316 407816 244322
rect 407764 244258 407816 244264
rect 407578 242992 407634 243001
rect 407578 242927 407634 242936
rect 407592 233102 407620 242927
rect 407580 233096 407632 233102
rect 407580 233038 407632 233044
rect 407776 155922 407804 244258
rect 407868 167822 407896 276791
rect 407856 167816 407908 167822
rect 407856 167758 407908 167764
rect 407960 157282 407988 302631
rect 407948 157276 408000 157282
rect 407948 157218 408000 157224
rect 407764 155916 407816 155922
rect 407764 155858 407816 155864
rect 407396 155848 407448 155854
rect 407396 155790 407448 155796
rect 408052 152930 408080 312831
rect 408144 153814 408172 335271
rect 408236 159322 408264 466375
rect 408328 160070 408356 501191
rect 408420 319025 408448 667111
rect 408972 578105 409000 680818
rect 408958 578096 409014 578105
rect 408958 578031 409014 578040
rect 409064 510105 409092 685238
rect 409156 570625 409184 685306
rect 454224 685296 454276 685302
rect 445114 685264 445170 685273
rect 436100 685228 436152 685234
rect 454224 685238 454276 685244
rect 445114 685199 445170 685208
rect 436100 685170 436152 685176
rect 409696 685160 409748 685166
rect 409696 685102 409748 685108
rect 409236 684956 409288 684962
rect 409236 684898 409288 684904
rect 409142 570616 409198 570625
rect 409142 570551 409198 570560
rect 409144 522980 409196 522986
rect 409144 522922 409196 522928
rect 409050 510096 409106 510105
rect 409050 510031 409106 510040
rect 408500 376780 408552 376786
rect 408500 376722 408552 376728
rect 408406 319016 408462 319025
rect 408406 318951 408462 318960
rect 408406 293992 408462 294001
rect 408406 293927 408462 293936
rect 408420 276826 408448 293927
rect 408408 276820 408460 276826
rect 408408 276762 408460 276768
rect 408406 259992 408462 260001
rect 408406 259927 408462 259936
rect 408420 239873 408448 259927
rect 408512 244322 408540 376722
rect 409156 285025 409184 522922
rect 409248 479505 409276 684898
rect 409512 684752 409564 684758
rect 409512 684694 409564 684700
rect 409328 683868 409380 683874
rect 409328 683810 409380 683816
rect 409234 479496 409290 479505
rect 409234 479431 409290 479440
rect 409340 476785 409368 683810
rect 409420 680468 409472 680474
rect 409420 680410 409472 680416
rect 409326 476776 409382 476785
rect 409326 476711 409382 476720
rect 409234 472016 409290 472025
rect 409234 471951 409290 471960
rect 409248 307086 409276 471951
rect 409432 428505 409460 680410
rect 409524 430545 409552 684694
rect 409604 679720 409656 679726
rect 409604 679662 409656 679668
rect 409616 459785 409644 679662
rect 409602 459776 409658 459785
rect 409602 459711 409658 459720
rect 409602 452976 409658 452985
rect 409602 452911 409658 452920
rect 409510 430536 409566 430545
rect 409510 430471 409566 430480
rect 409418 428496 409474 428505
rect 409418 428431 409474 428440
rect 409510 412176 409566 412185
rect 409510 412111 409566 412120
rect 409328 378820 409380 378826
rect 409328 378762 409380 378768
rect 409236 307080 409288 307086
rect 409236 307022 409288 307028
rect 409142 285016 409198 285025
rect 409142 284951 409198 284960
rect 409144 276820 409196 276826
rect 409144 276762 409196 276768
rect 408972 245614 409000 245645
rect 408960 245608 409012 245614
rect 408958 245576 408960 245585
rect 409012 245576 409014 245585
rect 408958 245511 409014 245520
rect 408500 244316 408552 244322
rect 408500 244258 408552 244264
rect 408868 243568 408920 243574
rect 408868 243510 408920 243516
rect 408406 239864 408462 239873
rect 408406 239799 408462 239808
rect 408880 238754 408908 243510
rect 408972 239766 409000 245511
rect 409052 244316 409104 244322
rect 409052 244258 409104 244264
rect 408960 239760 409012 239766
rect 408960 239702 409012 239708
rect 409064 239698 409092 244258
rect 409052 239692 409104 239698
rect 409052 239634 409104 239640
rect 408880 238726 409000 238754
rect 408316 160064 408368 160070
rect 408316 160006 408368 160012
rect 408224 159316 408276 159322
rect 408224 159258 408276 159264
rect 408132 153808 408184 153814
rect 408132 153750 408184 153756
rect 408040 152924 408092 152930
rect 408040 152866 408092 152872
rect 408972 150958 409000 238726
rect 409050 152416 409106 152425
rect 409050 152351 409106 152360
rect 408960 150952 409012 150958
rect 408960 150894 409012 150900
rect 403164 149932 403216 149938
rect 370964 149874 371016 149880
rect 407316 149926 408434 149954
rect 409064 149940 409092 152351
rect 409156 152318 409184 276762
rect 409236 253224 409288 253230
rect 409236 253166 409288 253172
rect 409248 159526 409276 253166
rect 409340 238338 409368 378762
rect 409418 318336 409474 318345
rect 409418 318271 409474 318280
rect 409432 244322 409460 318271
rect 409420 244316 409472 244322
rect 409420 244258 409472 244264
rect 409524 244202 409552 412111
rect 409432 244174 409552 244202
rect 409432 239630 409460 244174
rect 409510 241224 409566 241233
rect 409510 241159 409566 241168
rect 409524 241126 409552 241159
rect 409512 241120 409564 241126
rect 409512 241062 409564 241068
rect 409510 240816 409566 240825
rect 409510 240751 409566 240760
rect 409524 240650 409552 240751
rect 409512 240644 409564 240650
rect 409512 240586 409564 240592
rect 409420 239624 409472 239630
rect 409420 239566 409472 239572
rect 409328 238332 409380 238338
rect 409328 238274 409380 238280
rect 409236 159520 409288 159526
rect 409236 159462 409288 159468
rect 409616 152726 409644 452911
rect 409708 364585 409736 685102
rect 416134 684992 416190 685001
rect 416134 684927 416190 684936
rect 409788 684072 409840 684078
rect 409788 684014 409840 684020
rect 409694 364576 409750 364585
rect 409694 364511 409750 364520
rect 409694 342816 409750 342825
rect 409694 342751 409750 342760
rect 409708 233782 409736 342751
rect 409800 334665 409828 684014
rect 413558 683496 413614 683505
rect 413558 683431 413614 683440
rect 412914 682000 412970 682009
rect 412914 681935 412970 681944
rect 409880 680944 409932 680950
rect 409880 680886 409932 680892
rect 409892 665145 409920 680886
rect 411626 680368 411682 680377
rect 411626 680303 411682 680312
rect 411640 679946 411668 680303
rect 412928 679946 412956 681935
rect 413572 679946 413600 683431
rect 416148 679946 416176 684927
rect 425794 684856 425850 684865
rect 425794 684791 425850 684800
rect 423862 683768 423918 683777
rect 423862 683703 423918 683712
rect 422392 683664 422444 683670
rect 422392 683606 422444 683612
rect 416688 683256 416740 683262
rect 416688 683198 416740 683204
rect 416700 679946 416728 683198
rect 411640 679918 411976 679946
rect 412928 679918 413264 679946
rect 413572 679918 413908 679946
rect 415840 679918 416176 679946
rect 416484 679918 416728 679946
rect 419998 679960 420054 679969
rect 420054 679918 420348 679946
rect 419998 679895 420054 679904
rect 411260 679856 411312 679862
rect 411260 679798 411312 679804
rect 421472 679856 421524 679862
rect 422404 679810 422432 683606
rect 423876 679946 423904 683703
rect 424508 680468 424560 680474
rect 424508 680410 424560 680416
rect 424520 679946 424548 680410
rect 425808 679946 425836 684791
rect 435456 684616 435508 684622
rect 435456 684558 435508 684564
rect 429660 682168 429712 682174
rect 429660 682110 429712 682116
rect 428370 681864 428426 681873
rect 428370 681799 428426 681808
rect 427912 680400 427964 680406
rect 427912 680342 427964 680348
rect 423876 679918 424212 679946
rect 424520 679918 424856 679946
rect 425500 679918 425836 679946
rect 427924 679946 427952 680342
rect 428384 679946 428412 681799
rect 429672 679946 429700 682110
rect 432052 681012 432104 681018
rect 432052 680954 432104 680960
rect 434628 681012 434680 681018
rect 434628 680954 434680 680960
rect 427924 679918 428076 679946
rect 428384 679918 428720 679946
rect 429672 679918 430008 679946
rect 432064 679810 432092 680954
rect 433522 679960 433578 679969
rect 434640 679946 434668 680954
rect 435468 679946 435496 684558
rect 433578 679918 433872 679946
rect 434516 679918 434668 679946
rect 435160 679918 435496 679946
rect 435824 679992 435876 679998
rect 435824 679934 435876 679940
rect 436112 679946 436140 685170
rect 442538 684584 442594 684593
rect 442538 684519 442594 684528
rect 437572 683732 437624 683738
rect 437572 683674 437624 683680
rect 437584 679946 437612 683674
rect 441252 683664 441304 683670
rect 441252 683606 441304 683612
rect 438676 683596 438728 683602
rect 438676 683538 438728 683544
rect 437940 680128 437992 680134
rect 437940 680070 437992 680076
rect 433522 679895 433578 679904
rect 421472 679798 421524 679804
rect 411272 679522 411300 679798
rect 413744 679788 413796 679794
rect 413744 679730 413796 679736
rect 415216 679788 415268 679794
rect 415216 679730 415268 679736
rect 413756 679522 413784 679730
rect 415228 679590 415256 679730
rect 415492 679720 415544 679726
rect 415366 679668 415492 679674
rect 415366 679662 415544 679668
rect 415366 679658 415532 679662
rect 415354 679652 415532 679658
rect 415406 679646 415532 679652
rect 415354 679594 415406 679600
rect 415216 679584 415268 679590
rect 415216 679526 415268 679532
rect 421484 679522 421512 679798
rect 422280 679782 422432 679810
rect 431940 679782 432092 679810
rect 432696 679584 432748 679590
rect 432584 679532 432696 679538
rect 432584 679526 432748 679532
rect 411260 679516 411312 679522
rect 411260 679458 411312 679464
rect 413744 679516 413796 679522
rect 413744 679458 413796 679464
rect 421472 679516 421524 679522
rect 432584 679510 432736 679526
rect 432800 679522 433012 679538
rect 435836 679522 435864 679934
rect 436112 679918 436448 679946
rect 437584 679918 437736 679946
rect 437952 679522 437980 680070
rect 438688 679810 438716 683538
rect 439964 682304 440016 682310
rect 439964 682246 440016 682252
rect 439320 680400 439372 680406
rect 439320 680342 439372 680348
rect 439332 679946 439360 680342
rect 439024 679918 439360 679946
rect 438380 679782 438716 679810
rect 439976 679810 440004 682246
rect 441264 679946 441292 683606
rect 441896 682508 441948 682514
rect 441896 682450 441948 682456
rect 441804 680060 441856 680066
rect 441804 680002 441856 680008
rect 440956 679918 441292 679946
rect 441712 679924 441764 679930
rect 441712 679866 441764 679872
rect 439976 679782 440312 679810
rect 441724 679522 441752 679866
rect 441816 679522 441844 680002
rect 441908 679946 441936 682450
rect 442552 679946 442580 684519
rect 443000 682168 443052 682174
rect 443000 682110 443052 682116
rect 443012 681154 443040 682110
rect 443000 681148 443052 681154
rect 443000 681090 443052 681096
rect 445128 679946 445156 685199
rect 450268 685160 450320 685166
rect 450268 685102 450320 685108
rect 449900 684072 449952 684078
rect 449900 684014 449952 684020
rect 447690 682408 447746 682417
rect 447690 682343 447746 682352
rect 447140 682304 447192 682310
rect 447140 682246 447192 682252
rect 446862 681184 446918 681193
rect 446862 681119 446918 681128
rect 446220 680128 446272 680134
rect 446220 680070 446272 680076
rect 445760 680060 445812 680066
rect 445760 680002 445812 680008
rect 441908 679918 442244 679946
rect 442552 679918 442888 679946
rect 445128 679918 445464 679946
rect 442356 679788 442408 679794
rect 442356 679730 442408 679736
rect 442368 679522 442396 679730
rect 443920 679720 443972 679726
rect 443920 679662 443972 679668
rect 443932 679522 443960 679662
rect 445772 679522 445800 680002
rect 445944 679924 445996 679930
rect 445944 679866 445996 679872
rect 445956 679522 445984 679866
rect 446232 679590 446260 680070
rect 446876 679946 446904 681119
rect 447152 681086 447180 682246
rect 447140 681080 447192 681086
rect 447140 681022 447192 681028
rect 446752 679918 446904 679946
rect 446956 679992 447008 679998
rect 446956 679934 447008 679940
rect 447704 679946 447732 682343
rect 449912 680218 449940 684014
rect 449912 680190 449986 680218
rect 446220 679584 446272 679590
rect 446220 679526 446272 679532
rect 432788 679516 433024 679522
rect 421472 679458 421524 679464
rect 432840 679510 432972 679516
rect 432788 679458 432840 679464
rect 432972 679458 433024 679464
rect 435824 679516 435876 679522
rect 435824 679458 435876 679464
rect 437940 679516 437992 679522
rect 437940 679458 437992 679464
rect 441712 679516 441764 679522
rect 441712 679458 441764 679464
rect 441804 679516 441856 679522
rect 441804 679458 441856 679464
rect 442356 679516 442408 679522
rect 442356 679458 442408 679464
rect 443920 679516 443972 679522
rect 443920 679458 443972 679464
rect 445760 679516 445812 679522
rect 445760 679458 445812 679464
rect 445944 679516 445996 679522
rect 446968 679504 446996 679934
rect 447704 679918 448040 679946
rect 449958 679932 449986 680190
rect 450280 679946 450308 685102
rect 453854 684584 453910 684593
rect 453854 684519 453910 684528
rect 453868 680218 453896 684519
rect 453822 680190 453896 680218
rect 450280 679918 450616 679946
rect 453822 679932 453850 680190
rect 454236 679946 454264 685238
rect 454774 685128 454830 685137
rect 454774 685063 454830 685072
rect 454788 679946 454816 685063
rect 456892 685024 456944 685030
rect 456892 684966 456944 684972
rect 456904 679946 456932 684966
rect 457364 679946 457392 687278
rect 476580 686112 476632 686118
rect 476580 686054 476632 686060
rect 470876 685364 470928 685370
rect 470876 685306 470928 685312
rect 467012 684888 467064 684894
rect 467012 684830 467064 684836
rect 458640 682440 458692 682446
rect 458640 682382 458692 682388
rect 458456 682168 458508 682174
rect 458456 682110 458508 682116
rect 454236 679918 454480 679946
rect 454788 679918 455124 679946
rect 456904 679918 457056 679946
rect 457364 679918 457700 679946
rect 458468 679674 458496 682110
rect 458652 679946 458680 682382
rect 463792 682372 463844 682378
rect 463792 682314 463844 682320
rect 462502 682272 462558 682281
rect 462502 682207 462558 682216
rect 461216 681216 461268 681222
rect 461216 681158 461268 681164
rect 461228 679946 461256 681158
rect 462516 679946 462544 682207
rect 463804 679946 463832 682314
rect 467024 679946 467052 684830
rect 470692 684140 470744 684146
rect 470692 684082 470744 684088
rect 468392 684004 468444 684010
rect 468392 683946 468444 683952
rect 468300 683732 468352 683738
rect 468300 683674 468352 683680
rect 468312 679946 468340 683674
rect 458652 679918 458988 679946
rect 461228 679918 461564 679946
rect 462516 679918 462852 679946
rect 463804 679918 464140 679946
rect 465540 679924 465592 679930
rect 466716 679918 467052 679946
rect 467104 679924 467156 679930
rect 465540 679866 465592 679872
rect 468004 679918 468340 679946
rect 468404 679946 468432 683946
rect 468404 679918 468648 679946
rect 467104 679866 467156 679872
rect 462412 679788 462464 679794
rect 462412 679730 462464 679736
rect 458344 679646 458496 679674
rect 462424 679522 462452 679730
rect 465552 679522 465580 679866
rect 466184 679856 466236 679862
rect 466184 679798 466236 679804
rect 466196 679522 466224 679798
rect 467116 679522 467144 679866
rect 470704 679810 470732 684082
rect 470888 679946 470916 685306
rect 472808 685024 472860 685030
rect 472808 684966 472860 684972
rect 472820 679946 472848 684966
rect 476120 683936 476172 683942
rect 476120 683878 476172 683884
rect 470888 679918 471224 679946
rect 472512 679918 472848 679946
rect 476132 679946 476160 683878
rect 476592 679946 476620 686054
rect 477512 682446 477540 702406
rect 484400 700732 484452 700738
rect 484400 700674 484452 700680
rect 484412 692774 484440 700674
rect 527192 700670 527220 703520
rect 543476 700738 543504 703520
rect 543464 700732 543516 700738
rect 543464 700674 543516 700680
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 559668 700602 559696 703520
rect 559656 700596 559708 700602
rect 559656 700538 559708 700544
rect 551376 700528 551428 700534
rect 551376 700470 551428 700476
rect 550272 698964 550324 698970
rect 550272 698906 550324 698912
rect 498200 694816 498252 694822
rect 498200 694758 498252 694764
rect 484412 692746 484992 692774
rect 480534 683632 480590 683641
rect 480534 683567 480590 683576
rect 477500 682440 477552 682446
rect 477500 682382 477552 682388
rect 480352 682236 480404 682242
rect 480352 682178 480404 682184
rect 476132 679918 476376 679946
rect 476592 679918 477020 679946
rect 480364 679810 480392 682178
rect 480548 679946 480576 683567
rect 484860 681080 484912 681086
rect 484860 681022 484912 681028
rect 484872 679946 484900 681022
rect 480548 679918 480884 679946
rect 484748 679918 484900 679946
rect 484964 679946 484992 692746
rect 487618 685264 487674 685273
rect 487618 685199 487674 685208
rect 487632 679946 487660 685199
rect 489550 685128 489606 685137
rect 489550 685063 489606 685072
rect 490012 685092 490064 685098
rect 488722 681048 488778 681057
rect 488722 680983 488778 680992
rect 484964 679918 485392 679946
rect 487324 679918 487660 679946
rect 467564 679788 467616 679794
rect 470580 679782 470732 679810
rect 480240 679782 480392 679810
rect 467564 679730 467616 679736
rect 467196 679652 467248 679658
rect 467196 679594 467248 679600
rect 467208 679538 467236 679594
rect 467208 679522 467512 679538
rect 467576 679522 467604 679730
rect 488736 679674 488764 680983
rect 489564 679946 489592 685063
rect 490012 685034 490064 685040
rect 489256 679918 489592 679946
rect 490024 679810 490052 685034
rect 497280 683868 497332 683874
rect 497280 683810 497332 683816
rect 496636 681148 496688 681154
rect 496636 681090 496688 681096
rect 495162 680504 495218 680513
rect 495162 680439 495218 680448
rect 495176 679946 495204 680439
rect 496648 679946 496676 681090
rect 495052 679918 495204 679946
rect 496340 679918 496676 679946
rect 497292 679946 497320 683810
rect 498212 680218 498240 694758
rect 550088 692096 550140 692102
rect 550088 692038 550140 692044
rect 538220 688016 538272 688022
rect 538220 687958 538272 687964
rect 504270 687304 504326 687313
rect 504270 687239 504326 687248
rect 499856 683800 499908 683806
rect 499856 683742 499908 683748
rect 499212 681760 499264 681766
rect 499212 681702 499264 681708
rect 498212 680190 498286 680218
rect 497292 679918 497628 679946
rect 498258 679932 498286 680190
rect 499224 679946 499252 681702
rect 498916 679918 499252 679946
rect 499868 679946 499896 683742
rect 502522 683360 502578 683369
rect 502522 683295 502578 683304
rect 502248 682372 502300 682378
rect 502248 682314 502300 682320
rect 500498 682136 500554 682145
rect 500498 682071 500554 682080
rect 500512 679946 500540 682071
rect 501788 681216 501840 681222
rect 501788 681158 501840 681164
rect 501800 679946 501828 681158
rect 502260 679946 502288 682314
rect 499868 679918 500204 679946
rect 500512 679918 500848 679946
rect 501492 679918 501828 679946
rect 502136 679918 502288 679946
rect 502536 679946 502564 683295
rect 504284 679946 504312 687239
rect 528836 685976 528888 685982
rect 528836 685918 528888 685924
rect 510528 685092 510580 685098
rect 510528 685034 510580 685040
rect 509514 683224 509570 683233
rect 509514 683159 509570 683168
rect 507584 682508 507636 682514
rect 507584 682450 507636 682456
rect 505098 680912 505154 680921
rect 505098 680847 505154 680856
rect 505112 679946 505140 680847
rect 507596 679946 507624 682450
rect 509332 682304 509384 682310
rect 509332 682246 509384 682252
rect 502536 679918 502780 679946
rect 504284 679918 504712 679946
rect 505112 679918 505356 679946
rect 507288 679918 507624 679946
rect 509344 679810 509372 682246
rect 509528 679946 509556 683159
rect 510540 680218 510568 685034
rect 523040 684956 523092 684962
rect 523040 684898 523092 684904
rect 521844 684820 521896 684826
rect 521844 684762 521896 684768
rect 517244 682304 517296 682310
rect 517244 682246 517296 682252
rect 512736 682236 512788 682242
rect 512736 682178 512788 682184
rect 511446 680912 511502 680921
rect 511446 680847 511502 680856
rect 510494 680190 510568 680218
rect 509528 679918 509864 679946
rect 510494 679932 510522 680190
rect 511460 679946 511488 680847
rect 512748 679946 512776 682178
rect 514758 681320 514814 681329
rect 514758 681255 514814 681264
rect 511152 679918 511488 679946
rect 512440 679918 512776 679946
rect 514772 679946 514800 681255
rect 517256 679946 517284 682246
rect 517520 681760 517572 681766
rect 517520 681702 517572 681708
rect 517532 681290 517560 681702
rect 517520 681284 517572 681290
rect 517520 681226 517572 681232
rect 518990 680776 519046 680785
rect 518990 680711 519046 680720
rect 514772 679918 515016 679946
rect 516948 679918 517284 679946
rect 519004 679810 519032 680711
rect 521856 679946 521884 684762
rect 523052 679946 523080 684898
rect 524880 683800 524932 683806
rect 524880 683742 524932 683748
rect 524892 679946 524920 683742
rect 526258 682408 526314 682417
rect 526258 682343 526314 682352
rect 524972 682100 525024 682106
rect 524972 682042 525024 682048
rect 521856 679918 522100 679946
rect 523052 679918 523388 679946
rect 524676 679918 524920 679946
rect 524984 679946 525012 682042
rect 526272 679946 526300 682343
rect 528742 682272 528798 682281
rect 528742 682207 528798 682216
rect 528756 679946 528784 682207
rect 524984 679918 525320 679946
rect 525964 679918 526300 679946
rect 528540 679918 528784 679946
rect 528848 679946 528876 685918
rect 535460 684752 535512 684758
rect 535460 684694 535512 684700
rect 529664 682780 529716 682786
rect 529664 682722 529716 682728
rect 528848 679918 529184 679946
rect 489900 679782 490052 679810
rect 509220 679782 509372 679810
rect 518880 679782 519032 679810
rect 473464 679658 473800 679674
rect 473452 679652 473800 679658
rect 473504 679646 473800 679652
rect 488612 679646 488764 679674
rect 529676 679674 529704 682722
rect 530122 682544 530178 682553
rect 530122 682479 530178 682488
rect 530136 679946 530164 682479
rect 531226 682136 531282 682145
rect 531226 682071 531282 682080
rect 531240 679946 531268 682071
rect 534080 681964 534132 681970
rect 534080 681906 534132 681912
rect 535276 681964 535328 681970
rect 535276 681906 535328 681912
rect 532698 681456 532754 681465
rect 532698 681391 532754 681400
rect 530136 679918 530472 679946
rect 531116 679918 531268 679946
rect 532712 679946 532740 681391
rect 534092 679946 534120 681906
rect 535288 679946 535316 681906
rect 532712 679918 533048 679946
rect 534092 679918 534336 679946
rect 534980 679918 535316 679946
rect 535472 679946 535500 684694
rect 537852 681828 537904 681834
rect 537852 681770 537904 681776
rect 537864 679946 537892 681770
rect 538232 680218 538260 687958
rect 545578 684720 545634 684729
rect 539140 684684 539192 684690
rect 545578 684655 545634 684664
rect 539140 684626 539192 684632
rect 535472 679918 535624 679946
rect 537556 679918 537892 679946
rect 538186 680190 538260 680218
rect 538186 679932 538214 680190
rect 539152 679946 539180 684626
rect 545118 682680 545174 682689
rect 545118 682615 545174 682624
rect 541716 681760 541768 681766
rect 541716 681702 541768 681708
rect 541728 679946 541756 681702
rect 539152 679918 539488 679946
rect 541420 679918 541756 679946
rect 545132 679946 545160 682615
rect 545592 679946 545620 684655
rect 546960 682644 547012 682650
rect 546960 682586 547012 682592
rect 546866 682000 546922 682009
rect 546866 681935 546922 681944
rect 546880 679946 546908 681935
rect 545132 679918 545284 679946
rect 545592 679918 545928 679946
rect 546572 679918 546908 679946
rect 546972 679946 547000 682586
rect 549444 682100 549496 682106
rect 549444 682042 549496 682048
rect 548798 681864 548854 681873
rect 548798 681799 548854 681808
rect 548812 679946 548840 681799
rect 549456 679946 549484 682042
rect 549996 682032 550048 682038
rect 549996 681974 550048 681980
rect 550008 679946 550036 681974
rect 546972 679918 547216 679946
rect 548504 679918 548840 679946
rect 549148 679918 549484 679946
rect 549792 679918 550036 679946
rect 529676 679646 529828 679674
rect 473452 679594 473504 679600
rect 447094 679516 447146 679522
rect 446968 679476 447094 679504
rect 445944 679458 445996 679464
rect 447094 679458 447146 679464
rect 462412 679516 462464 679522
rect 462412 679458 462464 679464
rect 465540 679516 465592 679522
rect 465540 679458 465592 679464
rect 466184 679516 466236 679522
rect 466184 679458 466236 679464
rect 467104 679516 467156 679522
rect 467208 679516 467524 679522
rect 467208 679510 467472 679516
rect 467104 679458 467156 679464
rect 467472 679458 467524 679464
rect 467564 679516 467616 679522
rect 467564 679458 467616 679464
rect 409878 665136 409934 665145
rect 409878 665071 409934 665080
rect 550100 378865 550128 692038
rect 550180 682576 550232 682582
rect 550180 682518 550232 682524
rect 550192 564505 550220 682518
rect 550178 564496 550234 564505
rect 550178 564431 550234 564440
rect 550178 459776 550234 459785
rect 550178 459711 550234 459720
rect 550086 378856 550142 378865
rect 550086 378791 550142 378800
rect 409786 334656 409842 334665
rect 409786 334591 409842 334600
rect 409878 319696 409934 319705
rect 409878 319631 409934 319640
rect 409786 316976 409842 316985
rect 409786 316911 409842 316920
rect 409696 233776 409748 233782
rect 409696 233718 409748 233724
rect 409800 156466 409828 316911
rect 409892 203658 409920 319631
rect 550086 297936 550142 297945
rect 550086 297871 550142 297880
rect 410156 240644 410208 240650
rect 410156 240586 410208 240592
rect 537668 240644 537720 240650
rect 537668 240586 537720 240592
rect 410030 239850 410058 240108
rect 410030 239822 410104 239850
rect 409972 233844 410024 233850
rect 409972 233786 410024 233792
rect 409880 203652 409932 203658
rect 409880 203594 409932 203600
rect 409984 187202 410012 233786
rect 410076 204950 410104 239822
rect 410064 204944 410116 204950
rect 410064 204886 410116 204892
rect 409972 187196 410024 187202
rect 409972 187138 410024 187144
rect 410168 162042 410196 240586
rect 410338 240408 410394 240417
rect 410260 240366 410338 240394
rect 410260 230353 410288 240366
rect 410338 240343 410394 240352
rect 410352 240094 410688 240122
rect 410352 233850 410380 240094
rect 411318 239850 411346 240108
rect 412620 240094 412772 240122
rect 413264 240094 413600 240122
rect 414552 240094 414888 240122
rect 416484 240094 416728 240122
rect 411318 239822 411392 239850
rect 410340 233844 410392 233850
rect 410340 233786 410392 233792
rect 410246 230344 410302 230353
rect 410246 230279 410302 230288
rect 411364 202162 411392 239822
rect 411628 227384 411680 227390
rect 411628 227326 411680 227332
rect 411352 202156 411404 202162
rect 411352 202098 411404 202104
rect 410156 162036 410208 162042
rect 410156 161978 410208 161984
rect 409788 156460 409840 156466
rect 409788 156402 409840 156408
rect 409604 152720 409656 152726
rect 409604 152662 409656 152668
rect 410340 152380 410392 152386
rect 410340 152322 410392 152328
rect 409144 152312 409196 152318
rect 409144 152254 409196 152260
rect 410352 149940 410380 152322
rect 411640 149940 411668 227326
rect 412744 198393 412772 240094
rect 413572 237454 413600 240094
rect 414860 238066 414888 240094
rect 416700 238542 416728 240094
rect 416976 240094 417128 240122
rect 420012 240094 420348 240122
rect 420992 240094 421328 240122
rect 416688 238536 416740 238542
rect 416688 238478 416740 238484
rect 414848 238060 414900 238066
rect 414848 238002 414900 238008
rect 416700 237998 416728 238478
rect 416688 237992 416740 237998
rect 416688 237934 416740 237940
rect 413560 237448 413612 237454
rect 413560 237390 413612 237396
rect 414020 237448 414072 237454
rect 414020 237390 414072 237396
rect 413560 229628 413612 229634
rect 413560 229570 413612 229576
rect 412730 198384 412786 198393
rect 412730 198319 412786 198328
rect 412730 195392 412786 195401
rect 412730 195327 412786 195336
rect 412744 149954 412772 195327
rect 412744 149926 412942 149954
rect 413572 149940 413600 229570
rect 414032 151366 414060 237390
rect 416780 232484 416832 232490
rect 416780 232426 416832 232432
rect 414664 202904 414716 202910
rect 414664 202846 414716 202852
rect 414676 161974 414704 202846
rect 414664 161968 414716 161974
rect 414664 161910 414716 161916
rect 414848 152448 414900 152454
rect 414848 152390 414900 152396
rect 414020 151360 414072 151366
rect 414020 151302 414072 151308
rect 414860 149940 414888 152390
rect 416792 149940 416820 232426
rect 416976 210458 417004 240094
rect 417424 236700 417476 236706
rect 417424 236642 417476 236648
rect 416964 210452 417016 210458
rect 416964 210394 417016 210400
rect 417436 149940 417464 236642
rect 420012 233850 420040 240094
rect 421300 238134 421328 240094
rect 422588 240094 422924 240122
rect 423048 240094 423568 240122
rect 426452 240094 426788 240122
rect 426912 240094 427432 240122
rect 427832 240094 428076 240122
rect 428384 240094 428720 240122
rect 431940 240094 432092 240122
rect 422588 238202 422616 240094
rect 422576 238196 422628 238202
rect 422576 238138 422628 238144
rect 421288 238128 421340 238134
rect 421288 238070 421340 238076
rect 418804 233844 418856 233850
rect 418804 233786 418856 233792
rect 420000 233844 420052 233850
rect 420000 233786 420052 233792
rect 418068 225684 418120 225690
rect 418068 225626 418120 225632
rect 418080 149940 418108 225626
rect 418816 204270 418844 233786
rect 421932 231124 421984 231130
rect 421932 231066 421984 231072
rect 418804 204264 418856 204270
rect 418804 204206 418856 204212
rect 420000 161968 420052 161974
rect 420000 161910 420052 161916
rect 419356 152312 419408 152318
rect 419356 152254 419408 152260
rect 419368 149940 419396 152254
rect 420012 149940 420040 161910
rect 421944 149940 421972 231066
rect 423048 219434 423076 240094
rect 423588 238196 423640 238202
rect 423588 238138 423640 238144
rect 423600 237930 423628 238138
rect 423588 237924 423640 237930
rect 423588 237866 423640 237872
rect 422312 219406 423076 219434
rect 422312 198529 422340 219406
rect 422298 198520 422354 198529
rect 422298 198455 422354 198464
rect 426452 159254 426480 240094
rect 426912 219434 426940 240094
rect 427832 238814 427860 240094
rect 427820 238808 427872 238814
rect 427820 238750 427872 238756
rect 428384 238270 428412 240094
rect 428372 238264 428424 238270
rect 428372 238206 428424 238212
rect 430304 235544 430356 235550
rect 430304 235486 430356 235492
rect 429200 231192 429252 231198
rect 429200 231134 429252 231140
rect 426544 219406 426940 219434
rect 426544 188358 426572 219406
rect 426532 188352 426584 188358
rect 426532 188294 426584 188300
rect 427082 187096 427138 187105
rect 427082 187031 427138 187040
rect 426440 159248 426492 159254
rect 426440 159190 426492 159196
rect 425152 153128 425204 153134
rect 425152 153070 425204 153076
rect 425164 149940 425192 153070
rect 427096 149940 427124 187031
rect 429212 149954 429240 231134
rect 429212 149926 429686 149954
rect 430316 149940 430344 235486
rect 431224 212560 431276 212566
rect 431224 212502 431276 212508
rect 431236 177478 431264 212502
rect 431224 177472 431276 177478
rect 431224 177414 431276 177420
rect 432064 170406 432092 240094
rect 432248 240094 432584 240122
rect 433352 240094 434516 240122
rect 436448 240094 436784 240122
rect 432248 238474 432276 240094
rect 432236 238468 432288 238474
rect 432236 238410 432288 238416
rect 433352 211818 433380 240094
rect 436756 238814 436784 240094
rect 438872 240094 439024 240122
rect 436744 238808 436796 238814
rect 436744 238750 436796 238756
rect 436744 234524 436796 234530
rect 436744 234466 436796 234472
rect 435456 225752 435508 225758
rect 435456 225694 435508 225700
rect 433340 211812 433392 211818
rect 433340 211754 433392 211760
rect 432052 170400 432104 170406
rect 432052 170342 432104 170348
rect 434168 153196 434220 153202
rect 434168 153138 434220 153144
rect 434180 149940 434208 153138
rect 435468 149940 435496 225694
rect 436756 149940 436784 234466
rect 438676 217388 438728 217394
rect 438676 217330 438728 217336
rect 438688 149940 438716 217330
rect 438872 167890 438900 240094
rect 440298 239850 440326 240108
rect 440252 239822 440326 239850
rect 442552 240094 442888 240122
rect 443656 240094 444176 240122
rect 444820 240094 445156 240122
rect 446752 240094 447088 240122
rect 440252 238610 440280 239822
rect 440240 238604 440292 238610
rect 440240 238546 440292 238552
rect 442552 238338 442580 240094
rect 442540 238332 442592 238338
rect 442540 238274 442592 238280
rect 443656 219434 443684 240094
rect 445128 238474 445156 240094
rect 447060 238610 447088 240094
rect 449912 240094 450616 240122
rect 451384 240094 451904 240122
rect 447048 238604 447100 238610
rect 447048 238546 447100 238552
rect 445116 238468 445168 238474
rect 445116 238410 445168 238416
rect 444472 231260 444524 231266
rect 444472 231202 444524 231208
rect 443012 219406 443684 219434
rect 441620 210520 441672 210526
rect 441620 210462 441672 210468
rect 439320 169176 439372 169182
rect 439320 169118 439372 169124
rect 438860 167884 438912 167890
rect 438860 167826 438912 167832
rect 439332 149940 439360 169118
rect 440606 155680 440662 155689
rect 440606 155615 440662 155624
rect 440620 149940 440648 155615
rect 441632 149954 441660 210462
rect 443012 184210 443040 219406
rect 443000 184204 443052 184210
rect 443000 184146 443052 184152
rect 443184 176112 443236 176118
rect 443184 176054 443236 176060
rect 441632 149926 441922 149954
rect 443196 149940 443224 176054
rect 444484 149940 444512 231202
rect 448336 227316 448388 227322
rect 448336 227258 448388 227264
rect 445760 222896 445812 222902
rect 445760 222838 445812 222844
rect 445772 149954 445800 222838
rect 447690 153096 447746 153105
rect 447690 153031 447746 153040
rect 445772 149926 446430 149954
rect 447704 149940 447732 153031
rect 448348 149940 448376 227258
rect 449912 194138 449940 240094
rect 451384 219434 451412 240094
rect 452534 239850 452562 240108
rect 453192 240094 453528 240122
rect 452534 239822 452608 239850
rect 452580 232490 452608 239822
rect 453500 234598 453528 240094
rect 454144 240094 454480 240122
rect 454604 240094 455124 240122
rect 456412 240094 456748 240122
rect 457056 240094 457392 240122
rect 454144 238406 454172 240094
rect 454132 238400 454184 238406
rect 454132 238342 454184 238348
rect 453488 234592 453540 234598
rect 453488 234534 453540 234540
rect 452568 232484 452620 232490
rect 452568 232426 452620 232432
rect 454604 219434 454632 240094
rect 456720 234462 456748 240094
rect 457364 238406 457392 240094
rect 458192 240094 458344 240122
rect 457444 239012 457496 239018
rect 457444 238954 457496 238960
rect 457352 238400 457404 238406
rect 457352 238342 457404 238348
rect 456708 234456 456760 234462
rect 456708 234398 456760 234404
rect 451292 219406 451412 219434
rect 454144 219406 454632 219434
rect 449900 194132 449952 194138
rect 449900 194074 449952 194080
rect 451292 153746 451320 219406
rect 452842 195256 452898 195265
rect 452842 195191 452898 195200
rect 451280 153740 451332 153746
rect 451280 153682 451332 153688
rect 448980 153060 449032 153066
rect 448980 153002 449032 153008
rect 448992 149940 449020 153002
rect 452856 149940 452884 195191
rect 453486 192672 453542 192681
rect 453486 192607 453542 192616
rect 453500 149940 453528 192607
rect 454144 159662 454172 219406
rect 454132 159656 454184 159662
rect 454132 159598 454184 159604
rect 457456 152454 457484 238954
rect 458192 238513 458220 240094
rect 459618 239850 459646 240108
rect 459572 239822 459646 239850
rect 460906 239850 460934 240108
rect 461044 240094 461564 240122
rect 462332 240094 462852 240122
rect 463160 240094 463496 240122
rect 463712 240094 464140 240122
rect 465092 240094 465428 240122
rect 467852 240094 468004 240122
rect 468128 240094 468648 240122
rect 460906 239822 460980 239850
rect 458178 238504 458234 238513
rect 458178 238439 458234 238448
rect 458178 185736 458234 185745
rect 458178 185671 458234 185680
rect 457444 152448 457496 152454
rect 457444 152390 457496 152396
rect 458192 149954 458220 185671
rect 458192 149926 458666 149954
rect 459572 149938 459600 239822
rect 460952 232422 460980 239822
rect 460940 232416 460992 232422
rect 460940 232358 460992 232364
rect 459928 227248 459980 227254
rect 459928 227190 459980 227196
rect 459940 149940 459968 227190
rect 461044 219434 461072 240094
rect 461216 233844 461268 233850
rect 461216 233786 461268 233792
rect 460952 219406 461072 219434
rect 460570 184376 460626 184385
rect 460570 184311 460626 184320
rect 460584 149940 460612 184311
rect 460952 151230 460980 219406
rect 460940 151224 460992 151230
rect 460940 151166 460992 151172
rect 461228 149940 461256 233786
rect 462332 170406 462360 240094
rect 463160 238950 463188 240094
rect 463148 238944 463200 238950
rect 463148 238886 463200 238892
rect 463712 197130 463740 240094
rect 463700 197124 463752 197130
rect 463700 197066 463752 197072
rect 465092 195906 465120 240094
rect 465080 195900 465132 195906
rect 465080 195842 465132 195848
rect 462320 170400 462372 170406
rect 462320 170342 462372 170348
rect 467852 169250 467880 240094
rect 468128 219434 468156 240094
rect 469278 239850 469306 240108
rect 467944 219406 468156 219434
rect 469232 239822 469306 239850
rect 470566 239850 470594 240108
rect 470704 240094 471224 240122
rect 472512 240094 472664 240122
rect 470566 239822 470640 239850
rect 467944 198830 467972 219406
rect 467932 198824 467984 198830
rect 467932 198766 467984 198772
rect 468300 179376 468352 179382
rect 468300 179318 468352 179324
rect 467840 169244 467892 169250
rect 467840 169186 467892 169192
rect 463790 152960 463846 152969
rect 463790 152895 463846 152904
rect 463804 149940 463832 152895
rect 468312 149940 468340 179318
rect 469232 163674 469260 239822
rect 470612 238338 470640 239822
rect 470600 238332 470652 238338
rect 470600 238274 470652 238280
rect 470704 219434 470732 240094
rect 472636 238270 472664 240094
rect 472728 240094 473156 240122
rect 474444 240094 474688 240122
rect 472624 238264 472676 238270
rect 472624 238206 472676 238212
rect 472072 228404 472124 228410
rect 472072 228346 472124 228352
rect 470612 219406 470732 219434
rect 470612 187134 470640 219406
rect 470600 187128 470652 187134
rect 470600 187070 470652 187076
rect 470232 163804 470284 163810
rect 470232 163746 470284 163752
rect 469220 163668 469272 163674
rect 469220 163610 469272 163616
rect 470244 149940 470272 163746
rect 472084 149954 472112 228346
rect 472728 219434 472756 240094
rect 474660 235822 474688 240094
rect 474752 240094 475088 240122
rect 474648 235816 474700 235822
rect 474648 235758 474700 235764
rect 472808 233708 472860 233714
rect 472808 233650 472860 233656
rect 472176 219406 472756 219434
rect 472176 164898 472204 219406
rect 472164 164892 472216 164898
rect 472164 164834 472216 164840
rect 459560 149932 459612 149938
rect 403164 149874 403216 149880
rect 472084 149926 472190 149954
rect 472820 149940 472848 233650
rect 474648 150068 474700 150074
rect 474648 150010 474700 150016
rect 474660 149938 474688 150010
rect 474752 149938 474780 240094
rect 476362 239850 476390 240108
rect 476500 240094 477020 240122
rect 476362 239822 476436 239850
rect 476408 238202 476436 239822
rect 476396 238196 476448 238202
rect 476396 238138 476448 238144
rect 476500 219434 476528 240094
rect 477650 239850 477678 240108
rect 478938 239850 478966 240108
rect 480240 240094 480392 240122
rect 477604 239822 477678 239850
rect 478892 239822 478966 239850
rect 476672 224324 476724 224330
rect 476672 224266 476724 224272
rect 476224 219406 476528 219434
rect 476028 202156 476080 202162
rect 476028 202098 476080 202104
rect 476040 149940 476068 202098
rect 476224 197198 476252 219406
rect 476212 197192 476264 197198
rect 476212 197134 476264 197140
rect 476684 149940 476712 224266
rect 477604 217394 477632 239822
rect 478604 236564 478656 236570
rect 478604 236506 478656 236512
rect 477960 222964 478012 222970
rect 477960 222906 478012 222912
rect 477592 217388 477644 217394
rect 477592 217330 477644 217336
rect 477972 149940 478000 222906
rect 478616 149940 478644 236506
rect 478892 193050 478920 239822
rect 478880 193044 478932 193050
rect 478880 192986 478932 192992
rect 480364 190262 480392 240094
rect 481514 239850 481542 240108
rect 483124 240094 483460 240122
rect 483768 240094 484104 240122
rect 484872 240094 485392 240122
rect 487448 240094 487968 240122
rect 481514 239822 481588 239850
rect 481560 235754 481588 239822
rect 482928 237924 482980 237930
rect 482928 237866 482980 237872
rect 482940 237454 482968 237866
rect 482928 237448 482980 237454
rect 482928 237390 482980 237396
rect 481548 235748 481600 235754
rect 481548 235690 481600 235696
rect 481180 218748 481232 218754
rect 481180 218690 481232 218696
rect 480352 190256 480404 190262
rect 480352 190198 480404 190204
rect 480536 175976 480588 175982
rect 480536 175918 480588 175924
rect 480076 150068 480128 150074
rect 480076 150010 480128 150016
rect 480088 149938 480116 150010
rect 480548 149940 480576 175918
rect 481192 149940 481220 218690
rect 481824 156596 481876 156602
rect 481824 156538 481876 156544
rect 481836 149940 481864 156538
rect 482940 153066 482968 237390
rect 483124 159458 483152 240094
rect 483768 237454 483796 240094
rect 483756 237448 483808 237454
rect 483756 237390 483808 237396
rect 484872 219434 484900 240094
rect 486976 231124 487028 231130
rect 486976 231066 487028 231072
rect 485044 224392 485096 224398
rect 485044 224334 485096 224340
rect 484412 219406 484900 219434
rect 483112 159452 483164 159458
rect 483112 159394 483164 159400
rect 484412 158438 484440 219406
rect 484400 158432 484452 158438
rect 484400 158374 484452 158380
rect 482928 153060 482980 153066
rect 482928 153002 482980 153008
rect 482466 152824 482522 152833
rect 482466 152759 482522 152768
rect 482480 149940 482508 152759
rect 485056 149940 485084 224334
rect 486988 149940 487016 231066
rect 487448 219434 487476 240094
rect 488598 239850 488626 240108
rect 488736 240094 489256 240122
rect 488598 239822 488672 239850
rect 488644 235142 488672 239822
rect 488632 235136 488684 235142
rect 488632 235078 488684 235084
rect 488736 219434 488764 240094
rect 490530 239850 490558 240108
rect 491174 239850 491202 240108
rect 492048 240094 492476 240122
rect 496832 240094 496984 240122
rect 497628 240094 497964 240122
rect 490530 239822 490604 239850
rect 491174 239822 491248 239850
rect 490576 237998 490604 239822
rect 490564 237992 490616 237998
rect 490564 237934 490616 237940
rect 491116 237992 491168 237998
rect 491116 237934 491168 237940
rect 491128 232354 491156 237934
rect 491220 235074 491248 239822
rect 491208 235068 491260 235074
rect 491208 235010 491260 235016
rect 491300 233776 491352 233782
rect 491300 233718 491352 233724
rect 491116 232348 491168 232354
rect 491116 232290 491168 232296
rect 487172 219406 487476 219434
rect 488552 219406 488764 219434
rect 487172 197742 487200 219406
rect 487160 197736 487212 197742
rect 487160 197678 487212 197684
rect 488552 155553 488580 219406
rect 488906 167648 488962 167657
rect 488906 167583 488962 167592
rect 488538 155544 488594 155553
rect 488538 155479 488594 155488
rect 488920 149940 488948 167583
rect 490194 164928 490250 164937
rect 490194 164863 490250 164872
rect 490208 149940 490236 164863
rect 491312 153134 491340 233718
rect 492048 219434 492076 240094
rect 493416 235204 493468 235210
rect 493416 235146 493468 235152
rect 491404 219406 492076 219434
rect 491404 198422 491432 219406
rect 491392 198416 491444 198422
rect 491392 198358 491444 198364
rect 492770 180296 492826 180305
rect 492770 180231 492826 180240
rect 491300 153128 491352 153134
rect 491300 153070 491352 153076
rect 492128 153128 492180 153134
rect 492128 153070 492180 153076
rect 492140 149940 492168 153070
rect 492784 149940 492812 180231
rect 493428 149940 493456 235146
rect 496832 231130 496860 240094
rect 497936 238542 497964 240094
rect 498212 240094 498916 240122
rect 500328 240094 500848 240122
rect 501492 240094 501828 240122
rect 497924 238536 497976 238542
rect 497924 238478 497976 238484
rect 496820 231124 496872 231130
rect 496820 231066 496872 231072
rect 494060 220108 494112 220114
rect 494060 220050 494112 220056
rect 494072 149940 494100 220050
rect 497924 207664 497976 207670
rect 497924 207606 497976 207612
rect 497278 182880 497334 182889
rect 497278 182815 497334 182824
rect 495440 173188 495492 173194
rect 495440 173130 495492 173136
rect 495452 150278 495480 173130
rect 495440 150272 495492 150278
rect 495440 150214 495492 150220
rect 496636 150272 496688 150278
rect 496636 150214 496688 150220
rect 496648 149940 496676 150214
rect 497292 149940 497320 182815
rect 497936 149940 497964 207606
rect 498212 153134 498240 240094
rect 499212 236496 499264 236502
rect 499212 236438 499264 236444
rect 498200 153128 498252 153134
rect 498200 153070 498252 153076
rect 498566 152688 498622 152697
rect 498566 152623 498622 152632
rect 498580 149940 498608 152623
rect 499224 149940 499252 236438
rect 500328 219434 500356 240094
rect 501800 237998 501828 240094
rect 504376 240094 504712 240122
rect 505356 240094 505692 240122
rect 504376 238882 504404 240094
rect 505664 238882 505692 240094
rect 506630 239850 506658 240108
rect 506768 240094 507288 240122
rect 506630 239822 506704 239850
rect 506676 238950 506704 239822
rect 506664 238944 506716 238950
rect 506664 238886 506716 238892
rect 504364 238876 504416 238882
rect 504364 238818 504416 238824
rect 505652 238876 505704 238882
rect 505652 238818 505704 238824
rect 501788 237992 501840 237998
rect 501788 237934 501840 237940
rect 506768 219434 506796 240094
rect 507918 239850 507946 240108
rect 499592 219406 500356 219434
rect 506492 219406 506796 219434
rect 507872 239822 507946 239850
rect 509206 239850 509234 240108
rect 509344 240094 509864 240122
rect 514772 240094 515016 240122
rect 515324 240094 515660 240122
rect 509206 239822 509280 239850
rect 499592 152386 499620 219406
rect 500224 204944 500276 204950
rect 500224 204886 500276 204892
rect 500236 153202 500264 204886
rect 503720 203652 503772 203658
rect 503720 203594 503772 203600
rect 502430 162072 502486 162081
rect 502430 162007 502486 162016
rect 500224 153196 500276 153202
rect 500224 153138 500276 153144
rect 499856 152448 499908 152454
rect 499856 152390 499908 152396
rect 499580 152380 499632 152386
rect 499580 152322 499632 152328
rect 499868 149940 499896 152390
rect 502444 149940 502472 162007
rect 503076 152448 503128 152454
rect 503076 152390 503128 152396
rect 503088 149940 503116 152390
rect 503732 149940 503760 203594
rect 506492 192506 506520 219406
rect 507872 200802 507900 239822
rect 509252 238785 509280 239822
rect 509238 238776 509294 238785
rect 509238 238711 509294 238720
rect 509344 229634 509372 240094
rect 514772 236638 514800 240094
rect 515324 237862 515352 240094
rect 518866 239850 518894 240108
rect 519096 240094 519524 240122
rect 518866 239822 518940 239850
rect 515312 237856 515364 237862
rect 515312 237798 515364 237804
rect 514760 236632 514812 236638
rect 514760 236574 514812 236580
rect 511448 235612 511500 235618
rect 511448 235554 511500 235560
rect 509332 229628 509384 229634
rect 509332 229570 509384 229576
rect 508504 227248 508556 227254
rect 508504 227190 508556 227196
rect 507860 200796 507912 200802
rect 507860 200738 507912 200744
rect 506480 192500 506532 192506
rect 506480 192442 506532 192448
rect 508228 184204 508280 184210
rect 508228 184146 508280 184152
rect 506940 173324 506992 173330
rect 506940 173266 506992 173272
rect 506296 156936 506348 156942
rect 506296 156878 506348 156884
rect 505652 152312 505704 152318
rect 505652 152254 505704 152260
rect 505664 149940 505692 152254
rect 506308 149940 506336 156878
rect 506952 149940 506980 173266
rect 507584 153196 507636 153202
rect 507584 153138 507636 153144
rect 507676 153196 507728 153202
rect 507676 153138 507728 153144
rect 507596 149940 507624 153138
rect 507688 152386 507716 153138
rect 507676 152380 507728 152386
rect 507676 152322 507728 152328
rect 508240 149940 508268 184146
rect 508516 152318 508544 227190
rect 510160 161016 510212 161022
rect 510160 160958 510212 160964
rect 508504 152312 508556 152318
rect 508504 152254 508556 152260
rect 510172 149940 510200 160958
rect 511460 149940 511488 235554
rect 512092 214600 512144 214606
rect 512092 214542 512144 214548
rect 512104 149940 512132 214542
rect 514024 177472 514076 177478
rect 514024 177414 514076 177420
rect 514036 149940 514064 177414
rect 518912 153678 518940 239822
rect 519096 194410 519124 240094
rect 520154 239850 520182 240108
rect 524032 240094 524368 240122
rect 525320 240094 525656 240122
rect 527896 240094 528232 240122
rect 528540 240094 528784 240122
rect 520154 239822 520228 239850
rect 520200 238377 520228 239822
rect 520186 238368 520242 238377
rect 520186 238303 520242 238312
rect 524340 235618 524368 240094
rect 525628 238513 525656 240094
rect 525614 238504 525670 238513
rect 525614 238439 525670 238448
rect 528204 237930 528232 240094
rect 528192 237924 528244 237930
rect 528192 237866 528244 237872
rect 528756 235686 528784 240094
rect 528848 240094 529184 240122
rect 528848 238678 528876 240094
rect 529814 239850 529842 240108
rect 529952 240094 531116 240122
rect 531884 240094 532404 240122
rect 532712 240094 533048 240122
rect 534980 240094 535316 240122
rect 529814 239822 529888 239850
rect 528836 238672 528888 238678
rect 528836 238614 528888 238620
rect 529860 237658 529888 239822
rect 529848 237652 529900 237658
rect 529848 237594 529900 237600
rect 527548 235680 527600 235686
rect 527548 235622 527600 235628
rect 528744 235680 528796 235686
rect 528744 235622 528796 235628
rect 524328 235612 524380 235618
rect 524328 235554 524380 235560
rect 525800 225616 525852 225622
rect 525800 225558 525852 225564
rect 521660 221468 521712 221474
rect 521660 221410 521712 221416
rect 519176 207732 519228 207738
rect 519176 207674 519228 207680
rect 519084 194404 519136 194410
rect 519084 194346 519136 194352
rect 518900 153672 518952 153678
rect 518900 153614 518952 153620
rect 515036 150068 515088 150074
rect 515036 150010 515088 150016
rect 515048 149938 515076 150010
rect 519188 149940 519216 207674
rect 519820 182844 519872 182850
rect 519820 182786 519872 182792
rect 519832 149940 519860 182786
rect 521672 149954 521700 221410
rect 524972 213308 525024 213314
rect 524972 213250 525024 213256
rect 523038 206272 523094 206281
rect 523038 206207 523094 206216
rect 474648 149932 474700 149938
rect 459560 149874 459612 149880
rect 474648 149874 474700 149880
rect 474740 149932 474792 149938
rect 474740 149874 474792 149880
rect 480076 149932 480128 149938
rect 480076 149874 480128 149880
rect 515036 149932 515088 149938
rect 521672 149926 521778 149954
rect 523052 149940 523080 206207
rect 524984 149940 525012 213250
rect 525812 149954 525840 225558
rect 525812 149926 526286 149954
rect 527560 149940 527588 235622
rect 529952 192982 529980 240094
rect 531884 219434 531912 240094
rect 532056 238672 532108 238678
rect 532056 238614 532108 238620
rect 531332 219406 531912 219434
rect 531332 193225 531360 219406
rect 531318 193216 531374 193225
rect 531318 193151 531374 193160
rect 529940 192976 529992 192982
rect 529940 192918 529992 192924
rect 528836 169040 528888 169046
rect 528836 168982 528888 168988
rect 528848 149940 528876 168982
rect 529940 158024 529992 158030
rect 529940 157966 529992 157972
rect 529204 152992 529256 152998
rect 529204 152934 529256 152940
rect 529216 152454 529244 152934
rect 529204 152448 529256 152454
rect 529204 152390 529256 152396
rect 529952 149954 529980 157966
rect 531412 152992 531464 152998
rect 531412 152934 531464 152940
rect 529952 149926 530150 149954
rect 531424 149940 531452 152934
rect 532068 149940 532096 238614
rect 532712 236774 532740 240094
rect 535288 239018 535316 240094
rect 536898 239850 536926 240108
rect 536852 239822 536926 239850
rect 535276 239012 535328 239018
rect 535276 238954 535328 238960
rect 532700 236768 532752 236774
rect 532700 236710 532752 236716
rect 536852 229294 536880 239822
rect 537482 239456 537538 239465
rect 537482 239391 537538 239400
rect 534724 229288 534776 229294
rect 534724 229230 534776 229236
rect 536840 229288 536892 229294
rect 536840 229230 536892 229236
rect 534736 152998 534764 229230
rect 535920 213240 535972 213246
rect 535920 213182 535972 213188
rect 534724 152992 534776 152998
rect 534724 152934 534776 152940
rect 534632 152448 534684 152454
rect 534632 152390 534684 152396
rect 534644 149940 534672 152390
rect 535932 149940 535960 213182
rect 536104 207120 536156 207126
rect 536104 207062 536156 207068
rect 536116 151230 536144 207062
rect 536840 159860 536892 159866
rect 536840 159802 536892 159808
rect 536852 152386 536880 159802
rect 537496 152454 537524 239391
rect 537574 237960 537630 237969
rect 537574 237895 537630 237904
rect 537588 152998 537616 237895
rect 537576 152992 537628 152998
rect 537576 152934 537628 152940
rect 537484 152448 537536 152454
rect 537484 152390 537536 152396
rect 536840 152380 536892 152386
rect 536840 152322 536892 152328
rect 537680 151366 537708 240586
rect 549996 240304 550048 240310
rect 549996 240246 550048 240252
rect 549260 240236 549312 240242
rect 549260 240178 549312 240184
rect 542372 240094 543352 240122
rect 543996 240094 544240 240122
rect 541164 238060 541216 238066
rect 541164 238002 541216 238008
rect 540242 234288 540298 234297
rect 540242 234223 540298 234232
rect 538864 232960 538916 232966
rect 538864 232902 538916 232908
rect 537760 203584 537812 203590
rect 537760 203526 537812 203532
rect 537668 151360 537720 151366
rect 537668 151302 537720 151308
rect 536104 151224 536156 151230
rect 536104 151166 536156 151172
rect 537772 150006 537800 203526
rect 537852 162512 537904 162518
rect 537852 162454 537904 162460
rect 537864 152454 537892 162454
rect 537942 158672 537998 158681
rect 537942 158607 537998 158616
rect 537852 152448 537904 152454
rect 537852 152390 537904 152396
rect 537956 150074 537984 158607
rect 538876 150482 538904 232902
rect 538956 180124 539008 180130
rect 538956 180066 539008 180072
rect 538864 150476 538916 150482
rect 538864 150418 538916 150424
rect 538862 150376 538918 150385
rect 538862 150311 538918 150320
rect 537944 150068 537996 150074
rect 537944 150010 537996 150016
rect 537760 150000 537812 150006
rect 537760 149942 537812 149948
rect 538876 149938 538904 150311
rect 538968 149938 538996 180066
rect 539968 177404 540020 177410
rect 539968 177346 540020 177352
rect 539782 173224 539838 173233
rect 539782 173159 539838 173168
rect 539048 162240 539100 162246
rect 539048 162182 539100 162188
rect 539060 150414 539088 162182
rect 539232 162104 539284 162110
rect 539232 162046 539284 162052
rect 539048 150408 539100 150414
rect 539048 150350 539100 150356
rect 539244 150249 539272 162046
rect 539324 162036 539376 162042
rect 539324 161978 539376 161984
rect 539230 150240 539286 150249
rect 539230 150175 539286 150184
rect 539336 150142 539364 161978
rect 539324 150136 539376 150142
rect 539324 150078 539376 150084
rect 539796 149940 539824 173159
rect 538864 149932 538916 149938
rect 515036 149874 515088 149880
rect 538864 149874 538916 149880
rect 538956 149932 539008 149938
rect 538956 149874 539008 149880
rect 59648 132466 59768 132494
rect 59188 131158 59400 131186
rect 59636 131164 59688 131170
rect 58992 126948 59044 126954
rect 58992 126890 59044 126896
rect 58900 124160 58952 124166
rect 58900 124102 58952 124108
rect 58992 121644 59044 121650
rect 58992 121586 59044 121592
rect 58900 111852 58952 111858
rect 58900 111794 58952 111800
rect 58808 108248 58860 108254
rect 58808 108190 58860 108196
rect 58808 97980 58860 97986
rect 58808 97922 58860 97928
rect 58716 21276 58768 21282
rect 58716 21218 58768 21224
rect 58820 17406 58848 97922
rect 58912 18562 58940 111794
rect 59004 19310 59032 121586
rect 59188 120222 59216 131158
rect 59636 131106 59688 131112
rect 59360 126948 59412 126954
rect 59360 126890 59412 126896
rect 59268 124500 59320 124506
rect 59268 124442 59320 124448
rect 59280 121530 59308 124442
rect 59372 121650 59400 126890
rect 59452 124160 59504 124166
rect 59452 124102 59504 124108
rect 59360 121644 59412 121650
rect 59360 121586 59412 121592
rect 59280 121502 59400 121530
rect 59176 120216 59228 120222
rect 59176 120158 59228 120164
rect 59268 120148 59320 120154
rect 59268 120090 59320 120096
rect 59176 117972 59228 117978
rect 59176 117914 59228 117920
rect 59188 111874 59216 117914
rect 59280 111994 59308 120090
rect 59372 117978 59400 121502
rect 59464 120154 59492 124102
rect 59452 120148 59504 120154
rect 59452 120090 59504 120096
rect 59648 119406 59676 131106
rect 59636 119400 59688 119406
rect 59636 119342 59688 119348
rect 59544 118720 59596 118726
rect 59544 118662 59596 118668
rect 59360 117972 59412 117978
rect 59360 117914 59412 117920
rect 59268 111988 59320 111994
rect 59268 111930 59320 111936
rect 59188 111846 59400 111874
rect 59556 111858 59584 118662
rect 59740 118182 59768 132466
rect 59832 132466 59952 132494
rect 59832 124506 59860 132466
rect 59820 124500 59872 124506
rect 59820 124442 59872 124448
rect 59820 120216 59872 120222
rect 59820 120158 59872 120164
rect 59728 118176 59780 118182
rect 59728 118118 59780 118124
rect 59728 118040 59780 118046
rect 59728 117982 59780 117988
rect 59636 112124 59688 112130
rect 59636 112066 59688 112072
rect 59372 110378 59400 111846
rect 59544 111852 59596 111858
rect 59544 111794 59596 111800
rect 59648 110673 59676 112066
rect 59634 110664 59690 110673
rect 59634 110599 59690 110608
rect 59636 110492 59688 110498
rect 59636 110434 59688 110440
rect 59280 110350 59400 110378
rect 59280 89842 59308 110350
rect 59280 89814 59400 89842
rect 59372 67538 59400 89814
rect 59280 67510 59400 67538
rect 58992 19304 59044 19310
rect 58992 19246 59044 19252
rect 58900 18556 58952 18562
rect 58900 18498 58952 18504
rect 58808 17400 58860 17406
rect 58622 17368 58678 17377
rect 58808 17342 58860 17348
rect 58622 17303 58678 17312
rect 55956 17264 56008 17270
rect 55956 17206 56008 17212
rect 59280 17066 59308 67510
rect 59648 17542 59676 110434
rect 59740 98054 59768 117982
rect 59832 112130 59860 120158
rect 59820 112124 59872 112130
rect 59820 112066 59872 112072
rect 59820 111988 59872 111994
rect 59820 111930 59872 111936
rect 59728 98048 59780 98054
rect 59728 97990 59780 97996
rect 59728 97912 59780 97918
rect 59728 97854 59780 97860
rect 59740 25838 59768 97854
rect 59728 25832 59780 25838
rect 59728 25774 59780 25780
rect 59832 20058 59860 111930
rect 539980 46889 540008 177346
rect 540060 155916 540112 155922
rect 540060 155858 540112 155864
rect 539966 46880 540022 46889
rect 539966 46815 540022 46824
rect 59910 30560 59966 30569
rect 59966 30518 60030 30546
rect 59910 30495 59966 30504
rect 59910 29880 59966 29889
rect 59910 29815 59966 29824
rect 59924 29209 59952 29815
rect 61304 29617 61332 30124
rect 61290 29608 61346 29617
rect 61290 29543 61346 29552
rect 59910 29200 59966 29209
rect 59910 29135 59966 29144
rect 62592 27538 62620 30124
rect 63236 29578 63264 30124
rect 63224 29572 63276 29578
rect 63224 29514 63276 29520
rect 62580 27532 62632 27538
rect 62580 27474 62632 27480
rect 65168 27441 65196 30124
rect 65812 27577 65840 30124
rect 66456 29889 66484 30124
rect 66442 29880 66498 29889
rect 66442 29815 66498 29824
rect 67744 28898 67772 30124
rect 69048 29866 69076 30124
rect 69032 29838 69076 29866
rect 69032 29646 69060 29838
rect 69020 29640 69072 29646
rect 69020 29582 69072 29588
rect 69676 29510 69704 30124
rect 69664 29504 69716 29510
rect 69664 29446 69716 29452
rect 67732 28892 67784 28898
rect 67732 28834 67784 28840
rect 67638 28248 67694 28257
rect 67638 28183 67694 28192
rect 69570 28248 69626 28257
rect 69570 28183 69626 28192
rect 65798 27568 65854 27577
rect 65798 27503 65854 27512
rect 65154 27432 65210 27441
rect 65154 27367 65210 27376
rect 59820 20052 59872 20058
rect 59820 19994 59872 20000
rect 59636 17536 59688 17542
rect 59636 17478 59688 17484
rect 59268 17060 59320 17066
rect 59268 17002 59320 17008
rect 50172 16546 50292 16574
rect 52472 16546 53328 16574
rect 48780 4004 48832 4010
rect 48780 3946 48832 3952
rect 48228 3868 48280 3874
rect 48228 3810 48280 3816
rect 50158 3496 50214 3505
rect 50158 3431 50214 3440
rect 50172 480 50200 3431
rect 50264 3330 50292 16546
rect 50252 3324 50304 3330
rect 50252 3266 50304 3272
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 56784 11756 56836 11762
rect 56784 11698 56836 11704
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 11698
rect 64326 4856 64382 4865
rect 64326 4791 64382 4800
rect 60830 3496 60886 3505
rect 60830 3431 60886 3440
rect 60844 480 60872 3431
rect 64340 480 64368 4791
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 28183
rect 69584 22098 69612 28183
rect 69756 28144 69808 28150
rect 69756 28086 69808 28092
rect 69768 23458 69796 28086
rect 70320 27606 70348 30124
rect 70964 28966 70992 30124
rect 71608 29442 71636 30124
rect 72912 29866 72940 30124
rect 72896 29838 72940 29866
rect 71596 29436 71648 29442
rect 71596 29378 71648 29384
rect 70952 28960 71004 28966
rect 70952 28902 71004 28908
rect 72516 28348 72568 28354
rect 72516 28290 72568 28296
rect 70308 27600 70360 27606
rect 70308 27542 70360 27548
rect 71778 27568 71834 27577
rect 71778 27503 71834 27512
rect 71792 27010 71820 27503
rect 71608 26982 71820 27010
rect 71608 26761 71636 26982
rect 71780 26920 71832 26926
rect 71780 26862 71832 26868
rect 71792 26761 71820 26862
rect 71594 26752 71650 26761
rect 71594 26687 71650 26696
rect 71778 26752 71834 26761
rect 71778 26687 71834 26696
rect 70398 25936 70454 25945
rect 70398 25871 70454 25880
rect 69756 23452 69808 23458
rect 69756 23394 69808 23400
rect 69572 22092 69624 22098
rect 69572 22034 69624 22040
rect 70412 16574 70440 25871
rect 72528 19242 72556 28290
rect 72896 27577 72924 29838
rect 73540 28558 73568 30124
rect 73528 28552 73580 28558
rect 73528 28494 73580 28500
rect 74632 28552 74684 28558
rect 74632 28494 74684 28500
rect 72882 27568 72938 27577
rect 72882 27503 72938 27512
rect 74538 25800 74594 25809
rect 74538 25735 74594 25744
rect 72516 19236 72568 19242
rect 72516 19178 72568 19184
rect 74552 16574 74580 25735
rect 74644 22001 74672 28494
rect 78048 26234 78076 30124
rect 82556 28830 82584 30124
rect 82818 29744 82874 29753
rect 82818 29679 82874 29688
rect 82832 28830 82860 29679
rect 82544 28824 82596 28830
rect 82544 28766 82596 28772
rect 82820 28824 82872 28830
rect 82820 28766 82872 28772
rect 84488 26234 84516 30124
rect 85792 29866 85820 30124
rect 85776 29838 85820 29866
rect 85776 27305 85804 29838
rect 87708 28286 87736 30124
rect 89656 29866 89684 30124
rect 89640 29838 89684 29866
rect 89640 28422 89668 29838
rect 89628 28416 89680 28422
rect 89628 28358 89680 28364
rect 89720 28416 89772 28422
rect 89720 28358 89772 28364
rect 87696 28280 87748 28286
rect 87696 28222 87748 28228
rect 89076 28280 89128 28286
rect 89732 28234 89760 28358
rect 89076 28222 89128 28228
rect 88984 27668 89036 27674
rect 88984 27610 89036 27616
rect 85762 27296 85818 27305
rect 85762 27231 85818 27240
rect 77404 26206 78076 26234
rect 84212 26206 84516 26234
rect 77300 25356 77352 25362
rect 77300 25298 77352 25304
rect 74630 21992 74686 22001
rect 74630 21927 74686 21936
rect 77312 16574 77340 25298
rect 77404 24449 77432 26206
rect 81440 25424 81492 25430
rect 81440 25366 81492 25372
rect 77390 24440 77446 24449
rect 77390 24375 77446 24384
rect 81452 16574 81480 25366
rect 84212 17921 84240 26206
rect 85578 25664 85634 25673
rect 85578 25599 85634 25608
rect 84198 17912 84254 17921
rect 84198 17847 84254 17856
rect 85592 16574 85620 25599
rect 88338 25528 88394 25537
rect 88338 25463 88394 25472
rect 88352 16574 88380 25463
rect 88996 19310 89024 27610
rect 88984 19304 89036 19310
rect 88984 19246 89036 19252
rect 89088 18562 89116 28222
rect 89640 28206 89760 28234
rect 89640 27674 89668 28206
rect 89628 27668 89680 27674
rect 89628 27610 89680 27616
rect 91572 26234 91600 30124
rect 92216 27946 92244 30124
rect 95436 28234 95464 30124
rect 95344 28206 95464 28234
rect 92204 27940 92256 27946
rect 92204 27882 92256 27888
rect 91204 26206 91600 26234
rect 91204 24857 91232 26206
rect 91190 24848 91246 24857
rect 91190 24783 91246 24792
rect 95344 23934 95372 28206
rect 96080 26234 96108 30124
rect 98656 26234 98684 30124
rect 99300 28121 99328 30124
rect 99286 28112 99342 28121
rect 99286 28047 99342 28056
rect 100588 26994 100616 30124
rect 100576 26988 100628 26994
rect 100576 26930 100628 26936
rect 101232 26234 101260 30124
rect 103164 26234 103192 30124
rect 103808 28626 103836 30124
rect 103796 28620 103848 28626
rect 103796 28562 103848 28568
rect 105096 28490 105124 30124
rect 105636 28620 105688 28626
rect 105636 28562 105688 28568
rect 105084 28484 105136 28490
rect 105084 28426 105136 28432
rect 105544 28484 105596 28490
rect 105544 28426 105596 28432
rect 95436 26206 96108 26234
rect 98012 26206 98684 26234
rect 100772 26206 101260 26234
rect 102152 26206 103192 26234
rect 95332 23928 95384 23934
rect 95332 23870 95384 23876
rect 95240 19780 95292 19786
rect 95240 19722 95292 19728
rect 89076 18556 89128 18562
rect 89076 18498 89128 18504
rect 95252 16574 95280 19722
rect 95436 19009 95464 26206
rect 98012 25498 98040 26206
rect 100772 25566 100800 26206
rect 100760 25560 100812 25566
rect 100760 25502 100812 25508
rect 98000 25492 98052 25498
rect 98000 25434 98052 25440
rect 102152 22642 102180 26206
rect 102140 22636 102192 22642
rect 102140 22578 102192 22584
rect 99378 19952 99434 19961
rect 99378 19887 99434 19896
rect 95422 19000 95478 19009
rect 95422 18935 95478 18944
rect 99392 16574 99420 19887
rect 105556 17066 105584 28426
rect 105648 18630 105676 28562
rect 107028 26234 107056 30124
rect 106384 26206 107056 26234
rect 107672 26234 107700 30124
rect 108960 26234 108988 30124
rect 109604 29034 109632 30124
rect 109592 29028 109644 29034
rect 109592 28970 109644 28976
rect 107672 26206 107792 26234
rect 105636 18624 105688 18630
rect 105636 18566 105688 18572
rect 106278 18592 106334 18601
rect 106278 18527 106334 18536
rect 105544 17060 105596 17066
rect 105544 17002 105596 17008
rect 106292 16574 106320 18527
rect 106384 17785 106412 26206
rect 107764 23225 107792 26206
rect 107948 26206 108988 26234
rect 107948 23225 107976 26206
rect 107750 23216 107806 23225
rect 107750 23151 107806 23160
rect 107934 23216 107990 23225
rect 107934 23151 107990 23160
rect 116044 22710 116072 30124
rect 116688 27266 116716 30124
rect 117976 28937 118004 30124
rect 117962 28928 118018 28937
rect 117962 28863 118018 28872
rect 120552 28150 120580 30124
rect 120540 28144 120592 28150
rect 120540 28086 120592 28092
rect 123772 27470 123800 30124
rect 124416 28218 124444 30124
rect 125704 28234 125732 30124
rect 124404 28212 124456 28218
rect 124404 28154 124456 28160
rect 125612 28206 125732 28234
rect 123760 27464 123812 27470
rect 123760 27406 123812 27412
rect 116676 27260 116728 27266
rect 116676 27202 116728 27208
rect 116032 22704 116084 22710
rect 116032 22646 116084 22652
rect 124218 22672 124274 22681
rect 124218 22607 124274 22616
rect 113178 18728 113234 18737
rect 113178 18663 113234 18672
rect 106370 17776 106426 17785
rect 106370 17711 106426 17720
rect 113192 16574 113220 18663
rect 117320 17128 117372 17134
rect 117320 17070 117372 17076
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 77312 16546 78168 16574
rect 81452 16546 81664 16574
rect 85592 16546 85712 16574
rect 88352 16546 89208 16574
rect 95252 16546 95832 16574
rect 99392 16546 99880 16574
rect 106292 16546 106504 16574
rect 113192 16546 114048 16574
rect 71516 480 71544 16546
rect 75012 480 75040 16546
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 85684 480 85712 16546
rect 89180 480 89208 16546
rect 92478 15872 92534 15881
rect 92478 15807 92534 15816
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 15807
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 16546
rect 99852 480 99880 16546
rect 103334 3360 103390 3369
rect 103334 3295 103390 3304
rect 103348 480 103376 3295
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 110512 3324 110564 3330
rect 110512 3266 110564 3272
rect 110524 480 110552 3266
rect 114020 480 114048 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 17070
rect 124232 16574 124260 22607
rect 125612 19854 125640 28206
rect 126348 26234 126376 30124
rect 127652 29866 127680 30124
rect 127636 29838 127680 29866
rect 127636 27946 127664 29838
rect 128924 28082 128952 30124
rect 128912 28076 128964 28082
rect 128912 28018 128964 28024
rect 127624 27940 127676 27946
rect 127624 27882 127676 27888
rect 129568 26234 129596 30124
rect 131516 29866 131544 30124
rect 125704 26206 126376 26234
rect 128464 26206 129596 26234
rect 131132 29838 131544 29866
rect 125704 21593 125732 26206
rect 125690 21584 125746 21593
rect 125690 21519 125746 21528
rect 128358 21312 128414 21321
rect 128464 21282 128492 26206
rect 131132 22574 131160 29838
rect 132144 26234 132172 30124
rect 138584 26234 138612 30124
rect 139888 29866 139916 30124
rect 131224 26206 132172 26234
rect 138032 26206 138612 26234
rect 139412 29838 139916 29866
rect 131224 25634 131252 26206
rect 131212 25628 131264 25634
rect 131212 25570 131264 25576
rect 138032 23458 138060 26206
rect 138020 23452 138072 23458
rect 138020 23394 138072 23400
rect 131120 22568 131172 22574
rect 131120 22510 131172 22516
rect 139412 21418 139440 29838
rect 141804 26234 141832 30124
rect 143092 26234 143120 30124
rect 140792 26206 141832 26234
rect 142172 26206 143120 26234
rect 139400 21412 139452 21418
rect 139400 21354 139452 21360
rect 140792 21350 140820 26206
rect 142172 24002 142200 26206
rect 142160 23996 142212 24002
rect 142160 23938 142212 23944
rect 140780 21344 140832 21350
rect 140780 21286 140832 21292
rect 128358 21247 128414 21256
rect 128452 21276 128504 21282
rect 125600 19848 125652 19854
rect 125600 19790 125652 19796
rect 128372 16574 128400 21247
rect 128452 21218 128504 21224
rect 135260 20732 135312 20738
rect 135260 20674 135312 20680
rect 124232 16546 124720 16574
rect 128372 16546 128952 16574
rect 120632 15904 120684 15910
rect 120632 15846 120684 15852
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 15846
rect 124692 480 124720 16546
rect 125876 4140 125928 4146
rect 125876 4082 125928 4088
rect 125888 480 125916 4082
rect 126978 3360 127034 3369
rect 126978 3295 127034 3304
rect 126992 480 127020 3295
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 132960 11824 133012 11830
rect 132960 11766 133012 11772
rect 130568 3392 130620 3398
rect 130568 3334 130620 3340
rect 130580 480 130608 3334
rect 132972 480 133000 11766
rect 134156 4072 134208 4078
rect 134156 4014 134208 4020
rect 134168 480 134196 4014
rect 135272 3398 135300 20674
rect 139398 20088 139454 20097
rect 139398 20023 139454 20032
rect 136638 17232 136694 17241
rect 136638 17167 136694 17176
rect 136652 16574 136680 17167
rect 139412 16574 139440 20023
rect 146312 18766 146340 30124
rect 148888 28218 148916 30124
rect 147680 28212 147732 28218
rect 147680 28154 147732 28160
rect 148876 28212 148928 28218
rect 148876 28154 148928 28160
rect 147692 21554 147720 28154
rect 149532 26234 149560 30124
rect 151464 26234 151492 30124
rect 154684 26234 154712 30124
rect 155972 28234 156000 30124
rect 157276 29866 157304 30124
rect 157260 29838 157304 29866
rect 155972 28206 156092 28234
rect 155960 28144 156012 28150
rect 155960 28086 156012 28092
rect 149072 26206 149560 26234
rect 150452 26206 151492 26234
rect 154592 26206 154712 26234
rect 147680 21548 147732 21554
rect 147680 21490 147732 21496
rect 146390 21448 146446 21457
rect 146390 21383 146446 21392
rect 146300 18760 146352 18766
rect 146300 18702 146352 18708
rect 146404 16574 146432 21383
rect 149072 19922 149100 26206
rect 149060 19916 149112 19922
rect 149060 19858 149112 19864
rect 150452 18834 150480 26206
rect 150440 18828 150492 18834
rect 150440 18770 150492 18776
rect 154592 18698 154620 26206
rect 155972 21486 156000 28086
rect 156064 25702 156092 28206
rect 157260 28150 157288 29838
rect 158548 29034 158576 30124
rect 159836 29374 159864 30124
rect 161140 29866 161168 30124
rect 160112 29838 161168 29866
rect 159824 29368 159876 29374
rect 159824 29310 159876 29316
rect 158536 29028 158588 29034
rect 158536 28970 158588 28976
rect 157248 28144 157300 28150
rect 157248 28086 157300 28092
rect 156052 25696 156104 25702
rect 156052 25638 156104 25644
rect 155960 21480 156012 21486
rect 155960 21422 156012 21428
rect 154580 18692 154632 18698
rect 154580 18634 154632 18640
rect 160112 18426 160140 29838
rect 162412 26234 162440 30124
rect 161492 26206 162440 26234
rect 161492 24070 161520 26206
rect 164238 24168 164294 24177
rect 164238 24103 164294 24112
rect 161480 24064 161532 24070
rect 161480 24006 161532 24012
rect 161480 20800 161532 20806
rect 161480 20742 161532 20748
rect 160100 18420 160152 18426
rect 160100 18362 160152 18368
rect 153198 17504 153254 17513
rect 153198 17439 153254 17448
rect 147680 17196 147732 17202
rect 147680 17138 147732 17144
rect 147692 16574 147720 17138
rect 153212 16574 153240 17439
rect 161492 16574 161520 20742
rect 164252 16574 164280 24103
rect 164344 18494 164372 30124
rect 165648 29866 165676 30124
rect 165648 29838 165752 29866
rect 165620 28212 165672 28218
rect 165620 28154 165672 28160
rect 165632 23769 165660 28154
rect 165724 25770 165752 29838
rect 166276 28218 166304 30124
rect 166920 28393 166948 30124
rect 166906 28384 166962 28393
rect 166906 28319 166962 28328
rect 168208 28218 168236 30124
rect 169512 29918 169540 30124
rect 168380 29912 168432 29918
rect 168380 29854 168432 29860
rect 169500 29912 169552 29918
rect 169500 29854 169552 29860
rect 166264 28212 166316 28218
rect 166264 28154 166316 28160
rect 167000 28212 167052 28218
rect 167000 28154 167052 28160
rect 168196 28212 168248 28218
rect 168196 28154 168248 28160
rect 165712 25764 165764 25770
rect 165712 25706 165764 25712
rect 165618 23760 165674 23769
rect 165618 23695 165674 23704
rect 167012 19990 167040 28154
rect 167000 19984 167052 19990
rect 167000 19926 167052 19932
rect 168392 19145 168420 29854
rect 170784 29306 170812 30124
rect 170772 29300 170824 29306
rect 170772 29242 170824 29248
rect 171428 26234 171456 30124
rect 174020 29866 174048 30124
rect 174004 29838 174048 29866
rect 174004 28665 174032 29838
rect 173990 28656 174046 28665
rect 173990 28591 174046 28600
rect 174648 27470 174676 30124
rect 175292 27985 175320 30124
rect 175278 27976 175334 27985
rect 175278 27911 175334 27920
rect 174636 27464 174688 27470
rect 174636 27406 174688 27412
rect 178512 26234 178540 30124
rect 179800 26234 179828 30124
rect 181088 26234 181116 30124
rect 182392 29866 182420 30124
rect 182376 29838 182420 29866
rect 182376 29209 182404 29838
rect 182362 29200 182418 29209
rect 182362 29135 182418 29144
rect 183020 26234 183048 30124
rect 183664 26234 183692 30124
rect 171152 26206 171456 26234
rect 178144 26206 178540 26234
rect 179432 26206 179828 26234
rect 180812 26206 181116 26234
rect 182192 26206 183048 26234
rect 183572 26206 183692 26234
rect 184952 26234 184980 30124
rect 186256 29866 186284 30124
rect 186240 29838 186284 29866
rect 186240 28257 186268 29838
rect 187528 29170 187556 30124
rect 187516 29164 187568 29170
rect 187516 29106 187568 29112
rect 188816 28529 188844 30124
rect 188802 28520 188858 28529
rect 188802 28455 188858 28464
rect 186226 28248 186282 28257
rect 186226 28183 186282 28192
rect 189460 26234 189488 30124
rect 190764 29866 190792 30124
rect 190748 29838 190792 29866
rect 190748 28558 190776 29838
rect 190736 28552 190788 28558
rect 190736 28494 190788 28500
rect 191392 26234 191420 30124
rect 191840 28212 191892 28218
rect 191840 28154 191892 28160
rect 184952 26206 185072 26234
rect 171152 24002 171180 26206
rect 171140 23996 171192 24002
rect 171140 23938 171192 23944
rect 178038 22672 178094 22681
rect 178038 22607 178094 22616
rect 176660 21412 176712 21418
rect 176660 21354 176712 21360
rect 168378 19136 168434 19145
rect 168378 19071 168434 19080
rect 164332 18488 164384 18494
rect 164332 18430 164384 18436
rect 165620 17264 165672 17270
rect 165620 17206 165672 17212
rect 165632 16574 165660 17206
rect 136652 16546 137232 16574
rect 139412 16546 139624 16574
rect 146404 16546 147168 16574
rect 147692 16546 147904 16574
rect 153212 16546 153792 16574
rect 161492 16546 162072 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 136468 480 136496 3334
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 144734 16008 144790 16017
rect 144734 15943 144790 15952
rect 143540 13116 143592 13122
rect 143540 13058 143592 13064
rect 141240 10328 141292 10334
rect 141240 10270 141292 10276
rect 141252 480 141280 10270
rect 143552 480 143580 13058
rect 144748 480 144776 15943
rect 147140 480 147168 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 151820 4004 151872 4010
rect 151820 3946 151872 3952
rect 150622 3496 150678 3505
rect 150622 3431 150678 3440
rect 150636 480 150664 3431
rect 151832 480 151860 3946
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155406 4992 155462 5001
rect 155406 4927 155462 4936
rect 155420 480 155448 4927
rect 158904 3936 158956 3942
rect 158904 3878 158956 3884
rect 157798 3632 157854 3641
rect 157798 3567 157854 3576
rect 157812 480 157840 3567
rect 158916 480 158944 3878
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 161308 480 161336 3402
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 175464 14544 175516 14550
rect 175464 14486 175516 14492
rect 171968 14476 172020 14482
rect 171968 14418 172020 14424
rect 169574 3768 169630 3777
rect 169574 3703 169630 3712
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 168392 480 168420 3402
rect 169588 480 169616 3703
rect 171980 480 172008 14418
rect 173164 3868 173216 3874
rect 173164 3810 173216 3816
rect 173176 480 173204 3810
rect 175476 480 175504 14486
rect 176672 480 176700 21354
rect 178052 16574 178080 22607
rect 178144 17649 178172 26206
rect 179432 21622 179460 26206
rect 179420 21616 179472 21622
rect 179420 21558 179472 21564
rect 179420 20868 179472 20874
rect 179420 20810 179472 20816
rect 178130 17640 178186 17649
rect 178130 17575 178186 17584
rect 179432 16574 179460 20810
rect 180812 17105 180840 26206
rect 182192 22778 182220 26206
rect 183572 22846 183600 26206
rect 184938 25528 184994 25537
rect 184938 25463 184994 25472
rect 183560 22840 183612 22846
rect 183560 22782 183612 22788
rect 182180 22772 182232 22778
rect 182180 22714 182232 22720
rect 183558 21584 183614 21593
rect 183558 21519 183614 21528
rect 180798 17096 180854 17105
rect 180798 17031 180854 17040
rect 183572 16574 183600 21519
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 183572 16546 183784 16574
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 182546 3224 182602 3233
rect 182546 3159 182602 3168
rect 182560 480 182588 3159
rect 183756 480 183784 16546
rect 184952 3534 184980 25463
rect 185044 23390 185072 26206
rect 189092 26206 189488 26234
rect 190564 26206 191420 26234
rect 185032 23384 185084 23390
rect 185032 23326 185084 23332
rect 189092 18902 189120 26206
rect 189080 18896 189132 18902
rect 189080 18838 189132 18844
rect 190564 17882 190592 26206
rect 190552 17876 190604 17882
rect 190552 17818 190604 17824
rect 191852 17338 191880 28154
rect 192036 26234 192064 30124
rect 192680 28218 192708 30124
rect 192668 28212 192720 28218
rect 192668 28154 192720 28160
rect 193324 26234 193352 30124
rect 195256 28694 195284 30124
rect 195244 28688 195296 28694
rect 195244 28630 195296 28636
rect 195900 28218 195928 30124
rect 194692 28212 194744 28218
rect 194692 28154 194744 28160
rect 195888 28212 195940 28218
rect 195888 28154 195940 28160
rect 191944 26206 192064 26234
rect 193232 26206 193352 26234
rect 191944 24818 191972 26206
rect 191932 24812 191984 24818
rect 191932 24754 191984 24760
rect 193232 22506 193260 26206
rect 193220 22500 193272 22506
rect 193220 22442 193272 22448
rect 194704 18970 194732 28154
rect 197832 26234 197860 30124
rect 199764 29238 199792 30124
rect 199752 29232 199804 29238
rect 199752 29174 199804 29180
rect 201696 26234 201724 30124
rect 203628 26234 203656 30124
rect 204916 28762 204944 30124
rect 205560 29102 205588 30124
rect 205548 29096 205600 29102
rect 205548 29038 205600 29044
rect 204904 28756 204956 28762
rect 204904 28698 204956 28704
rect 206204 26234 206232 30124
rect 208136 26234 208164 30124
rect 210068 26234 210096 30124
rect 211372 29866 211400 30124
rect 211356 29838 211400 29866
rect 211356 28626 211384 29838
rect 211344 28620 211396 28626
rect 211344 28562 211396 28568
rect 212000 26234 212028 30124
rect 197372 26206 197860 26234
rect 201512 26206 201724 26234
rect 202892 26206 203656 26234
rect 205652 26206 206232 26234
rect 207032 26206 208164 26234
rect 209792 26206 210096 26234
rect 211264 26206 212028 26234
rect 197372 24138 197400 26206
rect 197360 24132 197412 24138
rect 197360 24074 197412 24080
rect 194692 18964 194744 18970
rect 194692 18906 194744 18912
rect 191840 17332 191892 17338
rect 191840 17274 191892 17280
rect 201512 16998 201540 26206
rect 202892 20126 202920 26206
rect 205652 21690 205680 26206
rect 207032 21729 207060 26206
rect 207110 24304 207166 24313
rect 207110 24239 207166 24248
rect 207018 21720 207074 21729
rect 205640 21684 205692 21690
rect 207018 21655 207074 21664
rect 205640 21626 205692 21632
rect 202880 20120 202932 20126
rect 202880 20062 202932 20068
rect 201592 19372 201644 19378
rect 201592 19314 201644 19320
rect 201500 16992 201552 16998
rect 201500 16934 201552 16940
rect 194416 11892 194468 11898
rect 194416 11834 194468 11840
rect 189724 3800 189776 3806
rect 189724 3742 189776 3748
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 186136 3528 186188 3534
rect 186136 3470 186188 3476
rect 186148 480 186176 3470
rect 187332 3392 187384 3398
rect 187332 3334 187384 3340
rect 187344 480 187372 3334
rect 189736 480 189764 3742
rect 193220 3732 193272 3738
rect 193220 3674 193272 3680
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 190840 480 190868 3470
rect 193232 480 193260 3674
rect 194428 480 194456 11834
rect 201604 6914 201632 19314
rect 203430 14920 203486 14929
rect 203430 14855 203486 14864
rect 201512 6886 201632 6914
rect 197910 4040 197966 4049
rect 197910 3975 197966 3984
rect 196808 3664 196860 3670
rect 196808 3606 196860 3612
rect 196820 480 196848 3606
rect 197924 480 197952 3975
rect 200302 3904 200358 3913
rect 200302 3839 200358 3848
rect 200316 480 200344 3839
rect 201512 480 201540 6886
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 14855
rect 205086 10296 205142 10305
rect 205086 10231 205142 10240
rect 205100 480 205128 10231
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 24239
rect 209792 24206 209820 26206
rect 211264 25838 211292 26206
rect 211252 25832 211304 25838
rect 211252 25774 211304 25780
rect 209780 24200 209832 24206
rect 209780 24142 209832 24148
rect 209872 24132 209924 24138
rect 209872 24074 209924 24080
rect 209884 16574 209912 24074
rect 212644 17513 212672 30124
rect 213288 28286 213316 30124
rect 213276 28280 213328 28286
rect 213276 28222 213328 28228
rect 213932 25906 213960 30124
rect 216508 28218 216536 30124
rect 215300 28212 215352 28218
rect 215300 28154 215352 28160
rect 216496 28212 216548 28218
rect 216496 28154 216548 28160
rect 213920 25900 213972 25906
rect 213920 25842 213972 25848
rect 215312 19106 215340 28154
rect 217152 26234 217180 30124
rect 217796 28014 217824 30124
rect 219744 29866 219772 30124
rect 219452 29838 219772 29866
rect 217784 28008 217836 28014
rect 217784 27950 217836 27956
rect 216784 26206 217180 26234
rect 216784 20058 216812 26206
rect 219452 24342 219480 29838
rect 220372 26234 220400 30124
rect 221016 26234 221044 30124
rect 222948 26234 222976 30124
rect 224252 29866 224280 30124
rect 228116 29866 228144 30124
rect 224236 29838 224280 29866
rect 227732 29838 228144 29866
rect 224236 27266 224264 29838
rect 224224 27260 224276 27266
rect 224224 27202 224276 27208
rect 219544 26206 220400 26234
rect 220924 26206 221044 26234
rect 222212 26206 222976 26234
rect 219440 24336 219492 24342
rect 219440 24278 219492 24284
rect 219544 24274 219572 26206
rect 219532 24268 219584 24274
rect 219532 24210 219584 24216
rect 220820 24200 220872 24206
rect 220820 24142 220872 24148
rect 216772 20052 216824 20058
rect 216772 19994 216824 20000
rect 215300 19100 215352 19106
rect 215300 19042 215352 19048
rect 212630 17504 212686 17513
rect 212630 17439 212686 17448
rect 209884 16546 211016 16574
rect 208582 13016 208638 13025
rect 208582 12951 208638 12960
rect 208596 480 208624 12951
rect 210988 480 211016 16546
rect 214470 14648 214526 14657
rect 214470 14583 214526 14592
rect 212172 3596 212224 3602
rect 212172 3538 212224 3544
rect 212184 480 212212 3538
rect 214484 480 214512 14583
rect 218058 11656 218114 11665
rect 218058 11591 218114 11600
rect 218072 3602 218100 11591
rect 220832 6914 220860 24142
rect 220924 15162 220952 26206
rect 222212 17377 222240 26206
rect 224958 24440 225014 24449
rect 224958 24375 225014 24384
rect 222198 17368 222254 17377
rect 222198 17303 222254 17312
rect 224972 16574 225000 24375
rect 227732 17406 227760 29838
rect 230032 26234 230060 30124
rect 232624 29866 232652 30124
rect 229112 26206 230060 26234
rect 231964 29838 232652 29866
rect 229112 21758 229140 26206
rect 231858 25664 231914 25673
rect 231858 25599 231914 25608
rect 229100 21752 229152 21758
rect 229100 21694 229152 21700
rect 229100 21480 229152 21486
rect 229100 21422 229152 21428
rect 227720 17400 227772 17406
rect 227720 17342 227772 17348
rect 229112 16574 229140 21422
rect 224972 16546 225184 16574
rect 229112 16546 229416 16574
rect 220912 15156 220964 15162
rect 220912 15098 220964 15104
rect 222750 11792 222806 11801
rect 222750 11727 222806 11736
rect 220832 6886 221136 6914
rect 218152 3732 218204 3738
rect 218152 3674 218204 3680
rect 218060 3596 218112 3602
rect 218060 3538 218112 3544
rect 215668 3392 215720 3398
rect 215668 3334 215720 3340
rect 215680 480 215708 3334
rect 218164 1850 218192 3674
rect 219256 3596 219308 3602
rect 219256 3538 219308 3544
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 218072 1822 218192 1850
rect 218072 480 218100 1822
rect 219268 480 219296 3538
rect 219360 3398 219388 3538
rect 219348 3392 219400 3398
rect 219348 3334 219400 3340
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 6886
rect 222764 480 222792 11727
rect 225156 480 225184 16546
rect 226338 14784 226394 14793
rect 226338 14719 226394 14728
rect 226352 480 226380 14719
rect 228272 11960 228324 11966
rect 228272 11902 228324 11908
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 11902
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 25599
rect 231964 13705 231992 29838
rect 233252 13802 233280 30124
rect 234540 28529 234568 30124
rect 234526 28520 234582 28529
rect 234526 28455 234582 28464
rect 235184 26234 235212 30124
rect 237116 26234 237144 30124
rect 238404 26234 238432 30124
rect 243556 26234 243584 30124
rect 244200 27130 244228 30124
rect 244188 27124 244240 27130
rect 244188 27066 244240 27072
rect 246776 26234 246804 30124
rect 247420 28966 247448 30124
rect 247408 28960 247460 28966
rect 247408 28902 247460 28908
rect 249996 28830 250024 30124
rect 249984 28824 250036 28830
rect 249984 28766 250036 28772
rect 251284 28234 251312 30124
rect 234632 26206 235212 26234
rect 236012 26206 237144 26234
rect 237392 26206 238432 26234
rect 243004 26206 243584 26234
rect 245764 26206 246804 26234
rect 251192 28206 251312 28234
rect 234632 17474 234660 26206
rect 236012 17746 236040 26206
rect 236000 17740 236052 17746
rect 236000 17682 236052 17688
rect 234620 17468 234672 17474
rect 234620 17410 234672 17416
rect 234620 17264 234672 17270
rect 234620 17206 234672 17212
rect 233424 14680 233476 14686
rect 233424 14622 233476 14628
rect 233240 13796 233292 13802
rect 233240 13738 233292 13744
rect 231950 13696 232006 13705
rect 231950 13631 232006 13640
rect 233436 480 233464 14622
rect 234632 3398 234660 17206
rect 237392 16930 237420 26206
rect 237380 16924 237432 16930
rect 237380 16866 237432 16872
rect 243004 16561 243032 26206
rect 245660 24268 245712 24274
rect 245660 24210 245712 24216
rect 245672 16574 245700 24210
rect 245764 17610 245792 26206
rect 249800 21548 249852 21554
rect 249800 21490 249852 21496
rect 245752 17604 245804 17610
rect 245752 17546 245804 17552
rect 249812 16574 249840 21490
rect 251192 17542 251220 28206
rect 251928 26234 251956 30124
rect 252572 28354 252600 30124
rect 252560 28348 252612 28354
rect 252560 28290 252612 28296
rect 256436 26234 256464 30124
rect 257740 29866 257768 30124
rect 251284 26206 251956 26234
rect 255332 26206 256464 26234
rect 256712 29838 257768 29866
rect 251284 17610 251312 26206
rect 255332 24721 255360 26206
rect 255318 24712 255374 24721
rect 255318 24647 255374 24656
rect 256712 24410 256740 29838
rect 259012 28422 259040 30124
rect 259000 28416 259052 28422
rect 259000 28358 259052 28364
rect 256700 24404 256752 24410
rect 256700 24346 256752 24352
rect 260838 19000 260894 19009
rect 260838 18935 260894 18944
rect 251272 17604 251324 17610
rect 251272 17546 251324 17552
rect 251180 17536 251232 17542
rect 251180 17478 251232 17484
rect 259460 17400 259512 17406
rect 259460 17342 259512 17348
rect 256700 17332 256752 17338
rect 256700 17274 256752 17280
rect 242990 16552 243046 16561
rect 245672 16546 245976 16574
rect 249812 16546 250024 16574
rect 242990 16487 243046 16496
rect 242898 11928 242954 11937
rect 242898 11863 242954 11872
rect 240506 6352 240562 6361
rect 240506 6287 240562 6296
rect 239312 3868 239364 3874
rect 239312 3810 239364 3816
rect 237012 3732 237064 3738
rect 237012 3674 237064 3680
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 235828 480 235856 3334
rect 237024 480 237052 3674
rect 239324 480 239352 3810
rect 240520 480 240548 6287
rect 242912 480 242940 11863
rect 244096 3800 244148 3806
rect 244096 3742 244148 3748
rect 244108 480 244136 3742
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247592 14816 247644 14822
rect 247592 14758 247644 14764
rect 247604 480 247632 14758
rect 249996 480 250024 16546
rect 251178 15056 251234 15065
rect 251178 14991 251234 15000
rect 251192 480 251220 14991
rect 254216 14884 254268 14890
rect 254216 14826 254268 14832
rect 253480 14612 253532 14618
rect 253480 14554 253532 14560
rect 253492 480 253520 14554
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 14826
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 17274
rect 258264 8968 258316 8974
rect 258264 8910 258316 8916
rect 258276 480 258304 8910
rect 259472 3398 259500 17342
rect 260852 16574 260880 18935
rect 260944 17542 260972 30124
rect 266112 29866 266140 30124
rect 266096 29838 266140 29866
rect 266096 28422 266124 29838
rect 266084 28416 266136 28422
rect 266084 28358 266136 28364
rect 266740 26234 266768 30124
rect 268028 28354 268056 30124
rect 268016 28348 268068 28354
rect 268016 28290 268068 28296
rect 268672 27130 268700 30124
rect 270620 29866 270648 30124
rect 270512 29838 270648 29866
rect 268660 27124 268712 27130
rect 268660 27066 268712 27072
rect 266372 26206 266768 26234
rect 266372 24478 266400 26206
rect 266360 24472 266412 24478
rect 266360 24414 266412 24420
rect 270512 21826 270540 29838
rect 271248 28558 271276 30124
rect 271236 28552 271288 28558
rect 271236 28494 271288 28500
rect 272536 28490 272564 30124
rect 272524 28484 272576 28490
rect 272524 28426 272576 28432
rect 275112 26234 275140 30124
rect 275756 28762 275784 30124
rect 275744 28756 275796 28762
rect 275744 28698 275796 28704
rect 276400 26234 276428 30124
rect 280264 26234 280292 30124
rect 284128 29481 284156 30124
rect 284114 29472 284170 29481
rect 284114 29407 284170 29416
rect 286060 26234 286088 30124
rect 287364 29866 287392 30124
rect 287348 29838 287392 29866
rect 287348 29102 287376 29838
rect 287336 29096 287388 29102
rect 287336 29038 287388 29044
rect 289280 26234 289308 30124
rect 291228 29866 291256 30124
rect 291228 29838 291332 29866
rect 291200 28144 291252 28150
rect 291200 28086 291252 28092
rect 274652 26206 275140 26234
rect 276032 26206 276428 26234
rect 280172 26206 280292 26234
rect 285692 26206 286088 26234
rect 288452 26206 289308 26234
rect 274652 24721 274680 26206
rect 274638 24712 274694 24721
rect 274638 24647 274694 24656
rect 270500 21820 270552 21826
rect 270500 21762 270552 21768
rect 271880 19984 271932 19990
rect 271880 19926 271932 19932
rect 267740 18624 267792 18630
rect 267740 18566 267792 18572
rect 260932 17536 260984 17542
rect 260932 17478 260984 17484
rect 267752 16574 267780 18566
rect 271892 16574 271920 19926
rect 260852 16546 261800 16574
rect 267752 16546 268424 16574
rect 271892 16546 272472 16574
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 260668 480 260696 3334
rect 261772 480 261800 16546
rect 264980 14748 265032 14754
rect 264980 14690 265032 14696
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 14690
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 272444 480 272472 16546
rect 276032 10985 276060 26206
rect 280172 25906 280200 26206
rect 280160 25900 280212 25906
rect 280160 25842 280212 25848
rect 285692 24614 285720 26206
rect 285680 24608 285732 24614
rect 285680 24550 285732 24556
rect 278778 18864 278834 18873
rect 278778 18799 278834 18808
rect 276112 18692 276164 18698
rect 276112 18634 276164 18640
rect 276018 10976 276074 10985
rect 276018 10911 276074 10920
rect 276124 6914 276152 18634
rect 278792 16574 278820 18799
rect 282918 17368 282974 17377
rect 282918 17303 282974 17312
rect 282932 16574 282960 17303
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 276032 6886 276152 6914
rect 276032 480 276060 6886
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 283116 480 283144 16546
rect 288452 5506 288480 26206
rect 289818 19136 289874 19145
rect 291212 19106 291240 28086
rect 291304 24546 291332 29838
rect 291856 28150 291884 30124
rect 291844 28144 291896 28150
rect 291844 28086 291896 28092
rect 293144 27062 293172 30124
rect 293132 27056 293184 27062
rect 293132 26998 293184 27004
rect 294432 26234 294460 30124
rect 295736 29866 295764 30124
rect 295720 29838 295764 29866
rect 295720 28490 295748 29838
rect 295708 28484 295760 28490
rect 295708 28426 295760 28432
rect 297008 26234 297036 30124
rect 299600 29866 299628 30124
rect 293972 26206 294460 26234
rect 296732 26206 297036 26234
rect 299492 29838 299628 29866
rect 291292 24540 291344 24546
rect 291292 24482 291344 24488
rect 289818 19071 289874 19080
rect 291200 19100 291252 19106
rect 288440 5500 288492 5506
rect 288440 5442 288492 5448
rect 286600 3936 286652 3942
rect 286600 3878 286652 3884
rect 286612 480 286640 3878
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 19071
rect 291200 19042 291252 19048
rect 293972 19038 294000 26206
rect 296732 22914 296760 26206
rect 296720 22908 296772 22914
rect 296720 22850 296772 22856
rect 296720 20052 296772 20058
rect 296720 19994 296772 20000
rect 293960 19032 294012 19038
rect 293960 18974 294012 18980
rect 296732 16574 296760 19994
rect 299492 17474 299520 29838
rect 300872 29345 300900 30124
rect 300858 29336 300914 29345
rect 300858 29271 300914 29280
rect 302160 28218 302188 30124
rect 304108 29866 304136 30124
rect 303632 29838 304136 29866
rect 300860 28212 300912 28218
rect 300860 28154 300912 28160
rect 302148 28212 302200 28218
rect 302148 28154 302200 28160
rect 299480 17468 299532 17474
rect 299480 17410 299532 17416
rect 296732 16546 297312 16574
rect 293224 15972 293276 15978
rect 293224 15914 293276 15920
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 15914
rect 297284 480 297312 16546
rect 300872 15706 300900 28154
rect 303632 24041 303660 29838
rect 306024 26234 306052 30124
rect 306668 26234 306696 30124
rect 308600 26234 308628 30124
rect 311176 26234 311204 30124
rect 312480 29866 312508 30124
rect 305012 26206 306052 26234
rect 306392 26206 306696 26234
rect 307772 26206 308628 26234
rect 310624 26206 311204 26234
rect 311912 29838 312508 29866
rect 305012 24585 305040 26206
rect 304998 24576 305054 24585
rect 304998 24511 305054 24520
rect 303618 24032 303674 24041
rect 303618 23967 303674 23976
rect 306392 23118 306420 26206
rect 306380 23112 306432 23118
rect 306380 23054 306432 23060
rect 307772 23050 307800 26206
rect 307760 23044 307812 23050
rect 307760 22986 307812 22992
rect 310518 20088 310574 20097
rect 310518 20023 310574 20032
rect 307760 18760 307812 18766
rect 307760 18702 307812 18708
rect 307772 16574 307800 18702
rect 307772 16546 307984 16574
rect 300860 15700 300912 15706
rect 300860 15642 300912 15648
rect 303894 13152 303950 13161
rect 303894 13087 303950 13096
rect 299480 12028 299532 12034
rect 299480 11970 299532 11976
rect 299492 3398 299520 11970
rect 299480 3392 299532 3398
rect 299480 3334 299532 3340
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 13087
rect 307956 480 307984 16546
rect 310532 6914 310560 20023
rect 310624 16522 310652 26206
rect 311912 20194 311940 29838
rect 313752 26234 313780 30124
rect 314396 29345 314424 30124
rect 314382 29336 314438 29345
rect 314382 29271 314438 29280
rect 315040 26234 315068 30124
rect 318904 28234 318932 30124
rect 313292 26206 313780 26234
rect 314672 26206 315068 26234
rect 318812 28206 318932 28234
rect 311900 20188 311952 20194
rect 311900 20130 311952 20136
rect 310612 16516 310664 16522
rect 310612 16458 310664 16464
rect 313292 12374 313320 26206
rect 313280 12368 313332 12374
rect 313280 12310 313332 12316
rect 314672 11014 314700 26206
rect 318812 21865 318840 28206
rect 319548 26234 319576 30124
rect 321480 28218 321508 30124
rect 322124 28626 322152 30124
rect 322112 28620 322164 28626
rect 322112 28562 322164 28568
rect 322768 28218 322796 30124
rect 320180 28212 320232 28218
rect 320180 28154 320232 28160
rect 321468 28212 321520 28218
rect 321468 28154 321520 28160
rect 321560 28212 321612 28218
rect 321560 28154 321612 28160
rect 322756 28212 322808 28218
rect 322756 28154 322808 28160
rect 318904 26206 319576 26234
rect 318904 22953 318932 26206
rect 318890 22944 318946 22953
rect 318890 22879 318946 22888
rect 318798 21856 318854 21865
rect 318798 21791 318854 21800
rect 314752 18828 314804 18834
rect 314752 18770 314804 18776
rect 314660 11008 314712 11014
rect 314660 10950 314712 10956
rect 310532 6886 311480 6914
rect 311452 480 311480 6886
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314764 354 314792 18770
rect 320192 13734 320220 28154
rect 321572 23905 321600 28154
rect 323412 26234 323440 30124
rect 324716 29866 324744 30124
rect 322952 26206 323440 26234
rect 324332 29838 324744 29866
rect 322952 25838 322980 26206
rect 322940 25832 322992 25838
rect 322940 25774 322992 25780
rect 321558 23896 321614 23905
rect 321558 23831 321614 23840
rect 324332 22982 324360 29838
rect 325344 26234 325372 30124
rect 325988 28234 326016 30124
rect 324424 26206 325372 26234
rect 325712 28206 326016 28234
rect 324320 22976 324372 22982
rect 324320 22918 324372 22924
rect 324318 20224 324374 20233
rect 324318 20159 324374 20168
rect 321560 18896 321612 18902
rect 321560 18838 321612 18844
rect 321572 16574 321600 18838
rect 321572 16546 322152 16574
rect 320180 13728 320232 13734
rect 320180 13670 320232 13676
rect 318524 4820 318576 4826
rect 318524 4762 318576 4768
rect 318536 480 318564 4762
rect 322124 480 322152 16546
rect 324332 2106 324360 20159
rect 324424 15094 324452 26206
rect 325712 24682 325740 28206
rect 326632 26234 326660 30124
rect 327276 27062 327304 30124
rect 329224 29866 329252 30124
rect 328472 29838 329252 29866
rect 327264 27056 327316 27062
rect 327264 26998 327316 27004
rect 325804 26206 326660 26234
rect 325804 25770 325832 26206
rect 325792 25764 325844 25770
rect 325792 25706 325844 25712
rect 325700 24676 325752 24682
rect 325700 24618 325752 24624
rect 324412 15088 324464 15094
rect 324412 15030 324464 15036
rect 328472 10946 328500 29838
rect 331140 28218 331168 30124
rect 333716 28393 333744 30124
rect 333702 28384 333758 28393
rect 333702 28319 333758 28328
rect 329840 28212 329892 28218
rect 329840 28154 329892 28160
rect 331128 28212 331180 28218
rect 331128 28154 331180 28160
rect 329852 18465 329880 28154
rect 334360 26234 334388 30124
rect 336292 26234 336320 30124
rect 337596 29866 337624 30124
rect 333992 26206 334388 26234
rect 335464 26206 336320 26234
rect 336752 29838 337624 29866
rect 333992 20262 334020 26206
rect 333980 20256 334032 20262
rect 333980 20198 334032 20204
rect 329838 18456 329894 18465
rect 329838 18391 329894 18400
rect 335358 18456 335414 18465
rect 335358 18391 335414 18400
rect 328734 12064 328790 12073
rect 328734 11999 328790 12008
rect 328460 10940 328512 10946
rect 328460 10882 328512 10888
rect 324320 2100 324372 2106
rect 324320 2042 324372 2048
rect 325608 2100 325660 2106
rect 325608 2042 325660 2048
rect 325620 480 325648 2042
rect 314998 354 315110 480
rect 314764 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 11999
rect 335372 6914 335400 18391
rect 335464 12306 335492 26206
rect 336752 19174 336780 29838
rect 338224 26234 338252 30124
rect 338132 26206 338252 26234
rect 336740 19168 336792 19174
rect 336740 19110 336792 19116
rect 335452 12300 335504 12306
rect 335452 12242 335504 12248
rect 338132 10878 338160 26206
rect 338120 10872 338172 10878
rect 338120 10814 338172 10820
rect 339512 10810 339540 30124
rect 342104 29918 342132 30124
rect 340880 29912 340932 29918
rect 340880 29854 340932 29860
rect 342092 29912 342144 29918
rect 342092 29854 342144 29860
rect 339592 18964 339644 18970
rect 339592 18906 339644 18912
rect 339500 10804 339552 10810
rect 339500 10746 339552 10752
rect 335372 6886 336320 6914
rect 332692 6180 332744 6186
rect 332692 6122 332744 6128
rect 332704 480 332732 6122
rect 336292 480 336320 6886
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339604 354 339632 18906
rect 340892 13666 340920 29854
rect 343376 26234 343404 30124
rect 344020 26994 344048 30124
rect 344008 26988 344060 26994
rect 344008 26930 344060 26936
rect 347240 26234 347268 30124
rect 347780 28212 347832 28218
rect 347780 28154 347832 28160
rect 342272 26206 343404 26234
rect 346412 26206 347268 26234
rect 342272 20330 342300 26206
rect 342260 20324 342312 20330
rect 342260 20266 342312 20272
rect 342904 16040 342956 16046
rect 342904 15982 342956 15988
rect 340880 13660 340932 13666
rect 340880 13602 340932 13608
rect 339838 354 339950 480
rect 339604 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 15982
rect 346412 10742 346440 26206
rect 346952 16108 347004 16114
rect 346952 16050 347004 16056
rect 346400 10736 346452 10742
rect 346400 10678 346452 10684
rect 346964 480 346992 16050
rect 347792 12238 347820 28154
rect 347884 24041 347912 30124
rect 348528 28218 348556 30124
rect 348516 28212 348568 28218
rect 348516 28154 348568 28160
rect 352392 26234 352420 30124
rect 354968 28234 354996 30124
rect 351932 26206 352420 26234
rect 354692 28206 354996 28234
rect 347870 24032 347926 24041
rect 347870 23967 347926 23976
rect 349160 16244 349212 16250
rect 349160 16186 349212 16192
rect 347780 12232 347832 12238
rect 347780 12174 347832 12180
rect 349172 3398 349200 16186
rect 351932 13598 351960 26206
rect 354692 20398 354720 28206
rect 355612 26234 355640 30124
rect 356256 26234 356284 30124
rect 356900 29170 356928 30124
rect 356888 29164 356940 29170
rect 356888 29106 356940 29112
rect 357544 26234 357572 30124
rect 358848 29866 358876 30124
rect 354784 26206 355640 26234
rect 356072 26206 356284 26234
rect 357452 26206 357572 26234
rect 358832 29838 358876 29866
rect 354784 25945 354812 26206
rect 354770 25936 354826 25945
rect 354770 25871 354826 25880
rect 356072 20466 356100 26206
rect 356060 20460 356112 20466
rect 356060 20402 356112 20408
rect 354680 20392 354732 20398
rect 354680 20334 354732 20340
rect 353300 19032 353352 19038
rect 353300 18974 353352 18980
rect 353312 16574 353340 18974
rect 353312 16546 353616 16574
rect 351920 13592 351972 13598
rect 351920 13534 351972 13540
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 357452 13530 357480 26206
rect 358832 22953 358860 29838
rect 359476 28257 359504 30124
rect 359462 28248 359518 28257
rect 359462 28183 359518 28192
rect 360120 28014 360148 30124
rect 362712 29918 362740 30124
rect 361580 29912 361632 29918
rect 361580 29854 361632 29860
rect 362700 29912 362752 29918
rect 362700 29854 362752 29860
rect 360108 28008 360160 28014
rect 360108 27950 360160 27956
rect 361592 23118 361620 29854
rect 363340 26234 363368 30124
rect 363984 27198 364012 30124
rect 364628 28234 364656 30124
rect 364352 28206 364656 28234
rect 363972 27192 364024 27198
rect 363972 27134 364024 27140
rect 363064 26206 363368 26234
rect 361580 23112 361632 23118
rect 361580 23054 361632 23060
rect 358818 22944 358874 22953
rect 358818 22879 358874 22888
rect 360200 22772 360252 22778
rect 360200 22714 360252 22720
rect 360212 16574 360240 22714
rect 360212 16546 361160 16574
rect 357532 16176 357584 16182
rect 357532 16118 357584 16124
rect 357440 13524 357492 13530
rect 357440 13466 357492 13472
rect 357544 480 357572 16118
rect 361132 480 361160 16546
rect 363064 13462 363092 26206
rect 364352 18358 364380 28206
rect 365272 26234 365300 30124
rect 365916 27198 365944 30124
rect 367220 29866 367248 30124
rect 367112 29838 367248 29866
rect 365904 27192 365956 27198
rect 365904 27134 365956 27140
rect 364444 26206 365300 26234
rect 364444 20534 364472 26206
rect 364432 20528 364484 20534
rect 364432 20470 364484 20476
rect 367112 19281 367140 29838
rect 367848 26234 367876 30124
rect 368480 28212 368532 28218
rect 368480 28154 368532 28160
rect 367204 26206 367876 26234
rect 367204 26081 367232 26206
rect 367190 26072 367246 26081
rect 367190 26007 367246 26016
rect 368492 23186 368520 28154
rect 369136 26897 369164 30124
rect 369780 28218 369808 30124
rect 373000 29238 373028 30124
rect 372988 29232 373040 29238
rect 372988 29174 373040 29180
rect 369768 28212 369820 28218
rect 369768 28154 369820 28160
rect 373644 27033 373672 30124
rect 375592 29866 375620 30124
rect 375392 29838 375620 29866
rect 373630 27024 373686 27033
rect 373630 26959 373686 26968
rect 369122 26888 369178 26897
rect 369122 26823 369178 26832
rect 368480 23180 368532 23186
rect 368480 23122 368532 23128
rect 367098 19272 367154 19281
rect 367098 19207 367154 19216
rect 364340 18352 364392 18358
rect 364340 18294 364392 18300
rect 375392 17678 375420 29838
rect 377508 26234 377536 30124
rect 378152 28234 378180 30124
rect 379456 29866 379484 30124
rect 379440 29838 379484 29866
rect 378152 28206 378272 28234
rect 378140 28144 378192 28150
rect 378140 28086 378192 28092
rect 376772 26206 377536 26234
rect 376772 23186 376800 26206
rect 376760 23180 376812 23186
rect 376760 23122 376812 23128
rect 375380 17672 375432 17678
rect 375380 17614 375432 17620
rect 364616 16312 364668 16318
rect 364616 16254 364668 16260
rect 363052 13456 363104 13462
rect 363052 13398 363104 13404
rect 364628 480 364656 16254
rect 367744 14952 367796 14958
rect 367744 14894 367796 14900
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 14894
rect 378152 13394 378180 28086
rect 378244 26081 378272 28206
rect 379440 28150 379468 29838
rect 381372 28898 381400 30124
rect 381360 28892 381412 28898
rect 381360 28834 381412 28840
rect 379428 28144 379480 28150
rect 379428 28086 379480 28092
rect 382016 26234 382044 30124
rect 382660 26234 382688 30124
rect 384592 26234 384620 30124
rect 385236 27169 385264 30124
rect 385222 27160 385278 27169
rect 385222 27095 385278 27104
rect 385880 26234 385908 30124
rect 386524 26234 386552 30124
rect 387828 29866 387856 30124
rect 387812 29838 387856 29866
rect 387064 28756 387116 28762
rect 387064 28698 387116 28704
rect 380912 26206 382044 26234
rect 382292 26206 382688 26234
rect 383672 26206 384620 26234
rect 385144 26206 385908 26234
rect 386432 26206 386552 26234
rect 378230 26072 378286 26081
rect 378230 26007 378286 26016
rect 378414 16144 378470 16153
rect 378414 16079 378470 16088
rect 378140 13388 378192 13394
rect 378140 13330 378192 13336
rect 371700 9036 371752 9042
rect 371700 8978 371752 8984
rect 371712 480 371740 8978
rect 375288 4888 375340 4894
rect 375288 4830 375340 4836
rect 375300 480 375328 4830
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16079
rect 380912 15026 380940 26206
rect 382292 23254 382320 26206
rect 383672 23254 383700 26206
rect 385038 25800 385094 25809
rect 385038 25735 385094 25744
rect 382280 23248 382332 23254
rect 382280 23190 382332 23196
rect 383660 23248 383712 23254
rect 383660 23190 383712 23196
rect 385052 16574 385080 25735
rect 385144 24682 385172 26206
rect 385132 24676 385184 24682
rect 385132 24618 385184 24624
rect 385052 16546 386000 16574
rect 382372 16380 382424 16386
rect 382372 16322 382424 16328
rect 380900 15020 380952 15026
rect 380900 14962 380952 14968
rect 382384 480 382412 16322
rect 385972 480 386000 16546
rect 386432 13258 386460 26206
rect 386420 13252 386472 13258
rect 386420 13194 386472 13200
rect 387076 10674 387104 28698
rect 387812 25974 387840 29838
rect 389100 27878 389128 30124
rect 389088 27872 389140 27878
rect 389088 27814 389140 27820
rect 389744 27334 389772 30124
rect 389732 27328 389784 27334
rect 389732 27270 389784 27276
rect 390388 26234 390416 30124
rect 392964 26234 392992 30124
rect 394252 26234 394280 30124
rect 398116 26234 398144 30124
rect 398760 27334 398788 30124
rect 398748 27328 398800 27334
rect 398748 27270 398800 27276
rect 399404 26234 399432 30124
rect 401336 26234 401364 30124
rect 403268 26234 403296 30124
rect 404572 29866 404600 30124
rect 409080 29866 409108 30124
rect 389284 26206 390416 26234
rect 391952 26206 392992 26234
rect 393332 26206 394280 26234
rect 397472 26206 398144 26234
rect 398852 26206 399432 26234
rect 400232 26206 401364 26234
rect 403084 26206 403296 26234
rect 404372 29838 404600 29866
rect 408512 29838 409108 29866
rect 389284 25974 389312 26206
rect 391952 26042 391980 26206
rect 391940 26036 391992 26042
rect 391940 25978 391992 25984
rect 387800 25968 387852 25974
rect 387800 25910 387852 25916
rect 389272 25968 389324 25974
rect 389272 25910 389324 25916
rect 389180 22840 389232 22846
rect 389180 22782 389232 22788
rect 391938 22808 391994 22817
rect 389192 16574 389220 22782
rect 391938 22743 391994 22752
rect 391952 16574 391980 22743
rect 389192 16546 389496 16574
rect 391952 16546 392624 16574
rect 387064 10668 387116 10674
rect 387064 10610 387116 10616
rect 389468 480 389496 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 393332 13054 393360 26206
rect 396080 25560 396132 25566
rect 396080 25502 396132 25508
rect 393320 13048 393372 13054
rect 393320 12990 393372 12996
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 25502
rect 397472 24750 397500 26206
rect 397460 24744 397512 24750
rect 397460 24686 397512 24692
rect 398852 12170 398880 26206
rect 400232 21894 400260 26206
rect 400220 21888 400272 21894
rect 400220 21830 400272 21836
rect 403084 16454 403112 26206
rect 403072 16448 403124 16454
rect 403072 16390 403124 16396
rect 403624 15836 403676 15842
rect 403624 15778 403676 15784
rect 398932 13184 398984 13190
rect 398932 13126 398984 13132
rect 398840 12164 398892 12170
rect 398840 12106 398892 12112
rect 398944 3398 398972 13126
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 403636 480 403664 15778
rect 404372 13326 404400 29838
rect 408512 23089 408540 29838
rect 409708 26790 409736 30124
rect 410352 26926 410380 30124
rect 410340 26920 410392 26926
rect 410340 26862 410392 26868
rect 409696 26784 409748 26790
rect 409696 26726 409748 26732
rect 410996 26234 411024 30124
rect 411640 26234 411668 30124
rect 416148 29073 416176 30124
rect 417452 29866 417480 30124
rect 417436 29838 417480 29866
rect 416134 29064 416190 29073
rect 416134 28999 416190 29008
rect 417436 26858 417464 29838
rect 417424 26852 417476 26858
rect 417424 26794 417476 26800
rect 420012 26234 420040 30124
rect 421316 29866 421344 30124
rect 409892 26206 411024 26234
rect 411272 26206 411668 26234
rect 419552 26206 420040 26234
rect 420932 29838 421344 29866
rect 409892 24750 409920 26206
rect 409880 24744 409932 24750
rect 409880 24686 409932 24692
rect 408498 23080 408554 23089
rect 408498 23015 408554 23024
rect 411272 21962 411300 26206
rect 411260 21956 411312 21962
rect 411260 21898 411312 21904
rect 419552 21894 419580 26206
rect 420932 21962 420960 29838
rect 421944 27169 421972 30124
rect 421930 27160 421986 27169
rect 421930 27095 421986 27104
rect 423876 26234 423904 30124
rect 426440 28212 426492 28218
rect 426440 28154 426492 28160
rect 423692 26206 423904 26234
rect 423692 26042 423720 26206
rect 423680 26036 423732 26042
rect 423680 25978 423732 25984
rect 420920 21956 420972 21962
rect 420920 21898 420972 21904
rect 419540 21888 419592 21894
rect 419540 21830 419592 21836
rect 416780 21684 416832 21690
rect 416780 21626 416832 21632
rect 407120 21616 407172 21622
rect 407120 21558 407172 21564
rect 407132 16574 407160 21558
rect 416792 16574 416820 21626
rect 426452 19242 426480 28154
rect 427096 26234 427124 30124
rect 427740 28218 427768 30124
rect 429028 28218 429056 30124
rect 427728 28212 427780 28218
rect 427728 28154 427780 28160
rect 427820 28212 427872 28218
rect 427820 28154 427872 28160
rect 429016 28212 429068 28218
rect 429016 28154 429068 28160
rect 426544 26206 427124 26234
rect 426544 23322 426572 26206
rect 426532 23316 426584 23322
rect 426532 23258 426584 23264
rect 426440 19236 426492 19242
rect 426440 19178 426492 19184
rect 427832 17814 427860 28154
rect 431604 26234 431632 30124
rect 432248 26234 432276 30124
rect 434196 29866 434224 30124
rect 430592 26206 431632 26234
rect 431972 26206 432276 26234
rect 433352 29838 434224 29866
rect 430592 25702 430620 26206
rect 430580 25696 430632 25702
rect 430580 25638 430632 25644
rect 427912 20120 427964 20126
rect 427912 20062 427964 20068
rect 427820 17808 427872 17814
rect 427820 17750 427872 17756
rect 427924 16574 427952 20062
rect 407132 16546 407252 16574
rect 416792 16546 417464 16574
rect 427924 16546 428504 16574
rect 404360 13320 404412 13326
rect 404360 13262 404412 13268
rect 407224 480 407252 16546
rect 414296 14408 414348 14414
rect 414296 14350 414348 14356
rect 410800 12980 410852 12986
rect 410800 12922 410852 12928
rect 410812 480 410840 12922
rect 414308 480 414336 14350
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 421380 7608 421432 7614
rect 421380 7550 421432 7556
rect 421392 480 421420 7550
rect 424968 4004 425020 4010
rect 424968 3946 425020 3952
rect 424980 480 425008 3946
rect 428476 480 428504 16546
rect 431972 16425 432000 26206
rect 431958 16416 432014 16425
rect 431958 16351 432014 16360
rect 433352 15774 433380 29838
rect 435468 26234 435496 30124
rect 437400 28218 437428 30124
rect 436100 28212 436152 28218
rect 436100 28154 436152 28160
rect 437388 28212 437440 28218
rect 437388 28154 437440 28160
rect 434824 26206 435496 26234
rect 434824 23322 434852 26206
rect 434812 23316 434864 23322
rect 434812 23258 434864 23264
rect 434720 22908 434772 22914
rect 434720 22850 434772 22856
rect 434732 16574 434760 22850
rect 436112 20369 436140 28154
rect 439332 26234 439360 30124
rect 440620 26234 440648 30124
rect 441264 27402 441292 30124
rect 443196 29306 443224 30124
rect 443184 29300 443236 29306
rect 443184 29242 443236 29248
rect 444380 28212 444432 28218
rect 444380 28154 444432 28160
rect 441252 27396 441304 27402
rect 441252 27338 441304 27344
rect 438872 26206 439360 26234
rect 440344 26206 440648 26234
rect 436098 20360 436154 20369
rect 436098 20295 436154 20304
rect 438872 17678 438900 26206
rect 440344 18562 440372 26206
rect 440332 18556 440384 18562
rect 440332 18498 440384 18504
rect 444392 17950 444420 28154
rect 444484 23089 444512 30124
rect 445128 28218 445156 30124
rect 445116 28212 445168 28218
rect 445116 28154 445168 28160
rect 444470 23080 444526 23089
rect 444470 23015 444526 23024
rect 445772 17950 445800 30124
rect 447076 29918 447104 30124
rect 445852 29912 445904 29918
rect 445852 29854 445904 29860
rect 447064 29912 447116 29918
rect 447064 29854 447116 29860
rect 445864 22250 445892 29854
rect 448348 28218 448376 30124
rect 448992 28234 449020 30124
rect 447140 28212 447192 28218
rect 447140 28154 447192 28160
rect 448336 28212 448388 28218
rect 448336 28154 448388 28160
rect 448532 28206 449020 28234
rect 447152 23050 447180 28154
rect 447140 23044 447192 23050
rect 447140 22986 447192 22992
rect 445864 22222 446076 22250
rect 445850 19816 445906 19825
rect 445850 19751 445906 19760
rect 445864 19378 445892 19751
rect 446048 19689 446076 22222
rect 446034 19680 446090 19689
rect 446034 19615 446090 19624
rect 445852 19372 445904 19378
rect 445852 19314 445904 19320
rect 444380 17944 444432 17950
rect 444380 17886 444432 17892
rect 445760 17944 445812 17950
rect 445760 17886 445812 17892
rect 448532 17814 448560 28206
rect 449636 26234 449664 30124
rect 450940 29866 450968 30124
rect 448624 26206 449664 26234
rect 449912 29838 450968 29866
rect 448624 22030 448652 26206
rect 448612 22024 448664 22030
rect 448612 21966 448664 21972
rect 449912 20534 449940 29838
rect 451568 28830 451596 30124
rect 451556 28824 451608 28830
rect 451556 28766 451608 28772
rect 452856 27033 452884 30124
rect 459312 29918 459340 30124
rect 458180 29912 458232 29918
rect 458180 29854 458232 29860
rect 459300 29912 459352 29918
rect 459300 29854 459352 29860
rect 452842 27024 452898 27033
rect 452842 26959 452898 26968
rect 458192 20670 458220 29854
rect 459940 26738 459968 30124
rect 459572 26710 459968 26738
rect 458180 20664 458232 20670
rect 458180 20606 458232 20612
rect 449900 20528 449952 20534
rect 449900 20470 449952 20476
rect 459572 20466 459600 26710
rect 460584 26234 460612 30124
rect 461228 28234 461256 30124
rect 459664 26206 460612 26234
rect 460952 28206 461256 28234
rect 459664 21185 459692 26206
rect 459650 21176 459706 21185
rect 459650 21111 459706 21120
rect 459560 20460 459612 20466
rect 459560 20402 459612 20408
rect 452660 20188 452712 20194
rect 452660 20130 452712 20136
rect 448520 17808 448572 17814
rect 448520 17750 448572 17756
rect 438860 17672 438912 17678
rect 438860 17614 438912 17620
rect 452672 16574 452700 20130
rect 460952 17202 460980 28206
rect 461872 26234 461900 30124
rect 462516 26234 462544 30124
rect 463820 29866 463848 30124
rect 463804 29838 463848 29866
rect 463700 28212 463752 28218
rect 463700 28154 463752 28160
rect 461044 26206 461900 26234
rect 462332 26206 462544 26234
rect 461044 19786 461072 26206
rect 462332 20602 462360 26206
rect 462320 20596 462372 20602
rect 462320 20538 462372 20544
rect 463712 20330 463740 28154
rect 463804 21865 463832 29838
rect 464448 28218 464476 30124
rect 464436 28212 464488 28218
rect 464436 28154 464488 28160
rect 463790 21856 463846 21865
rect 463790 21791 463846 21800
rect 463700 20324 463752 20330
rect 463700 20266 463752 20272
rect 461032 19780 461084 19786
rect 461032 19722 461084 19728
rect 465092 19174 465120 30124
rect 465736 28234 465764 30124
rect 465184 28206 465764 28234
rect 465184 24614 465212 28206
rect 466380 26234 466408 30124
rect 465276 26206 466408 26234
rect 465172 24608 465224 24614
rect 465172 24550 465224 24556
rect 465276 24478 465304 26206
rect 465264 24472 465316 24478
rect 465264 24414 465316 24420
rect 468956 23361 468984 30124
rect 468942 23352 468998 23361
rect 468942 23287 468998 23296
rect 469600 22094 469628 30124
rect 470888 26110 470916 30124
rect 473464 26722 473492 30124
rect 474752 30002 474780 30124
rect 474660 29974 474780 30002
rect 474660 29578 474688 29974
rect 476056 29918 476084 30124
rect 474740 29912 474792 29918
rect 474740 29854 474792 29860
rect 476044 29912 476096 29918
rect 476044 29854 476096 29860
rect 474648 29572 474700 29578
rect 474648 29514 474700 29520
rect 474004 28552 474056 28558
rect 474004 28494 474056 28500
rect 473452 26716 473504 26722
rect 473452 26658 473504 26664
rect 470876 26104 470928 26110
rect 470876 26046 470928 26052
rect 469232 22066 469628 22094
rect 469232 20602 469260 22066
rect 470600 21752 470652 21758
rect 470600 21694 470652 21700
rect 469220 20596 469272 20602
rect 469220 20538 469272 20544
rect 465080 19168 465132 19174
rect 465080 19110 465132 19116
rect 460940 17196 460992 17202
rect 460940 17138 460992 17144
rect 434732 16546 435128 16574
rect 452672 16546 453344 16574
rect 433340 15768 433392 15774
rect 433340 15710 433392 15716
rect 432052 6248 432104 6254
rect 432052 6190 432104 6196
rect 432064 480 432092 6190
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 446220 6520 446272 6526
rect 446220 6462 446272 6468
rect 442632 6384 442684 6390
rect 442632 6326 442684 6332
rect 439136 6316 439188 6322
rect 439136 6258 439188 6264
rect 439148 480 439176 6258
rect 442644 480 442672 6326
rect 446232 480 446260 6462
rect 449808 6452 449860 6458
rect 449808 6394 449860 6400
rect 449820 480 449848 6394
rect 453316 480 453344 16546
rect 456892 12912 456944 12918
rect 456892 12854 456944 12860
rect 456904 480 456932 12854
rect 467472 12096 467524 12102
rect 467472 12038 467524 12044
rect 460388 6724 460440 6730
rect 460388 6666 460440 6672
rect 460400 480 460428 6666
rect 463976 6588 464028 6594
rect 463976 6530 464028 6536
rect 463988 480 464016 6530
rect 467484 480 467512 12038
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 21694
rect 474016 14346 474044 28494
rect 474752 20262 474780 29854
rect 474832 29572 474884 29578
rect 474832 29514 474884 29520
rect 474844 28218 474872 29514
rect 476684 28234 476712 30124
rect 474832 28212 474884 28218
rect 474832 28154 474884 28160
rect 476132 28206 476712 28234
rect 476132 21729 476160 28206
rect 477328 26234 477356 30124
rect 478616 26234 478644 30124
rect 479260 28801 479288 30124
rect 480564 29866 480592 30124
rect 480272 29838 480592 29866
rect 479246 28792 479302 28801
rect 479246 28727 479302 28736
rect 476224 26206 477356 26234
rect 477604 26206 478644 26234
rect 480272 26217 480300 29838
rect 481836 29073 481864 30124
rect 481822 29064 481878 29073
rect 481822 28999 481878 29008
rect 483124 28082 483152 30124
rect 484428 29866 484456 30124
rect 484428 29838 484624 29866
rect 484400 28280 484452 28286
rect 484400 28222 484452 28228
rect 483112 28076 483164 28082
rect 483112 28018 483164 28024
rect 480258 26208 480314 26217
rect 476224 26110 476252 26206
rect 476212 26104 476264 26110
rect 476212 26046 476264 26052
rect 477500 25628 477552 25634
rect 477500 25570 477552 25576
rect 476118 21720 476174 21729
rect 476118 21655 476174 21664
rect 474740 20256 474792 20262
rect 474740 20198 474792 20204
rect 477512 16574 477540 25570
rect 477604 20398 477632 26206
rect 480258 26143 480314 26152
rect 484412 21185 484440 28222
rect 484492 28144 484544 28150
rect 484492 28086 484544 28092
rect 484504 22982 484532 28086
rect 484596 25401 484624 29838
rect 485056 28286 485084 30124
rect 485044 28280 485096 28286
rect 485044 28222 485096 28228
rect 485700 28150 485728 30124
rect 487632 28801 487660 30124
rect 487618 28792 487674 28801
rect 487618 28727 487674 28736
rect 485688 28144 485740 28150
rect 485688 28086 485740 28092
rect 489564 26234 489592 30124
rect 491496 26234 491524 30124
rect 492800 29866 492828 30124
rect 492784 29838 492828 29866
rect 492784 27538 492812 29838
rect 493428 28558 493456 30124
rect 493416 28552 493468 28558
rect 493416 28494 493468 28500
rect 492772 27532 492824 27538
rect 492772 27474 492824 27480
rect 488552 26206 489592 26234
rect 491312 26206 491524 26234
rect 484582 25392 484638 25401
rect 484582 25327 484638 25336
rect 484492 22976 484544 22982
rect 484492 22918 484544 22924
rect 488552 22030 488580 26206
rect 491312 22545 491340 26206
rect 494072 26178 494100 30124
rect 499224 26234 499252 30124
rect 502340 27804 502392 27810
rect 502340 27746 502392 27752
rect 498212 26206 499252 26234
rect 494060 26172 494112 26178
rect 494060 26114 494112 26120
rect 498212 22710 498240 26206
rect 498200 22704 498252 22710
rect 498200 22646 498252 22652
rect 491298 22536 491354 22545
rect 491298 22471 491354 22480
rect 488540 22024 488592 22030
rect 488540 21966 488592 21972
rect 484398 21176 484454 21185
rect 484398 21111 484454 21120
rect 477592 20392 477644 20398
rect 477592 20334 477644 20340
rect 502352 16574 502380 27746
rect 502444 24342 502472 30124
rect 503088 26234 503116 30124
rect 504376 28778 504404 30124
rect 505680 29866 505708 30124
rect 502536 26206 503116 26234
rect 503732 28750 504404 28778
rect 505664 29838 505708 29866
rect 502536 24546 502564 26206
rect 502524 24540 502576 24546
rect 502524 24482 502576 24488
rect 503732 24410 503760 28750
rect 504180 28620 504232 28626
rect 504180 28562 504232 28568
rect 503720 24404 503772 24410
rect 503720 24346 503772 24352
rect 502432 24336 502484 24342
rect 502432 24278 502484 24284
rect 503732 23526 503760 24346
rect 503720 23520 503772 23526
rect 503720 23462 503772 23468
rect 504192 19922 504220 28562
rect 505664 28286 505692 29838
rect 505652 28280 505704 28286
rect 505652 28222 505704 28228
rect 506308 28150 506336 30124
rect 506952 29374 506980 30124
rect 509544 29866 509572 30124
rect 509528 29838 509572 29866
rect 509528 29442 509556 29838
rect 509516 29436 509568 29442
rect 509516 29378 509568 29384
rect 506940 29368 506992 29374
rect 506940 29310 506992 29316
rect 505100 28144 505152 28150
rect 505100 28086 505152 28092
rect 506296 28144 506348 28150
rect 506296 28086 506348 28092
rect 506388 28144 506440 28150
rect 506388 28086 506440 28092
rect 504364 23520 504416 23526
rect 504364 23462 504416 23468
rect 504180 19916 504232 19922
rect 504180 19858 504232 19864
rect 477512 16546 478184 16574
rect 502352 16546 503024 16574
rect 474004 14340 474056 14346
rect 474004 14282 474056 14288
rect 474554 6624 474610 6633
rect 474554 6559 474610 6568
rect 474568 480 474596 6559
rect 478156 480 478184 16546
rect 499396 6792 499448 6798
rect 499396 6734 499448 6740
rect 485228 6656 485280 6662
rect 485228 6598 485280 6604
rect 481730 6488 481786 6497
rect 481730 6423 481786 6432
rect 481744 480 481772 6423
rect 485240 480 485268 6598
rect 492312 4140 492364 4146
rect 492312 4082 492364 4088
rect 488816 4072 488868 4078
rect 488816 4014 488868 4020
rect 488828 480 488856 4014
rect 492324 480 492352 4082
rect 495900 3392 495952 3398
rect 495900 3334 495952 3340
rect 495912 480 495940 3334
rect 499408 480 499436 6734
rect 502996 480 503024 16546
rect 504376 11830 504404 23462
rect 505112 21214 505140 28086
rect 506400 27810 506428 28086
rect 506388 27804 506440 27810
rect 506388 27746 506440 27752
rect 510172 26234 510200 30124
rect 510816 26234 510844 30124
rect 511264 28960 511316 28966
rect 511264 28902 511316 28908
rect 509252 26206 510200 26234
rect 510632 26206 510844 26234
rect 509252 26178 509280 26206
rect 509240 26172 509292 26178
rect 509240 26114 509292 26120
rect 510632 24070 510660 26206
rect 510620 24064 510672 24070
rect 510620 24006 510672 24012
rect 505100 21208 505152 21214
rect 505100 21150 505152 21156
rect 511276 17134 511304 28902
rect 511460 27402 511488 30124
rect 512104 28626 512132 30124
rect 514052 29866 514080 30124
rect 514036 29838 514080 29866
rect 514036 29510 514064 29838
rect 515968 29578 515996 30124
rect 515956 29572 516008 29578
rect 515956 29514 516008 29520
rect 514024 29504 514076 29510
rect 514024 29446 514076 29452
rect 512092 28620 512144 28626
rect 512092 28562 512144 28568
rect 511448 27396 511500 27402
rect 511448 27338 511500 27344
rect 516612 26722 516640 30124
rect 519188 29481 519216 30124
rect 519174 29472 519230 29481
rect 519174 29407 519230 29416
rect 516600 26716 516652 26722
rect 516600 26658 516652 26664
rect 519832 26234 519860 30124
rect 520476 26654 520504 30124
rect 521120 29617 521148 30124
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 523052 28694 523080 30124
rect 523040 28688 523092 28694
rect 523040 28630 523092 28636
rect 522304 28416 522356 28422
rect 522304 28358 522356 28364
rect 520464 26648 520516 26654
rect 520464 26590 520516 26596
rect 518912 26206 519860 26234
rect 513380 25492 513432 25498
rect 513380 25434 513432 25440
rect 511264 17128 511316 17134
rect 511264 17070 511316 17076
rect 504364 11824 504416 11830
rect 504364 11766 504416 11772
rect 506480 6860 506532 6866
rect 506480 6802 506532 6808
rect 506492 480 506520 6802
rect 510068 3324 510120 3330
rect 510068 3266 510120 3272
rect 510080 480 510108 3266
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 25434
rect 516140 25356 516192 25362
rect 516140 25298 516192 25304
rect 516152 16574 516180 25298
rect 518912 23361 518940 26206
rect 520280 25424 520332 25430
rect 520280 25366 520332 25372
rect 518898 23352 518954 23361
rect 518898 23287 518954 23296
rect 516152 16546 517192 16574
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 25366
rect 522316 16590 522344 28358
rect 523040 26240 523092 26246
rect 523696 26234 523724 30124
rect 524340 26625 524368 30124
rect 525628 27577 525656 30124
rect 526932 29918 526960 30124
rect 525800 29912 525852 29918
rect 525800 29854 525852 29860
rect 526920 29912 526972 29918
rect 526920 29854 526972 29860
rect 525614 27568 525670 27577
rect 525614 27503 525670 27512
rect 524326 26616 524382 26625
rect 524326 26551 524382 26560
rect 523092 26206 523724 26234
rect 523040 26182 523092 26188
rect 523040 21820 523092 21826
rect 523040 21762 523092 21768
rect 522304 16584 522356 16590
rect 523052 16574 523080 21762
rect 525812 20505 525840 29854
rect 527178 28520 527234 28529
rect 527178 28455 527234 28464
rect 527824 28484 527876 28490
rect 527192 28422 527220 28455
rect 527824 28426 527876 28432
rect 527180 28416 527232 28422
rect 527180 28358 527232 28364
rect 527180 28008 527232 28014
rect 527180 27950 527232 27956
rect 527192 20670 527220 27950
rect 527180 20664 527232 20670
rect 527180 20606 527232 20612
rect 525798 20496 525854 20505
rect 525798 20431 525854 20440
rect 527836 19310 527864 28426
rect 528204 27606 528232 30124
rect 528848 28529 528876 30124
rect 528834 28520 528890 28529
rect 529492 28490 529520 30124
rect 531424 29646 531452 30124
rect 531412 29640 531464 29646
rect 531412 29582 531464 29588
rect 531228 29028 531280 29034
rect 531228 28970 531280 28976
rect 531240 28762 531268 28970
rect 531228 28756 531280 28762
rect 531228 28698 531280 28704
rect 528834 28455 528890 28464
rect 529480 28484 529532 28490
rect 529480 28426 529532 28432
rect 528560 28348 528612 28354
rect 528560 28290 528612 28296
rect 528192 27600 528244 27606
rect 528192 27542 528244 27548
rect 528572 22001 528600 28290
rect 532068 27305 532096 30124
rect 534816 29640 534868 29646
rect 534816 29582 534868 29588
rect 535460 29640 535512 29646
rect 535460 29582 535512 29588
rect 534828 29102 534856 29582
rect 535472 29238 535500 29582
rect 535460 29232 535512 29238
rect 535460 29174 535512 29180
rect 534816 29096 534868 29102
rect 534816 29038 534868 29044
rect 536576 27985 536604 30124
rect 536840 29708 536892 29714
rect 536840 29650 536892 29656
rect 536852 28082 536880 29650
rect 537220 28422 537248 30124
rect 537864 29238 537892 30124
rect 539168 29866 539196 30124
rect 538324 29838 539196 29866
rect 539506 29880 539562 29889
rect 537852 29232 537904 29238
rect 537852 29174 537904 29180
rect 537208 28416 537260 28422
rect 537208 28358 537260 28364
rect 536840 28076 536892 28082
rect 536840 28018 536892 28024
rect 536562 27976 536618 27985
rect 536562 27911 536618 27920
rect 534724 27872 534776 27878
rect 534724 27814 534776 27820
rect 532054 27296 532110 27305
rect 532054 27231 532110 27240
rect 534736 24818 534764 27814
rect 538220 26240 538272 26246
rect 538220 26182 538272 26188
rect 534724 24812 534776 24818
rect 534724 24754 534776 24760
rect 528558 21992 528614 22001
rect 528558 21927 528614 21936
rect 533344 19848 533396 19854
rect 533344 19790 533396 19796
rect 527824 19304 527876 19310
rect 527824 19246 527876 19252
rect 523052 16546 523816 16574
rect 522304 16526 522356 16532
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 531318 3904 531374 3913
rect 533356 3874 533384 19790
rect 531318 3839 531374 3848
rect 533344 3868 533396 3874
rect 527824 3188 527876 3194
rect 527824 3130 527876 3136
rect 527836 480 527864 3130
rect 531332 480 531360 3839
rect 533344 3810 533396 3816
rect 534908 3868 534960 3874
rect 534908 3810 534960 3816
rect 534920 480 534948 3810
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 26182
rect 538324 20641 538352 29838
rect 539506 29815 539562 29824
rect 539520 29034 539548 29815
rect 539508 29028 539560 29034
rect 539508 28970 539560 28976
rect 539506 28928 539562 28937
rect 539506 28863 539562 28872
rect 539520 28354 539548 28863
rect 539508 28348 539560 28354
rect 539508 28290 539560 28296
rect 538310 20632 538366 20641
rect 538310 20567 538366 20576
rect 540072 20330 540100 155858
rect 540152 149932 540204 149938
rect 540152 149874 540204 149880
rect 540164 149841 540192 149874
rect 540150 149832 540206 149841
rect 540150 149767 540206 149776
rect 540256 149161 540284 234223
rect 540428 233164 540480 233170
rect 540428 233106 540480 233112
rect 540336 230444 540388 230450
rect 540336 230386 540388 230392
rect 540348 154714 540376 230386
rect 540440 160970 540468 233106
rect 540520 230104 540572 230110
rect 540520 230046 540572 230052
rect 540532 171134 540560 230046
rect 540532 171106 540836 171134
rect 540440 160942 540652 160970
rect 540624 154834 540652 160942
rect 540808 157334 540836 171106
rect 541072 159724 541124 159730
rect 541072 159666 541124 159672
rect 540808 157306 540928 157334
rect 540612 154828 540664 154834
rect 540612 154770 540664 154776
rect 540348 154686 540744 154714
rect 540612 154624 540664 154630
rect 540612 154566 540664 154572
rect 540520 154556 540572 154562
rect 540520 154498 540572 154504
rect 540336 152448 540388 152454
rect 540336 152390 540388 152396
rect 540242 149152 540298 149161
rect 540242 149087 540298 149096
rect 540150 147384 540206 147393
rect 540150 147319 540206 147328
rect 540164 144906 540192 147319
rect 540348 147257 540376 152390
rect 540428 150068 540480 150074
rect 540428 150010 540480 150016
rect 540440 149297 540468 150010
rect 540426 149288 540482 149297
rect 540426 149223 540482 149232
rect 540426 147656 540482 147665
rect 540426 147591 540482 147600
rect 540334 147248 540390 147257
rect 540334 147183 540390 147192
rect 540334 146976 540390 146985
rect 540334 146911 540390 146920
rect 540152 144900 540204 144906
rect 540152 144842 540204 144848
rect 540348 139641 540376 146911
rect 540334 139632 540390 139641
rect 540334 139567 540390 139576
rect 540440 137358 540468 147591
rect 540532 146130 540560 154498
rect 540624 150346 540652 154566
rect 540612 150340 540664 150346
rect 540612 150282 540664 150288
rect 540610 150104 540666 150113
rect 540610 150039 540666 150048
rect 540520 146124 540572 146130
rect 540520 146066 540572 146072
rect 540520 144220 540572 144226
rect 540520 144162 540572 144168
rect 540428 137352 540480 137358
rect 540428 137294 540480 137300
rect 540244 137284 540296 137290
rect 540244 137226 540296 137232
rect 540150 122768 540206 122777
rect 540150 122703 540206 122712
rect 540164 114209 540192 122703
rect 540150 114200 540206 114209
rect 540150 114135 540206 114144
rect 540152 79348 540204 79354
rect 540152 79290 540204 79296
rect 540060 20324 540112 20330
rect 540060 20266 540112 20272
rect 540164 10810 540192 79290
rect 540256 14346 540284 137226
rect 540336 126268 540388 126274
rect 540336 126210 540388 126216
rect 540348 19038 540376 126210
rect 540532 114374 540560 144162
rect 540624 143410 540652 150039
rect 540716 146946 540744 154686
rect 540796 153808 540848 153814
rect 540796 153750 540848 153756
rect 540704 146940 540756 146946
rect 540704 146882 540756 146888
rect 540704 146260 540756 146266
rect 540704 146202 540756 146208
rect 540612 143404 540664 143410
rect 540612 143346 540664 143352
rect 540612 139528 540664 139534
rect 540612 139470 540664 139476
rect 540624 122834 540652 139470
rect 540716 130898 540744 146202
rect 540808 143478 540836 153750
rect 540900 147674 540928 157306
rect 540980 150476 541032 150482
rect 540980 150418 541032 150424
rect 540992 150249 541020 150418
rect 540978 150240 541034 150249
rect 540978 150175 541034 150184
rect 540900 147646 541020 147674
rect 540992 146266 541020 147646
rect 540980 146260 541032 146266
rect 540980 146202 541032 146208
rect 540888 143540 540940 143546
rect 540888 143482 540940 143488
rect 540796 143472 540848 143478
rect 540796 143414 540848 143420
rect 540796 139596 540848 139602
rect 540796 139538 540848 139544
rect 540808 135153 540836 139538
rect 540900 139534 540928 143482
rect 540888 139528 540940 139534
rect 540888 139470 540940 139476
rect 540978 139496 541034 139505
rect 540978 139431 541034 139440
rect 540992 137442 541020 139431
rect 540900 137414 541020 137442
rect 540794 135144 540850 135153
rect 540794 135079 540850 135088
rect 540796 131096 540848 131102
rect 540796 131038 540848 131044
rect 540704 130892 540756 130898
rect 540704 130834 540756 130840
rect 540808 125662 540836 131038
rect 540900 129849 540928 137414
rect 540980 137352 541032 137358
rect 540980 137294 541032 137300
rect 540992 131170 541020 137294
rect 540980 131164 541032 131170
rect 540980 131106 541032 131112
rect 540886 129840 540942 129849
rect 540886 129775 540942 129784
rect 540980 127628 541032 127634
rect 540980 127570 541032 127576
rect 540796 125656 540848 125662
rect 540796 125598 540848 125604
rect 540992 125474 541020 127570
rect 540900 125446 541020 125474
rect 540624 122806 540836 122834
rect 540704 117564 540756 117570
rect 540704 117506 540756 117512
rect 540520 114368 540572 114374
rect 540520 114310 540572 114316
rect 540612 114028 540664 114034
rect 540612 113970 540664 113976
rect 540520 98048 540572 98054
rect 540520 97990 540572 97996
rect 540426 86864 540482 86873
rect 540426 86799 540482 86808
rect 540440 79354 540468 86799
rect 540532 85814 540560 97990
rect 540624 90001 540652 113970
rect 540716 98870 540744 117506
rect 540808 107642 540836 122806
rect 540900 120154 540928 125446
rect 540888 120148 540940 120154
rect 540888 120090 540940 120096
rect 540888 110560 540940 110566
rect 540888 110502 540940 110508
rect 540796 107636 540848 107642
rect 540796 107578 540848 107584
rect 540796 107500 540848 107506
rect 540796 107442 540848 107448
rect 540704 98864 540756 98870
rect 540704 98806 540756 98812
rect 540610 89992 540666 90001
rect 540610 89927 540666 89936
rect 540612 88324 540664 88330
rect 540612 88266 540664 88272
rect 540520 85808 540572 85814
rect 540520 85750 540572 85756
rect 540520 82952 540572 82958
rect 540520 82894 540572 82900
rect 540428 79348 540480 79354
rect 540428 79290 540480 79296
rect 540532 64874 540560 82894
rect 540624 75886 540652 88266
rect 540808 85542 540836 107442
rect 540900 102338 540928 110502
rect 540888 102332 540940 102338
rect 540888 102274 540940 102280
rect 540980 100020 541032 100026
rect 540980 99962 541032 99968
rect 540888 89820 540940 89826
rect 540888 89762 540940 89768
rect 540796 85536 540848 85542
rect 540796 85478 540848 85484
rect 540612 75880 540664 75886
rect 540612 75822 540664 75828
rect 540900 69018 540928 89762
rect 540888 69012 540940 69018
rect 540888 68954 540940 68960
rect 540612 66700 540664 66706
rect 540612 66642 540664 66648
rect 540440 64846 540560 64874
rect 540336 19032 540388 19038
rect 540336 18974 540388 18980
rect 540244 14340 540296 14346
rect 540244 14282 540296 14288
rect 540152 10804 540204 10810
rect 540152 10746 540204 10752
rect 540440 10674 540468 64846
rect 540624 45554 540652 66642
rect 540532 45526 540652 45554
rect 540532 14890 540560 45526
rect 540888 36780 540940 36786
rect 540888 36722 540940 36728
rect 540900 31657 540928 36722
rect 540886 31648 540942 31657
rect 540886 31583 540942 31592
rect 540888 31136 540940 31142
rect 540888 31078 540940 31084
rect 540704 31068 540756 31074
rect 540704 31010 540756 31016
rect 540612 30320 540664 30326
rect 540612 30262 540664 30268
rect 540520 14884 540572 14890
rect 540520 14826 540572 14832
rect 540624 10878 540652 30262
rect 540716 25702 540744 31010
rect 540900 26790 540928 31078
rect 540888 26784 540940 26790
rect 540888 26726 540940 26732
rect 540704 25696 540756 25702
rect 540704 25638 540756 25644
rect 540612 10872 540664 10878
rect 540612 10814 540664 10820
rect 540428 10668 540480 10674
rect 540428 10610 540480 10616
rect 540992 6914 541020 99962
rect 541084 24478 541112 159666
rect 541176 144226 541204 238002
rect 541900 237516 541952 237522
rect 541900 237458 541952 237464
rect 541624 235816 541676 235822
rect 541624 235758 541676 235764
rect 541254 235512 541310 235521
rect 541254 235447 541310 235456
rect 541268 151745 541296 235447
rect 541440 233980 541492 233986
rect 541440 233922 541492 233928
rect 541348 157344 541400 157350
rect 541348 157286 541400 157292
rect 541254 151736 541310 151745
rect 541254 151671 541310 151680
rect 541256 146668 541308 146674
rect 541256 146610 541308 146616
rect 541164 144220 541216 144226
rect 541164 144162 541216 144168
rect 541164 142180 541216 142186
rect 541164 142122 541216 142128
rect 541176 139466 541204 142122
rect 541268 139534 541296 146610
rect 541256 139528 541308 139534
rect 541256 139470 541308 139476
rect 541164 139460 541216 139466
rect 541164 139402 541216 139408
rect 541164 107636 541216 107642
rect 541164 107578 541216 107584
rect 541072 24472 541124 24478
rect 541072 24414 541124 24420
rect 541176 16318 541204 107578
rect 541360 101561 541388 157286
rect 541452 133521 541480 233922
rect 541530 147928 541586 147937
rect 541530 147863 541586 147872
rect 541544 147558 541572 147863
rect 541532 147552 541584 147558
rect 541532 147494 541584 147500
rect 541636 144838 541664 235758
rect 541716 234388 541768 234394
rect 541716 234330 541768 234336
rect 541728 147694 541756 234330
rect 541808 230172 541860 230178
rect 541808 230114 541860 230120
rect 541716 147688 541768 147694
rect 541716 147630 541768 147636
rect 541820 146334 541848 230114
rect 541912 198898 541940 237458
rect 541900 198892 541952 198898
rect 541900 198834 541952 198840
rect 542372 197334 542400 240094
rect 543924 238128 543976 238134
rect 543924 238070 543976 238076
rect 544014 238096 544070 238105
rect 543832 233980 543884 233986
rect 543832 233922 543884 233928
rect 542544 233028 542596 233034
rect 542544 232970 542596 232976
rect 542452 224256 542504 224262
rect 542452 224198 542504 224204
rect 542360 197328 542412 197334
rect 542360 197270 542412 197276
rect 542268 152584 542320 152590
rect 542268 152526 542320 152532
rect 541992 152380 542044 152386
rect 541992 152322 542044 152328
rect 541900 151020 541952 151026
rect 541900 150962 541952 150968
rect 541808 146328 541860 146334
rect 541808 146270 541860 146276
rect 541716 145580 541768 145586
rect 541716 145522 541768 145528
rect 541624 144832 541676 144838
rect 541624 144774 541676 144780
rect 541532 140888 541584 140894
rect 541532 140830 541584 140836
rect 541438 133512 541494 133521
rect 541438 133447 541494 133456
rect 541440 115456 541492 115462
rect 541440 115398 541492 115404
rect 541346 101552 541402 101561
rect 541346 101487 541402 101496
rect 541452 98734 541480 115398
rect 541544 104786 541572 140830
rect 541728 139602 541756 145522
rect 541716 139596 541768 139602
rect 541716 139538 541768 139544
rect 541808 139460 541860 139466
rect 541808 139402 541860 139408
rect 541716 131300 541768 131306
rect 541716 131242 541768 131248
rect 541624 126880 541676 126886
rect 541624 126822 541676 126828
rect 541532 104780 541584 104786
rect 541532 104722 541584 104728
rect 541440 98728 541492 98734
rect 541440 98670 541492 98676
rect 541254 89856 541310 89865
rect 541254 89791 541310 89800
rect 541268 75857 541296 89791
rect 541254 75848 541310 75857
rect 541254 75783 541310 75792
rect 541164 16312 541216 16318
rect 541164 16254 541216 16260
rect 540992 6886 541572 6914
rect 541544 3482 541572 6886
rect 541636 6730 541664 126822
rect 541728 30569 541756 131242
rect 541820 116618 541848 139402
rect 541912 126954 541940 150962
rect 542004 143342 542032 152322
rect 542280 146282 542308 152526
rect 542176 146260 542228 146266
rect 542280 146254 542400 146282
rect 542176 146202 542228 146208
rect 542084 143948 542136 143954
rect 542084 143890 542136 143896
rect 541992 143336 542044 143342
rect 541992 143278 542044 143284
rect 541990 138136 542046 138145
rect 541990 138071 542046 138080
rect 542004 137426 542032 138071
rect 541992 137420 542044 137426
rect 541992 137362 542044 137368
rect 541992 131232 542044 131238
rect 541992 131174 542044 131180
rect 542004 127650 542032 131174
rect 542096 128246 542124 143890
rect 542188 141166 542216 146202
rect 542176 141160 542228 141166
rect 542176 141102 542228 141108
rect 542268 140820 542320 140826
rect 542268 140762 542320 140768
rect 542176 138032 542228 138038
rect 542176 137974 542228 137980
rect 542188 131170 542216 137974
rect 542280 133890 542308 140762
rect 542268 133884 542320 133890
rect 542268 133826 542320 133832
rect 542268 133748 542320 133754
rect 542268 133690 542320 133696
rect 542176 131164 542228 131170
rect 542176 131106 542228 131112
rect 542084 128240 542136 128246
rect 542084 128182 542136 128188
rect 542004 127622 542216 127650
rect 541900 126948 541952 126954
rect 541900 126890 541952 126896
rect 541992 125656 542044 125662
rect 541992 125598 542044 125604
rect 541808 116612 541860 116618
rect 541808 116554 541860 116560
rect 541808 115932 541860 115938
rect 541808 115874 541860 115880
rect 541714 30560 541770 30569
rect 541714 30495 541770 30504
rect 541820 17678 541848 115874
rect 542004 115530 542032 125598
rect 542084 125588 542136 125594
rect 542084 125530 542136 125536
rect 541992 115524 542044 115530
rect 541992 115466 542044 115472
rect 542096 114510 542124 125530
rect 542084 114504 542136 114510
rect 542084 114446 542136 114452
rect 542188 108390 542216 127622
rect 542280 125730 542308 133690
rect 542268 125724 542320 125730
rect 542268 125666 542320 125672
rect 542372 115462 542400 146254
rect 542360 115456 542412 115462
rect 542360 115398 542412 115404
rect 542360 114504 542412 114510
rect 542360 114446 542412 114452
rect 542268 113144 542320 113150
rect 542268 113086 542320 113092
rect 542280 109002 542308 113086
rect 542268 108996 542320 109002
rect 542268 108938 542320 108944
rect 542176 108384 542228 108390
rect 542176 108326 542228 108332
rect 542176 108248 542228 108254
rect 542176 108190 542228 108196
rect 541900 104168 541952 104174
rect 541900 104110 541952 104116
rect 541808 17672 541860 17678
rect 541808 17614 541860 17620
rect 541912 15842 541940 104110
rect 542188 102270 542216 108190
rect 542372 104922 542400 114446
rect 542360 104916 542412 104922
rect 542360 104858 542412 104864
rect 542176 102264 542228 102270
rect 542176 102206 542228 102212
rect 542268 102196 542320 102202
rect 542268 102138 542320 102144
rect 542176 102128 542228 102134
rect 542176 102070 542228 102076
rect 541992 98728 542044 98734
rect 541992 98670 542044 98676
rect 541900 15836 541952 15842
rect 541900 15778 541952 15784
rect 542004 12306 542032 98670
rect 542188 98054 542216 102070
rect 542176 98048 542228 98054
rect 542176 97990 542228 97996
rect 542280 95198 542308 102138
rect 542360 98864 542412 98870
rect 542360 98806 542412 98812
rect 542268 95192 542320 95198
rect 542268 95134 542320 95140
rect 542372 93854 542400 98806
rect 542464 95441 542492 224198
rect 542556 147014 542584 232970
rect 543096 230036 543148 230042
rect 543096 229978 543148 229984
rect 543004 227180 543056 227186
rect 543004 227122 543056 227128
rect 542820 215960 542872 215966
rect 542820 215902 542872 215908
rect 542636 156528 542688 156534
rect 542636 156470 542688 156476
rect 542544 147008 542596 147014
rect 542544 146950 542596 146956
rect 542542 144800 542598 144809
rect 542542 144735 542598 144744
rect 542556 140865 542584 144735
rect 542542 140856 542598 140865
rect 542542 140791 542598 140800
rect 542544 133884 542596 133890
rect 542544 133826 542596 133832
rect 542450 95432 542506 95441
rect 542450 95367 542506 95376
rect 542280 93826 542400 93854
rect 542280 90914 542308 93826
rect 542268 90908 542320 90914
rect 542268 90850 542320 90856
rect 542360 84652 542412 84658
rect 542360 84594 542412 84600
rect 542372 84561 542400 84594
rect 542358 84552 542414 84561
rect 542358 84487 542414 84496
rect 542452 75880 542504 75886
rect 542452 75822 542504 75828
rect 542176 73228 542228 73234
rect 542176 73170 542228 73176
rect 542084 70644 542136 70650
rect 542084 70586 542136 70592
rect 542096 15094 542124 70586
rect 542188 17406 542216 73170
rect 542358 42392 542414 42401
rect 542358 42327 542360 42336
rect 542412 42327 542414 42336
rect 542360 42298 542412 42304
rect 542358 37632 542414 37641
rect 542358 37567 542414 37576
rect 542372 26761 542400 37567
rect 542358 26752 542414 26761
rect 542358 26687 542414 26696
rect 542176 17400 542228 17406
rect 542176 17342 542228 17348
rect 542084 15088 542136 15094
rect 542084 15030 542136 15036
rect 542464 13258 542492 75822
rect 542556 36786 542584 133826
rect 542648 107681 542676 156470
rect 542728 154284 542780 154290
rect 542728 154226 542780 154232
rect 542634 107672 542690 107681
rect 542634 107607 542690 107616
rect 542636 89752 542688 89758
rect 542636 89694 542688 89700
rect 542648 69902 542676 89694
rect 542740 75041 542768 154226
rect 542832 147098 542860 215902
rect 542912 159180 542964 159186
rect 542912 159122 542964 159128
rect 542924 147354 542952 159122
rect 543016 147370 543044 227122
rect 543108 147801 543136 229978
rect 543844 227254 543872 233922
rect 543832 227248 543884 227254
rect 543832 227190 543884 227196
rect 543936 151814 543964 238070
rect 544014 238031 544070 238040
rect 543844 151786 543964 151814
rect 543188 151700 543240 151706
rect 543188 151642 543240 151648
rect 543094 147792 543150 147801
rect 543094 147727 543150 147736
rect 542912 147348 542964 147354
rect 543016 147342 543136 147370
rect 542912 147290 542964 147296
rect 542832 147070 543044 147098
rect 542820 147008 542872 147014
rect 542820 146950 542872 146956
rect 542912 147008 542964 147014
rect 542912 146950 542964 146956
rect 542832 143546 542860 146950
rect 542820 143540 542872 143546
rect 542820 143482 542872 143488
rect 542820 143404 542872 143410
rect 542820 143346 542872 143352
rect 542832 137358 542860 143346
rect 542820 137352 542872 137358
rect 542820 137294 542872 137300
rect 542818 129976 542874 129985
rect 542818 129911 542874 129920
rect 542832 115938 542860 129911
rect 542820 115932 542872 115938
rect 542820 115874 542872 115880
rect 542820 108384 542872 108390
rect 542820 108326 542872 108332
rect 542832 102202 542860 108326
rect 542820 102196 542872 102202
rect 542820 102138 542872 102144
rect 542726 75032 542782 75041
rect 542726 74967 542782 74976
rect 542820 71052 542872 71058
rect 542820 70994 542872 71000
rect 542636 69896 542688 69902
rect 542636 69838 542688 69844
rect 542636 69012 542688 69018
rect 542636 68954 542688 68960
rect 542544 36780 542596 36786
rect 542544 36722 542596 36728
rect 542452 13252 542504 13258
rect 542452 13194 542504 13200
rect 542648 12374 542676 68954
rect 542832 65521 542860 70994
rect 542818 65512 542874 65521
rect 542818 65447 542874 65456
rect 542924 17202 542952 146950
rect 543016 145761 543044 147070
rect 543108 146198 543136 147342
rect 543096 146192 543148 146198
rect 543096 146134 543148 146140
rect 543002 145752 543058 145761
rect 543002 145687 543058 145696
rect 543200 144770 543228 151642
rect 543648 149116 543700 149122
rect 543648 149058 543700 149064
rect 543556 147620 543608 147626
rect 543556 147562 543608 147568
rect 543568 146441 543596 147562
rect 543554 146432 543610 146441
rect 543554 146367 543610 146376
rect 543556 146328 543608 146334
rect 543556 146270 543608 146276
rect 543464 146124 543516 146130
rect 543464 146066 543516 146072
rect 543280 144900 543332 144906
rect 543280 144842 543332 144848
rect 543188 144764 543240 144770
rect 543188 144706 543240 144712
rect 543004 143608 543056 143614
rect 543004 143550 543056 143556
rect 543016 113558 543044 143550
rect 543188 143540 543240 143546
rect 543188 143482 543240 143488
rect 543096 143200 543148 143206
rect 543096 143142 543148 143148
rect 543108 143041 543136 143142
rect 543094 143032 543150 143041
rect 543094 142967 543150 142976
rect 543200 142361 543228 143482
rect 543186 142352 543242 142361
rect 543186 142287 543242 142296
rect 543292 142154 543320 144842
rect 543108 142126 543320 142154
rect 543108 127673 543136 142126
rect 543188 141704 543240 141710
rect 543186 141672 543188 141681
rect 543240 141672 543242 141681
rect 543186 141607 543242 141616
rect 543280 141160 543332 141166
rect 543280 141102 543332 141108
rect 543292 133890 543320 141102
rect 543280 133884 543332 133890
rect 543280 133826 543332 133832
rect 543094 127664 543150 127673
rect 543094 127599 543150 127608
rect 543188 126948 543240 126954
rect 543188 126890 543240 126896
rect 543200 121310 543228 126890
rect 543476 126886 543504 146066
rect 543568 140826 543596 146270
rect 543660 144906 543688 149058
rect 543740 147688 543792 147694
rect 543740 147630 543792 147636
rect 543648 144900 543700 144906
rect 543648 144842 543700 144848
rect 543752 143614 543780 147630
rect 543740 143608 543792 143614
rect 543740 143550 543792 143556
rect 543648 142112 543700 142118
rect 543648 142054 543700 142060
rect 543660 141001 543688 142054
rect 543646 140992 543702 141001
rect 543646 140927 543702 140936
rect 543844 140894 543872 151786
rect 543924 147552 543976 147558
rect 543924 147494 543976 147500
rect 543936 144809 543964 147494
rect 543922 144800 543978 144809
rect 543922 144735 543978 144744
rect 544028 143954 544056 238031
rect 544212 237794 544240 240094
rect 544304 240094 544640 240122
rect 545592 240094 545928 240122
rect 544200 237788 544252 237794
rect 544200 237730 544252 237736
rect 544304 233986 544332 240094
rect 544474 239320 544530 239329
rect 544474 239255 544530 239264
rect 544384 234184 544436 234190
rect 544384 234126 544436 234132
rect 544292 233980 544344 233986
rect 544292 233922 544344 233928
rect 544108 227044 544160 227050
rect 544108 226986 544160 226992
rect 544120 146266 544148 226986
rect 544200 207052 544252 207058
rect 544200 206994 544252 207000
rect 544108 146260 544160 146266
rect 544108 146202 544160 146208
rect 544016 143948 544068 143954
rect 544016 143890 544068 143896
rect 543924 143472 543976 143478
rect 543924 143414 543976 143420
rect 543832 140888 543884 140894
rect 543832 140830 543884 140836
rect 543556 140820 543608 140826
rect 543556 140762 543608 140768
rect 543556 139392 543608 139398
rect 543556 139334 543608 139340
rect 543568 138281 543596 139334
rect 543554 138272 543610 138281
rect 543554 138207 543610 138216
rect 543830 137320 543886 137329
rect 543830 137255 543886 137264
rect 543556 136604 543608 136610
rect 543556 136546 543608 136552
rect 543568 136241 543596 136546
rect 543648 136536 543700 136542
rect 543648 136478 543700 136484
rect 543554 136232 543610 136241
rect 543554 136167 543610 136176
rect 543660 135561 543688 136478
rect 543646 135552 543702 135561
rect 543646 135487 543702 135496
rect 543648 135448 543700 135454
rect 543648 135390 543700 135396
rect 543556 135244 543608 135250
rect 543556 135186 543608 135192
rect 543568 134201 543596 135186
rect 543554 134192 543610 134201
rect 543554 134127 543610 134136
rect 543556 132456 543608 132462
rect 543556 132398 543608 132404
rect 543568 131481 543596 132398
rect 543660 131510 543688 135390
rect 543648 131504 543700 131510
rect 543554 131472 543610 131481
rect 543648 131446 543700 131452
rect 543554 131407 543610 131416
rect 543740 131164 543792 131170
rect 543740 131106 543792 131112
rect 543556 131096 543608 131102
rect 543556 131038 543608 131044
rect 543568 130801 543596 131038
rect 543554 130792 543610 130801
rect 543554 130727 543610 130736
rect 543752 128330 543780 131106
rect 543556 128308 543608 128314
rect 543556 128250 543608 128256
rect 543660 128302 543780 128330
rect 543568 128081 543596 128250
rect 543554 128072 543610 128081
rect 543554 128007 543610 128016
rect 543464 126880 543516 126886
rect 543464 126822 543516 126828
rect 543556 125588 543608 125594
rect 543556 125530 543608 125536
rect 543568 125361 543596 125530
rect 543660 125474 543688 128302
rect 543844 125746 543872 137255
rect 543752 125718 543872 125746
rect 543752 125662 543780 125718
rect 543740 125656 543792 125662
rect 543740 125598 543792 125604
rect 543830 125624 543886 125633
rect 543830 125559 543886 125568
rect 543660 125446 543780 125474
rect 543554 125352 543610 125361
rect 543554 125287 543610 125296
rect 543372 123412 543424 123418
rect 543372 123354 543424 123360
rect 543188 121304 543240 121310
rect 543188 121246 543240 121252
rect 543096 120148 543148 120154
rect 543096 120090 543148 120096
rect 543004 113552 543056 113558
rect 543004 113494 543056 113500
rect 543108 110634 543136 120090
rect 543384 117994 543412 123354
rect 543556 122800 543608 122806
rect 543556 122742 543608 122748
rect 543568 121961 543596 122742
rect 543554 121952 543610 121961
rect 543554 121887 543610 121896
rect 543556 121440 543608 121446
rect 543556 121382 543608 121388
rect 543568 120601 543596 121382
rect 543554 120592 543610 120601
rect 543554 120527 543610 120536
rect 543200 117966 543412 117994
rect 543096 110628 543148 110634
rect 543096 110570 543148 110576
rect 543004 110492 543056 110498
rect 543004 110434 543056 110440
rect 542912 17196 542964 17202
rect 542912 17138 542964 17144
rect 543016 16250 543044 110434
rect 543200 109750 543228 117966
rect 543556 117292 543608 117298
rect 543556 117234 543608 117240
rect 543568 116521 543596 117234
rect 543554 116512 543610 116521
rect 543554 116447 543610 116456
rect 543556 115864 543608 115870
rect 543554 115832 543556 115841
rect 543608 115832 543610 115841
rect 543554 115767 543610 115776
rect 543556 114504 543608 114510
rect 543554 114472 543556 114481
rect 543608 114472 543610 114481
rect 543554 114407 543610 114416
rect 543648 114436 543700 114442
rect 543648 114378 543700 114384
rect 543660 113801 543688 114378
rect 543646 113792 543702 113801
rect 543646 113727 543702 113736
rect 543752 113642 543780 125446
rect 543384 113614 543780 113642
rect 543384 110566 543412 113614
rect 543844 113540 543872 125559
rect 543660 113512 543872 113540
rect 543372 110560 543424 110566
rect 543372 110502 543424 110508
rect 543556 110424 543608 110430
rect 543554 110392 543556 110401
rect 543608 110392 543610 110401
rect 543554 110327 543610 110336
rect 543188 109744 543240 109750
rect 543188 109686 543240 109692
rect 543096 108996 543148 109002
rect 543096 108938 543148 108944
rect 543108 101862 543136 108938
rect 543660 108866 543688 113512
rect 543832 110628 543884 110634
rect 543832 110570 543884 110576
rect 543648 108860 543700 108866
rect 543648 108802 543700 108808
rect 543740 108452 543792 108458
rect 543740 108394 543792 108400
rect 543188 107908 543240 107914
rect 543188 107850 543240 107856
rect 543096 101856 543148 101862
rect 543096 101798 543148 101804
rect 543096 97300 543148 97306
rect 543096 97242 543148 97248
rect 543004 16244 543056 16250
rect 543004 16186 543056 16192
rect 542636 12368 542688 12374
rect 542636 12310 542688 12316
rect 541992 12300 542044 12306
rect 541992 12242 542044 12248
rect 541624 6724 541676 6730
rect 541624 6666 541676 6672
rect 543108 6526 543136 97242
rect 543200 20126 543228 107850
rect 543280 107636 543332 107642
rect 543280 107578 543332 107584
rect 543292 106321 543320 107578
rect 543278 106312 543334 106321
rect 543278 106247 543334 106256
rect 543752 106026 543780 108394
rect 543844 107710 543872 110570
rect 543832 107704 543884 107710
rect 543832 107646 543884 107652
rect 543660 105998 543780 106026
rect 543464 104236 543516 104242
rect 543464 104178 543516 104184
rect 543372 95192 543424 95198
rect 543372 95134 543424 95140
rect 543280 94104 543332 94110
rect 543280 94046 543332 94052
rect 543188 20120 543240 20126
rect 543188 20062 543240 20068
rect 543292 17474 543320 94046
rect 543384 88482 543412 95134
rect 543476 90574 543504 104178
rect 543660 102354 543688 105998
rect 543832 104848 543884 104854
rect 543832 104790 543884 104796
rect 543568 102326 543688 102354
rect 543568 98666 543596 102326
rect 543648 102264 543700 102270
rect 543648 102206 543700 102212
rect 543556 98660 543608 98666
rect 543556 98602 543608 98608
rect 543556 97980 543608 97986
rect 543556 97922 543608 97928
rect 543568 97481 543596 97922
rect 543554 97472 543610 97481
rect 543554 97407 543610 97416
rect 543556 96620 543608 96626
rect 543556 96562 543608 96568
rect 543568 96121 543596 96562
rect 543554 96112 543610 96121
rect 543554 96047 543610 96056
rect 543556 95192 543608 95198
rect 543556 95134 543608 95140
rect 543568 94081 543596 95134
rect 543554 94072 543610 94081
rect 543554 94007 543610 94016
rect 543556 93968 543608 93974
rect 543556 93910 543608 93916
rect 543568 92154 543596 93910
rect 543660 93854 543688 102206
rect 543660 93826 543780 93854
rect 543568 92126 543688 92154
rect 543554 92032 543610 92041
rect 543554 91967 543610 91976
rect 543568 91254 543596 91967
rect 543556 91248 543608 91254
rect 543556 91190 543608 91196
rect 543464 90568 543516 90574
rect 543464 90510 543516 90516
rect 543556 89684 543608 89690
rect 543556 89626 543608 89632
rect 543568 88641 543596 89626
rect 543554 88632 543610 88641
rect 543554 88567 543610 88576
rect 543384 88454 543596 88482
rect 543464 87644 543516 87650
rect 543464 87586 543516 87592
rect 543476 85898 543504 87586
rect 543568 86850 543596 88454
rect 543660 88210 543688 92126
rect 543752 89826 543780 93826
rect 543740 89820 543792 89826
rect 543740 89762 543792 89768
rect 543844 88330 543872 104790
rect 543832 88324 543884 88330
rect 543832 88266 543884 88272
rect 543660 88182 543872 88210
rect 543568 86822 543780 86850
rect 543384 85870 543504 85898
rect 543280 17468 543332 17474
rect 543280 17410 543332 17416
rect 543384 17338 543412 85870
rect 543464 85808 543516 85814
rect 543464 85750 543516 85756
rect 543476 72570 543504 85750
rect 543556 84176 543608 84182
rect 543556 84118 543608 84124
rect 543568 83881 543596 84118
rect 543752 83978 543780 86822
rect 543844 85814 543872 88182
rect 543832 85808 543884 85814
rect 543832 85750 543884 85756
rect 543740 83972 543792 83978
rect 543740 83914 543792 83920
rect 543554 83872 543610 83881
rect 543554 83807 543610 83816
rect 543556 82816 543608 82822
rect 543556 82758 543608 82764
rect 543568 82521 543596 82758
rect 543554 82512 543610 82521
rect 543554 82447 543610 82456
rect 543648 78668 543700 78674
rect 543648 78610 543700 78616
rect 543556 78600 543608 78606
rect 543556 78542 543608 78548
rect 543568 78441 543596 78542
rect 543554 78432 543610 78441
rect 543554 78367 543610 78376
rect 543660 77761 543688 78610
rect 543646 77752 543702 77761
rect 543646 77687 543702 77696
rect 543556 77240 543608 77246
rect 543556 77182 543608 77188
rect 543568 76401 543596 77182
rect 543554 76392 543610 76401
rect 543554 76327 543610 76336
rect 543554 75712 543610 75721
rect 543554 75647 543610 75656
rect 543568 75274 543596 75647
rect 543556 75268 543608 75274
rect 543556 75210 543608 75216
rect 543476 72542 543780 72570
rect 543556 72480 543608 72486
rect 543556 72422 543608 72428
rect 543568 71641 543596 72422
rect 543554 71632 543610 71641
rect 543554 71567 543610 71576
rect 543556 70372 543608 70378
rect 543556 70314 543608 70320
rect 543568 70281 543596 70314
rect 543554 70272 543610 70281
rect 543554 70207 543610 70216
rect 543752 69698 543780 72542
rect 543740 69692 543792 69698
rect 543740 69634 543792 69640
rect 543556 66224 543608 66230
rect 543554 66192 543556 66201
rect 543608 66192 543610 66201
rect 543554 66127 543610 66136
rect 543554 64152 543610 64161
rect 543554 64087 543610 64096
rect 543568 64054 543596 64087
rect 543556 64048 543608 64054
rect 543556 63990 543608 63996
rect 543554 62112 543610 62121
rect 543554 62047 543556 62056
rect 543608 62047 543610 62056
rect 543556 62018 543608 62024
rect 543648 62008 543700 62014
rect 543648 61950 543700 61956
rect 543660 60761 543688 61950
rect 543646 60752 543702 60761
rect 543646 60687 543702 60696
rect 543556 57928 543608 57934
rect 543556 57870 543608 57876
rect 543568 56681 543596 57870
rect 543554 56672 543610 56681
rect 543554 56607 543610 56616
rect 543556 53780 543608 53786
rect 543556 53722 543608 53728
rect 543568 52601 543596 53722
rect 543554 52592 543610 52601
rect 543554 52527 543610 52536
rect 543464 50856 543516 50862
rect 543464 50798 543516 50804
rect 543476 49881 543504 50798
rect 543462 49872 543518 49881
rect 543462 49807 543518 49816
rect 543556 49700 543608 49706
rect 543556 49642 543608 49648
rect 543568 48521 543596 49642
rect 543554 48512 543610 48521
rect 543554 48447 543610 48456
rect 543556 48272 543608 48278
rect 543556 48214 543608 48220
rect 543568 47841 543596 48214
rect 543554 47832 543610 47841
rect 543554 47767 543610 47776
rect 543556 45552 543608 45558
rect 543556 45494 543608 45500
rect 543568 45121 543596 45494
rect 543648 45484 543700 45490
rect 543648 45426 543700 45432
rect 543554 45112 543610 45121
rect 543554 45047 543610 45056
rect 543660 44441 543688 45426
rect 543646 44432 543702 44441
rect 543646 44367 543702 44376
rect 543556 44124 543608 44130
rect 543556 44066 543608 44072
rect 543568 43761 543596 44066
rect 543554 43752 543610 43761
rect 543554 43687 543610 43696
rect 543556 41404 543608 41410
rect 543556 41346 543608 41352
rect 543568 41041 543596 41346
rect 543554 41032 543610 41041
rect 543554 40967 543610 40976
rect 543556 37256 543608 37262
rect 543556 37198 543608 37204
rect 543568 36281 543596 37198
rect 543554 36272 543610 36281
rect 543554 36207 543610 36216
rect 543556 35896 543608 35902
rect 543556 35838 543608 35844
rect 543568 35601 543596 35838
rect 543554 35592 543610 35601
rect 543554 35527 543610 35536
rect 543556 31748 543608 31754
rect 543556 31690 543608 31696
rect 543568 30841 543596 31690
rect 543554 30832 543610 30841
rect 543554 30767 543610 30776
rect 543936 21894 543964 143414
rect 544212 142186 544240 206994
rect 544396 149734 544424 234126
rect 544488 167686 544516 239255
rect 545592 238746 545620 240094
rect 547846 239850 547874 240108
rect 548168 240094 548504 240122
rect 547846 239822 547920 239850
rect 547788 239488 547840 239494
rect 547788 239430 547840 239436
rect 547236 239420 547288 239426
rect 547236 239362 547288 239368
rect 547420 239420 547472 239426
rect 547420 239362 547472 239368
rect 545580 238740 545632 238746
rect 545580 238682 545632 238688
rect 546222 238504 546278 238513
rect 546222 238439 546278 238448
rect 545486 237280 545542 237289
rect 545486 237215 545542 237224
rect 545500 236881 545528 237215
rect 545762 237144 545818 237153
rect 545762 237079 545818 237088
rect 545486 236872 545542 236881
rect 545486 236807 545542 236816
rect 545212 234320 545264 234326
rect 545212 234262 545264 234268
rect 544844 234252 544896 234258
rect 544844 234194 544896 234200
rect 544660 230240 544712 230246
rect 544660 230182 544712 230188
rect 544476 167680 544528 167686
rect 544476 167622 544528 167628
rect 544384 149728 544436 149734
rect 544384 149670 544436 149676
rect 544474 148880 544530 148889
rect 544474 148815 544530 148824
rect 544384 144832 544436 144838
rect 544384 144774 544436 144780
rect 544292 144764 544344 144770
rect 544292 144706 544344 144712
rect 544200 142180 544252 142186
rect 544200 142122 544252 142128
rect 544106 130112 544162 130121
rect 544106 130047 544162 130056
rect 544016 128240 544068 128246
rect 544016 128182 544068 128188
rect 544028 110498 544056 128182
rect 544120 122874 544148 130047
rect 544108 122868 544160 122874
rect 544108 122810 544160 122816
rect 544016 110492 544068 110498
rect 544016 110434 544068 110440
rect 544200 108860 544252 108866
rect 544200 108802 544252 108808
rect 544016 104780 544068 104786
rect 544016 104722 544068 104728
rect 544028 24818 544056 104722
rect 544108 90568 544160 90574
rect 544108 90510 544160 90516
rect 544120 73234 544148 90510
rect 544212 89758 544240 108802
rect 544200 89752 544252 89758
rect 544200 89694 544252 89700
rect 544108 73228 544160 73234
rect 544108 73170 544160 73176
rect 544108 69896 544160 69902
rect 544108 69838 544160 69844
rect 544016 24812 544068 24818
rect 544016 24754 544068 24760
rect 543924 21888 543976 21894
rect 543924 21830 543976 21836
rect 544120 18562 544148 69838
rect 544200 42356 544252 42362
rect 544200 42298 544252 42304
rect 544108 18556 544160 18562
rect 544108 18498 544160 18504
rect 543372 17332 543424 17338
rect 543372 17274 543424 17280
rect 544212 12442 544240 42298
rect 544304 20466 544332 144706
rect 544396 124166 544424 144774
rect 544488 144158 544516 148815
rect 544672 146674 544700 230182
rect 544660 146668 544712 146674
rect 544660 146610 544712 146616
rect 544752 144900 544804 144906
rect 544752 144842 544804 144848
rect 544476 144152 544528 144158
rect 544476 144094 544528 144100
rect 544764 137562 544792 144842
rect 544752 137556 544804 137562
rect 544752 137498 544804 137504
rect 544752 137420 544804 137426
rect 544752 137362 544804 137368
rect 544660 137352 544712 137358
rect 544660 137294 544712 137300
rect 544672 130830 544700 137294
rect 544764 130966 544792 137362
rect 544752 130960 544804 130966
rect 544752 130902 544804 130908
rect 544660 130824 544712 130830
rect 544660 130766 544712 130772
rect 544476 130076 544528 130082
rect 544476 130018 544528 130024
rect 544384 124160 544436 124166
rect 544384 124102 544436 124108
rect 544384 115048 544436 115054
rect 544384 114990 544436 114996
rect 544292 20460 544344 20466
rect 544292 20402 544344 20408
rect 544396 13530 544424 114990
rect 544488 108254 544516 130018
rect 544568 125724 544620 125730
rect 544568 125666 544620 125672
rect 544476 108248 544528 108254
rect 544476 108190 544528 108196
rect 544476 100768 544528 100774
rect 544476 100710 544528 100716
rect 544488 30326 544516 100710
rect 544580 94110 544608 125666
rect 544658 117328 544714 117337
rect 544658 117263 544714 117272
rect 544672 110537 544700 117263
rect 544658 110528 544714 110537
rect 544658 110463 544714 110472
rect 544568 94104 544620 94110
rect 544568 94046 544620 94052
rect 544568 83020 544620 83026
rect 544568 82962 544620 82968
rect 544476 30320 544528 30326
rect 544476 30262 544528 30268
rect 544580 14686 544608 82962
rect 544658 82920 544714 82929
rect 544658 82855 544714 82864
rect 544672 19922 544700 82855
rect 544660 19916 544712 19922
rect 544660 19858 544712 19864
rect 544568 14680 544620 14686
rect 544568 14622 544620 14628
rect 544856 13734 544884 234194
rect 545028 208412 545080 208418
rect 545028 208354 545080 208360
rect 544936 154012 544988 154018
rect 544936 153954 544988 153960
rect 544948 84658 544976 153954
rect 545040 143206 545068 208354
rect 545120 152652 545172 152658
rect 545120 152594 545172 152600
rect 545028 143200 545080 143206
rect 545028 143142 545080 143148
rect 545132 142154 545160 152594
rect 545224 149122 545252 234262
rect 545672 159928 545724 159934
rect 545672 159870 545724 159876
rect 545304 151156 545356 151162
rect 545304 151098 545356 151104
rect 545212 149116 545264 149122
rect 545212 149058 545264 149064
rect 545212 146192 545264 146198
rect 545212 146134 545264 146140
rect 545040 142126 545160 142154
rect 545040 135318 545068 142126
rect 545120 140072 545172 140078
rect 545120 140014 545172 140020
rect 545028 135312 545080 135318
rect 545028 135254 545080 135260
rect 545026 135144 545082 135153
rect 545026 135079 545082 135088
rect 545040 131073 545068 135079
rect 545132 133958 545160 140014
rect 545224 138038 545252 146134
rect 545212 138032 545264 138038
rect 545212 137974 545264 137980
rect 545120 133952 545172 133958
rect 545120 133894 545172 133900
rect 545026 131064 545082 131073
rect 545026 130999 545082 131008
rect 545028 130960 545080 130966
rect 545028 130902 545080 130908
rect 545040 127634 545068 130902
rect 545028 127628 545080 127634
rect 545028 127570 545080 127576
rect 545120 121508 545172 121514
rect 545120 121450 545172 121456
rect 545132 120170 545160 121450
rect 545040 120142 545160 120170
rect 545040 117230 545068 120142
rect 545028 117224 545080 117230
rect 545028 117166 545080 117172
rect 545120 114640 545172 114646
rect 545120 114582 545172 114588
rect 545132 113218 545160 114582
rect 545120 113212 545172 113218
rect 545120 113154 545172 113160
rect 545028 108384 545080 108390
rect 545028 108326 545080 108332
rect 545040 104242 545068 108326
rect 545028 104236 545080 104242
rect 545028 104178 545080 104184
rect 545028 102332 545080 102338
rect 545028 102274 545080 102280
rect 545040 102082 545068 102274
rect 545040 102054 545160 102082
rect 545132 93974 545160 102054
rect 545120 93968 545172 93974
rect 545120 93910 545172 93916
rect 545028 88324 545080 88330
rect 545028 88266 545080 88272
rect 544936 84652 544988 84658
rect 544936 84594 544988 84600
rect 545040 83910 545068 88266
rect 545028 83904 545080 83910
rect 545028 83846 545080 83852
rect 545120 72276 545172 72282
rect 545120 72218 545172 72224
rect 545132 66706 545160 72218
rect 545120 66700 545172 66706
rect 545120 66642 545172 66648
rect 545316 27402 545344 151098
rect 545488 143336 545540 143342
rect 545488 143278 545540 143284
rect 545396 139528 545448 139534
rect 545396 139470 545448 139476
rect 545408 130082 545436 139470
rect 545396 130076 545448 130082
rect 545396 130018 545448 130024
rect 545396 124160 545448 124166
rect 545396 124102 545448 124108
rect 545304 27396 545356 27402
rect 545304 27338 545356 27344
rect 544844 13728 544896 13734
rect 544844 13670 544896 13676
rect 544384 13524 544436 13530
rect 544384 13466 544436 13472
rect 544200 12436 544252 12442
rect 544200 12378 544252 12384
rect 545408 12102 545436 124102
rect 545500 115054 545528 143278
rect 545580 133884 545632 133890
rect 545580 133826 545632 133832
rect 545488 115048 545540 115054
rect 545488 114990 545540 114996
rect 545488 114368 545540 114374
rect 545488 114310 545540 114316
rect 545396 12096 545448 12102
rect 545396 12038 545448 12044
rect 545500 11966 545528 114310
rect 545592 100774 545620 133826
rect 545580 100768 545632 100774
rect 545580 100710 545632 100716
rect 545684 22710 545712 159870
rect 545776 145586 545804 237079
rect 545856 230376 545908 230382
rect 545856 230318 545908 230324
rect 545764 145580 545816 145586
rect 545764 145522 545816 145528
rect 545868 145518 545896 230318
rect 546038 230208 546094 230217
rect 546038 230143 546094 230152
rect 545948 229696 546000 229702
rect 545948 229638 546000 229644
rect 545960 146266 545988 229638
rect 546052 149054 546080 230143
rect 546132 149796 546184 149802
rect 546132 149738 546184 149744
rect 546040 149048 546092 149054
rect 546040 148990 546092 148996
rect 545948 146260 546000 146266
rect 545948 146202 546000 146208
rect 546040 145648 546092 145654
rect 546040 145590 546092 145596
rect 545856 145512 545908 145518
rect 545856 145454 545908 145460
rect 545948 137556 546000 137562
rect 545948 137498 546000 137504
rect 545960 133142 545988 137498
rect 546052 135182 546080 145590
rect 546040 135176 546092 135182
rect 546040 135118 546092 135124
rect 545948 133136 546000 133142
rect 545948 133078 546000 133084
rect 545856 132796 545908 132802
rect 545856 132738 545908 132744
rect 545764 115932 545816 115938
rect 545764 115874 545816 115880
rect 545672 22704 545724 22710
rect 545672 22646 545724 22652
rect 545488 11960 545540 11966
rect 545488 11902 545540 11908
rect 543096 6520 543148 6526
rect 543096 6462 543148 6468
rect 545776 3806 545804 115874
rect 545868 29714 545896 132738
rect 546144 132394 546172 149738
rect 546132 132388 546184 132394
rect 546132 132330 546184 132336
rect 545948 131028 546000 131034
rect 545948 130970 546000 130976
rect 545960 120578 545988 130970
rect 546236 124137 546264 238439
rect 547144 237448 547196 237454
rect 547144 237390 547196 237396
rect 546958 234016 547014 234025
rect 546958 233951 547014 233960
rect 546776 159792 546828 159798
rect 546776 159734 546828 159740
rect 546316 154488 546368 154494
rect 546316 154430 546368 154436
rect 546222 124128 546278 124137
rect 546222 124063 546278 124072
rect 545960 120550 546264 120578
rect 546040 120420 546092 120426
rect 546040 120362 546092 120368
rect 545948 108112 546000 108118
rect 545948 108054 546000 108060
rect 545960 88330 545988 108054
rect 546052 106282 546080 120362
rect 546132 117360 546184 117366
rect 546132 117302 546184 117308
rect 546144 114034 546172 117302
rect 546132 114028 546184 114034
rect 546132 113970 546184 113976
rect 546236 108322 546264 120550
rect 546224 108316 546276 108322
rect 546224 108258 546276 108264
rect 546040 106276 546092 106282
rect 546040 106218 546092 106224
rect 546132 89616 546184 89622
rect 546132 89558 546184 89564
rect 545948 88324 546000 88330
rect 545948 88266 546000 88272
rect 546144 82958 546172 89558
rect 546132 82952 546184 82958
rect 546132 82894 546184 82900
rect 546040 82884 546092 82890
rect 546040 82826 546092 82832
rect 545948 74588 546000 74594
rect 545948 74530 546000 74536
rect 545856 29708 545908 29714
rect 545856 29650 545908 29656
rect 545960 13462 545988 74530
rect 546052 73234 546080 82826
rect 546040 73228 546092 73234
rect 546040 73170 546092 73176
rect 546040 67652 546092 67658
rect 546040 67594 546092 67600
rect 545948 13456 546000 13462
rect 545948 13398 546000 13404
rect 546052 10742 546080 67594
rect 546328 29238 546356 154430
rect 546592 154352 546644 154358
rect 546592 154294 546644 154300
rect 546500 150136 546552 150142
rect 546500 150078 546552 150084
rect 546408 146124 546460 146130
rect 546408 146066 546460 146072
rect 546420 133210 546448 146066
rect 546512 135454 546540 150078
rect 546604 141710 546632 154294
rect 546682 152416 546738 152425
rect 546682 152351 546738 152360
rect 546592 141704 546644 141710
rect 546592 141646 546644 141652
rect 546590 141264 546646 141273
rect 546590 141199 546646 141208
rect 546500 135448 546552 135454
rect 546500 135390 546552 135396
rect 546408 133204 546460 133210
rect 546408 133146 546460 133152
rect 546408 133068 546460 133074
rect 546408 133010 546460 133016
rect 546420 123026 546448 133010
rect 546604 131034 546632 141199
rect 546592 131028 546644 131034
rect 546592 130970 546644 130976
rect 546590 125488 546646 125497
rect 546590 125423 546646 125432
rect 546420 122998 546540 123026
rect 546408 122868 546460 122874
rect 546408 122810 546460 122816
rect 546420 117314 546448 122810
rect 546512 122738 546540 122998
rect 546500 122732 546552 122738
rect 546500 122674 546552 122680
rect 546604 117366 546632 125423
rect 546592 117360 546644 117366
rect 546420 117286 546540 117314
rect 546592 117302 546644 117308
rect 546408 111852 546460 111858
rect 546408 111794 546460 111800
rect 546420 89554 546448 111794
rect 546512 106185 546540 117286
rect 546592 117224 546644 117230
rect 546592 117166 546644 117172
rect 546604 108118 546632 117166
rect 546592 108112 546644 108118
rect 546592 108054 546644 108060
rect 546498 106176 546554 106185
rect 546498 106111 546554 106120
rect 546408 89548 546460 89554
rect 546408 89490 546460 89496
rect 546500 83904 546552 83910
rect 546500 83846 546552 83852
rect 546512 70650 546540 83846
rect 546500 70644 546552 70650
rect 546500 70586 546552 70592
rect 546500 70508 546552 70514
rect 546500 70450 546552 70456
rect 546512 67658 546540 70450
rect 546500 67652 546552 67658
rect 546500 67594 546552 67600
rect 546316 29232 546368 29238
rect 546316 29174 546368 29180
rect 546040 10736 546092 10742
rect 546040 10678 546092 10684
rect 545764 3800 545816 3806
rect 545764 3742 545816 3748
rect 541544 3454 542032 3482
rect 542004 480 542032 3454
rect 545488 3256 545540 3262
rect 545488 3198 545540 3204
rect 545500 480 545528 3198
rect 546696 3194 546724 152351
rect 546788 29442 546816 159734
rect 546868 154148 546920 154154
rect 546868 154090 546920 154096
rect 546776 29436 546828 29442
rect 546776 29378 546828 29384
rect 546880 28422 546908 154090
rect 546972 131238 547000 233951
rect 547052 151292 547104 151298
rect 547052 151234 547104 151240
rect 546960 131232 547012 131238
rect 546960 131174 547012 131180
rect 546960 130892 547012 130898
rect 546960 130834 547012 130840
rect 546972 117570 547000 130834
rect 546960 117564 547012 117570
rect 546960 117506 547012 117512
rect 546960 69692 547012 69698
rect 546960 69634 547012 69640
rect 546868 28416 546920 28422
rect 546868 28358 546920 28364
rect 546972 10946 547000 69634
rect 547064 50862 547092 151234
rect 547052 50856 547104 50862
rect 547052 50798 547104 50804
rect 546960 10940 547012 10946
rect 546960 10882 547012 10888
rect 547156 4826 547184 237390
rect 547248 151162 547276 239362
rect 547328 230512 547380 230518
rect 547328 230454 547380 230460
rect 547340 152590 547368 230454
rect 547432 167958 547460 239362
rect 547800 238746 547828 239430
rect 547788 238740 547840 238746
rect 547788 238682 547840 238688
rect 547604 237992 547656 237998
rect 547604 237934 547656 237940
rect 547512 236768 547564 236774
rect 547512 236710 547564 236716
rect 547524 186969 547552 236710
rect 547510 186960 547566 186969
rect 547510 186895 547566 186904
rect 547420 167952 547472 167958
rect 547420 167894 547472 167900
rect 547328 152584 547380 152590
rect 547328 152526 547380 152532
rect 547236 151156 547288 151162
rect 547236 151098 547288 151104
rect 547236 130824 547288 130830
rect 547236 130766 547288 130772
rect 547248 115938 547276 130766
rect 547510 128480 547566 128489
rect 547510 128415 547566 128424
rect 547524 126177 547552 128415
rect 547510 126168 547566 126177
rect 547510 126103 547566 126112
rect 547236 115932 547288 115938
rect 547236 115874 547288 115880
rect 547328 114572 547380 114578
rect 547328 114514 547380 114520
rect 547236 104168 547288 104174
rect 547236 104110 547288 104116
rect 547248 20670 547276 104110
rect 547340 97306 547368 114514
rect 547420 106276 547472 106282
rect 547420 106218 547472 106224
rect 547328 97300 547380 97306
rect 547328 97242 547380 97248
rect 547432 95334 547460 106218
rect 547420 95328 547472 95334
rect 547420 95270 547472 95276
rect 547328 95260 547380 95266
rect 547328 95202 547380 95208
rect 547340 86873 547368 95202
rect 547420 89480 547472 89486
rect 547420 89422 547472 89428
rect 547326 86864 547382 86873
rect 547326 86799 547382 86808
rect 547328 85536 547380 85542
rect 547328 85478 547380 85484
rect 547340 71738 547368 85478
rect 547432 82890 547460 89422
rect 547420 82884 547472 82890
rect 547420 82826 547472 82832
rect 547328 71732 547380 71738
rect 547328 71674 547380 71680
rect 547616 22778 547644 237934
rect 547696 237652 547748 237658
rect 547696 237594 547748 237600
rect 547708 25566 547736 237594
rect 547892 237454 547920 239822
rect 548168 238649 548196 240094
rect 549134 239850 549162 240108
rect 549134 239822 549208 239850
rect 549076 239556 549128 239562
rect 549076 239498 549128 239504
rect 548154 238640 548210 238649
rect 548154 238575 548210 238584
rect 547880 237448 547932 237454
rect 547880 237390 547932 237396
rect 548982 237280 549038 237289
rect 548982 237215 549038 237224
rect 548524 233096 548576 233102
rect 548524 233038 548576 233044
rect 548064 230308 548116 230314
rect 548064 230250 548116 230256
rect 547970 229936 548026 229945
rect 547970 229871 548026 229880
rect 547878 154048 547934 154057
rect 547878 153983 547934 153992
rect 547892 151298 547920 153983
rect 547880 151292 547932 151298
rect 547880 151234 547932 151240
rect 547880 149048 547932 149054
rect 547880 148990 547932 148996
rect 547892 131186 547920 148990
rect 547984 147121 548012 229871
rect 547970 147112 548026 147121
rect 547970 147047 548026 147056
rect 548076 146962 548104 230250
rect 548248 229968 548300 229974
rect 548248 229910 548300 229916
rect 548156 151360 548208 151366
rect 548156 151302 548208 151308
rect 547984 146934 548104 146962
rect 547984 146130 548012 146934
rect 548062 146840 548118 146849
rect 548062 146775 548118 146784
rect 547972 146124 548024 146130
rect 547972 146066 548024 146072
rect 547972 143608 548024 143614
rect 547972 143550 548024 143556
rect 547984 133074 548012 143550
rect 548076 140078 548104 146775
rect 548064 140072 548116 140078
rect 548064 140014 548116 140020
rect 547972 133068 548024 133074
rect 547972 133010 548024 133016
rect 548064 131504 548116 131510
rect 548064 131446 548116 131452
rect 547800 131158 547920 131186
rect 547800 126993 547828 131158
rect 547786 126984 547842 126993
rect 547786 126919 547842 126928
rect 547880 121304 547932 121310
rect 547880 121246 547932 121252
rect 547788 116680 547840 116686
rect 547788 116622 547840 116628
rect 547800 114918 547828 116622
rect 547788 114912 547840 114918
rect 547788 114854 547840 114860
rect 547892 114646 547920 121246
rect 547972 114912 548024 114918
rect 547972 114854 548024 114860
rect 547880 114640 547932 114646
rect 547880 114582 547932 114588
rect 547880 113552 547932 113558
rect 547880 113494 547932 113500
rect 547892 108934 547920 113494
rect 547984 113218 548012 114854
rect 548076 114578 548104 131446
rect 548064 114572 548116 114578
rect 548064 114514 548116 114520
rect 547972 113212 548024 113218
rect 547972 113154 548024 113160
rect 547970 109032 548026 109041
rect 547970 108967 548026 108976
rect 547880 108928 547932 108934
rect 547880 108870 547932 108876
rect 547880 95328 547932 95334
rect 547880 95270 547932 95276
rect 547892 89622 547920 95270
rect 547984 95266 548012 108967
rect 547972 95260 548024 95266
rect 547972 95202 548024 95208
rect 547880 89616 547932 89622
rect 547880 89558 547932 89564
rect 547972 89548 548024 89554
rect 547972 89490 548024 89496
rect 547880 83972 547932 83978
rect 547880 83914 547932 83920
rect 547892 72457 547920 83914
rect 547984 83026 548012 89490
rect 547972 83020 548024 83026
rect 547972 82962 548024 82968
rect 547878 72448 547934 72457
rect 547878 72383 547934 72392
rect 548168 29578 548196 151302
rect 548260 131306 548288 229910
rect 548340 163600 548392 163606
rect 548340 163542 548392 163548
rect 548248 131300 548300 131306
rect 548248 131242 548300 131248
rect 548248 73160 548300 73166
rect 548248 73102 548300 73108
rect 548156 29572 548208 29578
rect 548156 29514 548208 29520
rect 547696 25560 547748 25566
rect 547696 25502 547748 25508
rect 547604 22772 547656 22778
rect 547604 22714 547656 22720
rect 547236 20664 547288 20670
rect 547236 20606 547288 20612
rect 548260 11014 548288 73102
rect 548352 29510 548380 163542
rect 548432 151632 548484 151638
rect 548432 151574 548484 151580
rect 548340 29504 548392 29510
rect 548340 29446 548392 29452
rect 548444 24342 548472 151574
rect 548536 149802 548564 233038
rect 548996 229094 549024 237215
rect 549088 233866 549116 239498
rect 549180 238066 549208 239822
rect 549168 238060 549220 238066
rect 549168 238002 549220 238008
rect 549272 237425 549300 240178
rect 549536 240168 549588 240174
rect 549536 240110 549588 240116
rect 549258 237416 549314 237425
rect 549258 237351 549314 237360
rect 549088 233838 549208 233866
rect 548996 229066 549116 229094
rect 548892 153944 548944 153950
rect 548892 153886 548944 153892
rect 548706 149968 548762 149977
rect 548706 149903 548762 149912
rect 548524 149796 548576 149802
rect 548524 149738 548576 149744
rect 548720 138014 548748 149903
rect 548720 137986 548840 138014
rect 548524 133204 548576 133210
rect 548524 133146 548576 133152
rect 548536 121514 548564 133146
rect 548616 131028 548668 131034
rect 548616 130970 548668 130976
rect 548524 121508 548576 121514
rect 548524 121450 548576 121456
rect 548524 119400 548576 119406
rect 548524 119342 548576 119348
rect 548432 24336 548484 24342
rect 548432 24278 548484 24284
rect 548536 16386 548564 119342
rect 548628 27266 548656 130970
rect 548812 116686 548840 137986
rect 548800 116680 548852 116686
rect 548800 116622 548852 116628
rect 548800 115524 548852 115530
rect 548800 115466 548852 115472
rect 548708 105936 548760 105942
rect 548708 105878 548760 105884
rect 548616 27260 548668 27266
rect 548616 27202 548668 27208
rect 548524 16380 548576 16386
rect 548524 16322 548576 16328
rect 548720 13054 548748 105878
rect 548812 102134 548840 115466
rect 548800 102128 548852 102134
rect 548800 102070 548852 102076
rect 548800 94240 548852 94246
rect 548800 94182 548852 94188
rect 548708 13048 548760 13054
rect 548708 12990 548760 12996
rect 548248 11008 548300 11014
rect 548248 10950 548300 10956
rect 548812 6594 548840 94182
rect 548904 28286 548932 153886
rect 549088 150686 549116 229066
rect 549076 150680 549128 150686
rect 549076 150622 549128 150628
rect 548984 132388 549036 132394
rect 548984 132330 549036 132336
rect 548996 107914 549024 132330
rect 549076 122732 549128 122738
rect 549076 122674 549128 122680
rect 549088 117230 549116 122674
rect 549180 118833 549208 233838
rect 549442 230072 549498 230081
rect 549442 230007 549498 230016
rect 549352 229832 549404 229838
rect 549352 229774 549404 229780
rect 549260 162308 549312 162314
rect 549260 162250 549312 162256
rect 549272 143614 549300 162250
rect 549364 145654 549392 229774
rect 549456 147665 549484 230007
rect 549548 198762 549576 240110
rect 549640 240094 549792 240122
rect 549640 237522 549668 240094
rect 549628 237516 549680 237522
rect 549628 237458 549680 237464
rect 550008 235890 550036 240246
rect 549996 235884 550048 235890
rect 549996 235826 550048 235832
rect 549904 232688 549956 232694
rect 549904 232630 549956 232636
rect 549536 198756 549588 198762
rect 549536 198698 549588 198704
rect 549536 160880 549588 160886
rect 549536 160822 549588 160828
rect 549442 147656 549498 147665
rect 549442 147591 549498 147600
rect 549352 145648 549404 145654
rect 549352 145590 549404 145596
rect 549352 145512 549404 145518
rect 549352 145454 549404 145460
rect 549260 143608 549312 143614
rect 549260 143550 549312 143556
rect 549260 135176 549312 135182
rect 549260 135118 549312 135124
rect 549272 120426 549300 135118
rect 549260 120420 549312 120426
rect 549260 120362 549312 120368
rect 549166 118824 549222 118833
rect 549166 118759 549222 118768
rect 549076 117224 549128 117230
rect 549076 117166 549128 117172
rect 548984 107908 549036 107914
rect 548984 107850 549036 107856
rect 549260 85808 549312 85814
rect 549260 85750 549312 85756
rect 549272 70514 549300 85750
rect 549260 70508 549312 70514
rect 549260 70450 549312 70456
rect 548892 28280 548944 28286
rect 548892 28222 548944 28228
rect 549364 12238 549392 145454
rect 549444 144152 549496 144158
rect 549444 144094 549496 144100
rect 549456 135930 549484 144094
rect 549444 135924 549496 135930
rect 549444 135866 549496 135872
rect 549444 135312 549496 135318
rect 549444 135254 549496 135260
rect 549456 13394 549484 135254
rect 549548 64054 549576 160822
rect 549812 158160 549864 158166
rect 549812 158102 549864 158108
rect 549718 151056 549774 151065
rect 549718 150991 549774 151000
rect 549628 150408 549680 150414
rect 549628 150350 549680 150356
rect 549640 108458 549668 150350
rect 549628 108452 549680 108458
rect 549628 108394 549680 108400
rect 549628 101856 549680 101862
rect 549628 101798 549680 101804
rect 549640 89486 549668 101798
rect 549732 91254 549760 150991
rect 549824 146962 549852 158102
rect 549916 148442 549944 232630
rect 550100 186998 550128 297871
rect 550088 186992 550140 186998
rect 550088 186934 550140 186940
rect 550088 158296 550140 158302
rect 550088 158238 550140 158244
rect 550100 151814 550128 158238
rect 550008 151786 550128 151814
rect 549904 148436 549956 148442
rect 549904 148378 549956 148384
rect 550008 148374 550036 151786
rect 550088 149728 550140 149734
rect 550088 149670 550140 149676
rect 550100 149002 550128 149670
rect 550192 149161 550220 459711
rect 550284 431905 550312 698906
rect 551100 693456 551152 693462
rect 551100 693398 551152 693404
rect 550640 687948 550692 687954
rect 550640 687890 550692 687896
rect 550652 507385 550680 687890
rect 550732 681012 550784 681018
rect 550732 680954 550784 680960
rect 550638 507376 550694 507385
rect 550638 507311 550694 507320
rect 550362 495816 550418 495825
rect 550362 495751 550418 495760
rect 550270 431896 550326 431905
rect 550270 431831 550326 431840
rect 550376 248414 550404 495751
rect 550744 271425 550772 680954
rect 550916 680604 550968 680610
rect 550916 680546 550968 680552
rect 550824 679040 550876 679046
rect 550824 678982 550876 678988
rect 550836 600545 550864 678982
rect 550928 605985 550956 680546
rect 551008 680400 551060 680406
rect 551008 680342 551060 680348
rect 550914 605976 550970 605985
rect 550914 605911 550970 605920
rect 550822 600536 550878 600545
rect 550822 600471 550878 600480
rect 550822 596456 550878 596465
rect 550822 596391 550878 596400
rect 550730 271416 550786 271425
rect 550730 271351 550786 271360
rect 550730 268696 550786 268705
rect 550730 268631 550786 268640
rect 550376 248386 550496 248414
rect 550364 241528 550416 241534
rect 550364 241470 550416 241476
rect 550270 240816 550326 240825
rect 550270 240751 550326 240760
rect 550284 240174 550312 240751
rect 550272 240168 550324 240174
rect 550272 240110 550324 240116
rect 550376 234614 550404 241470
rect 550468 240310 550496 248386
rect 550638 247616 550694 247625
rect 550638 247551 550694 247560
rect 550548 240576 550600 240582
rect 550548 240518 550600 240524
rect 550456 240304 550508 240310
rect 550456 240246 550508 240252
rect 550456 240168 550508 240174
rect 550456 240110 550508 240116
rect 550468 239630 550496 240110
rect 550456 239624 550508 239630
rect 550456 239566 550508 239572
rect 550284 234586 550404 234614
rect 550178 149152 550234 149161
rect 550178 149087 550234 149096
rect 550100 148974 550220 149002
rect 549996 148368 550048 148374
rect 549996 148310 550048 148316
rect 549824 146934 550036 146962
rect 549812 146872 549864 146878
rect 549812 146814 549864 146820
rect 549904 146872 549956 146878
rect 549904 146814 549956 146820
rect 549824 137290 549852 146814
rect 549812 137284 549864 137290
rect 549812 137226 549864 137232
rect 549916 133929 549944 146814
rect 549902 133920 549958 133929
rect 549902 133855 549958 133864
rect 550008 122834 550036 146934
rect 550192 142050 550220 148974
rect 550180 142044 550232 142050
rect 550180 141986 550232 141992
rect 549824 122806 550036 122834
rect 549720 91248 549772 91254
rect 549720 91190 549772 91196
rect 549720 90908 549772 90914
rect 549720 90850 549772 90856
rect 549628 89480 549680 89486
rect 549628 89422 549680 89428
rect 549536 64048 549588 64054
rect 549536 63990 549588 63996
rect 549732 16590 549760 90850
rect 549824 74594 549852 122806
rect 549996 120148 550048 120154
rect 549996 120090 550048 120096
rect 549904 113144 549956 113150
rect 549904 113086 549956 113092
rect 549916 103154 549944 113086
rect 550008 111858 550036 120090
rect 549996 111852 550048 111858
rect 549996 111794 550048 111800
rect 550088 108928 550140 108934
rect 550088 108870 550140 108876
rect 549904 103148 549956 103154
rect 549904 103090 549956 103096
rect 549996 100768 550048 100774
rect 549996 100710 550048 100716
rect 549812 74588 549864 74594
rect 549812 74530 549864 74536
rect 549904 73228 549956 73234
rect 549904 73170 549956 73176
rect 549812 71732 549864 71738
rect 549812 71674 549864 71680
rect 549824 19310 549852 71674
rect 549812 19304 549864 19310
rect 549812 19246 549864 19252
rect 549720 16584 549772 16590
rect 549720 16526 549772 16532
rect 549916 13705 549944 73170
rect 550008 72282 550036 100710
rect 549996 72276 550048 72282
rect 549996 72218 550048 72224
rect 550100 19854 550128 108870
rect 550284 75274 550312 234586
rect 550560 219434 550588 240518
rect 550652 236706 550680 247551
rect 550640 236700 550692 236706
rect 550640 236642 550692 236648
rect 550468 219406 550588 219434
rect 550468 197266 550496 219406
rect 550456 197260 550508 197266
rect 550456 197202 550508 197208
rect 550744 182918 550772 268631
rect 550836 238270 550864 596391
rect 550914 562456 550970 562465
rect 550914 562391 550970 562400
rect 550824 238264 550876 238270
rect 550824 238206 550876 238212
rect 550928 236570 550956 562391
rect 551020 468625 551048 680342
rect 551112 555665 551140 693398
rect 551284 682780 551336 682786
rect 551284 682722 551336 682728
rect 551192 680808 551244 680814
rect 551192 680750 551244 680756
rect 551204 622985 551232 680750
rect 551296 667894 551324 682722
rect 551284 667888 551336 667894
rect 551284 667830 551336 667836
rect 551190 622976 551246 622985
rect 551190 622911 551246 622920
rect 551284 615936 551336 615942
rect 551284 615878 551336 615884
rect 551098 555656 551154 555665
rect 551098 555591 551154 555600
rect 551098 539336 551154 539345
rect 551098 539271 551154 539280
rect 551006 468616 551062 468625
rect 551006 468551 551062 468560
rect 551006 323776 551062 323785
rect 551006 323711 551062 323720
rect 550916 236564 550968 236570
rect 550916 236506 550968 236512
rect 550822 232792 550878 232801
rect 550822 232727 550878 232736
rect 550732 182912 550784 182918
rect 550732 182854 550784 182860
rect 550836 146878 550864 232727
rect 550916 162784 550968 162790
rect 550916 162726 550968 162732
rect 550824 146872 550876 146878
rect 550824 146814 550876 146820
rect 550364 146260 550416 146266
rect 550364 146202 550416 146208
rect 550272 75268 550324 75274
rect 550272 75210 550324 75216
rect 550088 19848 550140 19854
rect 550088 19790 550140 19796
rect 549902 13696 549958 13705
rect 549902 13631 549958 13640
rect 549444 13388 549496 13394
rect 549444 13330 549496 13336
rect 549352 12232 549404 12238
rect 549352 12174 549404 12180
rect 548800 6588 548852 6594
rect 548800 6530 548852 6536
rect 550376 5506 550404 146202
rect 550732 109744 550784 109750
rect 550732 109686 550784 109692
rect 550640 108316 550692 108322
rect 550640 108258 550692 108264
rect 550652 87650 550680 108258
rect 550744 100774 550772 109686
rect 550732 100768 550784 100774
rect 550732 100710 550784 100716
rect 550640 87644 550692 87650
rect 550640 87586 550692 87592
rect 550928 29102 550956 162726
rect 550916 29096 550968 29102
rect 550916 29038 550968 29044
rect 551020 12918 551048 323711
rect 551112 238814 551140 539271
rect 551190 333976 551246 333985
rect 551190 333911 551246 333920
rect 551100 238808 551152 238814
rect 551100 238750 551152 238756
rect 551098 238640 551154 238649
rect 551098 238575 551154 238584
rect 551112 192545 551140 238575
rect 551204 198354 551232 333911
rect 551296 238406 551324 615878
rect 551388 546514 551416 700470
rect 566004 700460 566056 700466
rect 566004 700402 566056 700408
rect 551468 700392 551520 700398
rect 551468 700334 551520 700340
rect 551480 565894 551508 700334
rect 552204 697604 552256 697610
rect 552204 697546 552256 697552
rect 552112 680876 552164 680882
rect 552112 680818 552164 680824
rect 552020 679584 552072 679590
rect 552020 679526 552072 679532
rect 552032 678978 552060 679526
rect 552020 678972 552072 678978
rect 552020 678914 552072 678920
rect 552124 678858 552152 680818
rect 552032 678830 552152 678858
rect 552032 678178 552060 678830
rect 552110 678736 552166 678745
rect 552110 678671 552166 678680
rect 551940 678150 552060 678178
rect 551940 677498 551968 678150
rect 552018 678056 552074 678065
rect 552018 677991 552074 678000
rect 552032 677618 552060 677991
rect 552124 677686 552152 678671
rect 552112 677680 552164 677686
rect 552112 677622 552164 677628
rect 552020 677612 552072 677618
rect 552020 677554 552072 677560
rect 551940 677470 552152 677498
rect 552018 676016 552074 676025
rect 552018 675951 552074 675960
rect 552032 674898 552060 675951
rect 552020 674892 552072 674898
rect 552020 674834 552072 674840
rect 552018 672480 552074 672489
rect 552018 672415 552074 672424
rect 552032 672110 552060 672415
rect 552020 672104 552072 672110
rect 552020 672046 552072 672052
rect 552124 671922 552152 677470
rect 552032 671894 552152 671922
rect 552032 661745 552060 671894
rect 552112 671832 552164 671838
rect 552112 671774 552164 671780
rect 552018 661736 552074 661745
rect 552018 661671 552074 661680
rect 552020 642252 552072 642258
rect 552020 642194 552072 642200
rect 552032 642025 552060 642194
rect 552018 642016 552074 642025
rect 552018 641951 552074 641960
rect 552018 637936 552074 637945
rect 552018 637871 552074 637880
rect 552032 637634 552060 637871
rect 552020 637628 552072 637634
rect 552020 637570 552072 637576
rect 552018 631816 552074 631825
rect 552018 631751 552020 631760
rect 552072 631751 552074 631760
rect 552020 631722 552072 631728
rect 552020 603968 552072 603974
rect 552018 603936 552020 603945
rect 552072 603936 552074 603945
rect 552018 603871 552074 603880
rect 552032 598505 552060 603871
rect 552018 598496 552074 598505
rect 552018 598431 552074 598440
rect 552018 591016 552074 591025
rect 552018 590951 552074 590960
rect 552032 590850 552060 590951
rect 552020 590844 552072 590850
rect 552020 590786 552072 590792
rect 552020 589008 552072 589014
rect 552018 588976 552020 588985
rect 552072 588976 552074 588985
rect 552018 588911 552074 588920
rect 552018 586936 552074 586945
rect 552018 586871 552074 586880
rect 552032 586566 552060 586871
rect 552020 586560 552072 586566
rect 552020 586502 552072 586508
rect 552018 585576 552074 585585
rect 552018 585511 552074 585520
rect 552032 585206 552060 585511
rect 552020 585200 552072 585206
rect 552020 585142 552072 585148
rect 552018 579456 552074 579465
rect 552018 579391 552074 579400
rect 552032 578270 552060 579391
rect 552020 578264 552072 578270
rect 552020 578206 552072 578212
rect 552018 578096 552074 578105
rect 552018 578031 552074 578040
rect 552032 577522 552060 578031
rect 552020 577516 552072 577522
rect 552020 577458 552072 577464
rect 552018 576056 552074 576065
rect 552018 575991 552074 576000
rect 552032 575550 552060 575991
rect 552020 575544 552072 575550
rect 552020 575486 552072 575492
rect 552018 574560 552074 574569
rect 552018 574495 552074 574504
rect 552032 574122 552060 574495
rect 552020 574116 552072 574122
rect 552020 574058 552072 574064
rect 552018 574016 552074 574025
rect 552018 573951 552074 573960
rect 552032 572762 552060 573951
rect 552020 572756 552072 572762
rect 552020 572698 552072 572704
rect 551468 565888 551520 565894
rect 551468 565830 551520 565836
rect 552020 553716 552072 553722
rect 552020 553658 552072 553664
rect 552032 553625 552060 553658
rect 552018 553616 552074 553625
rect 552018 553551 552074 553560
rect 552018 550896 552074 550905
rect 552018 550831 552020 550840
rect 552072 550831 552074 550840
rect 552020 550802 552072 550808
rect 552124 547505 552152 671774
rect 552110 547496 552166 547505
rect 552110 547431 552166 547440
rect 551376 546508 551428 546514
rect 551376 546450 551428 546456
rect 552020 546508 552072 546514
rect 552020 546450 552072 546456
rect 552032 522345 552060 546450
rect 552110 545456 552166 545465
rect 552110 545391 552166 545400
rect 552018 522336 552074 522345
rect 552018 522271 552074 522280
rect 552018 521656 552074 521665
rect 552018 521591 552074 521600
rect 552032 520334 552060 521591
rect 552020 520328 552072 520334
rect 552020 520270 552072 520276
rect 552018 519480 552074 519489
rect 552018 519415 552074 519424
rect 552032 519314 552060 519415
rect 552020 519308 552072 519314
rect 552020 519250 552072 519256
rect 552020 519036 552072 519042
rect 552020 518978 552072 518984
rect 552032 518945 552060 518978
rect 552018 518936 552074 518945
rect 552018 518871 552074 518880
rect 552018 516896 552074 516905
rect 552018 516831 552074 516840
rect 552032 516186 552060 516831
rect 552020 516180 552072 516186
rect 552020 516122 552072 516128
rect 552018 514856 552074 514865
rect 552018 514791 552020 514800
rect 552072 514791 552074 514800
rect 552020 514762 552072 514768
rect 551558 484936 551614 484945
rect 551558 484871 551614 484880
rect 551374 282296 551430 282305
rect 551374 282231 551430 282240
rect 551388 239018 551416 282231
rect 551376 239012 551428 239018
rect 551376 238954 551428 238960
rect 551284 238400 551336 238406
rect 551284 238342 551336 238348
rect 551284 235136 551336 235142
rect 551284 235078 551336 235084
rect 551192 198348 551244 198354
rect 551192 198290 551244 198296
rect 551098 192536 551154 192545
rect 551098 192471 551154 192480
rect 551190 160848 551246 160857
rect 551190 160783 551246 160792
rect 551100 149932 551152 149938
rect 551100 149874 551152 149880
rect 551112 20262 551140 149874
rect 551204 49706 551232 160783
rect 551296 131034 551324 235078
rect 551376 151088 551428 151094
rect 551376 151030 551428 151036
rect 551284 131028 551336 131034
rect 551284 130970 551336 130976
rect 551284 129668 551336 129674
rect 551284 129610 551336 129616
rect 551296 108390 551324 129610
rect 551388 110430 551416 151030
rect 551466 147520 551522 147529
rect 551466 147455 551522 147464
rect 551480 129742 551508 147455
rect 551468 129736 551520 129742
rect 551468 129678 551520 129684
rect 551376 110424 551428 110430
rect 551376 110366 551428 110372
rect 551284 108384 551336 108390
rect 551284 108326 551336 108332
rect 551284 98660 551336 98666
rect 551284 98602 551336 98608
rect 551192 49700 551244 49706
rect 551192 49642 551244 49648
rect 551100 20256 551152 20262
rect 551100 20198 551152 20204
rect 551296 13598 551324 98602
rect 551376 80096 551428 80102
rect 551376 80038 551428 80044
rect 551388 14822 551416 80038
rect 551376 14816 551428 14822
rect 551376 14758 551428 14764
rect 551284 13592 551336 13598
rect 551284 13534 551336 13540
rect 551008 12912 551060 12918
rect 551008 12854 551060 12860
rect 551572 11898 551600 484871
rect 552018 465896 552074 465905
rect 552018 465831 552074 465840
rect 552032 465118 552060 465831
rect 552020 465112 552072 465118
rect 552020 465054 552072 465060
rect 552018 464400 552074 464409
rect 552018 464335 552074 464344
rect 552032 463962 552060 464335
rect 552020 463956 552072 463962
rect 552020 463898 552072 463904
rect 552018 463176 552074 463185
rect 552018 463111 552074 463120
rect 552032 462398 552060 463111
rect 552020 462392 552072 462398
rect 552020 462334 552072 462340
rect 552018 460456 552074 460465
rect 552018 460391 552074 460400
rect 552032 459610 552060 460391
rect 552020 459604 552072 459610
rect 552020 459546 552072 459552
rect 552018 459096 552074 459105
rect 552018 459031 552020 459040
rect 552072 459031 552074 459040
rect 552020 459002 552072 459008
rect 552018 457736 552074 457745
rect 552018 457671 552074 457680
rect 552032 456822 552060 457671
rect 552020 456816 552072 456822
rect 552020 456758 552072 456764
rect 552018 456376 552074 456385
rect 552018 456311 552074 456320
rect 552032 456074 552060 456311
rect 552020 456068 552072 456074
rect 552020 456010 552072 456016
rect 552018 422376 552074 422385
rect 552018 422311 552074 422320
rect 552032 371385 552060 422311
rect 552018 371376 552074 371385
rect 552018 371311 552074 371320
rect 552020 368008 552072 368014
rect 552018 367976 552020 367985
rect 552072 367976 552074 367985
rect 552018 367911 552074 367920
rect 552018 365256 552074 365265
rect 552018 365191 552020 365200
rect 552072 365191 552074 365200
rect 552020 365162 552072 365168
rect 552020 342848 552072 342854
rect 552018 342816 552020 342825
rect 552072 342816 552074 342825
rect 552018 342751 552074 342760
rect 552018 322416 552074 322425
rect 552018 322351 552020 322360
rect 552072 322351 552074 322360
rect 552020 322322 552072 322328
rect 552020 307488 552072 307494
rect 552018 307456 552020 307465
rect 552072 307456 552074 307465
rect 552018 307391 552074 307400
rect 552018 293176 552074 293185
rect 552018 293111 552020 293120
rect 552072 293111 552074 293120
rect 552020 293082 552072 293088
rect 552018 291816 552074 291825
rect 552018 291751 552020 291760
rect 552072 291751 552074 291760
rect 552020 291722 552072 291728
rect 552124 267734 552152 545391
rect 552216 480185 552244 697546
rect 552848 696244 552900 696250
rect 552848 696186 552900 696192
rect 552296 683528 552348 683534
rect 552296 683470 552348 683476
rect 552308 525745 552336 683470
rect 552756 680740 552808 680746
rect 552756 680682 552808 680688
rect 552664 680536 552716 680542
rect 552664 680478 552716 680484
rect 552388 679516 552440 679522
rect 552388 679458 552440 679464
rect 552400 669314 552428 679458
rect 552478 679416 552534 679425
rect 552478 679351 552534 679360
rect 552492 679046 552520 679351
rect 552480 679040 552532 679046
rect 552480 678982 552532 678988
rect 552480 678904 552532 678910
rect 552480 678846 552532 678852
rect 552492 674665 552520 678846
rect 552478 674656 552534 674665
rect 552478 674591 552534 674600
rect 552572 674144 552624 674150
rect 552572 674086 552624 674092
rect 552400 669286 552520 669314
rect 552388 667888 552440 667894
rect 552388 667830 552440 667836
rect 552400 536625 552428 667830
rect 552492 640334 552520 669286
rect 552584 642705 552612 674086
rect 552676 654265 552704 680478
rect 552768 674150 552796 680682
rect 552756 674144 552808 674150
rect 552756 674086 552808 674092
rect 552754 670576 552810 670585
rect 552754 670511 552810 670520
rect 552768 669390 552796 670511
rect 552756 669384 552808 669390
rect 552756 669326 552808 669332
rect 552662 654256 552718 654265
rect 552662 654191 552718 654200
rect 552662 650176 552718 650185
rect 552662 650111 552718 650120
rect 552570 642696 552626 642705
rect 552570 642631 552626 642640
rect 552492 640306 552612 640334
rect 552478 638480 552534 638489
rect 552478 638415 552534 638424
rect 552492 637702 552520 638415
rect 552480 637696 552532 637702
rect 552480 637638 552532 637644
rect 552584 634545 552612 640306
rect 552570 634536 552626 634545
rect 552570 634471 552626 634480
rect 552676 615942 552704 650111
rect 552754 616176 552810 616185
rect 552754 616111 552810 616120
rect 552664 615936 552716 615942
rect 552664 615878 552716 615884
rect 552478 608696 552534 608705
rect 552478 608631 552480 608640
rect 552532 608631 552534 608640
rect 552480 608602 552532 608608
rect 552478 591424 552534 591433
rect 552478 591359 552534 591368
rect 552492 590714 552520 591359
rect 552480 590708 552532 590714
rect 552480 590650 552532 590656
rect 552480 565888 552532 565894
rect 552480 565830 552532 565836
rect 552386 536616 552442 536625
rect 552386 536551 552442 536560
rect 552388 532568 552440 532574
rect 552386 532536 552388 532545
rect 552440 532536 552442 532545
rect 552386 532471 552442 532480
rect 552388 530528 552440 530534
rect 552386 530496 552388 530505
rect 552440 530496 552442 530505
rect 552386 530431 552442 530440
rect 552386 526416 552442 526425
rect 552386 526351 552442 526360
rect 552400 526318 552428 526351
rect 552388 526312 552440 526318
rect 552388 526254 552440 526260
rect 552294 525736 552350 525745
rect 552294 525671 552350 525680
rect 552492 524385 552520 565830
rect 552570 544096 552626 544105
rect 552570 544031 552626 544040
rect 552584 543862 552612 544031
rect 552572 543856 552624 543862
rect 552572 543798 552624 543804
rect 552570 533896 552626 533905
rect 552570 533831 552626 533840
rect 552478 524376 552534 524385
rect 552478 524311 552534 524320
rect 552386 515536 552442 515545
rect 552386 515471 552442 515480
rect 552294 500576 552350 500585
rect 552294 500511 552350 500520
rect 552202 480176 552258 480185
rect 552202 480111 552258 480120
rect 552308 454345 552336 500511
rect 552294 454336 552350 454345
rect 552294 454271 552350 454280
rect 552202 451480 552258 451489
rect 552202 451415 552258 451424
rect 552216 432585 552244 451415
rect 552294 440736 552350 440745
rect 552294 440671 552350 440680
rect 552202 432576 552258 432585
rect 552202 432511 552258 432520
rect 552204 430228 552256 430234
rect 552204 430170 552256 430176
rect 552216 429865 552244 430170
rect 552202 429856 552258 429865
rect 552202 429791 552258 429800
rect 552204 421048 552256 421054
rect 552202 421016 552204 421025
rect 552256 421016 552258 421025
rect 552202 420951 552258 420960
rect 552202 393816 552258 393825
rect 552202 393751 552204 393760
rect 552256 393751 552258 393760
rect 552204 393722 552256 393728
rect 552202 372736 552258 372745
rect 552202 372671 552204 372680
rect 552256 372671 552258 372680
rect 552204 372642 552256 372648
rect 552202 369336 552258 369345
rect 552202 369271 552258 369280
rect 552216 368626 552244 369271
rect 552204 368620 552256 368626
rect 552204 368562 552256 368568
rect 552202 306096 552258 306105
rect 552202 306031 552258 306040
rect 552216 305522 552244 306031
rect 552204 305516 552256 305522
rect 552204 305458 552256 305464
rect 552124 267706 552244 267734
rect 552018 265296 552074 265305
rect 552018 265231 552020 265240
rect 552072 265231 552074 265240
rect 552020 265202 552072 265208
rect 552018 263256 552074 263265
rect 552018 263191 552020 263200
rect 552072 263191 552074 263200
rect 552020 263162 552072 263168
rect 552018 261896 552074 261905
rect 552018 261831 552074 261840
rect 552032 260914 552060 261831
rect 552020 260908 552072 260914
rect 552020 260850 552072 260856
rect 552110 260400 552166 260409
rect 552110 260335 552166 260344
rect 552018 259856 552074 259865
rect 552018 259791 552074 259800
rect 552032 259486 552060 259791
rect 552124 259554 552152 260335
rect 552112 259548 552164 259554
rect 552112 259490 552164 259496
rect 552020 259480 552072 259486
rect 552020 259422 552072 259428
rect 552110 259176 552166 259185
rect 552110 259111 552166 259120
rect 552018 258496 552074 258505
rect 552018 258431 552074 258440
rect 552032 258126 552060 258431
rect 552124 258194 552152 259111
rect 552112 258188 552164 258194
rect 552112 258130 552164 258136
rect 552020 258120 552072 258126
rect 552020 258062 552072 258068
rect 552018 257816 552074 257825
rect 552018 257751 552074 257760
rect 552032 256766 552060 257751
rect 552020 256760 552072 256766
rect 552020 256702 552072 256708
rect 552110 255096 552166 255105
rect 552110 255031 552166 255040
rect 552018 254416 552074 254425
rect 552018 254351 552074 254360
rect 552032 253978 552060 254351
rect 552124 254046 552152 255031
rect 552112 254040 552164 254046
rect 552112 253982 552164 253988
rect 552020 253972 552072 253978
rect 552020 253914 552072 253920
rect 552018 250336 552074 250345
rect 552018 250271 552074 250280
rect 552032 249830 552060 250271
rect 552020 249824 552072 249830
rect 552020 249766 552072 249772
rect 552216 248414 552244 267706
rect 552124 248386 552244 248414
rect 552018 242856 552074 242865
rect 552018 242791 552074 242800
rect 552032 239698 552060 242791
rect 552124 241534 552152 248386
rect 552202 246256 552258 246265
rect 552202 246191 552258 246200
rect 552216 245750 552244 246191
rect 552204 245744 552256 245750
rect 552204 245686 552256 245692
rect 552202 243400 552258 243409
rect 552202 243335 552258 243344
rect 552112 241528 552164 241534
rect 552112 241470 552164 241476
rect 552020 239692 552072 239698
rect 552020 239634 552072 239640
rect 552216 236842 552244 243335
rect 552204 236836 552256 236842
rect 552204 236778 552256 236784
rect 552112 235068 552164 235074
rect 552112 235010 552164 235016
rect 551650 162344 551706 162353
rect 551650 162279 551706 162288
rect 551664 24070 551692 162279
rect 551744 151496 551796 151502
rect 551744 151438 551796 151444
rect 551652 24064 551704 24070
rect 551652 24006 551704 24012
rect 551756 15774 551784 151438
rect 552020 133136 552072 133142
rect 552020 133078 552072 133084
rect 552032 129674 552060 133078
rect 552124 132802 552152 235010
rect 552308 177342 552336 440671
rect 552400 421705 552428 515471
rect 552584 492425 552612 533831
rect 552662 493776 552718 493785
rect 552662 493711 552718 493720
rect 552676 492726 552704 493711
rect 552664 492720 552716 492726
rect 552664 492662 552716 492668
rect 552570 492416 552626 492425
rect 552570 492351 552626 492360
rect 552662 484256 552718 484265
rect 552662 484191 552718 484200
rect 552676 483070 552704 484191
rect 552664 483064 552716 483070
rect 552664 483006 552716 483012
rect 552570 476096 552626 476105
rect 552570 476031 552626 476040
rect 552584 474842 552612 476031
rect 552572 474836 552624 474842
rect 552572 474778 552624 474784
rect 552570 449576 552626 449585
rect 552570 449511 552626 449520
rect 552584 448594 552612 449511
rect 552662 448896 552718 448905
rect 552662 448831 552718 448840
rect 552572 448588 552624 448594
rect 552572 448530 552624 448536
rect 552570 446856 552626 446865
rect 552570 446791 552626 446800
rect 552584 445806 552612 446791
rect 552572 445800 552624 445806
rect 552572 445742 552624 445748
rect 552570 445496 552626 445505
rect 552570 445431 552626 445440
rect 552584 444446 552612 445431
rect 552572 444440 552624 444446
rect 552572 444382 552624 444388
rect 552386 421696 552442 421705
rect 552386 421631 552442 421640
rect 552386 412856 552442 412865
rect 552386 412791 552388 412800
rect 552440 412791 552442 412800
rect 552388 412762 552440 412768
rect 552478 407416 552534 407425
rect 552478 407351 552534 407360
rect 552386 354376 552442 354385
rect 552386 354311 552442 354320
rect 552400 187066 552428 354311
rect 552492 240242 552520 407351
rect 552570 331256 552626 331265
rect 552570 331191 552626 331200
rect 552480 240236 552532 240242
rect 552480 240178 552532 240184
rect 552480 234116 552532 234122
rect 552480 234058 552532 234064
rect 552388 187060 552440 187066
rect 552388 187002 552440 187008
rect 552296 177336 552348 177342
rect 552296 177278 552348 177284
rect 552388 160744 552440 160750
rect 552388 160686 552440 160692
rect 552296 151224 552348 151230
rect 552296 151166 552348 151172
rect 552112 132796 552164 132802
rect 552112 132738 552164 132744
rect 552112 129736 552164 129742
rect 552112 129678 552164 129684
rect 552020 129668 552072 129674
rect 552020 129610 552072 129616
rect 552124 120154 552152 129678
rect 552112 120148 552164 120154
rect 552112 120090 552164 120096
rect 552112 117224 552164 117230
rect 552112 117166 552164 117172
rect 552124 105942 552152 117166
rect 552204 116612 552256 116618
rect 552204 116554 552256 116560
rect 552112 105936 552164 105942
rect 552112 105878 552164 105884
rect 552216 21962 552244 116554
rect 552308 70378 552336 151166
rect 552400 82822 552428 160686
rect 552492 123418 552520 234058
rect 552584 178702 552612 331191
rect 552676 252550 552704 448831
rect 552768 317626 552796 616111
rect 552860 597825 552888 696186
rect 554872 687268 554924 687274
rect 554872 687210 554924 687216
rect 554044 683664 554096 683670
rect 554044 683606 554096 683612
rect 553676 683460 553728 683466
rect 553676 683402 553728 683408
rect 553584 683392 553636 683398
rect 553584 683334 553636 683340
rect 553492 682712 553544 682718
rect 553492 682654 553544 682660
rect 553400 682508 553452 682514
rect 553400 682450 553452 682456
rect 552940 680944 552992 680950
rect 552940 680886 552992 680892
rect 552952 671838 552980 680886
rect 553122 679824 553178 679833
rect 553122 679759 553178 679768
rect 552940 671832 552992 671838
rect 552940 671774 552992 671780
rect 553136 665825 553164 679759
rect 553122 665816 553178 665825
rect 553122 665751 553178 665760
rect 553306 656976 553362 656985
rect 553306 656911 553308 656920
rect 553360 656911 553362 656920
rect 553308 656882 553360 656888
rect 553306 653576 553362 653585
rect 553306 653511 553362 653520
rect 553320 652798 553348 653511
rect 553308 652792 553360 652798
rect 553308 652734 553360 652740
rect 553306 648816 553362 648825
rect 553306 648751 553362 648760
rect 553320 648650 553348 648751
rect 553308 648644 553360 648650
rect 553308 648586 553360 648592
rect 552938 646776 552994 646785
rect 552938 646711 552994 646720
rect 552952 646202 552980 646711
rect 552940 646196 552992 646202
rect 552940 646138 552992 646144
rect 553306 645416 553362 645425
rect 553306 645351 553362 645360
rect 552938 644736 552994 644745
rect 552938 644671 552940 644680
rect 552992 644671 552994 644680
rect 552940 644642 552992 644648
rect 553320 644502 553348 645351
rect 553308 644496 553360 644502
rect 553308 644438 553360 644444
rect 553306 630456 553362 630465
rect 553306 630391 553362 630400
rect 553320 629338 553348 630391
rect 553308 629332 553360 629338
rect 553308 629274 553360 629280
rect 553306 624336 553362 624345
rect 553306 624271 553362 624280
rect 553320 623830 553348 624271
rect 553308 623824 553360 623830
rect 553308 623766 553360 623772
rect 553306 620256 553362 620265
rect 553306 620191 553362 620200
rect 553320 619682 553348 620191
rect 553308 619676 553360 619682
rect 553308 619618 553360 619624
rect 553306 617536 553362 617545
rect 553306 617471 553362 617480
rect 553320 616894 553348 617471
rect 553308 616888 553360 616894
rect 553308 616830 553360 616836
rect 553306 614816 553362 614825
rect 553306 614751 553362 614760
rect 553320 614174 553348 614751
rect 553308 614168 553360 614174
rect 553308 614110 553360 614116
rect 553306 613456 553362 613465
rect 553306 613391 553362 613400
rect 553320 612814 553348 613391
rect 553308 612808 553360 612814
rect 553308 612750 553360 612756
rect 553306 611416 553362 611425
rect 553306 611351 553308 611360
rect 553360 611351 553362 611360
rect 553308 611322 553360 611328
rect 553306 610736 553362 610745
rect 553306 610671 553362 610680
rect 553320 610026 553348 610671
rect 553308 610020 553360 610026
rect 553308 609962 553360 609968
rect 553306 607336 553362 607345
rect 553306 607271 553362 607280
rect 553320 607238 553348 607271
rect 553308 607232 553360 607238
rect 553308 607174 553360 607180
rect 553306 603256 553362 603265
rect 553306 603191 553362 603200
rect 553320 603158 553348 603191
rect 553308 603152 553360 603158
rect 553308 603094 553360 603100
rect 552846 597816 552902 597825
rect 552846 597751 552902 597760
rect 553214 584896 553270 584905
rect 553214 584831 553270 584840
rect 553122 568576 553178 568585
rect 553122 568511 553178 568520
rect 553136 567322 553164 568511
rect 553124 567316 553176 567322
rect 553124 567258 553176 567264
rect 553122 561096 553178 561105
rect 553122 561031 553178 561040
rect 553136 560318 553164 561031
rect 553124 560312 553176 560318
rect 553124 560254 553176 560260
rect 552938 558376 552994 558385
rect 552938 558311 552994 558320
rect 552952 558006 552980 558311
rect 552940 558000 552992 558006
rect 552940 557942 552992 557948
rect 553122 540696 553178 540705
rect 553122 540631 553178 540640
rect 553136 539646 553164 540631
rect 553124 539640 553176 539646
rect 553124 539582 553176 539588
rect 553122 493096 553178 493105
rect 553122 493031 553178 493040
rect 552846 453656 552902 453665
rect 552846 453591 552902 453600
rect 552860 452810 552888 453591
rect 552848 452804 552900 452810
rect 552848 452746 552900 452752
rect 553030 438696 553086 438705
rect 553030 438631 553086 438640
rect 553044 437442 553072 438631
rect 553032 437436 553084 437442
rect 553032 437378 553084 437384
rect 553030 437336 553086 437345
rect 553030 437271 553086 437280
rect 553044 436014 553072 437271
rect 553032 436008 553084 436014
rect 553032 435950 553084 435956
rect 553030 428496 553086 428505
rect 553030 428431 553086 428440
rect 553044 427854 553072 428431
rect 553032 427848 553084 427854
rect 553032 427790 553084 427796
rect 553032 426488 553084 426494
rect 553030 426456 553032 426465
rect 553084 426456 553086 426465
rect 553030 426391 553086 426400
rect 553032 425128 553084 425134
rect 553030 425096 553032 425105
rect 553084 425096 553086 425105
rect 553030 425031 553086 425040
rect 552938 424416 552994 424425
rect 552938 424351 552994 424360
rect 552952 423706 552980 424351
rect 553032 423768 553084 423774
rect 553030 423736 553032 423745
rect 553084 423736 553086 423745
rect 552940 423700 552992 423706
rect 553030 423671 553086 423680
rect 552940 423642 552992 423648
rect 553030 420336 553086 420345
rect 553030 420271 553086 420280
rect 553044 420170 553072 420271
rect 553032 420164 553084 420170
rect 553032 420106 553084 420112
rect 553030 416256 553086 416265
rect 553030 416191 553086 416200
rect 553044 416090 553072 416191
rect 553032 416084 553084 416090
rect 553032 416026 553084 416032
rect 553030 415576 553086 415585
rect 553030 415511 553086 415520
rect 553044 415478 553072 415511
rect 553032 415472 553084 415478
rect 553032 415414 553084 415420
rect 553030 413400 553086 413409
rect 553030 413335 553086 413344
rect 553044 412690 553072 413335
rect 553032 412684 553084 412690
rect 553032 412626 553084 412632
rect 553030 410816 553086 410825
rect 553030 410751 553086 410760
rect 553044 409902 553072 410751
rect 553032 409896 553084 409902
rect 553032 409838 553084 409844
rect 553032 405680 553084 405686
rect 553032 405622 553084 405628
rect 553044 405385 553072 405622
rect 553030 405376 553086 405385
rect 553030 405311 553086 405320
rect 553030 404016 553086 404025
rect 553030 403951 553086 403960
rect 553044 403714 553072 403951
rect 553032 403708 553084 403714
rect 553032 403650 553084 403656
rect 553030 403336 553086 403345
rect 553030 403271 553086 403280
rect 553044 403034 553072 403271
rect 553032 403028 553084 403034
rect 553032 402970 553084 402976
rect 553030 400480 553086 400489
rect 553030 400415 553086 400424
rect 553044 400246 553072 400415
rect 553032 400240 553084 400246
rect 553032 400182 553084 400188
rect 553030 395176 553086 395185
rect 553030 395111 553086 395120
rect 553044 394738 553072 395111
rect 553032 394732 553084 394738
rect 553032 394674 553084 394680
rect 553030 391776 553086 391785
rect 553030 391711 553086 391720
rect 553044 390658 553072 391711
rect 553032 390652 553084 390658
rect 553032 390594 553084 390600
rect 553030 390416 553086 390425
rect 553030 390351 553086 390360
rect 553044 389230 553072 390351
rect 553032 389224 553084 389230
rect 553032 389166 553084 389172
rect 553030 388376 553086 388385
rect 553030 388311 553086 388320
rect 553044 387870 553072 388311
rect 553032 387864 553084 387870
rect 553032 387806 553084 387812
rect 553030 387696 553086 387705
rect 553030 387631 553086 387640
rect 553044 386442 553072 387631
rect 553032 386436 553084 386442
rect 553032 386378 553084 386384
rect 553030 385656 553086 385665
rect 553030 385591 553086 385600
rect 553044 385082 553072 385591
rect 553032 385076 553084 385082
rect 553032 385018 553084 385024
rect 553030 381576 553086 381585
rect 553030 381511 553032 381520
rect 553084 381511 553086 381520
rect 553032 381482 553084 381488
rect 553032 378344 553084 378350
rect 553032 378286 553084 378292
rect 553044 378185 553072 378286
rect 553030 378176 553086 378185
rect 553030 378111 553086 378120
rect 553030 377496 553086 377505
rect 553030 377431 553086 377440
rect 553044 376786 553072 377431
rect 553032 376780 553084 376786
rect 553032 376722 553084 376728
rect 553030 370696 553086 370705
rect 553030 370631 553086 370640
rect 553044 369918 553072 370631
rect 553032 369912 553084 369918
rect 553032 369854 553084 369860
rect 553030 368656 553086 368665
rect 553030 368591 553086 368600
rect 553044 368558 553072 368591
rect 553032 368552 553084 368558
rect 553032 368494 553084 368500
rect 552938 366480 552994 366489
rect 552938 366415 552994 366424
rect 552952 365770 552980 366415
rect 553030 365936 553086 365945
rect 553030 365871 553086 365880
rect 553044 365838 553072 365871
rect 553032 365832 553084 365838
rect 553032 365774 553084 365780
rect 552940 365764 552992 365770
rect 552940 365706 552992 365712
rect 552938 361176 552994 361185
rect 552938 361111 552994 361120
rect 552952 360262 552980 361111
rect 553030 360496 553086 360505
rect 553030 360431 553032 360440
rect 553084 360431 553086 360440
rect 553032 360402 553084 360408
rect 552940 360256 552992 360262
rect 552940 360198 552992 360204
rect 553032 358760 553084 358766
rect 553032 358702 553084 358708
rect 552938 358456 552994 358465
rect 552938 358391 552994 358400
rect 552952 357474 552980 358391
rect 553044 357785 553072 358702
rect 553030 357776 553086 357785
rect 553030 357711 553086 357720
rect 552940 357468 552992 357474
rect 552940 357410 552992 357416
rect 553030 355736 553086 355745
rect 553030 355671 553086 355680
rect 553044 354754 553072 355671
rect 553032 354748 553084 354754
rect 553032 354690 553084 354696
rect 553030 353696 553086 353705
rect 553030 353631 553086 353640
rect 553044 353326 553072 353631
rect 553032 353320 553084 353326
rect 553032 353262 553084 353268
rect 552846 351656 552902 351665
rect 552846 351591 552902 351600
rect 552860 350606 552888 351591
rect 553136 351098 553164 493031
rect 552952 351070 553164 351098
rect 552848 350600 552900 350606
rect 552848 350542 552900 350548
rect 552952 340105 552980 351070
rect 553122 350976 553178 350985
rect 553122 350911 553124 350920
rect 553176 350911 553178 350920
rect 553124 350882 553176 350888
rect 553122 349480 553178 349489
rect 553122 349415 553178 349424
rect 553136 349178 553164 349415
rect 553124 349172 553176 349178
rect 553124 349114 553176 349120
rect 553030 347576 553086 347585
rect 553030 347511 553086 347520
rect 553044 346458 553072 347511
rect 553122 346896 553178 346905
rect 553122 346831 553178 346840
rect 553136 346526 553164 346831
rect 553124 346520 553176 346526
rect 553124 346462 553176 346468
rect 553032 346452 553084 346458
rect 553032 346394 553084 346400
rect 553030 343496 553086 343505
rect 553030 343431 553086 343440
rect 553044 343058 553072 343431
rect 553032 343052 553084 343058
rect 553032 342994 553084 343000
rect 552938 340096 552994 340105
rect 552938 340031 552994 340040
rect 553122 338736 553178 338745
rect 553122 338671 553178 338680
rect 553136 338162 553164 338671
rect 553124 338156 553176 338162
rect 553124 338098 553176 338104
rect 553030 336016 553086 336025
rect 553030 335951 553086 335960
rect 553044 335374 553072 335951
rect 553032 335368 553084 335374
rect 553032 335310 553084 335316
rect 553122 335336 553178 335345
rect 553122 335271 553124 335280
rect 553176 335271 553178 335280
rect 553124 335242 553176 335248
rect 552846 334656 552902 334665
rect 552846 334591 552902 334600
rect 552756 317620 552808 317626
rect 552756 317562 552808 317568
rect 552860 267734 552888 334591
rect 553030 327856 553086 327865
rect 553030 327791 553086 327800
rect 553044 327214 553072 327791
rect 553032 327208 553084 327214
rect 553032 327150 553084 327156
rect 553122 327176 553178 327185
rect 553122 327111 553124 327120
rect 553176 327111 553178 327120
rect 553124 327082 553176 327088
rect 553030 326496 553086 326505
rect 553030 326431 553086 326440
rect 553044 325786 553072 326431
rect 553122 325816 553178 325825
rect 553032 325780 553084 325786
rect 553122 325751 553178 325760
rect 553032 325722 553084 325728
rect 553136 325718 553164 325751
rect 553124 325712 553176 325718
rect 553124 325654 553176 325660
rect 553030 318336 553086 318345
rect 553030 318271 553086 318280
rect 553044 317490 553072 318271
rect 553122 317656 553178 317665
rect 553122 317591 553178 317600
rect 553136 317558 553164 317591
rect 553124 317552 553176 317558
rect 553124 317494 553176 317500
rect 553032 317484 553084 317490
rect 553032 317426 553084 317432
rect 553122 316296 553178 316305
rect 553122 316231 553178 316240
rect 553136 316062 553164 316231
rect 553124 316056 553176 316062
rect 553124 315998 553176 316004
rect 553122 314936 553178 314945
rect 553122 314871 553178 314880
rect 553136 314702 553164 314871
rect 553124 314696 553176 314702
rect 553124 314638 553176 314644
rect 553030 314256 553086 314265
rect 553030 314191 553086 314200
rect 553044 313342 553072 314191
rect 553032 313336 553084 313342
rect 553032 313278 553084 313284
rect 553124 313268 553176 313274
rect 553124 313210 553176 313216
rect 553136 312905 553164 313210
rect 553122 312896 553178 312905
rect 553122 312831 553178 312840
rect 553030 311400 553086 311409
rect 553030 311335 553086 311344
rect 553044 310554 553072 311335
rect 553122 310856 553178 310865
rect 553122 310791 553178 310800
rect 553136 310622 553164 310791
rect 553124 310616 553176 310622
rect 553124 310558 553176 310564
rect 553032 310548 553084 310554
rect 553032 310490 553084 310496
rect 553122 310176 553178 310185
rect 553122 310111 553178 310120
rect 553136 309194 553164 310111
rect 553124 309188 553176 309194
rect 553124 309130 553176 309136
rect 553122 308816 553178 308825
rect 553122 308751 553178 308760
rect 553136 307834 553164 308751
rect 553124 307828 553176 307834
rect 553124 307770 553176 307776
rect 553122 305416 553178 305425
rect 553122 305351 553178 305360
rect 553136 305046 553164 305351
rect 553124 305040 553176 305046
rect 553124 304982 553176 304988
rect 553030 302016 553086 302025
rect 553030 301951 553086 301960
rect 553044 300966 553072 301951
rect 553122 301336 553178 301345
rect 553122 301271 553178 301280
rect 553032 300960 553084 300966
rect 553032 300902 553084 300908
rect 553136 300898 553164 301271
rect 553124 300892 553176 300898
rect 553124 300834 553176 300840
rect 553122 300656 553178 300665
rect 553122 300591 553178 300600
rect 553136 299538 553164 300591
rect 553124 299532 553176 299538
rect 553124 299474 553176 299480
rect 553122 297256 553178 297265
rect 553122 297191 553178 297200
rect 553136 296750 553164 297191
rect 553124 296744 553176 296750
rect 553124 296686 553176 296692
rect 553122 292496 553178 292505
rect 553122 292431 553178 292440
rect 553136 291242 553164 292431
rect 553124 291236 553176 291242
rect 553124 291178 553176 291184
rect 553122 290456 553178 290465
rect 553122 290391 553178 290400
rect 553136 289882 553164 290391
rect 553124 289876 553176 289882
rect 553124 289818 553176 289824
rect 553030 289776 553086 289785
rect 553030 289711 553086 289720
rect 553044 288522 553072 289711
rect 553122 289096 553178 289105
rect 553122 289031 553178 289040
rect 553032 288516 553084 288522
rect 553032 288458 553084 288464
rect 553136 288454 553164 289031
rect 553124 288448 553176 288454
rect 553124 288390 553176 288396
rect 553122 287736 553178 287745
rect 553122 287671 553178 287680
rect 553136 287094 553164 287671
rect 553124 287088 553176 287094
rect 553124 287030 553176 287036
rect 553122 283656 553178 283665
rect 553122 283591 553124 283600
rect 553176 283591 553178 283600
rect 553124 283562 553176 283568
rect 553124 282872 553176 282878
rect 553124 282814 553176 282820
rect 553136 281625 553164 282814
rect 553122 281616 553178 281625
rect 553122 281551 553178 281560
rect 553030 280936 553086 280945
rect 553030 280871 553086 280880
rect 553044 280226 553072 280871
rect 553124 280288 553176 280294
rect 553122 280256 553124 280265
rect 553176 280256 553178 280265
rect 553032 280220 553084 280226
rect 553122 280191 553178 280200
rect 553032 280162 553084 280168
rect 553124 280152 553176 280158
rect 553124 280094 553176 280100
rect 553136 279585 553164 280094
rect 553122 279576 553178 279585
rect 553122 279511 553178 279520
rect 553122 278896 553178 278905
rect 553122 278831 553124 278840
rect 553176 278831 553178 278840
rect 553124 278802 553176 278808
rect 553122 277536 553178 277545
rect 553122 277471 553178 277480
rect 553136 277438 553164 277471
rect 553124 277432 553176 277438
rect 553124 277374 553176 277380
rect 553030 276176 553086 276185
rect 553030 276111 553032 276120
rect 553084 276111 553086 276120
rect 553032 276082 553084 276088
rect 553122 274816 553178 274825
rect 553122 274751 553178 274760
rect 553136 274718 553164 274751
rect 553124 274712 553176 274718
rect 553124 274654 553176 274660
rect 553122 273456 553178 273465
rect 553122 273391 553178 273400
rect 553136 273290 553164 273391
rect 553124 273284 553176 273290
rect 553124 273226 553176 273232
rect 553122 270736 553178 270745
rect 553122 270671 553178 270680
rect 553136 270570 553164 270671
rect 553124 270564 553176 270570
rect 553124 270506 553176 270512
rect 552860 267706 552980 267734
rect 552846 264616 552902 264625
rect 552846 264551 552902 264560
rect 552860 260438 552888 264551
rect 552952 260834 552980 267706
rect 553122 266656 553178 266665
rect 553122 266591 553178 266600
rect 553136 266422 553164 266591
rect 553124 266416 553176 266422
rect 553124 266358 553176 266364
rect 553122 263936 553178 263945
rect 553122 263871 553178 263880
rect 553136 263634 553164 263871
rect 553124 263628 553176 263634
rect 553124 263570 553176 263576
rect 552952 260806 553072 260834
rect 553044 260522 553072 260806
rect 552952 260494 553072 260522
rect 552848 260432 552900 260438
rect 552848 260374 552900 260380
rect 552664 252544 552716 252550
rect 552664 252486 552716 252492
rect 552664 249892 552716 249898
rect 552664 249834 552716 249840
rect 552572 178696 552624 178702
rect 552572 178638 552624 178644
rect 552572 160812 552624 160818
rect 552572 160754 552624 160760
rect 552480 123412 552532 123418
rect 552480 123354 552532 123360
rect 552480 103148 552532 103154
rect 552480 103090 552532 103096
rect 552388 82816 552440 82822
rect 552388 82758 552440 82764
rect 552492 80102 552520 103090
rect 552584 84182 552612 160754
rect 552572 84176 552624 84182
rect 552572 84118 552624 84124
rect 552480 80096 552532 80102
rect 552480 80038 552532 80044
rect 552296 70372 552348 70378
rect 552296 70314 552348 70320
rect 552676 28218 552704 249834
rect 552952 247722 552980 260494
rect 553032 260432 553084 260438
rect 553032 260374 553084 260380
rect 552940 247716 552992 247722
rect 552940 247658 552992 247664
rect 552756 239624 552808 239630
rect 552756 239566 552808 239572
rect 552768 200977 552796 239566
rect 552848 239488 552900 239494
rect 552848 239430 552900 239436
rect 552754 200968 552810 200977
rect 552754 200903 552810 200912
rect 552756 170400 552808 170406
rect 552756 170342 552808 170348
rect 552664 28212 552716 28218
rect 552664 28154 552716 28160
rect 552204 21956 552256 21962
rect 552204 21898 552256 21904
rect 551744 15768 551796 15774
rect 551744 15710 551796 15716
rect 551560 11892 551612 11898
rect 551560 11834 551612 11840
rect 550364 5500 550416 5506
rect 550364 5442 550416 5448
rect 547144 4820 547196 4826
rect 547144 4762 547196 4768
rect 549074 4040 549130 4049
rect 549074 3975 549130 3984
rect 546684 3188 546736 3194
rect 546684 3130 546736 3136
rect 549088 480 549116 3975
rect 552664 3800 552716 3806
rect 552664 3742 552716 3748
rect 552676 480 552704 3742
rect 552768 3058 552796 170342
rect 552860 167754 552888 239430
rect 553044 236881 553072 260374
rect 553122 253736 553178 253745
rect 553122 253671 553178 253680
rect 553136 252618 553164 253671
rect 553124 252612 553176 252618
rect 553124 252554 553176 252560
rect 553122 252376 553178 252385
rect 553122 252311 553178 252320
rect 553136 251258 553164 252311
rect 553124 251252 553176 251258
rect 553124 251194 553176 251200
rect 553122 248296 553178 248305
rect 553122 248231 553178 248240
rect 553136 247110 553164 248231
rect 553124 247104 553176 247110
rect 553124 247046 553176 247052
rect 553122 246936 553178 246945
rect 553122 246871 553178 246880
rect 553136 245682 553164 246871
rect 553124 245676 553176 245682
rect 553124 245618 553176 245624
rect 553122 244896 553178 244905
rect 553122 244831 553178 244840
rect 553136 244322 553164 244831
rect 553124 244316 553176 244322
rect 553124 244258 553176 244264
rect 553030 236872 553086 236881
rect 553030 236807 553086 236816
rect 553228 232529 553256 584831
rect 553306 567896 553362 567905
rect 553306 567831 553362 567840
rect 553320 567254 553348 567831
rect 553308 567248 553360 567254
rect 553308 567190 553360 567196
rect 553306 565176 553362 565185
rect 553306 565111 553362 565120
rect 553320 564466 553348 565111
rect 553308 564460 553360 564466
rect 553308 564402 553360 564408
rect 553306 560416 553362 560425
rect 553306 560351 553308 560360
rect 553360 560351 553362 560360
rect 553308 560322 553360 560328
rect 553306 557696 553362 557705
rect 553306 557631 553362 557640
rect 553320 557598 553348 557631
rect 553308 557592 553360 557598
rect 553308 557534 553360 557540
rect 553306 557016 553362 557025
rect 553306 556951 553362 556960
rect 553320 556578 553348 556951
rect 553308 556572 553360 556578
rect 553308 556514 553360 556520
rect 553306 556336 553362 556345
rect 553306 556271 553362 556280
rect 553320 556238 553348 556271
rect 553308 556232 553360 556238
rect 553308 556174 553360 556180
rect 553306 551576 553362 551585
rect 553306 551511 553362 551520
rect 553320 550662 553348 551511
rect 553308 550656 553360 550662
rect 553308 550598 553360 550604
rect 553306 549536 553362 549545
rect 553306 549471 553362 549480
rect 553320 549302 553348 549471
rect 553308 549296 553360 549302
rect 553308 549238 553360 549244
rect 553306 540016 553362 540025
rect 553306 539951 553362 539960
rect 553320 539714 553348 539951
rect 553308 539708 553360 539714
rect 553308 539650 553360 539656
rect 553306 535936 553362 535945
rect 553306 535871 553362 535880
rect 553320 535498 553348 535871
rect 553308 535492 553360 535498
rect 553308 535434 553360 535440
rect 553306 535256 553362 535265
rect 553306 535191 553362 535200
rect 553320 534138 553348 535191
rect 553308 534132 553360 534138
rect 553308 534074 553360 534080
rect 553306 531176 553362 531185
rect 553306 531111 553362 531120
rect 553320 530330 553348 531111
rect 553308 530324 553360 530330
rect 553308 530266 553360 530272
rect 553306 528456 553362 528465
rect 553306 528391 553362 528400
rect 553320 527202 553348 528391
rect 553308 527196 553360 527202
rect 553308 527138 553360 527144
rect 553306 510096 553362 510105
rect 553306 510031 553362 510040
rect 553320 509658 553348 510031
rect 553308 509652 553360 509658
rect 553308 509594 553360 509600
rect 553308 506456 553360 506462
rect 553308 506398 553360 506404
rect 553320 505345 553348 506398
rect 553306 505336 553362 505345
rect 553306 505271 553362 505280
rect 553306 504656 553362 504665
rect 553306 504591 553362 504600
rect 553320 503742 553348 504591
rect 553308 503736 553360 503742
rect 553308 503678 553360 503684
rect 553306 502480 553362 502489
rect 553306 502415 553308 502424
rect 553360 502415 553362 502424
rect 553308 502386 553360 502392
rect 553306 501936 553362 501945
rect 553306 501871 553362 501880
rect 553320 501362 553348 501871
rect 553308 501356 553360 501362
rect 553308 501298 553360 501304
rect 553306 501256 553362 501265
rect 553306 501191 553362 501200
rect 553320 501022 553348 501191
rect 553308 501016 553360 501022
rect 553308 500958 553360 500964
rect 553306 499896 553362 499905
rect 553306 499831 553308 499840
rect 553360 499831 553362 499840
rect 553308 499802 553360 499808
rect 553306 498536 553362 498545
rect 553306 498471 553308 498480
rect 553360 498471 553362 498480
rect 553308 498442 553360 498448
rect 553306 489016 553362 489025
rect 553306 488951 553362 488960
rect 553320 488918 553348 488951
rect 553308 488912 553360 488918
rect 553308 488854 553360 488860
rect 553306 488336 553362 488345
rect 553306 488271 553362 488280
rect 553320 487218 553348 488271
rect 553308 487212 553360 487218
rect 553308 487154 553360 487160
rect 553306 478816 553362 478825
rect 553306 478751 553362 478760
rect 553320 477562 553348 478751
rect 553308 477556 553360 477562
rect 553308 477498 553360 477504
rect 553306 475416 553362 475425
rect 553306 475351 553362 475360
rect 553320 474774 553348 475351
rect 553308 474768 553360 474774
rect 553308 474710 553360 474716
rect 553306 470656 553362 470665
rect 553306 470591 553308 470600
rect 553360 470591 553362 470600
rect 553308 470562 553360 470568
rect 553306 469976 553362 469985
rect 553306 469911 553362 469920
rect 553320 469266 553348 469911
rect 553308 469260 553360 469266
rect 553308 469202 553360 469208
rect 553306 466576 553362 466585
rect 553306 466511 553362 466520
rect 553320 466478 553348 466511
rect 553308 466472 553360 466478
rect 553308 466414 553360 466420
rect 553306 455016 553362 455025
rect 553306 454951 553362 454960
rect 553320 454102 553348 454951
rect 553308 454096 553360 454102
rect 553308 454038 553360 454044
rect 553306 450256 553362 450265
rect 553306 450191 553362 450200
rect 553320 449954 553348 450191
rect 553308 449948 553360 449954
rect 553308 449890 553360 449896
rect 553306 443456 553362 443465
rect 553306 443391 553362 443400
rect 553320 443018 553348 443391
rect 553308 443012 553360 443018
rect 553308 442954 553360 442960
rect 553306 438016 553362 438025
rect 553306 437951 553362 437960
rect 553320 437510 553348 437951
rect 553308 437504 553360 437510
rect 553308 437446 553360 437452
rect 553306 436656 553362 436665
rect 553306 436591 553362 436600
rect 553320 436150 553348 436591
rect 553308 436144 553360 436150
rect 553308 436086 553360 436092
rect 553308 436008 553360 436014
rect 553308 435950 553360 435956
rect 553214 232520 553270 232529
rect 553214 232455 553270 232464
rect 552848 167748 552900 167754
rect 552848 167690 552900 167696
rect 553320 159361 553348 435950
rect 553412 249898 553440 682450
rect 553504 496505 553532 682654
rect 553490 496496 553546 496505
rect 553490 496431 553546 496440
rect 553490 391096 553546 391105
rect 553490 391031 553546 391040
rect 553400 249892 553452 249898
rect 553400 249834 553452 249840
rect 553400 249756 553452 249762
rect 553400 249698 553452 249704
rect 553306 159352 553362 159361
rect 553306 159287 553362 159296
rect 553032 153876 553084 153882
rect 553032 153818 553084 153824
rect 552848 150000 552900 150006
rect 552848 149942 552900 149948
rect 552860 115161 552888 149942
rect 552846 115152 552902 115161
rect 552846 115087 552902 115096
rect 552940 83496 552992 83502
rect 552940 83438 552992 83444
rect 552848 82884 552900 82890
rect 552848 82826 552900 82832
rect 552860 3534 552888 82826
rect 552952 23118 552980 83438
rect 553044 27606 553072 153818
rect 553124 150884 553176 150890
rect 553124 150826 553176 150832
rect 553032 27600 553084 27606
rect 553032 27542 553084 27548
rect 553136 26110 553164 150826
rect 553124 26104 553176 26110
rect 553124 26046 553176 26052
rect 552940 23112 552992 23118
rect 552940 23054 552992 23060
rect 553412 13122 553440 249698
rect 553400 13116 553452 13122
rect 553400 13058 553452 13064
rect 553504 8974 553532 391031
rect 553596 363905 553624 683334
rect 553688 532574 553716 683402
rect 553768 679380 553820 679386
rect 553768 679322 553820 679328
rect 553676 532568 553728 532574
rect 553676 532510 553728 532516
rect 553780 530534 553808 679322
rect 553768 530528 553820 530534
rect 553768 530470 553820 530476
rect 553768 526312 553820 526318
rect 553768 526254 553820 526260
rect 553676 519308 553728 519314
rect 553676 519250 553728 519256
rect 553582 363896 553638 363905
rect 553582 363831 553638 363840
rect 553688 342854 553716 519250
rect 553780 368014 553808 526254
rect 553860 459060 553912 459066
rect 553860 459002 553912 459008
rect 553768 368008 553820 368014
rect 553768 367950 553820 367956
rect 553676 342848 553728 342854
rect 553676 342790 553728 342796
rect 553582 340776 553638 340785
rect 553582 340711 553638 340720
rect 553596 25537 553624 340711
rect 553676 322380 553728 322386
rect 553676 322322 553728 322328
rect 553582 25528 553638 25537
rect 553582 25463 553638 25472
rect 553688 9042 553716 322322
rect 553768 293140 553820 293146
rect 553768 293082 553820 293088
rect 553780 17270 553808 293082
rect 553872 198490 553900 459002
rect 553952 456068 554004 456074
rect 553952 456010 554004 456016
rect 553964 307494 553992 456010
rect 553952 307488 554004 307494
rect 553952 307430 554004 307436
rect 554056 293185 554084 683606
rect 554780 682168 554832 682174
rect 554780 682110 554832 682116
rect 554792 603974 554820 682110
rect 554780 603968 554832 603974
rect 554780 603910 554832 603916
rect 554884 589014 554912 687210
rect 554964 686044 555016 686050
rect 554964 685986 555016 685992
rect 554872 589008 554924 589014
rect 554872 588950 554924 588956
rect 554976 421054 555004 685986
rect 555148 684548 555200 684554
rect 555148 684490 555200 684496
rect 555056 680672 555108 680678
rect 555056 680614 555108 680620
rect 555068 430234 555096 680614
rect 555160 553722 555188 684490
rect 555240 683324 555292 683330
rect 555240 683266 555292 683272
rect 555252 642258 555280 683266
rect 560944 682372 560996 682378
rect 560944 682314 560996 682320
rect 557908 679448 557960 679454
rect 557908 679390 557960 679396
rect 556436 646196 556488 646202
rect 556436 646138 556488 646144
rect 555240 642252 555292 642258
rect 555240 642194 555292 642200
rect 555700 608660 555752 608666
rect 555700 608602 555752 608608
rect 555148 553716 555200 553722
rect 555148 553658 555200 553664
rect 555240 550860 555292 550866
rect 555240 550802 555292 550808
rect 555148 543856 555200 543862
rect 555148 543798 555200 543804
rect 555056 430228 555108 430234
rect 555056 430170 555108 430176
rect 554964 421048 555016 421054
rect 554964 420990 555016 420996
rect 554964 393780 555016 393786
rect 554964 393722 555016 393728
rect 554136 365220 554188 365226
rect 554136 365162 554188 365168
rect 554042 293176 554098 293185
rect 554042 293111 554098 293120
rect 554044 291780 554096 291786
rect 554044 291722 554096 291728
rect 553952 252544 554004 252550
rect 553952 252486 554004 252492
rect 553860 198484 553912 198490
rect 553860 198426 553912 198432
rect 553860 158364 553912 158370
rect 553860 158306 553912 158312
rect 553768 17264 553820 17270
rect 553768 17206 553820 17212
rect 553676 9036 553728 9042
rect 553676 8978 553728 8984
rect 553492 8968 553544 8974
rect 553492 8910 553544 8916
rect 553872 4146 553900 158306
rect 553964 28898 553992 252486
rect 554056 233918 554084 291722
rect 554148 240174 554176 365162
rect 554228 265260 554280 265266
rect 554228 265202 554280 265208
rect 554136 240168 554188 240174
rect 554136 240110 554188 240116
rect 554240 238474 554268 265202
rect 554780 263220 554832 263226
rect 554780 263162 554832 263168
rect 554228 238468 554280 238474
rect 554228 238410 554280 238416
rect 554792 238202 554820 263162
rect 554780 238196 554832 238202
rect 554780 238138 554832 238144
rect 554044 233912 554096 233918
rect 554044 233854 554096 233860
rect 554044 155372 554096 155378
rect 554044 155314 554096 155320
rect 553952 28892 554004 28898
rect 553952 28834 554004 28840
rect 554056 20398 554084 155314
rect 554136 152856 554188 152862
rect 554136 152798 554188 152804
rect 554148 149122 554176 152798
rect 554226 149288 554282 149297
rect 554226 149223 554282 149232
rect 554136 149116 554188 149122
rect 554136 149058 554188 149064
rect 554240 142154 554268 149223
rect 554148 142126 554268 142154
rect 554148 94246 554176 142126
rect 554228 142044 554280 142050
rect 554228 141986 554280 141992
rect 554240 133890 554268 141986
rect 554228 133884 554280 133890
rect 554228 133826 554280 133832
rect 554136 94240 554188 94246
rect 554136 94182 554188 94188
rect 554044 20392 554096 20398
rect 554044 20334 554096 20340
rect 554976 15978 555004 393722
rect 555056 372700 555108 372706
rect 555056 372642 555108 372648
rect 554964 15972 555016 15978
rect 554964 15914 555016 15920
rect 555068 13025 555096 372642
rect 555160 188698 555188 543798
rect 555252 235346 555280 550802
rect 555332 412820 555384 412826
rect 555332 412762 555384 412768
rect 555344 238950 555372 412762
rect 555424 368620 555476 368626
rect 555424 368562 555476 368568
rect 555332 238944 555384 238950
rect 555332 238886 555384 238892
rect 555436 236502 555464 368562
rect 555516 305516 555568 305522
rect 555516 305458 555568 305464
rect 555424 236496 555476 236502
rect 555424 236438 555476 236444
rect 555240 235340 555292 235346
rect 555240 235282 555292 235288
rect 555528 191146 555556 305458
rect 555608 232892 555660 232898
rect 555608 232834 555660 232840
rect 555516 191140 555568 191146
rect 555516 191082 555568 191088
rect 555148 188692 555200 188698
rect 555148 188634 555200 188640
rect 555238 162480 555294 162489
rect 555238 162415 555294 162424
rect 555148 152924 555200 152930
rect 555148 152866 555200 152872
rect 555054 13016 555110 13025
rect 555054 12951 555110 12960
rect 553860 4140 553912 4146
rect 553860 4082 553912 4088
rect 555160 4010 555188 152866
rect 555252 24410 555280 162415
rect 555516 157004 555568 157010
rect 555516 156946 555568 156952
rect 555332 152584 555384 152590
rect 555332 152526 555384 152532
rect 555344 27538 555372 152526
rect 555424 149116 555476 149122
rect 555424 149058 555476 149064
rect 555332 27532 555384 27538
rect 555332 27474 555384 27480
rect 555436 24750 555464 149058
rect 555528 95198 555556 156946
rect 555620 138718 555648 232834
rect 555608 138712 555660 138718
rect 555608 138654 555660 138660
rect 555516 95192 555568 95198
rect 555516 95134 555568 95140
rect 555712 26246 555740 608602
rect 555792 590844 555844 590850
rect 555792 590786 555844 590792
rect 555700 26240 555752 26246
rect 555700 26182 555752 26188
rect 555424 24744 555476 24750
rect 555424 24686 555476 24692
rect 555240 24404 555292 24410
rect 555240 24346 555292 24352
rect 555804 21622 555832 590786
rect 556160 577516 556212 577522
rect 556160 577458 556212 577464
rect 556172 21758 556200 577458
rect 556252 463956 556304 463962
rect 556252 463898 556304 463904
rect 556160 21752 556212 21758
rect 556160 21694 556212 21700
rect 555792 21616 555844 21622
rect 555792 21558 555844 21564
rect 556264 6186 556292 463898
rect 556344 452804 556396 452810
rect 556344 452746 556396 452752
rect 556356 22846 556384 452746
rect 556448 238338 556476 646138
rect 556804 644700 556856 644706
rect 556804 644642 556856 644648
rect 556816 632058 556844 644642
rect 556804 632052 556856 632058
rect 556804 631994 556856 632000
rect 556528 631780 556580 631786
rect 556528 631722 556580 631728
rect 556436 238332 556488 238338
rect 556436 238274 556488 238280
rect 556540 235414 556568 631722
rect 556620 558000 556672 558006
rect 556620 557942 556672 557948
rect 556528 235408 556580 235414
rect 556528 235350 556580 235356
rect 556632 195294 556660 557942
rect 557724 502444 557776 502450
rect 557724 502386 557776 502392
rect 557632 499860 557684 499866
rect 557632 499802 557684 499808
rect 557540 498500 557592 498506
rect 557540 498442 557592 498448
rect 556896 437436 556948 437442
rect 556896 437378 556948 437384
rect 556712 343052 556764 343058
rect 556712 342994 556764 343000
rect 556620 195288 556672 195294
rect 556620 195230 556672 195236
rect 556436 158228 556488 158234
rect 556436 158170 556488 158176
rect 556344 22840 556396 22846
rect 556344 22782 556396 22788
rect 556252 6180 556304 6186
rect 556252 6122 556304 6128
rect 555148 4004 555200 4010
rect 555148 3946 555200 3952
rect 552848 3528 552900 3534
rect 552848 3470 552900 3476
rect 556448 3398 556476 158170
rect 556528 155780 556580 155786
rect 556528 155722 556580 155728
rect 556540 26217 556568 155722
rect 556620 150680 556672 150686
rect 556620 150622 556672 150628
rect 556632 82890 556660 150622
rect 556620 82884 556672 82890
rect 556620 82826 556672 82832
rect 556526 26208 556582 26217
rect 556526 26143 556582 26152
rect 556724 19990 556752 342994
rect 556804 276140 556856 276146
rect 556804 276082 556856 276088
rect 556816 26926 556844 276082
rect 556908 238542 556936 437378
rect 557080 278860 557132 278866
rect 557080 278802 557132 278808
rect 556896 238536 556948 238542
rect 556896 238478 556948 238484
rect 556894 235376 556950 235385
rect 556894 235311 556950 235320
rect 556908 126274 556936 235311
rect 556988 232824 557040 232830
rect 556988 232766 557040 232772
rect 557000 134473 557028 232766
rect 557092 197810 557120 278802
rect 557080 197804 557132 197810
rect 557080 197746 557132 197752
rect 556986 134464 557042 134473
rect 556986 134399 557042 134408
rect 556988 133884 557040 133890
rect 556988 133826 557040 133832
rect 556896 126268 556948 126274
rect 556896 126210 556948 126216
rect 556894 112432 556950 112441
rect 556894 112367 556950 112376
rect 556908 73234 556936 112367
rect 557000 111110 557028 133826
rect 557078 126304 557134 126313
rect 557078 126239 557134 126248
rect 557092 113218 557120 126239
rect 557080 113212 557132 113218
rect 557080 113154 557132 113160
rect 556988 111104 557040 111110
rect 556988 111046 557040 111052
rect 556896 73228 556948 73234
rect 556896 73170 556948 73176
rect 556804 26920 556856 26926
rect 556804 26862 556856 26868
rect 556712 19984 556764 19990
rect 556712 19926 556764 19932
rect 557552 4894 557580 498442
rect 557644 13161 557672 499802
rect 557736 20194 557764 502386
rect 557816 403708 557868 403714
rect 557816 403650 557868 403656
rect 557828 21690 557856 403650
rect 557920 378350 557948 679390
rect 560392 652792 560444 652798
rect 560392 652734 560444 652740
rect 559288 567316 559340 567322
rect 559288 567258 559340 567264
rect 558000 530324 558052 530330
rect 558000 530266 558052 530272
rect 557908 378344 557960 378350
rect 557908 378286 557960 378292
rect 557908 360460 557960 360466
rect 557908 360402 557960 360408
rect 557816 21684 557868 21690
rect 557816 21626 557868 21632
rect 557724 20188 557776 20194
rect 557724 20130 557776 20136
rect 557630 13152 557686 13161
rect 557630 13087 557686 13096
rect 557920 10334 557948 360402
rect 558012 235210 558040 530266
rect 559196 501356 559248 501362
rect 559196 501298 559248 501304
rect 559104 488912 559156 488918
rect 559104 488854 559156 488860
rect 558092 381540 558144 381546
rect 558092 381482 558144 381488
rect 558000 235204 558052 235210
rect 558000 235146 558052 235152
rect 558104 190194 558132 381482
rect 558184 350940 558236 350946
rect 558184 350882 558236 350888
rect 558196 238678 558224 350882
rect 558184 238672 558236 238678
rect 558184 238614 558236 238620
rect 558184 232756 558236 232762
rect 558184 232698 558236 232704
rect 558092 190188 558144 190194
rect 558092 190130 558144 190136
rect 558000 154420 558052 154426
rect 558000 154362 558052 154368
rect 557908 10328 557960 10334
rect 557908 10270 557960 10276
rect 558012 6458 558040 154362
rect 558092 153060 558144 153066
rect 558092 153002 558144 153008
rect 558104 20534 558132 153002
rect 558196 137766 558224 232698
rect 558276 159316 558328 159322
rect 558276 159258 558328 159264
rect 558184 137760 558236 137766
rect 558184 137702 558236 137708
rect 558184 135924 558236 135930
rect 558184 135866 558236 135872
rect 558196 111926 558224 135866
rect 558288 115938 558316 159258
rect 559012 148436 559064 148442
rect 559012 148378 559064 148384
rect 559024 137358 559052 148378
rect 558368 137352 558420 137358
rect 558368 137294 558420 137300
rect 559012 137352 559064 137358
rect 559012 137294 559064 137300
rect 558276 115932 558328 115938
rect 558276 115874 558328 115880
rect 558276 113212 558328 113218
rect 558276 113154 558328 113160
rect 558184 111920 558236 111926
rect 558184 111862 558236 111868
rect 558288 89049 558316 113154
rect 558380 104242 558408 137294
rect 558368 104236 558420 104242
rect 558368 104178 558420 104184
rect 558274 89040 558330 89049
rect 558274 88975 558330 88984
rect 559116 22914 559144 488854
rect 559208 158098 559236 501298
rect 559300 234530 559328 567258
rect 559748 556572 559800 556578
rect 559748 556514 559800 556520
rect 559564 420164 559616 420170
rect 559564 420106 559616 420112
rect 559472 416084 559524 416090
rect 559472 416026 559524 416032
rect 559380 317620 559432 317626
rect 559380 317562 559432 317568
rect 559288 234524 559340 234530
rect 559288 234466 559340 234472
rect 559196 158092 559248 158098
rect 559196 158034 559248 158040
rect 559196 156460 559248 156466
rect 559196 156402 559248 156408
rect 559104 22908 559156 22914
rect 559104 22850 559156 22856
rect 558092 20528 558144 20534
rect 558092 20470 558144 20476
rect 559208 6914 559236 156402
rect 559288 151292 559340 151298
rect 559288 151234 559340 151240
rect 559300 16574 559328 151234
rect 559392 28257 559420 317562
rect 559484 195838 559512 416026
rect 559576 235278 559604 420106
rect 559564 235272 559616 235278
rect 559564 235214 559616 235220
rect 559472 195832 559524 195838
rect 559472 195774 559524 195780
rect 559564 160064 559616 160070
rect 559564 160006 559616 160012
rect 559472 159384 559524 159390
rect 559472 159326 559524 159332
rect 559484 139398 559512 159326
rect 559472 139392 559524 139398
rect 559472 139334 559524 139340
rect 559472 137760 559524 137766
rect 559472 137702 559524 137708
rect 559378 28248 559434 28257
rect 559378 28183 559434 28192
rect 559300 16546 559420 16574
rect 559208 6886 559328 6914
rect 558000 6452 558052 6458
rect 558000 6394 558052 6400
rect 557540 4888 557592 4894
rect 557540 4830 557592 4836
rect 556436 3392 556488 3398
rect 556436 3334 556488 3340
rect 552756 3052 552808 3058
rect 552756 2994 552808 3000
rect 556160 3052 556212 3058
rect 556160 2994 556212 3000
rect 556172 480 556200 2994
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 6886
rect 559392 6390 559420 16546
rect 559484 16114 559512 137702
rect 559576 114442 559604 160006
rect 559656 153196 559708 153202
rect 559656 153138 559708 153144
rect 559564 114436 559616 114442
rect 559564 114378 559616 114384
rect 559564 99408 559616 99414
rect 559564 99350 559616 99356
rect 559472 16108 559524 16114
rect 559472 16050 559524 16056
rect 559576 13666 559604 99350
rect 559668 77246 559696 153138
rect 559656 77240 559708 77246
rect 559656 77182 559708 77188
rect 559564 13660 559616 13666
rect 559564 13602 559616 13608
rect 559760 12986 559788 556514
rect 559840 509652 559892 509658
rect 559840 509594 559892 509600
rect 559748 12980 559800 12986
rect 559748 12922 559800 12928
rect 559852 7614 559880 509594
rect 560300 258188 560352 258194
rect 560300 258130 560352 258136
rect 560312 240786 560340 258130
rect 560300 240780 560352 240786
rect 560300 240722 560352 240728
rect 560404 239873 560432 652734
rect 560576 575544 560628 575550
rect 560576 575486 560628 575492
rect 560484 567248 560536 567254
rect 560484 567190 560536 567196
rect 560390 239864 560446 239873
rect 560390 239799 560446 239808
rect 560392 237924 560444 237930
rect 560392 237866 560444 237872
rect 560300 237788 560352 237794
rect 560300 237730 560352 237736
rect 560312 236842 560340 237730
rect 560300 236836 560352 236842
rect 560300 236778 560352 236784
rect 560300 149796 560352 149802
rect 560300 149738 560352 149744
rect 560312 137306 560340 149738
rect 560220 137278 560340 137306
rect 560220 100774 560248 137278
rect 560208 100768 560260 100774
rect 560208 100710 560260 100716
rect 560404 26858 560432 237866
rect 560496 178974 560524 567190
rect 560588 195974 560616 575486
rect 560760 535492 560812 535498
rect 560760 535434 560812 535440
rect 560668 369912 560720 369918
rect 560668 369854 560720 369860
rect 560576 195968 560628 195974
rect 560576 195910 560628 195916
rect 560484 178968 560536 178974
rect 560484 178910 560536 178916
rect 560484 156732 560536 156738
rect 560484 156674 560536 156680
rect 560496 44130 560524 156674
rect 560576 155576 560628 155582
rect 560576 155518 560628 155524
rect 560588 62014 560616 155518
rect 560576 62008 560628 62014
rect 560576 61950 560628 61956
rect 560484 44124 560536 44130
rect 560484 44066 560536 44072
rect 560680 27062 560708 369854
rect 560772 198801 560800 535434
rect 560852 459604 560904 459610
rect 560852 459546 560904 459552
rect 560758 198792 560814 198801
rect 560758 198727 560814 198736
rect 560864 196858 560892 459546
rect 560956 237454 560984 682314
rect 564622 682136 564678 682145
rect 564622 682071 564678 682080
rect 563980 669384 564032 669390
rect 563980 669326 564032 669332
rect 563336 656940 563388 656946
rect 563336 656882 563388 656888
rect 561864 648644 561916 648650
rect 561864 648586 561916 648592
rect 561128 474836 561180 474842
rect 561128 474778 561180 474784
rect 561036 386436 561088 386442
rect 561036 386378 561088 386384
rect 560944 237448 560996 237454
rect 560944 237390 560996 237396
rect 560944 236836 560996 236842
rect 560944 236778 560996 236784
rect 560852 196852 560904 196858
rect 560852 196794 560904 196800
rect 560852 165096 560904 165102
rect 560852 165038 560904 165044
rect 560760 155712 560812 155718
rect 560760 155654 560812 155660
rect 560772 62082 560800 155654
rect 560864 121446 560892 165038
rect 560852 121440 560904 121446
rect 560852 121382 560904 121388
rect 560852 100768 560904 100774
rect 560852 100710 560904 100716
rect 560760 62076 560812 62082
rect 560760 62018 560812 62024
rect 560668 27056 560720 27062
rect 560668 26998 560720 27004
rect 560392 26852 560444 26858
rect 560392 26794 560444 26800
rect 560298 20904 560354 20913
rect 560298 20839 560354 20848
rect 560312 20806 560340 20839
rect 560300 20800 560352 20806
rect 560300 20742 560352 20748
rect 560864 13326 560892 100710
rect 560956 29170 560984 236778
rect 561048 198966 561076 386378
rect 561036 198960 561088 198966
rect 561036 198902 561088 198908
rect 561036 159996 561088 160002
rect 561036 159938 561088 159944
rect 561048 78606 561076 159938
rect 561036 78600 561088 78606
rect 561036 78542 561088 78548
rect 560944 29164 560996 29170
rect 560944 29106 560996 29112
rect 561140 28830 561168 474778
rect 561680 251252 561732 251258
rect 561680 251194 561732 251200
rect 561692 248414 561720 251194
rect 561692 248386 561812 248414
rect 561680 247104 561732 247110
rect 561680 247046 561732 247052
rect 561692 239630 561720 247046
rect 561680 239624 561732 239630
rect 561680 239566 561732 239572
rect 561784 239329 561812 248386
rect 561770 239320 561826 239329
rect 561770 239255 561826 239264
rect 561772 237448 561824 237454
rect 561772 237390 561824 237396
rect 561680 111104 561732 111110
rect 561680 111046 561732 111052
rect 561692 99414 561720 111046
rect 561680 99408 561732 99414
rect 561680 99350 561732 99356
rect 561128 28824 561180 28830
rect 561128 28766 561180 28772
rect 561784 24614 561812 237390
rect 561876 147626 561904 648586
rect 562508 623824 562560 623830
rect 562508 623766 562560 623772
rect 562048 607232 562100 607238
rect 562048 607174 562100 607180
rect 561956 474768 562008 474774
rect 561956 474710 562008 474716
rect 561864 147620 561916 147626
rect 561864 147562 561916 147568
rect 561968 29306 561996 474710
rect 562060 190097 562088 607174
rect 562232 539708 562284 539714
rect 562232 539650 562284 539656
rect 562140 385076 562192 385082
rect 562140 385018 562192 385024
rect 562046 190088 562102 190097
rect 562046 190023 562102 190032
rect 562048 159588 562100 159594
rect 562048 159530 562100 159536
rect 562060 37262 562088 159530
rect 562048 37256 562100 37262
rect 562048 37198 562100 37204
rect 561956 29300 562008 29306
rect 561956 29242 562008 29248
rect 562152 26994 562180 385018
rect 562244 233850 562272 539650
rect 562416 477556 562468 477562
rect 562416 477498 562468 477504
rect 562428 437646 562456 477498
rect 562416 437640 562468 437646
rect 562416 437582 562468 437588
rect 562324 437504 562376 437510
rect 562324 437446 562376 437452
rect 562232 233844 562284 233850
rect 562232 233786 562284 233792
rect 562336 174758 562364 437446
rect 562324 174752 562376 174758
rect 562324 174694 562376 174700
rect 562324 162852 562376 162858
rect 562324 162794 562376 162800
rect 562232 150952 562284 150958
rect 562232 150894 562284 150900
rect 562140 26988 562192 26994
rect 562140 26930 562192 26936
rect 561772 24608 561824 24614
rect 561772 24550 561824 24556
rect 562244 19786 562272 150894
rect 562336 125594 562364 162794
rect 562416 155644 562468 155650
rect 562416 155586 562468 155592
rect 562324 125588 562376 125594
rect 562324 125530 562376 125536
rect 562324 124160 562376 124166
rect 562324 124102 562376 124108
rect 562232 19780 562284 19786
rect 562232 19722 562284 19728
rect 562336 16182 562364 124102
rect 562428 107642 562456 155586
rect 562416 107636 562468 107642
rect 562416 107578 562468 107584
rect 562520 72486 562548 623766
rect 563152 603152 563204 603158
rect 563152 603094 563204 603100
rect 562600 550656 562652 550662
rect 562600 550598 562652 550604
rect 562508 72480 562560 72486
rect 562508 72422 562560 72428
rect 562612 28393 562640 550598
rect 563060 155848 563112 155854
rect 563060 155790 563112 155796
rect 563072 128314 563100 155790
rect 563060 128308 563112 128314
rect 563060 128250 563112 128256
rect 563164 45490 563192 603094
rect 563244 437640 563296 437646
rect 563244 437582 563296 437588
rect 563152 45484 563204 45490
rect 563152 45426 563204 45432
rect 562598 28384 562654 28393
rect 562598 28319 562654 28328
rect 562324 16176 562376 16182
rect 562324 16118 562376 16124
rect 560852 13320 560904 13326
rect 560852 13262 560904 13268
rect 559840 7608 559892 7614
rect 559840 7550 559892 7556
rect 559380 6384 559432 6390
rect 559380 6326 559432 6332
rect 563256 480 563284 437582
rect 563348 143546 563376 656882
rect 563428 637696 563480 637702
rect 563428 637638 563480 637644
rect 563440 196654 563468 637638
rect 563612 578264 563664 578270
rect 563612 578206 563664 578212
rect 563520 574116 563572 574122
rect 563520 574058 563572 574064
rect 563428 196648 563480 196654
rect 563428 196590 563480 196596
rect 563532 171834 563560 574058
rect 563624 194041 563652 578206
rect 563704 564460 563756 564466
rect 563704 564402 563756 564408
rect 563610 194032 563666 194041
rect 563610 193967 563666 193976
rect 563716 189689 563744 564402
rect 563796 492720 563848 492726
rect 563796 492662 563848 492668
rect 563702 189680 563758 189689
rect 563702 189615 563758 189624
rect 563520 171828 563572 171834
rect 563520 171770 563572 171776
rect 563428 165232 563480 165238
rect 563428 165174 563480 165180
rect 563336 143540 563388 143546
rect 563336 143482 563388 143488
rect 563440 3330 563468 165174
rect 563808 163538 563836 492662
rect 563888 427848 563940 427854
rect 563888 427790 563940 427796
rect 563900 198014 563928 427790
rect 563888 198008 563940 198014
rect 563888 197950 563940 197956
rect 563796 163532 563848 163538
rect 563796 163474 563848 163480
rect 563610 156632 563666 156641
rect 563610 156567 563666 156576
rect 563520 151768 563572 151774
rect 563520 151710 563572 151716
rect 563532 6322 563560 151710
rect 563624 22982 563652 156567
rect 563888 152788 563940 152794
rect 563888 152730 563940 152736
rect 563794 150240 563850 150249
rect 563794 150175 563850 150184
rect 563704 140820 563756 140826
rect 563704 140762 563756 140768
rect 563612 22976 563664 22982
rect 563612 22918 563664 22924
rect 563716 20058 563744 140762
rect 563808 139534 563836 150175
rect 563796 139528 563848 139534
rect 563796 139470 563848 139476
rect 563796 138712 563848 138718
rect 563796 138654 563848 138660
rect 563808 104174 563836 138654
rect 563796 104168 563848 104174
rect 563796 104110 563848 104116
rect 563796 102196 563848 102202
rect 563796 102138 563848 102144
rect 563704 20052 563756 20058
rect 563704 19994 563756 20000
rect 563808 13802 563836 102138
rect 563900 41410 563928 152730
rect 563992 78674 564020 669326
rect 564532 637628 564584 637634
rect 564532 637570 564584 637576
rect 564440 263628 564492 263634
rect 564440 263570 564492 263576
rect 564452 239902 564480 263570
rect 564440 239896 564492 239902
rect 564440 239838 564492 239844
rect 563980 78668 564032 78674
rect 563980 78610 564032 78616
rect 563888 41404 563940 41410
rect 563888 41346 563940 41352
rect 564544 29481 564572 637570
rect 564636 197441 564664 682071
rect 565452 644496 565504 644502
rect 565452 644438 565504 644444
rect 564716 519036 564768 519042
rect 564716 518978 564768 518984
rect 564622 197432 564678 197441
rect 564622 197367 564678 197376
rect 564624 157276 564676 157282
rect 564624 157218 564676 157224
rect 564530 29472 564586 29481
rect 564530 29407 564586 29416
rect 564636 23322 564664 157218
rect 564728 136542 564756 518978
rect 564808 514820 564860 514826
rect 564808 514762 564860 514768
rect 564820 238746 564848 514762
rect 564992 288516 565044 288522
rect 564992 288458 565044 288464
rect 564900 245744 564952 245750
rect 564900 245686 564952 245692
rect 564808 238740 564860 238746
rect 564808 238682 564860 238688
rect 564808 232416 564860 232422
rect 564808 232358 564860 232364
rect 564716 136536 564768 136542
rect 564716 136478 564768 136484
rect 564714 124128 564770 124137
rect 564714 124063 564770 124072
rect 564624 23316 564676 23322
rect 564624 23258 564676 23264
rect 564728 15162 564756 124063
rect 564716 15156 564768 15162
rect 564716 15098 564768 15104
rect 564820 14482 564848 232358
rect 564912 24274 564940 245686
rect 565004 240553 565032 288458
rect 565084 274712 565136 274718
rect 565084 274654 565136 274660
rect 564990 240544 565046 240553
rect 564990 240479 565046 240488
rect 565096 239601 565124 274654
rect 565082 239592 565138 239601
rect 565082 239527 565138 239536
rect 564992 235612 565044 235618
rect 564992 235554 565044 235560
rect 564900 24268 564952 24274
rect 564900 24210 564952 24216
rect 565004 18426 565032 235554
rect 565176 235476 565228 235482
rect 565176 235418 565228 235424
rect 565084 154216 565136 154222
rect 565084 154158 565136 154164
rect 565096 23050 565124 154158
rect 565188 140826 565216 235418
rect 565360 149864 565412 149870
rect 565360 149806 565412 149812
rect 565176 140820 565228 140826
rect 565176 140762 565228 140768
rect 565176 139528 565228 139534
rect 565176 139470 565228 139476
rect 565268 139528 565320 139534
rect 565268 139470 565320 139476
rect 565188 83502 565216 139470
rect 565280 124166 565308 139470
rect 565372 139466 565400 149806
rect 565360 139460 565412 139466
rect 565360 139402 565412 139408
rect 565268 124160 565320 124166
rect 565268 124102 565320 124108
rect 565176 83496 565228 83502
rect 565176 83438 565228 83444
rect 565464 29073 565492 644438
rect 565912 454096 565964 454102
rect 565912 454038 565964 454044
rect 565820 256760 565872 256766
rect 565820 256702 565872 256708
rect 565832 239737 565860 256702
rect 565818 239728 565874 239737
rect 565818 239663 565874 239672
rect 565820 139460 565872 139466
rect 565820 139402 565872 139408
rect 565832 119406 565860 139402
rect 565820 119400 565872 119406
rect 565820 119342 565872 119348
rect 565820 111920 565872 111926
rect 565820 111862 565872 111868
rect 565832 102202 565860 111862
rect 565820 102196 565872 102202
rect 565820 102138 565872 102144
rect 565924 29374 565952 454038
rect 566016 282878 566044 700402
rect 566188 700324 566240 700330
rect 566188 700266 566240 700272
rect 566096 682440 566148 682446
rect 566096 682382 566148 682388
rect 566108 313274 566136 682382
rect 566200 335306 566228 700266
rect 579158 697232 579214 697241
rect 579158 697167 579214 697176
rect 576860 684616 576912 684622
rect 576860 684558 576912 684564
rect 567936 683596 567988 683602
rect 567936 683538 567988 683544
rect 566740 560380 566792 560386
rect 566740 560322 566792 560328
rect 566280 527196 566332 527202
rect 566280 527138 566332 527144
rect 566188 335300 566240 335306
rect 566188 335242 566240 335248
rect 566188 317552 566240 317558
rect 566188 317494 566240 317500
rect 566096 313268 566148 313274
rect 566096 313210 566148 313216
rect 566096 289876 566148 289882
rect 566096 289818 566148 289824
rect 566004 282872 566056 282878
rect 566004 282814 566056 282820
rect 566004 217320 566056 217326
rect 566004 217262 566056 217268
rect 565912 29368 565964 29374
rect 565912 29310 565964 29316
rect 565450 29064 565506 29073
rect 565450 28999 565506 29008
rect 565084 23044 565136 23050
rect 565084 22986 565136 22992
rect 564992 18420 565044 18426
rect 564992 18362 565044 18368
rect 564808 14476 564860 14482
rect 564808 14418 564860 14424
rect 563796 13796 563848 13802
rect 563796 13738 563848 13744
rect 563520 6316 563572 6322
rect 563520 6258 563572 6264
rect 565820 4004 565872 4010
rect 565820 3946 565872 3952
rect 565832 3466 565860 3946
rect 566016 3482 566044 217262
rect 566108 4010 566136 289818
rect 566200 283626 566228 317494
rect 566188 283620 566240 283626
rect 566188 283562 566240 283568
rect 566200 282946 566228 283562
rect 566188 282940 566240 282946
rect 566188 282882 566240 282888
rect 566292 280158 566320 527138
rect 566372 445800 566424 445806
rect 566372 445742 566424 445748
rect 566280 280152 566332 280158
rect 566280 280094 566332 280100
rect 566188 254040 566240 254046
rect 566188 253982 566240 253988
rect 566200 24138 566228 253982
rect 566384 240106 566412 445742
rect 566464 335368 566516 335374
rect 566464 335310 566516 335316
rect 566372 240100 566424 240106
rect 566372 240042 566424 240048
rect 566280 232348 566332 232354
rect 566280 232290 566332 232296
rect 566188 24132 566240 24138
rect 566188 24074 566240 24080
rect 566292 16522 566320 232290
rect 566476 193118 566504 335310
rect 566556 300960 566608 300966
rect 566556 300902 566608 300908
rect 566464 193112 566516 193118
rect 566464 193054 566516 193060
rect 566568 184249 566596 300902
rect 566648 282940 566700 282946
rect 566648 282882 566700 282888
rect 566660 239766 566688 282882
rect 566648 239760 566700 239766
rect 566648 239702 566700 239708
rect 566648 232620 566700 232626
rect 566648 232562 566700 232568
rect 566554 184240 566610 184249
rect 566554 184175 566610 184184
rect 566370 165064 566426 165073
rect 566370 164999 566426 165008
rect 566280 16516 566332 16522
rect 566280 16458 566332 16464
rect 566384 4078 566412 164999
rect 566464 155508 566516 155514
rect 566464 155450 566516 155456
rect 566476 6866 566504 155450
rect 566556 152720 566608 152726
rect 566556 152662 566608 152668
rect 566568 17814 566596 152662
rect 566660 139534 566688 232562
rect 566648 139528 566700 139534
rect 566648 139470 566700 139476
rect 566752 71058 566780 560322
rect 567292 539640 567344 539646
rect 567292 539582 567344 539588
rect 566832 280288 566884 280294
rect 566832 280230 566884 280236
rect 566844 193905 566872 280230
rect 567200 247716 567252 247722
rect 567200 247658 567252 247664
rect 567212 237114 567240 247658
rect 567200 237108 567252 237114
rect 567200 237050 567252 237056
rect 567304 236774 567332 539582
rect 567844 470620 567896 470626
rect 567844 470562 567896 470568
rect 567476 466472 567528 466478
rect 567476 466414 567528 466420
rect 567384 277432 567436 277438
rect 567384 277374 567436 277380
rect 567292 236768 567344 236774
rect 567292 236710 567344 236716
rect 566830 193896 566886 193905
rect 566830 193831 566886 193840
rect 567292 162716 567344 162722
rect 567292 162658 567344 162664
rect 566740 71052 566792 71058
rect 566740 70994 566792 71000
rect 566556 17808 566608 17814
rect 566556 17750 566608 17756
rect 566464 6860 566516 6866
rect 566464 6802 566516 6808
rect 567304 6662 567332 162658
rect 567396 18902 567424 277374
rect 567488 239834 567516 466414
rect 567568 365832 567620 365838
rect 567568 365774 567620 365780
rect 567476 239828 567528 239834
rect 567476 239770 567528 239776
rect 567580 194478 567608 365774
rect 567568 194472 567620 194478
rect 567568 194414 567620 194420
rect 567660 157140 567712 157146
rect 567660 157082 567712 157088
rect 567476 156868 567528 156874
rect 567476 156810 567528 156816
rect 567488 20602 567516 156810
rect 567568 148368 567620 148374
rect 567568 148310 567620 148316
rect 567476 20596 567528 20602
rect 567476 20538 567528 20544
rect 567384 18896 567436 18902
rect 567384 18838 567436 18844
rect 567580 15026 567608 148310
rect 567672 26042 567700 157082
rect 567752 151564 567804 151570
rect 567752 151506 567804 151512
rect 567764 31142 567792 151506
rect 567752 31136 567804 31142
rect 567752 31078 567804 31084
rect 567660 26036 567712 26042
rect 567660 25978 567712 25984
rect 567568 15020 567620 15026
rect 567568 14962 567620 14968
rect 567856 7614 567884 470562
rect 567948 139398 567976 683538
rect 571340 683256 571392 683262
rect 571340 683198 571392 683204
rect 570144 682032 570196 682038
rect 570144 681974 570196 681980
rect 568764 681964 568816 681970
rect 568764 681906 568816 681912
rect 568028 560312 568080 560318
rect 568028 560254 568080 560260
rect 568040 173874 568068 560254
rect 568672 557592 568724 557598
rect 568672 557534 568724 557540
rect 568120 354748 568172 354754
rect 568120 354690 568172 354696
rect 568028 173868 568080 173874
rect 568028 173810 568080 173816
rect 568028 153672 568080 153678
rect 568028 153614 568080 153620
rect 567936 139392 567988 139398
rect 567936 139334 567988 139340
rect 568040 117298 568068 153614
rect 568028 117292 568080 117298
rect 568028 117234 568080 117240
rect 568132 25362 568160 354690
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 568592 239970 568620 260850
rect 568580 239964 568632 239970
rect 568580 239906 568632 239912
rect 568580 162172 568632 162178
rect 568580 162114 568632 162120
rect 568592 135250 568620 162114
rect 568580 135244 568632 135250
rect 568580 135186 568632 135192
rect 568120 25356 568172 25362
rect 568120 25298 568172 25304
rect 568684 24206 568712 557534
rect 568776 239562 568804 681906
rect 569406 681864 569462 681873
rect 569406 681799 569462 681808
rect 569132 443012 569184 443018
rect 569132 442954 569184 442960
rect 569040 259548 569092 259554
rect 569040 259490 569092 259496
rect 568948 258120 569000 258126
rect 568948 258062 569000 258068
rect 568764 239556 568816 239562
rect 568764 239498 568816 239504
rect 568764 235680 568816 235686
rect 568764 235622 568816 235628
rect 568672 24200 568724 24206
rect 568672 24142 568724 24148
rect 568776 14550 568804 235622
rect 568856 156664 568908 156670
rect 568856 156606 568908 156612
rect 568868 31074 568896 156606
rect 568856 31068 568908 31074
rect 568856 31010 568908 31016
rect 568960 21554 568988 258062
rect 569052 25498 569080 259490
rect 569144 241194 569172 442954
rect 569224 338156 569276 338162
rect 569224 338098 569276 338104
rect 569132 241188 569184 241194
rect 569132 241130 569184 241136
rect 569236 237046 569264 338098
rect 569316 239420 569368 239426
rect 569316 239362 569368 239368
rect 569224 237040 569276 237046
rect 569224 236982 569276 236988
rect 569132 232484 569184 232490
rect 569132 232426 569184 232432
rect 569040 25492 569092 25498
rect 569040 25434 569092 25440
rect 568948 21548 569000 21554
rect 568948 21490 569000 21496
rect 569144 19106 569172 232426
rect 569328 191214 569356 239362
rect 569316 191208 569368 191214
rect 569316 191150 569368 191156
rect 569224 154080 569276 154086
rect 569224 154022 569276 154028
rect 569236 53786 569264 154022
rect 569224 53780 569276 53786
rect 569224 53722 569276 53728
rect 569132 19100 569184 19106
rect 569132 19042 569184 19048
rect 569420 18834 569448 681799
rect 570052 681080 570104 681086
rect 570052 681022 570104 681028
rect 569960 611380 570012 611386
rect 569960 611322 570012 611328
rect 569500 425128 569552 425134
rect 569500 425070 569552 425076
rect 569512 150385 569540 425070
rect 569498 150376 569554 150385
rect 569498 150311 569554 150320
rect 569972 28150 570000 611322
rect 570064 97986 570092 681022
rect 570156 100026 570184 681974
rect 570696 610020 570748 610026
rect 570696 609962 570748 609968
rect 570604 600976 570656 600982
rect 570604 600918 570656 600924
rect 570616 506462 570644 600918
rect 570708 525774 570736 609962
rect 570696 525768 570748 525774
rect 570696 525710 570748 525716
rect 570788 516180 570840 516186
rect 570788 516122 570840 516128
rect 570604 506456 570656 506462
rect 570604 506398 570656 506404
rect 570696 470620 570748 470626
rect 570696 470562 570748 470568
rect 570604 423768 570656 423774
rect 570604 423710 570656 423716
rect 570236 409896 570288 409902
rect 570236 409838 570288 409844
rect 570144 100020 570196 100026
rect 570144 99962 570196 99968
rect 570052 97980 570104 97986
rect 570052 97922 570104 97928
rect 569960 28144 570012 28150
rect 569960 28086 570012 28092
rect 569958 20904 570014 20913
rect 569958 20839 569960 20848
rect 570012 20839 570014 20848
rect 569960 20810 570012 20816
rect 569408 18828 569460 18834
rect 569408 18770 569460 18776
rect 568764 14544 568816 14550
rect 568764 14486 568816 14492
rect 567844 7608 567896 7614
rect 567844 7550 567896 7556
rect 567292 6656 567344 6662
rect 567292 6598 567344 6604
rect 566372 4072 566424 4078
rect 566372 4014 566424 4020
rect 566096 4004 566148 4010
rect 566096 3946 566148 3952
rect 570248 3505 570276 409838
rect 570420 389224 570472 389230
rect 570420 389166 570472 389172
rect 570328 287088 570380 287094
rect 570328 287030 570380 287036
rect 570340 18766 570368 287030
rect 570432 193186 570460 389166
rect 570512 327208 570564 327214
rect 570512 327150 570564 327156
rect 570524 238610 570552 327150
rect 570512 238604 570564 238610
rect 570512 238546 570564 238552
rect 570512 235748 570564 235754
rect 570512 235690 570564 235696
rect 570420 193180 570472 193186
rect 570420 193122 570472 193128
rect 570420 173868 570472 173874
rect 570420 173810 570472 173816
rect 570328 18760 570380 18766
rect 570328 18702 570380 18708
rect 570432 6914 570460 173810
rect 570524 14754 570552 235690
rect 570616 33114 570644 423710
rect 570708 238882 570736 470562
rect 570800 420238 570828 516122
rect 570788 420232 570840 420238
rect 570788 420174 570840 420180
rect 570788 252612 570840 252618
rect 570788 252554 570840 252560
rect 570696 238876 570748 238882
rect 570696 238818 570748 238824
rect 570800 198558 570828 252554
rect 570788 198552 570840 198558
rect 570788 198494 570840 198500
rect 570696 157072 570748 157078
rect 570696 157014 570748 157020
rect 570604 33108 570656 33114
rect 570604 33050 570656 33056
rect 570708 19242 570736 157014
rect 570696 19236 570748 19242
rect 570696 19178 570748 19184
rect 570512 14748 570564 14754
rect 570512 14690 570564 14696
rect 570340 6886 570460 6914
rect 570234 3496 570290 3505
rect 565820 3460 565872 3466
rect 566016 3454 566872 3482
rect 565820 3402 565872 3408
rect 563428 3324 563480 3330
rect 563428 3266 563480 3272
rect 566844 480 566872 3454
rect 570234 3431 570290 3440
rect 570340 480 570368 6886
rect 571352 4049 571380 683198
rect 574100 682304 574152 682310
rect 574100 682246 574152 682252
rect 571616 681828 571668 681834
rect 571616 681770 571668 681776
rect 571432 629332 571484 629338
rect 571432 629274 571484 629280
rect 571444 20890 571472 629274
rect 571524 520328 571576 520334
rect 571524 520270 571576 520276
rect 571536 25430 571564 520270
rect 571628 239465 571656 681770
rect 571984 681760 572036 681766
rect 571984 681702 572036 681708
rect 571708 672104 571760 672110
rect 571708 672046 571760 672052
rect 571720 241126 571748 672046
rect 571800 314696 571852 314702
rect 571800 314638 571852 314644
rect 571708 241120 571760 241126
rect 571708 241062 571760 241068
rect 571614 239456 571670 239465
rect 571812 239426 571840 314638
rect 571892 280220 571944 280226
rect 571892 280162 571944 280168
rect 571614 239391 571670 239400
rect 571800 239420 571852 239426
rect 571800 239362 571852 239368
rect 571616 234592 571668 234598
rect 571616 234534 571668 234540
rect 571524 25424 571576 25430
rect 571524 25366 571576 25372
rect 571444 20862 571564 20890
rect 571430 20768 571486 20777
rect 571430 20703 571432 20712
rect 571484 20703 571486 20712
rect 571432 20674 571484 20680
rect 571536 18698 571564 20862
rect 571524 18692 571576 18698
rect 571524 18634 571576 18640
rect 571338 4040 571394 4049
rect 571338 3975 571394 3984
rect 571628 3670 571656 234534
rect 571904 196994 571932 280162
rect 571892 196988 571944 196994
rect 571892 196930 571944 196936
rect 571996 193186 572024 681702
rect 572812 677680 572864 677686
rect 572812 677622 572864 677628
rect 572076 378208 572128 378214
rect 572076 378150 572128 378156
rect 572088 358766 572116 378150
rect 572076 358760 572128 358766
rect 572076 358702 572128 358708
rect 572076 310616 572128 310622
rect 572076 310558 572128 310564
rect 572088 240145 572116 310558
rect 572260 245676 572312 245682
rect 572260 245618 572312 245624
rect 572074 240136 572130 240145
rect 572074 240071 572130 240080
rect 572076 229628 572128 229634
rect 572076 229570 572128 229576
rect 571984 193180 572036 193186
rect 571984 193122 572036 193128
rect 571708 159520 571760 159526
rect 571708 159462 571760 159468
rect 571616 3664 571668 3670
rect 571616 3606 571668 3612
rect 571720 3262 571748 159462
rect 571982 156768 572038 156777
rect 571982 156703 572038 156712
rect 571892 155304 571944 155310
rect 571892 155246 571944 155252
rect 571904 6798 571932 155246
rect 571996 19174 572024 156703
rect 571984 19168 572036 19174
rect 571984 19110 572036 19116
rect 571892 6792 571944 6798
rect 571892 6734 571944 6740
rect 572088 3534 572116 229570
rect 572168 157208 572220 157214
rect 572168 157150 572220 157156
rect 572180 114510 572208 157150
rect 572168 114504 572220 114510
rect 572168 114446 572220 114452
rect 572272 17921 572300 245618
rect 572720 153128 572772 153134
rect 572720 153070 572772 153076
rect 572732 136610 572760 153070
rect 572824 151434 572852 677622
rect 573548 556232 573600 556238
rect 573548 556174 573600 556180
rect 572904 487212 572956 487218
rect 572904 487154 572956 487160
rect 572812 151428 572864 151434
rect 572812 151370 572864 151376
rect 572720 136604 572772 136610
rect 572720 136546 572772 136552
rect 572916 21418 572944 487154
rect 573088 462392 573140 462398
rect 573088 462334 573140 462340
rect 572996 368552 573048 368558
rect 572996 368494 573048 368500
rect 573008 25634 573036 368494
rect 573100 237318 573128 462334
rect 573272 357468 573324 357474
rect 573272 357410 573324 357416
rect 573180 253972 573232 253978
rect 573180 253914 573232 253920
rect 573088 237312 573140 237318
rect 573088 237254 573140 237260
rect 573086 233880 573142 233889
rect 573086 233815 573142 233824
rect 572996 25628 573048 25634
rect 572996 25570 573048 25576
rect 572904 21412 572956 21418
rect 572904 21354 572956 21360
rect 572258 17912 572314 17921
rect 572258 17847 572314 17856
rect 573100 3602 573128 233815
rect 573192 28558 573220 253914
rect 573284 235550 573312 357410
rect 573456 310548 573508 310554
rect 573456 310490 573508 310496
rect 573364 296744 573416 296750
rect 573364 296686 573416 296692
rect 573272 235544 573324 235550
rect 573272 235486 573324 235492
rect 573376 194546 573404 296686
rect 573468 240038 573496 310490
rect 573456 240032 573508 240038
rect 573456 239974 573508 239980
rect 573364 194540 573416 194546
rect 573364 194482 573416 194488
rect 573362 159488 573418 159497
rect 573362 159423 573418 159432
rect 573270 155136 573326 155145
rect 573270 155071 573326 155080
rect 573180 28552 573232 28558
rect 573180 28494 573232 28500
rect 573284 6254 573312 155071
rect 573376 20369 573404 159423
rect 573456 155440 573508 155446
rect 573456 155382 573508 155388
rect 573362 20360 573418 20369
rect 573362 20295 573418 20304
rect 573272 6248 573324 6254
rect 573272 6190 573324 6196
rect 573468 3874 573496 155382
rect 573560 18630 573588 556174
rect 574112 57934 574140 682246
rect 575572 682236 575624 682242
rect 575572 682178 575624 682184
rect 575480 681148 575532 681154
rect 575480 681090 575532 681096
rect 574284 674892 574336 674898
rect 574284 674834 574336 674840
rect 574192 549296 574244 549302
rect 574192 549238 574244 549244
rect 574100 57928 574152 57934
rect 574100 57870 574152 57876
rect 574204 18970 574232 549238
rect 574296 194342 574324 674834
rect 574560 503736 574612 503742
rect 574560 503678 574612 503684
rect 574376 483064 574428 483070
rect 574376 483006 574428 483012
rect 574284 194336 574336 194342
rect 574284 194278 574336 194284
rect 574284 153740 574336 153746
rect 574284 153682 574336 153688
rect 574192 18964 574244 18970
rect 574192 18906 574244 18912
rect 573548 18624 573600 18630
rect 573548 18566 573600 18572
rect 573456 3868 573508 3874
rect 573456 3810 573508 3816
rect 574296 3806 574324 153682
rect 574388 21486 574416 483006
rect 574468 300892 574520 300898
rect 574468 300834 574520 300840
rect 574376 21480 574428 21486
rect 574376 21422 574428 21428
rect 574480 11762 574508 300834
rect 574572 236910 574600 503678
rect 574928 501016 574980 501022
rect 574928 500958 574980 500964
rect 574836 423700 574888 423706
rect 574836 423642 574888 423648
rect 574744 360256 574796 360262
rect 574744 360198 574796 360204
rect 574652 266416 574704 266422
rect 574652 266358 574704 266364
rect 574560 236904 574612 236910
rect 574560 236846 574612 236852
rect 574560 162376 574612 162382
rect 574560 162318 574612 162324
rect 574572 26178 574600 162318
rect 574560 26172 574612 26178
rect 574560 26114 574612 26120
rect 574664 23254 574692 266358
rect 574756 60722 574784 360198
rect 574848 237017 574876 423642
rect 574940 325650 574968 500958
rect 574928 325644 574980 325650
rect 574928 325586 574980 325592
rect 575020 307828 575072 307834
rect 575020 307770 575072 307776
rect 574928 299532 574980 299538
rect 574928 299474 574980 299480
rect 574940 239358 574968 299474
rect 575032 273222 575060 307770
rect 575020 273216 575072 273222
rect 575020 273158 575072 273164
rect 574928 239352 574980 239358
rect 574928 239294 574980 239300
rect 574834 237008 574890 237017
rect 574834 236943 574890 236952
rect 574928 165028 574980 165034
rect 574928 164970 574980 164976
rect 574836 151156 574888 151162
rect 574836 151098 574888 151104
rect 574744 60716 574796 60722
rect 574744 60658 574796 60664
rect 574848 26722 574876 151098
rect 574940 122806 574968 164970
rect 574928 122800 574980 122806
rect 574928 122742 574980 122748
rect 575492 48278 575520 681090
rect 575584 96626 575612 682178
rect 576124 681216 576176 681222
rect 576124 681158 576176 681164
rect 575940 465112 575992 465118
rect 575940 465054 575992 465060
rect 575664 448588 575716 448594
rect 575664 448530 575716 448536
rect 575572 96620 575624 96626
rect 575572 96562 575624 96568
rect 575480 48272 575532 48278
rect 575480 48214 575532 48220
rect 574836 26716 574888 26722
rect 574836 26658 574888 26664
rect 574652 23248 574704 23254
rect 574652 23190 574704 23196
rect 575676 21826 575704 448530
rect 575848 353320 575900 353326
rect 575848 353262 575900 353268
rect 575756 346520 575808 346526
rect 575756 346462 575808 346468
rect 575664 21820 575716 21826
rect 575664 21762 575716 21768
rect 575768 16046 575796 346462
rect 575860 25906 575888 353262
rect 575952 191826 575980 465054
rect 576032 273284 576084 273290
rect 576032 273226 576084 273232
rect 575940 191820 575992 191826
rect 575940 191762 575992 191768
rect 575940 152992 575992 152998
rect 575940 152934 575992 152940
rect 575952 27577 575980 152934
rect 575938 27568 575994 27577
rect 575938 27503 575994 27512
rect 575848 25900 575900 25906
rect 575848 25842 575900 25848
rect 575756 16040 575808 16046
rect 575756 15982 575808 15988
rect 576044 15910 576072 273226
rect 576136 73166 576164 681158
rect 576216 456816 576268 456822
rect 576216 456758 576268 456764
rect 576228 113150 576256 456758
rect 576308 316056 576360 316062
rect 576308 315998 576360 316004
rect 576320 241262 576348 315998
rect 576308 241256 576360 241262
rect 576308 241198 576360 241204
rect 576308 229900 576360 229906
rect 576308 229842 576360 229848
rect 576216 113144 576268 113150
rect 576216 113086 576268 113092
rect 576124 73160 576176 73166
rect 576124 73102 576176 73108
rect 576032 15904 576084 15910
rect 576032 15846 576084 15852
rect 576320 13190 576348 229842
rect 576872 14618 576900 684558
rect 577044 682100 577096 682106
rect 577044 682042 577096 682048
rect 576950 680912 577006 680921
rect 576950 680847 577006 680856
rect 576964 23186 576992 680847
rect 577056 26081 577084 682042
rect 579068 679108 579120 679114
rect 579068 679050 579120 679056
rect 577504 619676 577556 619682
rect 577504 619618 577556 619624
rect 577228 585200 577280 585206
rect 577228 585142 577280 585148
rect 577136 426488 577188 426494
rect 577136 426430 577188 426436
rect 577042 26072 577098 26081
rect 577042 26007 577098 26016
rect 576952 23180 577004 23186
rect 576952 23122 577004 23128
rect 576860 14612 576912 14618
rect 576860 14554 576912 14560
rect 576308 13184 576360 13190
rect 576308 13126 576360 13132
rect 574468 11756 574520 11762
rect 574468 11698 574520 11704
rect 574284 3800 574336 3806
rect 574284 3742 574336 3748
rect 573088 3596 573140 3602
rect 573088 3538 573140 3544
rect 572076 3528 572128 3534
rect 572076 3470 572128 3476
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 571708 3256 571760 3262
rect 571708 3198 571760 3204
rect 573928 480 573956 3470
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577148 354 577176 426430
rect 577240 177313 577268 585142
rect 577320 469260 577372 469266
rect 577320 469202 577372 469208
rect 577226 177304 577282 177313
rect 577226 177239 577282 177248
rect 577226 162208 577282 162217
rect 577226 162143 577282 162152
rect 577240 17950 577268 162143
rect 577332 66230 577360 469202
rect 577412 309188 577464 309194
rect 577412 309130 577464 309136
rect 577320 66224 577372 66230
rect 577320 66166 577372 66172
rect 577424 28490 577452 309130
rect 577516 179382 577544 619618
rect 577596 616888 577648 616894
rect 577596 616830 577648 616836
rect 577608 431798 577636 616830
rect 578884 612808 578936 612814
rect 578884 612750 578936 612756
rect 578332 449948 578384 449954
rect 578332 449890 578384 449896
rect 577688 436144 577740 436150
rect 577688 436086 577740 436092
rect 577596 431792 577648 431798
rect 577596 431734 577648 431740
rect 577596 244316 577648 244322
rect 577596 244258 577648 244264
rect 577504 179376 577556 179382
rect 577504 179318 577556 179324
rect 577504 156800 577556 156806
rect 577504 156742 577556 156748
rect 577412 28484 577464 28490
rect 577412 28426 577464 28432
rect 577516 22030 577544 156742
rect 577504 22024 577556 22030
rect 577504 21966 577556 21972
rect 577228 17944 577280 17950
rect 577228 17886 577280 17892
rect 577608 17882 577636 244258
rect 577700 239494 577728 436086
rect 577688 239488 577740 239494
rect 577688 239430 577740 239436
rect 578240 155236 578292 155242
rect 578240 155178 578292 155184
rect 578252 131102 578280 155178
rect 578240 131096 578292 131102
rect 578240 131038 578292 131044
rect 578344 27470 578372 449890
rect 578424 365764 578476 365770
rect 578424 365706 578476 365712
rect 578332 27464 578384 27470
rect 578332 27406 578384 27412
rect 578436 25770 578464 365706
rect 578700 346452 578752 346458
rect 578700 346394 578752 346400
rect 578516 288448 578568 288454
rect 578516 288390 578568 288396
rect 578528 25838 578556 288390
rect 578608 270564 578660 270570
rect 578608 270506 578660 270512
rect 578620 27130 578648 270506
rect 578712 237182 578740 346394
rect 578792 327140 578844 327146
rect 578792 327082 578844 327088
rect 578804 240009 578832 327082
rect 578790 240000 578846 240009
rect 578790 239935 578846 239944
rect 578700 237176 578752 237182
rect 578700 237118 578752 237124
rect 578700 234048 578752 234054
rect 578700 233990 578752 233996
rect 578608 27124 578660 27130
rect 578608 27066 578660 27072
rect 578516 25832 578568 25838
rect 578516 25774 578568 25780
rect 578424 25764 578476 25770
rect 578424 25706 578476 25712
rect 578238 24032 578294 24041
rect 578238 23967 578240 23976
rect 578292 23967 578294 23976
rect 578240 23938 578292 23944
rect 577596 17876 577648 17882
rect 577596 17818 577648 17824
rect 578712 3942 578740 233990
rect 578792 160948 578844 160954
rect 578792 160890 578844 160896
rect 578804 132462 578832 160890
rect 578792 132456 578844 132462
rect 578792 132398 578844 132404
rect 578896 19825 578924 612750
rect 578976 586560 579028 586566
rect 578976 586502 579028 586508
rect 578882 19816 578938 19825
rect 578882 19751 578938 19760
rect 578700 3936 578752 3942
rect 578700 3878 578752 3884
rect 578988 3330 579016 586502
rect 579080 258913 579108 679050
rect 579172 405686 579200 697167
rect 580908 685908 580960 685914
rect 580908 685850 580960 685856
rect 579252 683732 579304 683738
rect 579252 683674 579304 683680
rect 579160 405680 579212 405686
rect 579160 405622 579212 405628
rect 579066 258904 579122 258913
rect 579066 258839 579122 258848
rect 579264 14414 579292 683674
rect 580356 683188 580408 683194
rect 580356 683130 580408 683136
rect 580264 681284 580316 681290
rect 580264 681226 580316 681232
rect 579620 677612 579672 677618
rect 579620 677554 579672 677560
rect 579632 25945 579660 677554
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 579896 431792 579948 431798
rect 579896 431734 579948 431740
rect 579908 431633 579936 431734
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579712 415472 579764 415478
rect 579712 415414 579764 415420
rect 579724 28694 579752 415414
rect 580080 412684 580132 412690
rect 580080 412626 580132 412632
rect 579896 403028 579948 403034
rect 579896 402970 579948 402976
rect 579804 387864 579856 387870
rect 579804 387806 579856 387812
rect 579816 35894 579844 387806
rect 579908 45558 579936 402970
rect 579988 317484 580040 317490
rect 579988 317426 580040 317432
rect 579896 45552 579948 45558
rect 579896 45494 579948 45500
rect 579816 35866 579936 35894
rect 579802 33144 579858 33153
rect 579802 33079 579804 33088
rect 579856 33079 579858 33088
rect 579804 33050 579856 33056
rect 579712 28688 579764 28694
rect 579712 28630 579764 28636
rect 579908 27198 579936 35866
rect 580000 27946 580028 317426
rect 580092 185774 580120 412626
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580172 232280 580224 232286
rect 580172 232222 580224 232228
rect 580080 185768 580132 185774
rect 580080 185710 580132 185716
rect 580080 179376 580132 179382
rect 580080 179318 580132 179324
rect 580092 179217 580120 179318
rect 580078 179208 580134 179217
rect 580078 179143 580134 179152
rect 580080 162444 580132 162450
rect 580080 162386 580132 162392
rect 579988 27940 580040 27946
rect 579988 27882 580040 27888
rect 579896 27192 579948 27198
rect 579896 27134 579948 27140
rect 580092 25974 580120 162386
rect 580080 25968 580132 25974
rect 579618 25936 579674 25945
rect 580080 25910 580132 25916
rect 579618 25871 579674 25880
rect 580184 17134 580212 232222
rect 580276 219065 580304 681226
rect 580368 484673 580396 683130
rect 580448 681896 580500 681902
rect 580448 681838 580500 681844
rect 580460 537849 580488 681838
rect 580724 681352 580776 681358
rect 580724 681294 580776 681300
rect 580630 680640 580686 680649
rect 580630 680575 580686 680584
rect 580540 679312 580592 679318
rect 580540 679254 580592 679260
rect 580552 564369 580580 679254
rect 580644 577697 580672 680575
rect 580736 591025 580764 681294
rect 580816 679176 580868 679182
rect 580816 679118 580868 679124
rect 580828 617545 580856 679118
rect 580920 670721 580948 685850
rect 581000 685092 581052 685098
rect 581000 685034 581052 685040
rect 580906 670712 580962 670721
rect 580906 670647 580962 670656
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580814 617536 580870 617545
rect 580814 617471 580870 617480
rect 580920 600982 580948 643991
rect 580908 600976 580960 600982
rect 580908 600918 580960 600924
rect 580722 591016 580778 591025
rect 580722 590951 580778 590960
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580538 564360 580594 564369
rect 580538 564295 580594 564304
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580354 484664 580410 484673
rect 580354 484599 580410 484608
rect 580448 420232 580500 420238
rect 580448 420174 580500 420180
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580368 235958 580396 418231
rect 580460 365129 580488 420174
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580446 312080 580502 312089
rect 580446 312015 580502 312024
rect 580460 237250 580488 312015
rect 580448 237244 580500 237250
rect 580448 237186 580500 237192
rect 580356 235952 580408 235958
rect 580356 235894 580408 235900
rect 580448 234456 580500 234462
rect 580448 234398 580500 234404
rect 580356 232552 580408 232558
rect 580356 232494 580408 232500
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 580264 193180 580316 193186
rect 580264 193122 580316 193128
rect 580276 192545 580304 193122
rect 580262 192536 580318 192545
rect 580262 192471 580318 192480
rect 580264 152516 580316 152522
rect 580264 152458 580316 152464
rect 580276 99521 580304 152458
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580264 73160 580316 73166
rect 580264 73102 580316 73108
rect 580276 73001 580304 73102
rect 580262 72992 580318 73001
rect 580262 72927 580318 72936
rect 580264 60716 580316 60722
rect 580264 60658 580316 60664
rect 580276 59673 580304 60658
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 580368 24682 580396 232494
rect 580460 232286 580488 234398
rect 580448 232280 580500 232286
rect 580448 232222 580500 232228
rect 580448 227112 580500 227118
rect 580448 227054 580500 227060
rect 580460 152697 580488 227054
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580448 139392 580500 139398
rect 580446 139360 580448 139369
rect 580500 139360 580502 139369
rect 580446 139295 580502 139304
rect 580448 113144 580500 113150
rect 580448 113086 580500 113092
rect 580460 112849 580488 113086
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580356 24676 580408 24682
rect 580356 24618 580408 24624
rect 580172 17128 580224 17134
rect 580172 17070 580224 17076
rect 581012 14958 581040 685034
rect 582380 685024 582432 685030
rect 582380 684966 582432 684972
rect 581184 614168 581236 614174
rect 581184 614110 581236 614116
rect 581092 590708 581144 590714
rect 581092 590650 581144 590656
rect 581104 23458 581132 590650
rect 581196 185638 581224 614110
rect 581460 534132 581512 534138
rect 581460 534074 581512 534080
rect 581276 444440 581328 444446
rect 581276 444382 581328 444388
rect 581184 185632 581236 185638
rect 581184 185574 581236 185580
rect 581184 162580 581236 162586
rect 581184 162522 581236 162528
rect 581092 23452 581144 23458
rect 581092 23394 581144 23400
rect 581000 14952 581052 14958
rect 581000 14894 581052 14900
rect 579252 14408 579304 14414
rect 579252 14350 579304 14356
rect 581196 12170 581224 162522
rect 581288 17542 581316 444382
rect 581368 325780 581420 325786
rect 581368 325722 581420 325728
rect 581380 23390 581408 325722
rect 581472 241330 581500 534074
rect 581736 394732 581788 394738
rect 581736 394674 581788 394680
rect 581644 390652 581696 390658
rect 581644 390594 581696 390600
rect 581460 241324 581512 241330
rect 581460 241266 581512 241272
rect 581550 229800 581606 229809
rect 581550 229735 581606 229744
rect 581460 211812 581512 211818
rect 581460 211754 581512 211760
rect 581368 23384 581420 23390
rect 581368 23326 581420 23332
rect 581276 17536 581328 17542
rect 581276 17478 581328 17484
rect 581184 12164 581236 12170
rect 581184 12106 581236 12112
rect 579804 7608 579856 7614
rect 579804 7550 579856 7556
rect 578976 3324 579028 3330
rect 578976 3266 579028 3272
rect 579816 480 579844 7550
rect 577382 354 577494 480
rect 577148 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 354 581082 480
rect 581472 354 581500 211754
rect 581564 3738 581592 229735
rect 581656 181490 581684 390594
rect 581748 189038 581776 394674
rect 581828 229764 581880 229770
rect 581828 229706 581880 229712
rect 581736 189032 581788 189038
rect 581736 188974 581788 188980
rect 581644 181484 581696 181490
rect 581644 181426 581696 181432
rect 581644 165164 581696 165170
rect 581644 165106 581696 165112
rect 581656 35902 581684 165106
rect 581736 164960 581788 164966
rect 581736 164902 581788 164908
rect 581748 89690 581776 164902
rect 581736 89684 581788 89690
rect 581736 89626 581788 89632
rect 581644 35896 581696 35902
rect 581644 35838 581696 35844
rect 581840 29646 581868 229706
rect 581828 29640 581880 29646
rect 581828 29582 581880 29588
rect 582392 15706 582420 684966
rect 582472 684888 582524 684894
rect 582472 684830 582524 684836
rect 582484 16454 582512 684830
rect 582564 683800 582616 683806
rect 582564 683742 582616 683748
rect 582576 30977 582604 683742
rect 582656 679040 582708 679046
rect 582656 678982 582708 678988
rect 582668 191758 582696 678982
rect 582932 572756 582984 572762
rect 582932 572698 582984 572704
rect 582748 400240 582800 400246
rect 582748 400182 582800 400188
rect 582656 191752 582708 191758
rect 582656 191694 582708 191700
rect 582656 162648 582708 162654
rect 582656 162590 582708 162596
rect 582562 30968 582618 30977
rect 582562 30903 582618 30912
rect 582668 24546 582696 162590
rect 582656 24540 582708 24546
rect 582656 24482 582708 24488
rect 582760 17746 582788 400182
rect 582840 376780 582892 376786
rect 582840 376722 582892 376728
rect 582852 27334 582880 376722
rect 582944 236978 582972 572698
rect 583024 350600 583076 350606
rect 583024 350542 583076 350548
rect 582932 236972 582984 236978
rect 582932 236914 582984 236920
rect 582932 210452 582984 210458
rect 582932 210394 582984 210400
rect 582840 27328 582892 27334
rect 582840 27270 582892 27276
rect 582748 17740 582800 17746
rect 582748 17682 582800 17688
rect 582944 16574 582972 210394
rect 583036 17610 583064 350542
rect 583484 349172 583536 349178
rect 583484 349114 583536 349120
rect 583116 313336 583168 313342
rect 583116 313278 583168 313284
rect 583128 28121 583156 313278
rect 583208 305040 583260 305046
rect 583208 304982 583260 304988
rect 583220 28626 583248 304982
rect 583300 291236 583352 291242
rect 583300 291178 583352 291184
rect 583312 31754 583340 291178
rect 583392 259480 583444 259486
rect 583392 259422 583444 259428
rect 583300 31748 583352 31754
rect 583300 31690 583352 31696
rect 583404 28762 583432 259422
rect 583496 237386 583524 349114
rect 583576 325712 583628 325718
rect 583576 325654 583628 325660
rect 583484 237380 583536 237386
rect 583484 237322 583536 237328
rect 583588 142118 583616 325654
rect 583668 238060 583720 238066
rect 583668 238002 583720 238008
rect 583576 142112 583628 142118
rect 583576 142054 583628 142060
rect 583392 28756 583444 28762
rect 583392 28698 583444 28704
rect 583208 28620 583260 28626
rect 583208 28562 583260 28568
rect 583114 28112 583170 28121
rect 583114 28047 583170 28056
rect 583024 17604 583076 17610
rect 583024 17546 583076 17552
rect 582944 16546 583432 16574
rect 582472 16448 582524 16454
rect 582472 16390 582524 16396
rect 582380 15700 582432 15706
rect 582380 15642 582432 15648
rect 581552 3732 581604 3738
rect 581552 3674 581604 3680
rect 582196 3324 582248 3330
rect 582196 3266 582248 3272
rect 582208 480 582236 3266
rect 583404 480 583432 16546
rect 583680 12034 583708 238002
rect 583668 12028 583720 12034
rect 583668 11970 583720 11976
rect 580970 326 581500 354
rect 580970 -960 581082 326
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 24306 700304 24362 700360
rect 21362 683304 21418 683360
rect 3238 566888 3294 566944
rect 3514 671200 3570 671256
rect 3606 658144 3662 658200
rect 3606 619112 3662 619168
rect 3698 606056 3754 606112
rect 3698 584296 3754 584352
rect 3422 553832 3478 553888
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3422 501744 3478 501800
rect 3146 449520 3202 449576
rect 2962 410488 3018 410544
rect 3146 358400 3202 358456
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 2962 201864 3018 201920
rect 3514 462576 3570 462632
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 345344 3570 345400
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 2962 194520 3018 194576
rect 2778 192480 2834 192536
rect 3146 136720 3202 136776
rect 2870 97552 2926 97608
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 84632 3570 84688
rect 3422 58520 3478 58576
rect 1674 7520 1730 7576
rect 3422 6432 3478 6488
rect 17866 19760 17922 19816
rect 20626 152632 20682 152688
rect 26882 683168 26938 683224
rect 24674 681400 24730 681456
rect 23386 587152 23442 587208
rect 22650 560904 22706 560960
rect 21638 151136 21694 151192
rect 22006 23296 22062 23352
rect 20534 20440 20590 20496
rect 19246 18944 19302 19000
rect 23294 29008 23350 29064
rect 24582 560768 24638 560824
rect 25962 561992 26018 562048
rect 26146 561856 26202 561912
rect 171782 681264 171838 681320
rect 165526 678136 165582 678192
rect 153106 677628 153108 677648
rect 153108 677628 153160 677648
rect 153160 677628 153162 677648
rect 153106 677592 153162 677628
rect 32862 628224 32918 628280
rect 31574 627952 31630 628008
rect 31390 625368 31446 625424
rect 28906 587288 28962 587344
rect 27526 562128 27582 562184
rect 27342 561312 27398 561368
rect 26882 253952 26938 254008
rect 27066 151000 27122 151056
rect 28078 198464 28134 198520
rect 27618 184456 27674 184512
rect 24766 17040 24822 17096
rect 28446 155216 28502 155272
rect 28262 151272 28318 151328
rect 31482 619656 31538 619712
rect 32770 622376 32826 622432
rect 31666 601704 31722 601760
rect 30102 561720 30158 561776
rect 29458 198328 29514 198384
rect 30010 561040 30066 561096
rect 30286 28872 30342 28928
rect 32678 600344 32734 600400
rect 33046 624144 33102 624200
rect 32954 621288 33010 621344
rect 32678 559952 32734 560008
rect 31390 193160 31446 193216
rect 19430 6160 19486 6216
rect 24214 3440 24270 3496
rect 31758 187176 31814 187232
rect 32402 186904 32458 186960
rect 35254 589872 35310 589928
rect 33046 198736 33102 198792
rect 32678 20576 32734 20632
rect 33690 184728 33746 184784
rect 34150 199144 34206 199200
rect 34242 152904 34298 152960
rect 35070 224168 35126 224224
rect 34978 211792 35034 211848
rect 34886 198600 34942 198656
rect 35254 17448 35310 17504
rect 35806 153040 35862 153096
rect 36542 199688 36598 199744
rect 50066 590552 50122 590608
rect 55862 590552 55918 590608
rect 60370 590552 60426 590608
rect 69018 590552 69074 590608
rect 74814 590552 74870 590608
rect 77850 590552 77906 590608
rect 42522 590008 42578 590064
rect 37646 201320 37702 201376
rect 37554 201048 37610 201104
rect 37186 199824 37242 199880
rect 38198 195744 38254 195800
rect 38382 197784 38438 197840
rect 38290 176024 38346 176080
rect 39762 195472 39818 195528
rect 39670 178880 39726 178936
rect 40314 183232 40370 183288
rect 41050 195608 41106 195664
rect 42246 560088 42302 560144
rect 42062 209480 42118 209536
rect 43350 558864 43406 558920
rect 43810 561176 43866 561232
rect 43626 292576 43682 292632
rect 43718 195336 43774 195392
rect 44730 321544 44786 321600
rect 45006 372952 45062 373008
rect 44914 283192 44970 283248
rect 44822 242936 44878 242992
rect 44730 241440 44786 241496
rect 45098 359352 45154 359408
rect 44730 152768 44786 152824
rect 44914 31048 44970 31104
rect 45282 339496 45338 339552
rect 45190 264696 45246 264752
rect 45190 237360 45246 237416
rect 46110 556552 46166 556608
rect 45926 556144 45982 556200
rect 45742 521736 45798 521792
rect 45650 520648 45706 520704
rect 45558 520396 45614 520432
rect 45558 520376 45560 520396
rect 45560 520376 45612 520396
rect 45612 520376 45614 520396
rect 45558 516568 45614 516624
rect 45558 515208 45614 515264
rect 45834 501336 45890 501392
rect 45834 497256 45890 497312
rect 45650 463800 45706 463856
rect 45650 425176 45706 425232
rect 45650 420980 45706 421016
rect 45650 420960 45652 420980
rect 45652 420960 45704 420980
rect 45704 420960 45706 420980
rect 45650 419620 45706 419656
rect 45650 419600 45652 419620
rect 45652 419600 45704 419620
rect 45704 419600 45706 419620
rect 45650 415540 45706 415576
rect 45650 415520 45652 415540
rect 45652 415520 45704 415540
rect 45704 415520 45706 415540
rect 45650 281580 45706 281616
rect 45650 281560 45652 281580
rect 45652 281560 45704 281580
rect 45704 281560 45706 281580
rect 45374 251776 45430 251832
rect 45558 232192 45614 232248
rect 45558 230560 45614 230616
rect 45558 227840 45614 227896
rect 45466 213968 45522 214024
rect 45558 211248 45614 211304
rect 46110 551248 46166 551304
rect 46110 550860 46166 550896
rect 46110 550840 46112 550860
rect 46112 550840 46164 550860
rect 46164 550840 46166 550860
rect 46110 549752 46166 549808
rect 46110 548256 46166 548312
rect 46110 544176 46166 544232
rect 46110 528944 46166 529000
rect 46294 526496 46350 526552
rect 46018 510856 46074 510912
rect 46018 494536 46074 494592
rect 46202 513848 46258 513904
rect 46110 474136 46166 474192
rect 46018 439592 46074 439648
rect 45926 429936 45982 429992
rect 45926 420008 45982 420064
rect 45926 418648 45982 418704
rect 45926 415928 45982 415984
rect 46110 392672 46166 392728
rect 46018 392128 46074 392184
rect 46110 385736 46166 385792
rect 46018 366016 46074 366072
rect 46110 310936 46166 310992
rect 46110 309188 46166 309224
rect 46110 309168 46112 309188
rect 46112 309168 46164 309188
rect 46164 309168 46166 309188
rect 46110 292576 46166 292632
rect 46018 258304 46074 258360
rect 45926 233416 45982 233472
rect 46018 230832 46074 230888
rect 46110 218592 46166 218648
rect 45558 207576 45614 207632
rect 45834 212608 45890 212664
rect 45650 206932 45652 206952
rect 45652 206932 45704 206952
rect 45704 206932 45706 206952
rect 45650 206896 45706 206932
rect 45650 205944 45706 206000
rect 46386 496032 46442 496088
rect 46386 489932 46442 489968
rect 46386 489912 46388 489932
rect 46388 489912 46440 489932
rect 46440 489912 46442 489932
rect 46294 318416 46350 318472
rect 46294 314744 46350 314800
rect 46294 310256 46350 310312
rect 46478 482296 46534 482352
rect 46754 545672 46810 545728
rect 46754 544312 46810 544368
rect 46754 541048 46810 541104
rect 46754 538056 46810 538112
rect 46754 533296 46810 533352
rect 46754 532072 46810 532128
rect 46754 529932 46756 529952
rect 46756 529932 46808 529952
rect 46808 529932 46810 529952
rect 46754 529896 46810 529932
rect 46754 525136 46810 525192
rect 46754 509496 46810 509552
rect 46754 505164 46810 505200
rect 46754 505144 46756 505164
rect 46756 505144 46808 505164
rect 46808 505144 46810 505164
rect 46754 500656 46810 500712
rect 46754 495896 46810 495952
rect 46754 495216 46810 495272
rect 46754 493176 46810 493232
rect 46754 490592 46810 490648
rect 46754 489812 46756 489832
rect 46756 489812 46808 489832
rect 46808 489812 46810 489832
rect 46754 489776 46810 489812
rect 46754 485852 46810 485888
rect 46754 485832 46756 485852
rect 46756 485832 46808 485852
rect 46808 485832 46810 485852
rect 46754 484744 46810 484800
rect 46754 483384 46810 483440
rect 46662 480256 46718 480312
rect 46570 475496 46626 475552
rect 46570 473456 46626 473512
rect 46570 468288 46626 468344
rect 46570 459856 46626 459912
rect 46754 476448 46810 476504
rect 46754 469648 46810 469704
rect 46754 468016 46810 468072
rect 46754 464208 46810 464264
rect 46754 463256 46810 463312
rect 46754 460964 46810 461000
rect 46754 460944 46756 460964
rect 46756 460944 46808 460964
rect 46808 460944 46810 460964
rect 46754 458244 46810 458280
rect 46754 458224 46756 458244
rect 46756 458224 46808 458244
rect 46808 458224 46810 458244
rect 46754 456456 46810 456512
rect 46754 450336 46810 450392
rect 46754 445848 46810 445904
rect 46754 445032 46810 445088
rect 46754 443264 46810 443320
rect 46662 442856 46718 442912
rect 46754 439048 46810 439104
rect 46754 436464 46810 436520
rect 46754 434732 46756 434752
rect 46756 434732 46808 434752
rect 46808 434732 46810 434752
rect 46754 434696 46810 434732
rect 46754 433608 46810 433664
rect 46754 431996 46810 432032
rect 46754 431976 46756 431996
rect 46756 431976 46808 431996
rect 46808 431976 46810 431996
rect 46662 428304 46718 428360
rect 46754 427896 46810 427952
rect 46662 425312 46718 425368
rect 46570 421232 46626 421288
rect 46478 390496 46534 390552
rect 46478 389272 46534 389328
rect 46478 386436 46534 386472
rect 46478 386416 46480 386436
rect 46480 386416 46532 386436
rect 46532 386416 46534 386436
rect 46478 385076 46534 385112
rect 46478 385056 46480 385076
rect 46480 385056 46532 385076
rect 46532 385056 46534 385076
rect 46478 383016 46534 383072
rect 46478 376216 46534 376272
rect 46478 354748 46534 354784
rect 46478 354728 46480 354748
rect 46480 354728 46532 354748
rect 46532 354728 46534 354748
rect 46478 353096 46534 353152
rect 46478 349172 46534 349208
rect 46478 349152 46480 349172
rect 46480 349152 46532 349172
rect 46532 349152 46534 349172
rect 46478 347112 46534 347168
rect 46478 345092 46534 345128
rect 46478 345072 46480 345092
rect 46480 345072 46532 345092
rect 46532 345072 46534 345092
rect 46478 336796 46534 336832
rect 46478 336776 46480 336796
rect 46480 336776 46532 336796
rect 46532 336776 46534 336796
rect 46478 330656 46534 330712
rect 46478 328888 46534 328944
rect 46478 325216 46534 325272
rect 46386 302912 46442 302968
rect 46294 302232 46350 302288
rect 46386 300892 46442 300928
rect 46386 300872 46388 300892
rect 46388 300872 46440 300892
rect 46440 300872 46442 300892
rect 46386 298172 46442 298208
rect 46386 298152 46388 298172
rect 46388 298152 46440 298172
rect 46440 298152 46442 298172
rect 46386 297064 46442 297120
rect 46386 292848 46442 292904
rect 46386 291488 46442 291544
rect 46386 285776 46442 285832
rect 46478 268232 46534 268288
rect 46386 267844 46442 267880
rect 46386 267824 46388 267844
rect 46388 267824 46440 267844
rect 46440 267824 46442 267844
rect 46478 256672 46534 256728
rect 46386 236000 46442 236056
rect 46294 226616 46350 226672
rect 46386 224848 46442 224904
rect 46294 217232 46350 217288
rect 46202 198056 46258 198112
rect 46386 202836 46442 202872
rect 46386 202816 46388 202836
rect 46388 202816 46440 202836
rect 46440 202816 46442 202836
rect 46386 201592 46442 201648
rect 46018 150456 46074 150512
rect 46018 100000 46074 100056
rect 46754 423700 46810 423736
rect 46754 423680 46756 423700
rect 46756 423680 46808 423700
rect 46808 423680 46810 423700
rect 46754 414044 46810 414080
rect 46754 414024 46756 414044
rect 46756 414024 46808 414044
rect 46808 414024 46810 414044
rect 46754 411324 46810 411360
rect 46754 411304 46756 411324
rect 46756 411304 46808 411324
rect 46808 411304 46810 411324
rect 46754 407632 46810 407688
rect 46754 403552 46810 403608
rect 46754 400288 46810 400344
rect 46754 399472 46810 399528
rect 46754 394732 46810 394768
rect 46754 394712 46756 394732
rect 46756 394712 46808 394732
rect 46808 394712 46810 394732
rect 46754 393488 46810 393544
rect 46662 247016 46718 247072
rect 46570 244296 46626 244352
rect 46662 238176 46718 238232
rect 46662 234660 46718 234696
rect 46662 234640 46664 234660
rect 46664 234640 46716 234660
rect 46716 234640 46718 234660
rect 46662 224032 46718 224088
rect 46662 222400 46718 222456
rect 46570 221312 46626 221368
rect 46662 221040 46718 221096
rect 46662 218320 46718 218376
rect 46662 216708 46718 216744
rect 46662 216688 46664 216708
rect 46664 216688 46716 216708
rect 46716 216688 46718 216708
rect 46662 215348 46718 215384
rect 46662 215328 46664 215348
rect 46664 215328 46716 215348
rect 46716 215328 46718 215348
rect 46662 203632 46718 203688
rect 47030 438776 47086 438832
rect 46846 380976 46902 381032
rect 46846 379752 46902 379808
rect 46846 372680 46902 372736
rect 46846 371456 46902 371512
rect 46846 368872 46902 368928
rect 46846 367512 46902 367568
rect 46846 363432 46902 363488
rect 46846 357856 46902 357912
rect 47030 335416 47086 335472
rect 46846 323040 46902 323096
rect 46846 321680 46902 321736
rect 46846 320204 46902 320240
rect 46846 320184 46848 320204
rect 46848 320184 46900 320204
rect 46900 320184 46902 320204
rect 46846 318980 46902 319016
rect 46846 318960 46848 318980
rect 46848 318960 46900 318980
rect 46900 318960 46902 318980
rect 46846 281832 46902 281888
rect 46846 277752 46902 277808
rect 46846 273672 46902 273728
rect 46846 253972 46902 254008
rect 46846 253952 46848 253972
rect 46848 253952 46900 253972
rect 46900 253952 46902 253972
rect 46846 247424 46902 247480
rect 46846 245792 46902 245848
rect 46754 200096 46810 200152
rect 46478 155896 46534 155952
rect 46938 210432 46994 210488
rect 46846 195200 46902 195256
rect 47398 524592 47454 524648
rect 47306 327936 47362 327992
rect 47306 304952 47362 305008
rect 47214 298016 47270 298072
rect 47490 504056 47546 504112
rect 47490 329840 47546 329896
rect 47398 282920 47454 282976
rect 47214 273264 47270 273320
rect 47122 270136 47178 270192
rect 47122 209616 47178 209672
rect 47398 220768 47454 220824
rect 47306 201184 47362 201240
rect 67638 589600 67694 589656
rect 51078 589464 51134 589520
rect 53838 589464 53894 589520
rect 60646 589464 60702 589520
rect 62210 589464 62266 589520
rect 47766 562264 47822 562320
rect 47766 558864 47822 558920
rect 47674 257896 47730 257952
rect 47582 229744 47638 229800
rect 47398 199008 47454 199064
rect 47766 200912 47822 200968
rect 47674 151408 47730 151464
rect 48962 562536 49018 562592
rect 51170 589328 51226 589384
rect 53746 589328 53802 589384
rect 53746 566344 53802 566400
rect 56690 589328 56746 589384
rect 57978 589328 58034 589384
rect 57978 562128 58034 562184
rect 57426 561992 57482 562048
rect 56690 560904 56746 560960
rect 60738 589328 60794 589384
rect 62118 589328 62174 589384
rect 59818 564440 59874 564496
rect 58530 561992 58586 562048
rect 58530 560088 58586 560144
rect 59910 561856 59966 561912
rect 60738 561856 60794 561912
rect 60738 561176 60794 561232
rect 63498 589328 63554 589384
rect 64786 589328 64842 589384
rect 65430 589328 65486 589384
rect 66258 589328 66314 589384
rect 67546 589328 67602 589384
rect 64786 566480 64842 566536
rect 63498 561040 63554 561096
rect 63222 560360 63278 560416
rect 72422 589464 72478 589520
rect 74538 589464 74594 589520
rect 67730 589328 67786 589384
rect 70306 589328 70362 589384
rect 71134 589328 71190 589384
rect 71778 589328 71834 589384
rect 71134 582936 71190 582992
rect 73158 589328 73214 589384
rect 72422 584432 72478 584488
rect 75182 590416 75238 590472
rect 77298 590416 77354 590472
rect 75182 589736 75238 589792
rect 75642 589328 75698 589384
rect 75918 589328 75974 589384
rect 78678 590416 78734 590472
rect 78678 589464 78734 589520
rect 77850 588512 77906 588568
rect 77942 564576 77998 564632
rect 99930 590552 99986 590608
rect 107566 590552 107622 590608
rect 127346 590552 127402 590608
rect 129738 590552 129794 590608
rect 92478 590416 92534 590472
rect 81346 589464 81402 589520
rect 82726 589464 82782 589520
rect 84198 589464 84254 589520
rect 88246 589464 88302 589520
rect 89626 589464 89682 589520
rect 91006 589464 91062 589520
rect 81438 589328 81494 589384
rect 82634 589328 82690 589384
rect 84106 589328 84162 589384
rect 85578 589328 85634 589384
rect 86958 589328 87014 589384
rect 85486 566752 85542 566808
rect 83094 563760 83150 563816
rect 89718 589328 89774 589384
rect 90914 589328 90970 589384
rect 90914 572056 90970 572112
rect 104898 589464 104954 589520
rect 122562 589736 122618 589792
rect 91098 589328 91154 589384
rect 93766 589328 93822 589384
rect 95146 589328 95202 589384
rect 103426 589328 103482 589384
rect 110326 589328 110382 589384
rect 113086 589328 113142 589384
rect 115846 589328 115902 589384
rect 117318 589328 117374 589384
rect 119986 589328 120042 589384
rect 89718 562400 89774 562456
rect 109590 566072 109646 566128
rect 106186 565936 106242 565992
rect 104346 562264 104402 562320
rect 137282 589600 137338 589656
rect 125506 589328 125562 589384
rect 132498 589328 132554 589384
rect 133878 589328 133934 589384
rect 140686 589328 140742 589384
rect 171230 671200 171286 671256
rect 157246 589328 157302 589384
rect 158626 589328 158682 589384
rect 130566 568792 130622 568848
rect 126058 568656 126114 568712
rect 121550 562672 121606 562728
rect 143446 566208 143502 566264
rect 171322 605648 171378 605704
rect 170770 561992 170826 562048
rect 172610 611360 172666 611416
rect 172518 606872 172574 606928
rect 173806 609728 173862 609784
rect 173806 608368 173862 608424
rect 325054 677592 325110 677648
rect 337566 677592 337622 677648
rect 325790 677048 325846 677104
rect 204166 628224 204222 628280
rect 203522 627952 203578 628008
rect 173898 561856 173954 561912
rect 180706 563352 180762 563408
rect 184846 561856 184902 561912
rect 190366 566616 190422 566672
rect 189446 562128 189502 562184
rect 195886 564712 195942 564768
rect 203062 601724 203118 601760
rect 203062 601704 203064 601724
rect 203064 601704 203116 601724
rect 203116 601704 203118 601724
rect 203614 625368 203670 625424
rect 204074 624144 204130 624200
rect 203982 622376 204038 622432
rect 203890 619656 203946 619712
rect 203798 599392 203854 599448
rect 201038 561992 201094 562048
rect 205546 621930 205602 621986
rect 204902 600344 204958 600400
rect 220818 590552 220874 590608
rect 223026 590552 223082 590608
rect 238390 590552 238446 590608
rect 241518 590552 241574 590608
rect 246670 590552 246726 590608
rect 252374 590552 252430 590608
rect 273258 590552 273314 590608
rect 289542 590552 289598 590608
rect 292118 590552 292174 590608
rect 207478 560904 207534 560960
rect 208766 562264 208822 562320
rect 223578 589328 223634 589384
rect 216862 567160 216918 567216
rect 225326 589328 225382 589384
rect 226614 589328 226670 589384
rect 240598 589736 240654 589792
rect 230202 589464 230258 589520
rect 230478 589464 230534 589520
rect 234526 589464 234582 589520
rect 235998 589464 236054 589520
rect 239954 589464 240010 589520
rect 229006 589328 229062 589384
rect 230386 589328 230442 589384
rect 231858 589328 231914 589384
rect 233238 589328 233294 589384
rect 234618 589328 234674 589384
rect 236090 589328 236146 589384
rect 237286 589328 237342 589384
rect 240046 589328 240102 589384
rect 242806 589464 242862 589520
rect 244278 589464 244334 589520
rect 248418 589464 248474 589520
rect 251178 589464 251234 589520
rect 240046 562400 240102 562456
rect 242898 589328 242954 589384
rect 244186 589328 244242 589384
rect 245566 589328 245622 589384
rect 247038 589328 247094 589384
rect 248326 589328 248382 589384
rect 256054 589736 256110 589792
rect 253938 589464 253994 589520
rect 248510 589328 248566 589384
rect 249798 589328 249854 589384
rect 251270 589328 251326 589384
rect 253846 589328 253902 589384
rect 248418 572192 248474 572248
rect 254122 589328 254178 589384
rect 257986 589464 258042 589520
rect 259458 589464 259514 589520
rect 260838 589464 260894 589520
rect 264886 589464 264942 589520
rect 266358 589464 266414 589520
rect 257894 589328 257950 589384
rect 253938 574776 253994 574832
rect 258078 589328 258134 589384
rect 259274 589328 259330 589384
rect 260746 589328 260802 589384
rect 262126 589328 262182 589384
rect 263506 589328 263562 589384
rect 264794 589328 264850 589384
rect 266266 589328 266322 589384
rect 270406 589328 270462 589384
rect 271878 589328 271934 589384
rect 266358 585656 266414 585712
rect 267922 561720 267978 561776
rect 278962 589600 279018 589656
rect 277306 589328 277362 589384
rect 282826 589328 282882 589384
rect 284298 589328 284354 589384
rect 273258 576000 273314 576056
rect 275006 564848 275062 564904
rect 274454 562672 274510 562728
rect 277030 563624 277086 563680
rect 293958 589464 294014 589520
rect 296718 589464 296774 589520
rect 299478 589464 299534 589520
rect 300858 589464 300914 589520
rect 284298 567840 284354 567896
rect 294326 563216 294382 563272
rect 297638 563216 297694 563272
rect 300858 574640 300914 574696
rect 298926 563488 298982 563544
rect 312082 590552 312138 590608
rect 306378 589464 306434 589520
rect 309138 589464 309194 589520
rect 329746 589600 329802 589656
rect 329654 589464 329710 589520
rect 309138 571920 309194 571976
rect 308310 567296 308366 567352
rect 311162 560768 311218 560824
rect 328366 560632 328422 560688
rect 330482 561312 330538 561368
rect 336186 563080 336242 563136
rect 343638 671200 343694 671256
rect 346306 611380 346362 611416
rect 346306 611360 346308 611380
rect 346308 611360 346360 611380
rect 346360 611360 346362 611380
rect 345018 609728 345074 609784
rect 345110 608368 345166 608424
rect 345570 606872 345626 606928
rect 345110 605648 345166 605704
rect 341982 561720 342038 561776
rect 340142 561040 340198 561096
rect 347778 471144 347834 471200
rect 347870 451424 347926 451480
rect 347870 445712 347926 445768
rect 347686 200368 347742 200424
rect 46662 14456 46718 14512
rect 43074 3440 43130 3496
rect 48778 188264 48834 188320
rect 48870 112376 48926 112432
rect 49974 198192 50030 198248
rect 49330 179152 49386 179208
rect 49330 29552 49386 29608
rect 49606 141344 49662 141400
rect 50618 138624 50674 138680
rect 50894 176568 50950 176624
rect 50802 139440 50858 139496
rect 50986 139440 51042 139496
rect 51630 178744 51686 178800
rect 50802 19216 50858 19272
rect 52458 171672 52514 171728
rect 53838 198600 53894 198656
rect 53194 197376 53250 197432
rect 54482 197376 54538 197432
rect 53378 132504 53434 132560
rect 54298 182960 54354 183016
rect 54390 106664 54446 106720
rect 58990 198600 59046 198656
rect 60278 197104 60334 197160
rect 55862 181328 55918 181384
rect 55494 147464 55550 147520
rect 54850 29688 54906 29744
rect 56046 119176 56102 119232
rect 56046 107480 56102 107536
rect 55954 98096 56010 98152
rect 56138 77016 56194 77072
rect 56782 189896 56838 189952
rect 56322 86536 56378 86592
rect 56230 55256 56286 55312
rect 57150 139576 57206 139632
rect 57058 131416 57114 131472
rect 57242 130736 57298 130792
rect 57242 128016 57298 128072
rect 57242 126656 57298 126712
rect 57242 125296 57298 125352
rect 57242 123256 57298 123312
rect 57058 81096 57114 81152
rect 56782 70216 56838 70272
rect 56690 67496 56746 67552
rect 56966 64096 57022 64152
rect 57058 46416 57114 46472
rect 57150 40296 57206 40352
rect 57334 120536 57390 120592
rect 57334 119856 57390 119912
rect 57334 117136 57390 117192
rect 57334 115776 57390 115832
rect 57426 113056 57482 113112
rect 57518 110336 57574 110392
rect 57518 108296 57574 108352
rect 57426 107616 57482 107672
rect 57518 104216 57574 104272
rect 57426 103536 57482 103592
rect 57518 102856 57574 102912
rect 57426 102176 57482 102232
rect 57518 99456 57574 99512
rect 57518 96736 57574 96792
rect 57334 30776 57390 30832
rect 57518 94016 57574 94072
rect 57794 168952 57850 169008
rect 57610 82456 57666 82512
rect 57610 75656 57666 75712
rect 57610 68176 57666 68232
rect 58346 195472 58402 195528
rect 57886 145696 57942 145752
rect 57886 141616 57942 141672
rect 57886 140256 57942 140312
rect 57886 137536 57942 137592
rect 57886 134816 57942 134872
rect 57886 132776 57942 132832
rect 57886 114280 57942 114336
rect 57886 92656 57942 92712
rect 57886 90616 57942 90672
rect 57886 89256 57942 89312
rect 57886 81776 57942 81832
rect 57886 64796 57942 64832
rect 57886 64776 57888 64796
rect 57888 64776 57940 64796
rect 57940 64776 57942 64796
rect 57702 63452 57704 63472
rect 57704 63452 57756 63472
rect 57756 63452 57758 63472
rect 57702 63416 57758 63452
rect 57702 62076 57758 62112
rect 57702 62056 57704 62076
rect 57704 62056 57756 62076
rect 57756 62056 57758 62076
rect 57794 59336 57850 59392
rect 57702 58656 57758 58712
rect 57702 57316 57758 57352
rect 57702 57296 57704 57316
rect 57704 57296 57756 57316
rect 57756 57296 57758 57316
rect 57886 55936 57942 55992
rect 57702 53216 57758 53272
rect 57702 47096 57758 47152
rect 58162 45736 58218 45792
rect 58438 138080 58494 138136
rect 58438 114416 58494 114472
rect 58530 89800 58586 89856
rect 58346 45056 58402 45112
rect 58254 41656 58310 41712
rect 57702 40976 57758 41032
rect 57702 39616 57758 39672
rect 57702 33496 57758 33552
rect 57702 32816 57758 32872
rect 57794 32136 57850 32192
rect 57702 31456 57758 31512
rect 58530 28464 58586 28520
rect 57610 19080 57666 19136
rect 59082 146512 59138 146568
rect 59358 140936 59414 140992
rect 61934 152496 61990 152552
rect 64510 159296 64566 159352
rect 67638 180104 67694 180160
rect 73342 175888 73398 175944
rect 72882 152360 72938 152416
rect 82818 197784 82874 197840
rect 84106 198872 84162 198928
rect 83462 197240 83518 197296
rect 87694 195608 87750 195664
rect 85670 190304 85726 190360
rect 81254 188536 81310 188592
rect 93122 198056 93178 198112
rect 94410 198056 94466 198112
rect 117318 151544 117374 151600
rect 122746 197920 122802 197976
rect 139398 192888 139454 192944
rect 129554 153040 129610 153096
rect 145654 152904 145710 152960
rect 147678 184048 147734 184104
rect 153658 198736 153714 198792
rect 158166 195880 158222 195936
rect 157890 189624 157946 189680
rect 153382 152632 153438 152688
rect 159178 181872 159234 181928
rect 172058 188808 172114 188864
rect 170126 152768 170182 152824
rect 179142 152632 179198 152688
rect 200026 195608 200082 195664
rect 197174 152768 197230 152824
rect 213918 152904 213974 152960
rect 227718 196832 227774 196888
rect 228362 195744 228418 195800
rect 237746 182008 237802 182064
rect 247038 198736 247094 198792
rect 257986 199552 258042 199608
rect 257894 199144 257950 199200
rect 270590 190032 270646 190088
rect 275742 188672 275798 188728
rect 296074 199416 296130 199472
rect 295338 199008 295394 199064
rect 292486 153040 292542 153096
rect 287702 152496 287758 152552
rect 291198 152496 291254 152552
rect 313094 175752 313150 175808
rect 317602 152224 317658 152280
rect 342350 196968 342406 197024
rect 347778 200252 347834 200288
rect 347778 200232 347780 200252
rect 347780 200232 347832 200252
rect 347832 200232 347834 200252
rect 347686 199280 347742 199336
rect 347778 199144 347834 199200
rect 348054 561584 348110 561640
rect 348054 511944 348110 512000
rect 347962 336504 348018 336560
rect 347962 331064 348018 331120
rect 348422 522960 348478 523016
rect 348330 477536 348386 477592
rect 348238 456456 348294 456512
rect 348146 410896 348202 410952
rect 348238 395868 348294 395924
rect 348146 391108 348202 391164
rect 348054 296384 348110 296440
rect 348054 262792 348110 262848
rect 348330 368668 348386 368724
rect 349158 541456 349214 541512
rect 349066 540912 349122 540968
rect 348606 511536 348662 511592
rect 348698 474952 348754 475008
rect 349066 469240 349122 469296
rect 349434 493856 349490 493912
rect 349434 465160 349490 465216
rect 349342 396616 349398 396672
rect 349250 346976 349306 347032
rect 349158 302232 349214 302288
rect 349250 288496 349306 288552
rect 349250 280472 349306 280528
rect 349618 455776 349674 455832
rect 350170 548936 350226 548992
rect 350262 547032 350318 547088
rect 350262 533432 350318 533488
rect 350262 523096 350318 523152
rect 349894 521736 349950 521792
rect 350170 520376 350226 520432
rect 350262 516568 350318 516624
rect 350262 513460 350318 513496
rect 350262 513440 350264 513460
rect 350264 513440 350316 513460
rect 350316 513440 350318 513460
rect 350262 505416 350318 505472
rect 349802 499976 349858 500032
rect 350262 491952 350318 492008
rect 350262 490184 350318 490240
rect 350170 489812 350172 489832
rect 350172 489812 350224 489832
rect 350224 489812 350226 489832
rect 350170 489776 350226 489812
rect 350262 487736 350318 487792
rect 349986 485152 350042 485208
rect 350262 483384 350318 483440
rect 350262 480664 350318 480720
rect 350170 476584 350226 476640
rect 349710 451016 349766 451072
rect 350262 476176 350318 476232
rect 350262 473456 350318 473512
rect 350262 465976 350318 466032
rect 350262 462848 350318 462904
rect 350262 461488 350318 461544
rect 350262 457272 350318 457328
rect 350262 446392 350318 446448
rect 350262 437824 350318 437880
rect 349802 433336 349858 433392
rect 350262 430888 350318 430944
rect 349986 421232 350042 421288
rect 350262 414432 350318 414488
rect 349526 409536 349582 409592
rect 349618 391312 349674 391368
rect 349434 295432 349490 295488
rect 349434 284280 349490 284336
rect 349342 202272 349398 202328
rect 349526 247696 349582 247752
rect 349618 245656 349674 245712
rect 349526 224984 349582 225040
rect 350078 381248 350134 381304
rect 349986 379480 350042 379536
rect 350078 376896 350134 376952
rect 350078 375808 350134 375864
rect 350078 370096 350134 370152
rect 350078 363296 350134 363352
rect 350078 349832 350134 349888
rect 350078 344392 350134 344448
rect 350078 311072 350134 311128
rect 349986 268776 350042 268832
rect 349894 257896 349950 257952
rect 349986 242936 350042 242992
rect 349986 219952 350042 220008
rect 350262 404912 350318 404968
rect 350262 394732 350318 394768
rect 350262 394712 350264 394732
rect 350264 394712 350316 394732
rect 350316 394712 350318 394732
rect 350262 389952 350318 390008
rect 350262 387096 350318 387152
rect 350262 382336 350318 382392
rect 350262 380976 350318 381032
rect 350262 377168 350318 377224
rect 350262 374856 350318 374912
rect 350262 372816 350318 372872
rect 350262 371320 350318 371376
rect 350262 358828 350318 358864
rect 350262 358808 350264 358828
rect 350264 358808 350316 358828
rect 350316 358808 350318 358828
rect 350262 358264 350318 358320
rect 350262 356632 350318 356688
rect 350262 355816 350318 355872
rect 350262 354748 350318 354784
rect 350262 354728 350264 354748
rect 350264 354728 350316 354748
rect 350316 354728 350318 354748
rect 350262 350648 350318 350704
rect 350262 349424 350318 349480
rect 350262 345752 350318 345808
rect 350262 343984 350318 344040
rect 350446 554376 350502 554432
rect 350446 551384 350502 551440
rect 350446 546644 350502 546680
rect 350446 546624 350448 546644
rect 350448 546624 350500 546644
rect 350500 546624 350502 546644
rect 350446 542952 350502 543008
rect 350446 538328 350502 538384
rect 350446 537104 350502 537160
rect 350446 534656 350502 534712
rect 350446 533024 350502 533080
rect 350446 532072 350502 532128
rect 350446 530712 350502 530768
rect 350446 527196 350502 527232
rect 350446 527176 350448 527196
rect 350448 527176 350500 527196
rect 350500 527176 350502 527196
rect 350446 526224 350502 526280
rect 350446 523232 350502 523288
rect 350446 517656 350502 517712
rect 350446 516180 350502 516216
rect 350446 516160 350448 516180
rect 350448 516160 350500 516180
rect 350500 516160 350502 516180
rect 350446 513712 350502 513768
rect 350446 508816 350502 508872
rect 350446 506912 350502 506968
rect 350446 505552 350502 505608
rect 350446 503784 350502 503840
rect 350446 500112 350502 500168
rect 350446 498228 350502 498264
rect 350446 498208 350448 498228
rect 350448 498208 350500 498228
rect 350500 498208 350502 498228
rect 350446 495508 350502 495544
rect 350446 495488 350448 495508
rect 350448 495488 350500 495508
rect 350500 495488 350502 495508
rect 350446 491408 350502 491464
rect 350446 490592 350502 490648
rect 350446 481652 350448 481672
rect 350448 481652 350500 481672
rect 350500 481652 350502 481672
rect 350446 481616 350502 481652
rect 350446 480276 350502 480312
rect 350446 480256 350448 480276
rect 350448 480256 350500 480276
rect 350500 480256 350502 480276
rect 350446 472232 350502 472288
rect 350446 466520 350502 466576
rect 350446 462576 350502 462632
rect 350446 461100 350502 461136
rect 350446 461080 350448 461100
rect 350448 461080 350500 461100
rect 350500 461080 350502 461100
rect 350446 459604 350502 459640
rect 350446 459584 350448 459604
rect 350448 459584 350500 459604
rect 350500 459584 350502 459604
rect 350446 456884 350502 456920
rect 350446 456864 350448 456884
rect 350448 456864 350500 456884
rect 350500 456864 350502 456884
rect 350446 454144 350502 454200
rect 350446 451832 350502 451888
rect 350446 449948 350502 449984
rect 350446 449928 350448 449948
rect 350448 449928 350500 449948
rect 350500 449928 350502 449948
rect 350446 447752 350502 447808
rect 350446 445576 350502 445632
rect 350446 440544 350502 440600
rect 350446 436736 350502 436792
rect 350446 434696 350502 434752
rect 350446 430652 350448 430672
rect 350448 430652 350500 430672
rect 350500 430652 350502 430672
rect 350446 430616 350502 430652
rect 350446 427896 350502 427952
rect 350446 426536 350502 426592
rect 350446 425312 350502 425368
rect 350446 422340 350502 422376
rect 350446 422320 350448 422340
rect 350448 422320 350500 422340
rect 350500 422320 350502 422340
rect 350446 420980 350502 421016
rect 350446 420960 350448 420980
rect 350448 420960 350500 420980
rect 350500 420960 350502 420980
rect 350446 419620 350502 419656
rect 350446 419600 350448 419620
rect 350448 419600 350500 419620
rect 350500 419600 350502 419620
rect 350446 418376 350502 418432
rect 350446 416880 350502 416936
rect 350446 414160 350502 414216
rect 350446 411324 350502 411360
rect 350446 411304 350448 411324
rect 350448 411304 350500 411324
rect 350500 411304 350502 411324
rect 350446 404388 350502 404424
rect 350446 404368 350448 404388
rect 350448 404368 350500 404388
rect 350500 404368 350502 404388
rect 350446 400288 350502 400344
rect 350446 399472 350502 399528
rect 350446 397568 350502 397624
rect 350446 396752 350502 396808
rect 350446 394612 350448 394632
rect 350448 394612 350500 394632
rect 350500 394612 350502 394632
rect 350446 394576 350502 394612
rect 350446 392264 350502 392320
rect 350446 389816 350502 389872
rect 350446 387812 350448 387832
rect 350448 387812 350500 387832
rect 350500 387812 350502 387832
rect 350446 387776 350502 387812
rect 350446 385056 350502 385112
rect 350354 334076 350410 334112
rect 350354 334056 350356 334076
rect 350356 334056 350408 334076
rect 350408 334056 350410 334076
rect 350354 332696 350410 332752
rect 350354 329860 350410 329896
rect 350354 329840 350356 329860
rect 350356 329840 350408 329860
rect 350408 329840 350410 329860
rect 350354 328888 350410 328944
rect 350354 325760 350410 325816
rect 350262 324536 350318 324592
rect 350354 321680 350410 321736
rect 350354 320592 350410 320648
rect 350354 319232 350410 319288
rect 350262 319096 350318 319152
rect 350354 317736 350410 317792
rect 350262 315152 350318 315208
rect 350354 315016 350410 315072
rect 350354 312296 350410 312352
rect 350354 308352 350410 308408
rect 350446 304272 350502 304328
rect 350446 302912 350502 302968
rect 350446 301008 350502 301064
rect 350446 300192 350502 300248
rect 350446 298832 350502 298888
rect 350446 296676 350502 296712
rect 350446 296656 350448 296676
rect 350448 296656 350500 296676
rect 350500 296656 350502 296676
rect 350446 295332 350448 295352
rect 350448 295332 350500 295352
rect 350500 295332 350502 295352
rect 350446 295296 350502 295332
rect 350446 293972 350448 293992
rect 350448 293972 350500 293992
rect 350500 293972 350502 293992
rect 350446 293936 350502 293972
rect 350446 288768 350502 288824
rect 350446 287156 350502 287192
rect 350446 287136 350448 287156
rect 350448 287136 350500 287156
rect 350500 287136 350502 287156
rect 350446 285776 350502 285832
rect 350354 285096 350410 285152
rect 350446 277480 350502 277536
rect 350446 275576 350502 275632
rect 350354 273808 350410 273864
rect 350446 273400 350502 273456
rect 350446 270136 350502 270192
rect 350446 268096 350502 268152
rect 350446 266736 350502 266792
rect 350446 263880 350502 263936
rect 350446 261296 350502 261352
rect 350446 258712 350502 258768
rect 350354 255992 350410 256048
rect 351366 560496 351422 560552
rect 351182 379752 351238 379808
rect 351090 365336 351146 365392
rect 351090 364520 351146 364576
rect 350998 342216 351054 342272
rect 350998 338136 351054 338192
rect 350722 279656 350778 279712
rect 350722 275984 350778 276040
rect 350630 262656 350686 262712
rect 350446 255332 350502 255368
rect 350446 255312 350448 255332
rect 350448 255312 350500 255332
rect 350500 255312 350502 255332
rect 350446 253972 350502 254008
rect 350446 253952 350448 253972
rect 350448 253952 350500 253972
rect 350500 253952 350502 253972
rect 350446 250144 350502 250200
rect 350446 248784 350502 248840
rect 350446 245928 350502 245984
rect 350538 244432 350594 244488
rect 350446 244316 350502 244352
rect 350446 244296 350448 244316
rect 350448 244296 350500 244316
rect 350500 244296 350502 244316
rect 350446 243208 350502 243264
rect 350446 239264 350502 239320
rect 350446 238856 350502 238912
rect 350446 236136 350502 236192
rect 350446 235048 350502 235104
rect 350446 232192 350502 232248
rect 350446 230560 350502 230616
rect 350446 229200 350502 229256
rect 350446 222536 350502 222592
rect 350446 221196 350502 221232
rect 350446 221176 350448 221196
rect 350448 221176 350500 221196
rect 350500 221176 350502 221196
rect 350446 218068 350502 218104
rect 350446 218048 350448 218068
rect 350448 218048 350500 218068
rect 350500 218048 350502 218068
rect 350446 217504 350502 217560
rect 350354 217096 350410 217152
rect 350446 215348 350502 215384
rect 350446 215328 350448 215348
rect 350448 215328 350500 215348
rect 350500 215328 350502 215348
rect 350446 213152 350502 213208
rect 350446 209908 350502 209944
rect 350446 209888 350448 209908
rect 350448 209888 350500 209908
rect 350500 209888 350502 209908
rect 350446 209072 350502 209128
rect 350446 207712 350502 207768
rect 350354 207304 350410 207360
rect 350446 206932 350448 206952
rect 350448 206932 350500 206952
rect 350500 206932 350502 206952
rect 350446 206896 350502 206932
rect 350354 204992 350410 205048
rect 350446 204212 350448 204232
rect 350448 204212 350500 204232
rect 350500 204212 350502 204232
rect 350446 204176 350502 204212
rect 350446 203224 350502 203280
rect 350446 201864 350502 201920
rect 349986 195472 350042 195528
rect 350814 272176 350870 272232
rect 351366 200368 351422 200424
rect 352654 214512 352710 214568
rect 353942 487192 353998 487248
rect 356702 562400 356758 562456
rect 356702 204856 356758 204912
rect 356978 199824 357034 199880
rect 358266 564712 358322 564768
rect 358542 237904 358598 237960
rect 358266 158344 358322 158400
rect 359462 562128 359518 562184
rect 359462 156848 359518 156904
rect 360382 563080 360438 563136
rect 360382 264968 360438 265024
rect 361762 560632 361818 560688
rect 360198 152224 360254 152280
rect 363878 240080 363934 240136
rect 364246 262928 364302 262984
rect 364706 184864 364762 184920
rect 363602 159568 363658 159624
rect 365994 562264 366050 562320
rect 365902 561856 365958 561912
rect 366086 180512 366142 180568
rect 366362 156712 366418 156768
rect 366546 190984 366602 191040
rect 366454 155896 366510 155952
rect 368570 185816 368626 185872
rect 369306 198872 369362 198928
rect 369490 181600 369546 181656
rect 365718 151408 365774 151464
rect 370594 153040 370650 153096
rect 373354 176160 373410 176216
rect 372342 167728 372398 167784
rect 375286 239944 375342 240000
rect 376206 563760 376262 563816
rect 376206 240488 376262 240544
rect 376850 158208 376906 158264
rect 377402 190304 377458 190360
rect 377034 181464 377090 181520
rect 377494 158208 377550 158264
rect 377586 155760 377642 155816
rect 379058 237224 379114 237280
rect 380346 563488 380402 563544
rect 380162 176296 380218 176352
rect 381818 237088 381874 237144
rect 382278 183640 382334 183696
rect 383106 229880 383162 229936
rect 384946 232600 385002 232656
rect 383014 174664 383070 174720
rect 384578 156576 384634 156632
rect 385774 563352 385830 563408
rect 385498 158480 385554 158536
rect 385958 230016 386014 230072
rect 386142 230152 386198 230208
rect 386326 236544 386382 236600
rect 386418 177656 386474 177712
rect 387246 238584 387302 238640
rect 387154 167728 387210 167784
rect 387706 239808 387762 239864
rect 388258 235184 388314 235240
rect 388626 562672 388682 562728
rect 388626 162288 388682 162344
rect 388442 162152 388498 162208
rect 388902 238040 388958 238096
rect 388994 150048 389050 150104
rect 389822 174800 389878 174856
rect 390466 232872 390522 232928
rect 393134 242256 393190 242312
rect 393226 238176 393282 238232
rect 394146 178608 394202 178664
rect 396630 233960 396686 234016
rect 396170 177384 396226 177440
rect 391846 151408 391902 151464
rect 397182 233824 397238 233880
rect 397090 174528 397146 174584
rect 398286 564576 398342 564632
rect 398286 152904 398342 152960
rect 399482 238720 399538 238776
rect 399942 150048 399998 150104
rect 402426 590280 402482 590336
rect 402610 587288 402666 587344
rect 402426 559952 402482 560008
rect 402794 234232 402850 234288
rect 404910 589872 404966 589928
rect 405186 590144 405242 590200
rect 405370 590008 405426 590064
rect 404174 165144 404230 165200
rect 406658 461080 406714 461136
rect 406382 437960 406438 438016
rect 406106 242392 406162 242448
rect 406658 433200 406714 433256
rect 406474 383016 406530 383072
rect 406750 377440 406806 377496
rect 406934 679632 406990 679688
rect 407118 678000 407174 678056
rect 407026 677592 407082 677648
rect 407118 670520 407174 670576
rect 407118 669160 407174 669216
rect 407118 667800 407174 667856
rect 407118 666440 407174 666496
rect 407118 663740 407174 663776
rect 407118 663720 407120 663740
rect 407120 663720 407172 663740
rect 407172 663720 407174 663740
rect 407210 662360 407266 662416
rect 407118 661680 407174 661736
rect 407118 654880 407174 654936
rect 407118 654200 407174 654256
rect 407118 652840 407174 652896
rect 407118 652160 407174 652216
rect 407302 650120 407358 650176
rect 407578 650120 407634 650176
rect 407210 649440 407266 649496
rect 407118 648760 407174 648816
rect 407118 644680 407174 644736
rect 407394 645360 407450 645416
rect 407210 644000 407266 644056
rect 407302 642096 407358 642152
rect 407210 641960 407266 642016
rect 407210 641280 407266 641336
rect 407486 638016 407542 638072
rect 407210 637200 407266 637256
rect 407210 633800 407266 633856
rect 407210 632440 407266 632496
rect 407210 631760 407266 631816
rect 407210 629040 407266 629096
rect 407394 625640 407450 625696
rect 407210 622920 407266 622976
rect 407210 618840 407266 618896
rect 407302 616800 407358 616856
rect 407302 614896 407358 614952
rect 407210 612756 407212 612776
rect 407212 612756 407264 612776
rect 407264 612756 407266 612776
rect 407210 612720 407266 612756
rect 407210 608660 407266 608696
rect 407210 608640 407212 608660
rect 407212 608640 407264 608660
rect 407264 608640 407266 608660
rect 407210 607280 407266 607336
rect 407670 614760 407726 614816
rect 407118 525680 407174 525736
rect 407118 522280 407174 522336
rect 407118 517556 407120 517576
rect 407120 517556 407172 517576
rect 407172 517556 407174 517576
rect 407118 517520 407174 517556
rect 407118 516196 407120 516216
rect 407120 516196 407172 516216
rect 407172 516196 407174 516216
rect 407118 516160 407174 516196
rect 407118 512760 407174 512816
rect 407118 512080 407174 512136
rect 407118 509360 407174 509416
rect 407118 500520 407174 500576
rect 407118 497120 407174 497176
rect 407118 495760 407174 495816
rect 407118 493040 407174 493096
rect 407118 491000 407174 491056
rect 407118 488960 407174 489016
rect 407118 487600 407174 487656
rect 407118 486920 407174 486976
rect 407026 485560 407082 485616
rect 407118 484880 407174 484936
rect 407118 484200 407174 484256
rect 407026 483520 407082 483576
rect 406934 478080 406990 478136
rect 406842 372000 406898 372056
rect 406842 356360 406898 356416
rect 406750 345208 406806 345264
rect 407118 482160 407174 482216
rect 407118 480120 407174 480176
rect 407118 475360 407174 475416
rect 407118 474000 407174 474056
rect 407118 469920 407174 469976
rect 407118 468152 407174 468208
rect 407118 465840 407174 465896
rect 407118 463800 407174 463856
rect 407118 462460 407174 462496
rect 407118 462440 407120 462460
rect 407120 462440 407172 462460
rect 407172 462440 407174 462460
rect 407118 461760 407174 461816
rect 407118 459040 407174 459096
rect 407118 457000 407174 457056
rect 407118 454280 407174 454336
rect 407118 453600 407174 453656
rect 407118 451308 407174 451344
rect 407118 451288 407120 451308
rect 407120 451288 407172 451308
rect 407172 451288 407174 451308
rect 407118 449520 407174 449576
rect 407118 446120 407174 446176
rect 407118 444760 407174 444816
rect 407118 442040 407174 442096
rect 407118 440000 407174 440056
rect 407118 437280 407174 437336
rect 407118 435920 407174 435976
rect 407670 602520 407726 602576
rect 407302 601840 407358 601896
rect 407762 601160 407818 601216
rect 407302 599120 407358 599176
rect 407302 597080 407358 597136
rect 407302 595040 407358 595096
rect 407302 593000 407358 593056
rect 407302 591096 407358 591152
rect 407302 588920 407358 588976
rect 407762 587152 407818 587208
rect 407302 586880 407358 586936
rect 407946 605920 408002 605976
rect 407946 594360 408002 594416
rect 407946 586200 408002 586256
rect 407670 585520 407726 585576
rect 407302 580080 407358 580136
rect 407302 577360 407358 577416
rect 407394 576680 407450 576736
rect 407302 572600 407358 572656
rect 407302 569880 407358 569936
rect 408038 573960 408094 574016
rect 407670 573280 407726 573336
rect 407394 567840 407450 567896
rect 407394 564460 407450 564496
rect 407394 564440 407396 564460
rect 407396 564440 407448 564460
rect 407448 564440 407450 564460
rect 407394 561040 407450 561096
rect 407670 556960 407726 557016
rect 407394 556280 407450 556336
rect 407486 552880 407542 552936
rect 407394 551520 407450 551576
rect 407394 550840 407450 550896
rect 407394 550160 407450 550216
rect 407486 548800 407542 548856
rect 407394 547440 407450 547496
rect 407394 544720 407450 544776
rect 407486 544040 407542 544096
rect 407394 542000 407450 542056
rect 407302 535200 407358 535256
rect 407302 533840 407358 533896
rect 407302 531800 407358 531856
rect 407302 525000 407358 525056
rect 407302 523640 407358 523696
rect 407394 522960 407450 523016
rect 407302 518200 407358 518256
rect 407302 516840 407358 516896
rect 407578 514800 407634 514856
rect 408038 559000 408094 559056
rect 407946 555600 408002 555656
rect 407762 508000 407818 508056
rect 407302 489640 407358 489696
rect 407302 476040 407358 476096
rect 407302 474680 407358 474736
rect 407302 467880 407358 467936
rect 407302 463120 407358 463176
rect 407302 455640 407358 455696
rect 407670 454960 407726 455016
rect 407302 447208 407358 447264
rect 407302 441360 407358 441416
rect 407486 438640 407542 438696
rect 407210 434560 407266 434616
rect 407118 429800 407174 429856
rect 407118 429120 407174 429176
rect 407210 427760 407266 427816
rect 407118 427080 407174 427136
rect 407946 425720 408002 425776
rect 407118 423700 407174 423736
rect 407118 423680 407120 423700
rect 407120 423680 407172 423700
rect 407172 423680 407174 423700
rect 407118 423000 407174 423056
rect 407854 421640 407910 421696
rect 407210 420280 407266 420336
rect 407118 419600 407174 419656
rect 407118 418920 407174 418976
rect 407118 416200 407174 416256
rect 407118 414840 407174 414896
rect 407118 411440 407174 411496
rect 407118 410760 407174 410816
rect 407118 408720 407174 408776
rect 407118 406000 407174 406056
rect 407210 404640 407266 404696
rect 407762 401920 407818 401976
rect 407486 400288 407542 400344
rect 407118 399200 407174 399256
rect 407118 397840 407174 397896
rect 407210 395800 407266 395856
rect 407118 395120 407174 395176
rect 407118 393760 407174 393816
rect 407578 393080 407634 393136
rect 407210 391720 407266 391776
rect 407118 391040 407174 391096
rect 407118 389680 407174 389736
rect 407118 385600 407174 385656
rect 407118 384920 407174 384976
rect 407118 382880 407174 382936
rect 407118 381520 407174 381576
rect 407118 378800 407174 378856
rect 407118 373360 407174 373416
rect 407118 370640 407174 370696
rect 407118 361120 407174 361176
rect 407118 360440 407174 360496
rect 407118 357040 407174 357096
rect 407118 353640 407174 353696
rect 407210 352960 407266 353016
rect 407118 352280 407174 352336
rect 407118 351600 407174 351656
rect 407118 349172 407174 349208
rect 407118 349152 407120 349172
rect 407120 349152 407172 349172
rect 407172 349152 407174 349172
rect 407118 346840 407174 346896
rect 407118 344800 407174 344856
rect 407118 343440 407174 343496
rect 407118 340720 407174 340776
rect 407118 339360 407174 339416
rect 407118 336676 407120 336696
rect 407120 336676 407172 336696
rect 407172 336676 407174 336696
rect 407118 336640 407174 336676
rect 407394 332560 407450 332616
rect 407118 330520 407174 330576
rect 407118 328500 407174 328536
rect 407118 328480 407120 328500
rect 407120 328480 407172 328500
rect 407172 328480 407174 328500
rect 407118 327800 407174 327856
rect 407118 325760 407174 325816
rect 407210 325080 407266 325136
rect 407210 323720 407266 323776
rect 407118 323040 407174 323096
rect 407210 322360 407266 322416
rect 407118 321680 407174 321736
rect 407302 321000 407358 321056
rect 407118 315560 407174 315616
rect 407210 311072 407266 311128
rect 407118 310800 407174 310856
rect 407118 310120 407174 310176
rect 407118 308080 407174 308136
rect 407118 306720 407174 306776
rect 407118 305360 407174 305416
rect 407118 304000 407174 304056
rect 407210 301960 407266 302016
rect 407118 301280 407174 301336
rect 407118 299920 407174 299976
rect 407118 295840 407174 295896
rect 407210 293800 407266 293856
rect 407118 292476 407120 292496
rect 407120 292476 407172 292496
rect 407172 292476 407174 292496
rect 407118 292440 407174 292476
rect 407210 291760 407266 291816
rect 407118 289720 407174 289776
rect 407302 289040 407358 289096
rect 407210 288360 407266 288416
rect 407118 287680 407174 287736
rect 407118 287000 407174 287056
rect 407118 284316 407120 284336
rect 407120 284316 407172 284336
rect 407172 284316 407174 284336
rect 407118 284280 407174 284316
rect 407210 283600 407266 283656
rect 407118 282940 407174 282976
rect 407118 282920 407120 282940
rect 407120 282920 407172 282940
rect 407172 282920 407174 282940
rect 407210 279520 407266 279576
rect 407118 278860 407174 278896
rect 407118 278840 407120 278860
rect 407120 278840 407172 278860
rect 407172 278840 407174 278860
rect 407118 276120 407174 276176
rect 407118 275440 407174 275496
rect 407118 271360 407174 271416
rect 407118 270000 407174 270056
rect 407118 267960 407174 268016
rect 407118 263880 407174 263936
rect 407118 262520 407174 262576
rect 407118 261840 407174 261896
rect 407118 259800 407174 259856
rect 407210 257760 407266 257816
rect 407118 257080 407174 257136
rect 407118 255040 407174 255096
rect 407118 251640 407174 251696
rect 407118 250960 407174 251016
rect 407210 250280 407266 250336
rect 407210 246880 407266 246936
rect 407118 246200 407174 246256
rect 407118 244840 407174 244896
rect 407118 242120 407174 242176
rect 407486 300600 407542 300656
rect 407578 298560 407634 298616
rect 408222 678272 408278 678328
rect 408866 680040 408922 680096
rect 408406 667120 408462 667176
rect 408314 565120 408370 565176
rect 408314 546080 408370 546136
rect 408314 501200 408370 501256
rect 408222 466520 408278 466576
rect 408222 466384 408278 466440
rect 408130 457680 408186 457736
rect 408130 433880 408186 433936
rect 408130 374040 408186 374096
rect 408038 362480 408094 362536
rect 408130 335280 408186 335336
rect 408038 312840 408094 312896
rect 407946 302640 408002 302696
rect 407854 276800 407910 276856
rect 407762 267280 407818 267336
rect 407486 254360 407542 254416
rect 407762 249600 407818 249656
rect 407578 242936 407634 242992
rect 408958 578040 409014 578096
rect 445114 685208 445170 685264
rect 409142 570560 409198 570616
rect 409050 510040 409106 510096
rect 408406 318960 408462 319016
rect 408406 293936 408462 293992
rect 408406 259936 408462 259992
rect 409234 479440 409290 479496
rect 409326 476720 409382 476776
rect 409234 471960 409290 472016
rect 409602 459720 409658 459776
rect 409602 452920 409658 452976
rect 409510 430480 409566 430536
rect 409418 428440 409474 428496
rect 409510 412120 409566 412176
rect 409142 284960 409198 285016
rect 408958 245556 408960 245576
rect 408960 245556 409012 245576
rect 409012 245556 409014 245576
rect 408958 245520 409014 245556
rect 408406 239808 408462 239864
rect 409050 152360 409106 152416
rect 409418 318280 409474 318336
rect 409510 241168 409566 241224
rect 409510 240760 409566 240816
rect 416134 684936 416190 684992
rect 409694 364520 409750 364576
rect 409694 342760 409750 342816
rect 413558 683440 413614 683496
rect 412914 681944 412970 682000
rect 411626 680312 411682 680368
rect 425794 684800 425850 684856
rect 423862 683712 423918 683768
rect 419998 679904 420054 679960
rect 428370 681808 428426 681864
rect 433522 679904 433578 679960
rect 442538 684528 442594 684584
rect 447690 682352 447746 682408
rect 446862 681128 446918 681184
rect 453854 684528 453910 684584
rect 454774 685072 454830 685128
rect 462502 682216 462558 682272
rect 480534 683576 480590 683632
rect 487618 685208 487674 685264
rect 489550 685072 489606 685128
rect 488722 680992 488778 681048
rect 495162 680448 495218 680504
rect 504270 687248 504326 687304
rect 502522 683304 502578 683360
rect 500498 682080 500554 682136
rect 509514 683168 509570 683224
rect 505098 680856 505154 680912
rect 511446 680856 511502 680912
rect 514758 681264 514814 681320
rect 518990 680720 519046 680776
rect 526258 682352 526314 682408
rect 528742 682216 528798 682272
rect 530122 682488 530178 682544
rect 531226 682080 531282 682136
rect 532698 681400 532754 681456
rect 545578 684664 545634 684720
rect 545118 682624 545174 682680
rect 546866 681944 546922 682000
rect 548798 681808 548854 681864
rect 409878 665080 409934 665136
rect 550178 564440 550234 564496
rect 550178 459720 550234 459776
rect 550086 378800 550142 378856
rect 409786 334600 409842 334656
rect 409878 319640 409934 319696
rect 409786 316920 409842 316976
rect 550086 297880 550142 297936
rect 410338 240352 410394 240408
rect 410246 230288 410302 230344
rect 412730 198328 412786 198384
rect 412730 195336 412786 195392
rect 422298 198464 422354 198520
rect 427082 187040 427138 187096
rect 440606 155624 440662 155680
rect 447690 153040 447746 153096
rect 452842 195200 452898 195256
rect 453486 192616 453542 192672
rect 458178 238448 458234 238504
rect 458178 185680 458234 185736
rect 460570 184320 460626 184376
rect 463790 152904 463846 152960
rect 482466 152768 482522 152824
rect 488906 167592 488962 167648
rect 488538 155488 488594 155544
rect 490194 164872 490250 164928
rect 492770 180240 492826 180296
rect 497278 182824 497334 182880
rect 498566 152632 498622 152688
rect 502430 162016 502486 162072
rect 509238 238720 509294 238776
rect 520186 238312 520242 238368
rect 525614 238448 525670 238504
rect 523038 206216 523094 206272
rect 531318 193160 531374 193216
rect 537482 239400 537538 239456
rect 537574 237904 537630 237960
rect 540242 234232 540298 234288
rect 537942 158616 537998 158672
rect 538862 150320 538918 150376
rect 539782 173168 539838 173224
rect 539230 150184 539286 150240
rect 59634 110608 59690 110664
rect 58622 17312 58678 17368
rect 539966 46824 540022 46880
rect 59910 30504 59966 30560
rect 59910 29824 59966 29880
rect 61290 29552 61346 29608
rect 59910 29144 59966 29200
rect 66442 29824 66498 29880
rect 67638 28192 67694 28248
rect 69570 28192 69626 28248
rect 65798 27512 65854 27568
rect 65154 27376 65210 27432
rect 50158 3440 50214 3496
rect 64326 4800 64382 4856
rect 60830 3440 60886 3496
rect 71778 27512 71834 27568
rect 71594 26696 71650 26752
rect 71778 26696 71834 26752
rect 70398 25880 70454 25936
rect 72882 27512 72938 27568
rect 74538 25744 74594 25800
rect 82818 29688 82874 29744
rect 85762 27240 85818 27296
rect 74630 21936 74686 21992
rect 77390 24384 77446 24440
rect 85578 25608 85634 25664
rect 84198 17856 84254 17912
rect 88338 25472 88394 25528
rect 91190 24792 91246 24848
rect 99286 28056 99342 28112
rect 99378 19896 99434 19952
rect 95422 18944 95478 19000
rect 106278 18536 106334 18592
rect 107750 23160 107806 23216
rect 107934 23160 107990 23216
rect 117962 28872 118018 28928
rect 124218 22616 124274 22672
rect 113178 18672 113234 18728
rect 106370 17720 106426 17776
rect 92478 15816 92534 15872
rect 103334 3304 103390 3360
rect 125690 21528 125746 21584
rect 128358 21256 128414 21312
rect 126978 3304 127034 3360
rect 139398 20032 139454 20088
rect 136638 17176 136694 17232
rect 146390 21392 146446 21448
rect 164238 24112 164294 24168
rect 153198 17448 153254 17504
rect 166906 28328 166962 28384
rect 165618 23704 165674 23760
rect 173990 28600 174046 28656
rect 175278 27920 175334 27976
rect 182362 29144 182418 29200
rect 188802 28464 188858 28520
rect 186226 28192 186282 28248
rect 178038 22616 178094 22672
rect 168378 19080 168434 19136
rect 144734 15952 144790 16008
rect 150622 3440 150678 3496
rect 155406 4936 155462 4992
rect 157798 3576 157854 3632
rect 169574 3712 169630 3768
rect 178130 17584 178186 17640
rect 184938 25472 184994 25528
rect 183558 21528 183614 21584
rect 180798 17040 180854 17096
rect 182546 3168 182602 3224
rect 207110 24248 207166 24304
rect 207018 21664 207074 21720
rect 203430 14864 203486 14920
rect 197910 3984 197966 4040
rect 200302 3848 200358 3904
rect 205086 10240 205142 10296
rect 212630 17448 212686 17504
rect 208582 12960 208638 13016
rect 214470 14592 214526 14648
rect 218058 11600 218114 11656
rect 224958 24384 225014 24440
rect 222198 17312 222254 17368
rect 231858 25608 231914 25664
rect 222750 11736 222806 11792
rect 226338 14728 226394 14784
rect 234526 28464 234582 28520
rect 231950 13640 232006 13696
rect 255318 24656 255374 24712
rect 260838 18944 260894 19000
rect 242990 16496 243046 16552
rect 242898 11872 242954 11928
rect 240506 6296 240562 6352
rect 251178 15000 251234 15056
rect 284114 29416 284170 29472
rect 274638 24656 274694 24712
rect 278778 18808 278834 18864
rect 276018 10920 276074 10976
rect 282918 17312 282974 17368
rect 289818 19080 289874 19136
rect 300858 29280 300914 29336
rect 304998 24520 305054 24576
rect 303618 23976 303674 24032
rect 310518 20032 310574 20088
rect 303894 13096 303950 13152
rect 314382 29280 314438 29336
rect 318890 22888 318946 22944
rect 318798 21800 318854 21856
rect 321558 23840 321614 23896
rect 324318 20168 324374 20224
rect 333702 28328 333758 28384
rect 329838 18400 329894 18456
rect 335358 18400 335414 18456
rect 328734 12008 328790 12064
rect 347870 23976 347926 24032
rect 354770 25880 354826 25936
rect 359462 28192 359518 28248
rect 358818 22888 358874 22944
rect 367190 26016 367246 26072
rect 373630 26968 373686 27024
rect 369122 26832 369178 26888
rect 367098 19216 367154 19272
rect 385222 27104 385278 27160
rect 378230 26016 378286 26072
rect 378414 16088 378470 16144
rect 385038 25744 385094 25800
rect 391938 22752 391994 22808
rect 416134 29008 416190 29064
rect 408498 23024 408554 23080
rect 421930 27104 421986 27160
rect 431958 16360 432014 16416
rect 436098 20304 436154 20360
rect 444470 23024 444526 23080
rect 445850 19760 445906 19816
rect 446034 19624 446090 19680
rect 452842 26968 452898 27024
rect 459650 21120 459706 21176
rect 463790 21800 463846 21856
rect 468942 23296 468998 23352
rect 479246 28736 479302 28792
rect 481822 29008 481878 29064
rect 476118 21664 476174 21720
rect 480258 26152 480314 26208
rect 487618 28736 487674 28792
rect 484582 25336 484638 25392
rect 491298 22480 491354 22536
rect 484398 21120 484454 21176
rect 474554 6568 474610 6624
rect 481730 6432 481786 6488
rect 519174 29416 519230 29472
rect 521106 29552 521162 29608
rect 518898 23296 518954 23352
rect 525614 27512 525670 27568
rect 524326 26560 524382 26616
rect 527178 28464 527234 28520
rect 525798 20440 525854 20496
rect 528834 28464 528890 28520
rect 536562 27920 536618 27976
rect 532054 27240 532110 27296
rect 528558 21936 528614 21992
rect 531318 3848 531374 3904
rect 539506 29824 539562 29880
rect 539506 28872 539562 28928
rect 538310 20576 538366 20632
rect 540150 149776 540206 149832
rect 540242 149096 540298 149152
rect 540150 147328 540206 147384
rect 540426 149232 540482 149288
rect 540426 147600 540482 147656
rect 540334 147192 540390 147248
rect 540334 146920 540390 146976
rect 540334 139576 540390 139632
rect 540610 150048 540666 150104
rect 540150 122712 540206 122768
rect 540150 114144 540206 114200
rect 540978 150184 541034 150240
rect 540978 139440 541034 139496
rect 540794 135088 540850 135144
rect 540886 129784 540942 129840
rect 540426 86808 540482 86864
rect 540610 89936 540666 89992
rect 540886 31592 540942 31648
rect 541254 235456 541310 235512
rect 541254 151680 541310 151736
rect 541530 147872 541586 147928
rect 541438 133456 541494 133512
rect 541346 101496 541402 101552
rect 541254 89800 541310 89856
rect 541254 75792 541310 75848
rect 541990 138080 542046 138136
rect 541714 30504 541770 30560
rect 542542 144744 542598 144800
rect 542542 140800 542598 140856
rect 542450 95376 542506 95432
rect 542358 84496 542414 84552
rect 542358 42356 542414 42392
rect 542358 42336 542360 42356
rect 542360 42336 542412 42356
rect 542412 42336 542414 42356
rect 542358 37576 542414 37632
rect 542358 26696 542414 26752
rect 542634 107616 542690 107672
rect 544014 238040 544070 238096
rect 543094 147736 543150 147792
rect 542818 129920 542874 129976
rect 542726 74976 542782 75032
rect 542818 65456 542874 65512
rect 543002 145696 543058 145752
rect 543554 146376 543610 146432
rect 543094 142976 543150 143032
rect 543186 142296 543242 142352
rect 543186 141652 543188 141672
rect 543188 141652 543240 141672
rect 543240 141652 543242 141672
rect 543186 141616 543242 141652
rect 543094 127608 543150 127664
rect 543646 140936 543702 140992
rect 543922 144744 543978 144800
rect 544474 239264 544530 239320
rect 543554 138216 543610 138272
rect 543830 137264 543886 137320
rect 543554 136176 543610 136232
rect 543646 135496 543702 135552
rect 543554 134136 543610 134192
rect 543554 131416 543610 131472
rect 543554 130736 543610 130792
rect 543554 128016 543610 128072
rect 543830 125568 543886 125624
rect 543554 125296 543610 125352
rect 543554 121896 543610 121952
rect 543554 120536 543610 120592
rect 543554 116456 543610 116512
rect 543554 115812 543556 115832
rect 543556 115812 543608 115832
rect 543608 115812 543610 115832
rect 543554 115776 543610 115812
rect 543554 114452 543556 114472
rect 543556 114452 543608 114472
rect 543608 114452 543610 114472
rect 543554 114416 543610 114452
rect 543646 113736 543702 113792
rect 543554 110372 543556 110392
rect 543556 110372 543608 110392
rect 543608 110372 543610 110392
rect 543554 110336 543610 110372
rect 543278 106256 543334 106312
rect 543554 97416 543610 97472
rect 543554 96056 543610 96112
rect 543554 94016 543610 94072
rect 543554 91976 543610 92032
rect 543554 88576 543610 88632
rect 543554 83816 543610 83872
rect 543554 82456 543610 82512
rect 543554 78376 543610 78432
rect 543646 77696 543702 77752
rect 543554 76336 543610 76392
rect 543554 75656 543610 75712
rect 543554 71576 543610 71632
rect 543554 70216 543610 70272
rect 543554 66172 543556 66192
rect 543556 66172 543608 66192
rect 543608 66172 543610 66192
rect 543554 66136 543610 66172
rect 543554 64096 543610 64152
rect 543554 62076 543610 62112
rect 543554 62056 543556 62076
rect 543556 62056 543608 62076
rect 543608 62056 543610 62076
rect 543646 60696 543702 60752
rect 543554 56616 543610 56672
rect 543554 52536 543610 52592
rect 543462 49816 543518 49872
rect 543554 48456 543610 48512
rect 543554 47776 543610 47832
rect 543554 45056 543610 45112
rect 543646 44376 543702 44432
rect 543554 43696 543610 43752
rect 543554 40976 543610 41032
rect 543554 36216 543610 36272
rect 543554 35536 543610 35592
rect 543554 30776 543610 30832
rect 546222 238448 546278 238504
rect 545486 237224 545542 237280
rect 545762 237088 545818 237144
rect 545486 236816 545542 236872
rect 544474 148824 544530 148880
rect 544106 130056 544162 130112
rect 544658 117272 544714 117328
rect 544658 110472 544714 110528
rect 544658 82864 544714 82920
rect 545026 135088 545082 135144
rect 545026 131008 545082 131064
rect 546038 230152 546094 230208
rect 546958 233960 547014 234016
rect 546222 124072 546278 124128
rect 546682 152360 546738 152416
rect 546590 141208 546646 141264
rect 546590 125432 546646 125488
rect 546498 106120 546554 106176
rect 547510 186904 547566 186960
rect 547510 128424 547566 128480
rect 547510 126112 547566 126168
rect 547326 86808 547382 86864
rect 548154 238584 548210 238640
rect 548982 237224 549038 237280
rect 547970 229880 548026 229936
rect 547878 153992 547934 154048
rect 547970 147056 548026 147112
rect 548062 146784 548118 146840
rect 547786 126928 547842 126984
rect 547970 108976 548026 109032
rect 547878 72392 547934 72448
rect 549258 237360 549314 237416
rect 548706 149912 548762 149968
rect 549442 230016 549498 230072
rect 549442 147600 549498 147656
rect 549166 118768 549222 118824
rect 549718 151000 549774 151056
rect 550638 507320 550694 507376
rect 550362 495760 550418 495816
rect 550270 431840 550326 431896
rect 550914 605920 550970 605976
rect 550822 600480 550878 600536
rect 550822 596400 550878 596456
rect 550730 271360 550786 271416
rect 550730 268640 550786 268696
rect 550270 240760 550326 240816
rect 550638 247560 550694 247616
rect 550178 149096 550234 149152
rect 549902 133864 549958 133920
rect 550914 562400 550970 562456
rect 551190 622920 551246 622976
rect 551098 555600 551154 555656
rect 551098 539280 551154 539336
rect 551006 468560 551062 468616
rect 551006 323720 551062 323776
rect 550822 232736 550878 232792
rect 549902 13640 549958 13696
rect 551190 333920 551246 333976
rect 551098 238584 551154 238640
rect 552110 678680 552166 678736
rect 552018 678000 552074 678056
rect 552018 675960 552074 676016
rect 552018 672424 552074 672480
rect 552018 661680 552074 661736
rect 552018 641960 552074 642016
rect 552018 637880 552074 637936
rect 552018 631780 552074 631816
rect 552018 631760 552020 631780
rect 552020 631760 552072 631780
rect 552072 631760 552074 631780
rect 552018 603916 552020 603936
rect 552020 603916 552072 603936
rect 552072 603916 552074 603936
rect 552018 603880 552074 603916
rect 552018 598440 552074 598496
rect 552018 590960 552074 591016
rect 552018 588956 552020 588976
rect 552020 588956 552072 588976
rect 552072 588956 552074 588976
rect 552018 588920 552074 588956
rect 552018 586880 552074 586936
rect 552018 585520 552074 585576
rect 552018 579400 552074 579456
rect 552018 578040 552074 578096
rect 552018 576000 552074 576056
rect 552018 574504 552074 574560
rect 552018 573960 552074 574016
rect 552018 553560 552074 553616
rect 552018 550860 552074 550896
rect 552018 550840 552020 550860
rect 552020 550840 552072 550860
rect 552072 550840 552074 550860
rect 552110 547440 552166 547496
rect 552110 545400 552166 545456
rect 552018 522280 552074 522336
rect 552018 521600 552074 521656
rect 552018 519424 552074 519480
rect 552018 518880 552074 518936
rect 552018 516840 552074 516896
rect 552018 514820 552074 514856
rect 552018 514800 552020 514820
rect 552020 514800 552072 514820
rect 552072 514800 552074 514820
rect 551558 484880 551614 484936
rect 551374 282240 551430 282296
rect 551098 192480 551154 192536
rect 551190 160792 551246 160848
rect 551466 147464 551522 147520
rect 552018 465840 552074 465896
rect 552018 464344 552074 464400
rect 552018 463120 552074 463176
rect 552018 460400 552074 460456
rect 552018 459060 552074 459096
rect 552018 459040 552020 459060
rect 552020 459040 552072 459060
rect 552072 459040 552074 459060
rect 552018 457680 552074 457736
rect 552018 456320 552074 456376
rect 552018 422320 552074 422376
rect 552018 371320 552074 371376
rect 552018 367956 552020 367976
rect 552020 367956 552072 367976
rect 552072 367956 552074 367976
rect 552018 367920 552074 367956
rect 552018 365220 552074 365256
rect 552018 365200 552020 365220
rect 552020 365200 552072 365220
rect 552072 365200 552074 365220
rect 552018 342796 552020 342816
rect 552020 342796 552072 342816
rect 552072 342796 552074 342816
rect 552018 342760 552074 342796
rect 552018 322380 552074 322416
rect 552018 322360 552020 322380
rect 552020 322360 552072 322380
rect 552072 322360 552074 322380
rect 552018 307436 552020 307456
rect 552020 307436 552072 307456
rect 552072 307436 552074 307456
rect 552018 307400 552074 307436
rect 552018 293140 552074 293176
rect 552018 293120 552020 293140
rect 552020 293120 552072 293140
rect 552072 293120 552074 293140
rect 552018 291780 552074 291816
rect 552018 291760 552020 291780
rect 552020 291760 552072 291780
rect 552072 291760 552074 291780
rect 552478 679360 552534 679416
rect 552478 674600 552534 674656
rect 552754 670520 552810 670576
rect 552662 654200 552718 654256
rect 552662 650120 552718 650176
rect 552570 642640 552626 642696
rect 552478 638424 552534 638480
rect 552570 634480 552626 634536
rect 552754 616120 552810 616176
rect 552478 608660 552534 608696
rect 552478 608640 552480 608660
rect 552480 608640 552532 608660
rect 552532 608640 552534 608660
rect 552478 591368 552534 591424
rect 552386 536560 552442 536616
rect 552386 532516 552388 532536
rect 552388 532516 552440 532536
rect 552440 532516 552442 532536
rect 552386 532480 552442 532516
rect 552386 530476 552388 530496
rect 552388 530476 552440 530496
rect 552440 530476 552442 530496
rect 552386 530440 552442 530476
rect 552386 526360 552442 526416
rect 552294 525680 552350 525736
rect 552570 544040 552626 544096
rect 552570 533840 552626 533896
rect 552478 524320 552534 524376
rect 552386 515480 552442 515536
rect 552294 500520 552350 500576
rect 552202 480120 552258 480176
rect 552294 454280 552350 454336
rect 552202 451424 552258 451480
rect 552294 440680 552350 440736
rect 552202 432520 552258 432576
rect 552202 429800 552258 429856
rect 552202 420996 552204 421016
rect 552204 420996 552256 421016
rect 552256 420996 552258 421016
rect 552202 420960 552258 420996
rect 552202 393780 552258 393816
rect 552202 393760 552204 393780
rect 552204 393760 552256 393780
rect 552256 393760 552258 393780
rect 552202 372700 552258 372736
rect 552202 372680 552204 372700
rect 552204 372680 552256 372700
rect 552256 372680 552258 372700
rect 552202 369280 552258 369336
rect 552202 306040 552258 306096
rect 552018 265260 552074 265296
rect 552018 265240 552020 265260
rect 552020 265240 552072 265260
rect 552072 265240 552074 265260
rect 552018 263220 552074 263256
rect 552018 263200 552020 263220
rect 552020 263200 552072 263220
rect 552072 263200 552074 263220
rect 552018 261840 552074 261896
rect 552110 260344 552166 260400
rect 552018 259800 552074 259856
rect 552110 259120 552166 259176
rect 552018 258440 552074 258496
rect 552018 257760 552074 257816
rect 552110 255040 552166 255096
rect 552018 254360 552074 254416
rect 552018 250280 552074 250336
rect 552018 242800 552074 242856
rect 552202 246200 552258 246256
rect 552202 243344 552258 243400
rect 551650 162288 551706 162344
rect 552662 493720 552718 493776
rect 552570 492360 552626 492416
rect 552662 484200 552718 484256
rect 552570 476040 552626 476096
rect 552570 449520 552626 449576
rect 552662 448840 552718 448896
rect 552570 446800 552626 446856
rect 552570 445440 552626 445496
rect 552386 421640 552442 421696
rect 552386 412820 552442 412856
rect 552386 412800 552388 412820
rect 552388 412800 552440 412820
rect 552440 412800 552442 412820
rect 552478 407360 552534 407416
rect 552386 354320 552442 354376
rect 552570 331200 552626 331256
rect 553122 679768 553178 679824
rect 553122 665760 553178 665816
rect 553306 656940 553362 656976
rect 553306 656920 553308 656940
rect 553308 656920 553360 656940
rect 553360 656920 553362 656940
rect 553306 653520 553362 653576
rect 553306 648760 553362 648816
rect 552938 646720 552994 646776
rect 553306 645360 553362 645416
rect 552938 644700 552994 644736
rect 552938 644680 552940 644700
rect 552940 644680 552992 644700
rect 552992 644680 552994 644700
rect 553306 630400 553362 630456
rect 553306 624280 553362 624336
rect 553306 620200 553362 620256
rect 553306 617480 553362 617536
rect 553306 614760 553362 614816
rect 553306 613400 553362 613456
rect 553306 611380 553362 611416
rect 553306 611360 553308 611380
rect 553308 611360 553360 611380
rect 553360 611360 553362 611380
rect 553306 610680 553362 610736
rect 553306 607280 553362 607336
rect 553306 603200 553362 603256
rect 552846 597760 552902 597816
rect 553214 584840 553270 584896
rect 553122 568520 553178 568576
rect 553122 561040 553178 561096
rect 552938 558320 552994 558376
rect 553122 540640 553178 540696
rect 553122 493040 553178 493096
rect 552846 453600 552902 453656
rect 553030 438640 553086 438696
rect 553030 437280 553086 437336
rect 553030 428440 553086 428496
rect 553030 426436 553032 426456
rect 553032 426436 553084 426456
rect 553084 426436 553086 426456
rect 553030 426400 553086 426436
rect 553030 425076 553032 425096
rect 553032 425076 553084 425096
rect 553084 425076 553086 425096
rect 553030 425040 553086 425076
rect 552938 424360 552994 424416
rect 553030 423716 553032 423736
rect 553032 423716 553084 423736
rect 553084 423716 553086 423736
rect 553030 423680 553086 423716
rect 553030 420280 553086 420336
rect 553030 416200 553086 416256
rect 553030 415520 553086 415576
rect 553030 413344 553086 413400
rect 553030 410760 553086 410816
rect 553030 405320 553086 405376
rect 553030 403960 553086 404016
rect 553030 403280 553086 403336
rect 553030 400424 553086 400480
rect 553030 395120 553086 395176
rect 553030 391720 553086 391776
rect 553030 390360 553086 390416
rect 553030 388320 553086 388376
rect 553030 387640 553086 387696
rect 553030 385600 553086 385656
rect 553030 381540 553086 381576
rect 553030 381520 553032 381540
rect 553032 381520 553084 381540
rect 553084 381520 553086 381540
rect 553030 378120 553086 378176
rect 553030 377440 553086 377496
rect 553030 370640 553086 370696
rect 553030 368600 553086 368656
rect 552938 366424 552994 366480
rect 553030 365880 553086 365936
rect 552938 361120 552994 361176
rect 553030 360460 553086 360496
rect 553030 360440 553032 360460
rect 553032 360440 553084 360460
rect 553084 360440 553086 360460
rect 552938 358400 552994 358456
rect 553030 357720 553086 357776
rect 553030 355680 553086 355736
rect 553030 353640 553086 353696
rect 552846 351600 552902 351656
rect 553122 350940 553178 350976
rect 553122 350920 553124 350940
rect 553124 350920 553176 350940
rect 553176 350920 553178 350940
rect 553122 349424 553178 349480
rect 553030 347520 553086 347576
rect 553122 346840 553178 346896
rect 553030 343440 553086 343496
rect 552938 340040 552994 340096
rect 553122 338680 553178 338736
rect 553030 335960 553086 336016
rect 553122 335300 553178 335336
rect 553122 335280 553124 335300
rect 553124 335280 553176 335300
rect 553176 335280 553178 335300
rect 552846 334600 552902 334656
rect 553030 327800 553086 327856
rect 553122 327140 553178 327176
rect 553122 327120 553124 327140
rect 553124 327120 553176 327140
rect 553176 327120 553178 327140
rect 553030 326440 553086 326496
rect 553122 325760 553178 325816
rect 553030 318280 553086 318336
rect 553122 317600 553178 317656
rect 553122 316240 553178 316296
rect 553122 314880 553178 314936
rect 553030 314200 553086 314256
rect 553122 312840 553178 312896
rect 553030 311344 553086 311400
rect 553122 310800 553178 310856
rect 553122 310120 553178 310176
rect 553122 308760 553178 308816
rect 553122 305360 553178 305416
rect 553030 301960 553086 302016
rect 553122 301280 553178 301336
rect 553122 300600 553178 300656
rect 553122 297200 553178 297256
rect 553122 292440 553178 292496
rect 553122 290400 553178 290456
rect 553030 289720 553086 289776
rect 553122 289040 553178 289096
rect 553122 287680 553178 287736
rect 553122 283620 553178 283656
rect 553122 283600 553124 283620
rect 553124 283600 553176 283620
rect 553176 283600 553178 283620
rect 553122 281560 553178 281616
rect 553030 280880 553086 280936
rect 553122 280236 553124 280256
rect 553124 280236 553176 280256
rect 553176 280236 553178 280256
rect 553122 280200 553178 280236
rect 553122 279520 553178 279576
rect 553122 278860 553178 278896
rect 553122 278840 553124 278860
rect 553124 278840 553176 278860
rect 553176 278840 553178 278860
rect 553122 277480 553178 277536
rect 553030 276140 553086 276176
rect 553030 276120 553032 276140
rect 553032 276120 553084 276140
rect 553084 276120 553086 276140
rect 553122 274760 553178 274816
rect 553122 273400 553178 273456
rect 553122 270680 553178 270736
rect 552846 264560 552902 264616
rect 553122 266600 553178 266656
rect 553122 263880 553178 263936
rect 552754 200912 552810 200968
rect 549074 3984 549130 4040
rect 553122 253680 553178 253736
rect 553122 252320 553178 252376
rect 553122 248240 553178 248296
rect 553122 246880 553178 246936
rect 553122 244840 553178 244896
rect 553030 236816 553086 236872
rect 553306 567840 553362 567896
rect 553306 565120 553362 565176
rect 553306 560380 553362 560416
rect 553306 560360 553308 560380
rect 553308 560360 553360 560380
rect 553360 560360 553362 560380
rect 553306 557640 553362 557696
rect 553306 556960 553362 557016
rect 553306 556280 553362 556336
rect 553306 551520 553362 551576
rect 553306 549480 553362 549536
rect 553306 539960 553362 540016
rect 553306 535880 553362 535936
rect 553306 535200 553362 535256
rect 553306 531120 553362 531176
rect 553306 528400 553362 528456
rect 553306 510040 553362 510096
rect 553306 505280 553362 505336
rect 553306 504600 553362 504656
rect 553306 502444 553362 502480
rect 553306 502424 553308 502444
rect 553308 502424 553360 502444
rect 553360 502424 553362 502444
rect 553306 501880 553362 501936
rect 553306 501200 553362 501256
rect 553306 499860 553362 499896
rect 553306 499840 553308 499860
rect 553308 499840 553360 499860
rect 553360 499840 553362 499860
rect 553306 498500 553362 498536
rect 553306 498480 553308 498500
rect 553308 498480 553360 498500
rect 553360 498480 553362 498500
rect 553306 488960 553362 489016
rect 553306 488280 553362 488336
rect 553306 478760 553362 478816
rect 553306 475360 553362 475416
rect 553306 470620 553362 470656
rect 553306 470600 553308 470620
rect 553308 470600 553360 470620
rect 553360 470600 553362 470620
rect 553306 469920 553362 469976
rect 553306 466520 553362 466576
rect 553306 454960 553362 455016
rect 553306 450200 553362 450256
rect 553306 443400 553362 443456
rect 553306 437960 553362 438016
rect 553306 436600 553362 436656
rect 553214 232464 553270 232520
rect 553490 496440 553546 496496
rect 553490 391040 553546 391096
rect 553306 159296 553362 159352
rect 552846 115096 552902 115152
rect 553582 363840 553638 363896
rect 553582 340720 553638 340776
rect 553582 25472 553638 25528
rect 554042 293120 554098 293176
rect 554226 149232 554282 149288
rect 555238 162424 555294 162480
rect 555054 12960 555110 13016
rect 556526 26152 556582 26208
rect 556894 235320 556950 235376
rect 556986 134408 557042 134464
rect 556894 112376 556950 112432
rect 557078 126248 557134 126304
rect 557630 13096 557686 13152
rect 558274 88984 558330 89040
rect 559378 28192 559434 28248
rect 560390 239808 560446 239864
rect 560758 198736 560814 198792
rect 564622 682080 564678 682136
rect 560298 20848 560354 20904
rect 561770 239264 561826 239320
rect 562046 190032 562102 190088
rect 562598 28328 562654 28384
rect 563610 193976 563666 194032
rect 563702 189624 563758 189680
rect 563610 156576 563666 156632
rect 563794 150184 563850 150240
rect 564622 197376 564678 197432
rect 564530 29416 564586 29472
rect 564714 124072 564770 124128
rect 564990 240488 565046 240544
rect 565082 239536 565138 239592
rect 565818 239672 565874 239728
rect 579158 697176 579214 697232
rect 565450 29008 565506 29064
rect 566554 184184 566610 184240
rect 566370 165008 566426 165064
rect 566830 193840 566886 193896
rect 569406 681808 569462 681864
rect 569498 150320 569554 150376
rect 569958 20868 570014 20904
rect 569958 20848 569960 20868
rect 569960 20848 570012 20868
rect 570012 20848 570014 20868
rect 570234 3440 570290 3496
rect 571614 239400 571670 239456
rect 571430 20732 571486 20768
rect 571430 20712 571432 20732
rect 571432 20712 571484 20732
rect 571484 20712 571486 20732
rect 571338 3984 571394 4040
rect 572074 240080 572130 240136
rect 571982 156712 572038 156768
rect 573086 233824 573142 233880
rect 572258 17856 572314 17912
rect 573362 159432 573418 159488
rect 573270 155080 573326 155136
rect 573362 20304 573418 20360
rect 574834 236952 574890 237008
rect 575938 27512 575994 27568
rect 576950 680856 577006 680912
rect 577042 26016 577098 26072
rect 577226 177248 577282 177304
rect 577226 162152 577282 162208
rect 578790 239944 578846 240000
rect 578238 23996 578294 24032
rect 578238 23976 578240 23996
rect 578240 23976 578292 23996
rect 578292 23976 578294 23996
rect 578882 19760 578938 19816
rect 579066 258848 579122 258904
rect 580170 630808 580226 630864
rect 580170 524456 580226 524512
rect 580170 471416 580226 471472
rect 579894 431568 579950 431624
rect 579802 33108 579858 33144
rect 579802 33088 579804 33108
rect 579804 33088 579856 33108
rect 579856 33088 579858 33108
rect 580170 378392 580226 378448
rect 580170 325216 580226 325272
rect 580170 272176 580226 272232
rect 580170 232328 580226 232384
rect 580078 179152 580134 179208
rect 579618 25880 579674 25936
rect 580630 680584 580686 680640
rect 580906 670656 580962 670712
rect 580906 644000 580962 644056
rect 580814 617480 580870 617536
rect 580722 590960 580778 591016
rect 580630 577632 580686 577688
rect 580538 564304 580594 564360
rect 580446 537784 580502 537840
rect 580354 484608 580410 484664
rect 580354 418240 580410 418296
rect 580446 365064 580502 365120
rect 580446 312024 580502 312080
rect 580262 219000 580318 219056
rect 580262 192480 580318 192536
rect 580262 99456 580318 99512
rect 580262 72936 580318 72992
rect 580262 59608 580318 59664
rect 580446 152632 580502 152688
rect 580446 139340 580448 139360
rect 580448 139340 580500 139360
rect 580500 139340 580502 139360
rect 580446 139304 580502 139340
rect 580446 112784 580502 112840
rect 581550 229744 581606 229800
rect 582562 30912 582618 30968
rect 583114 28056 583170 28112
<< metal3 >>
rect 24301 700362 24367 700365
rect 566038 700362 566044 700364
rect 24301 700360 566044 700362
rect 24301 700304 24306 700360
rect 24362 700304 566044 700360
rect 24301 700302 566044 700304
rect 24301 700299 24367 700302
rect 566038 700300 566044 700302
rect 566108 700300 566114 700364
rect -960 697220 480 697460
rect 579153 697234 579219 697237
rect 583520 697234 584960 697324
rect 579153 697232 584960 697234
rect 579153 697176 579158 697232
rect 579214 697176 584960 697232
rect 579153 697174 584960 697176
rect 579153 697171 579219 697174
rect 583520 697084 584960 697174
rect 359406 687244 359412 687308
rect 359476 687306 359482 687308
rect 504265 687306 504331 687309
rect 359476 687304 504331 687306
rect 359476 687248 504270 687304
rect 504326 687248 504331 687304
rect 359476 687246 504331 687248
rect 359476 687244 359482 687246
rect 504265 687243 504331 687246
rect 28206 685884 28212 685948
rect 28276 685946 28282 685948
rect 552054 685946 552060 685948
rect 28276 685886 552060 685946
rect 28276 685884 28282 685886
rect 552054 685884 552060 685886
rect 552124 685884 552130 685948
rect 382774 685204 382780 685268
rect 382844 685266 382850 685268
rect 445109 685266 445175 685269
rect 382844 685264 445175 685266
rect 382844 685208 445114 685264
rect 445170 685208 445175 685264
rect 382844 685206 445175 685208
rect 382844 685204 382850 685206
rect 445109 685203 445175 685206
rect 487613 685266 487679 685269
rect 575422 685266 575428 685268
rect 487613 685264 575428 685266
rect 487613 685208 487618 685264
rect 487674 685208 575428 685264
rect 487613 685206 575428 685208
rect 487613 685203 487679 685206
rect 575422 685204 575428 685206
rect 575492 685204 575498 685268
rect 355174 685068 355180 685132
rect 355244 685130 355250 685132
rect 454769 685130 454835 685133
rect 355244 685128 454835 685130
rect 355244 685072 454774 685128
rect 454830 685072 454835 685128
rect 355244 685070 454835 685072
rect 355244 685068 355250 685070
rect 454769 685067 454835 685070
rect 489545 685130 489611 685133
rect 579654 685130 579660 685132
rect 489545 685128 579660 685130
rect 489545 685072 489550 685128
rect 489606 685072 579660 685128
rect 489545 685070 579660 685072
rect 489545 685067 489611 685070
rect 579654 685068 579660 685070
rect 579724 685068 579730 685132
rect 416129 684994 416195 684997
rect 551686 684994 551692 684996
rect 416129 684992 551692 684994
rect 416129 684936 416134 684992
rect 416190 684936 551692 684992
rect 416129 684934 551692 684936
rect 416129 684931 416195 684934
rect 551686 684932 551692 684934
rect 551756 684932 551762 684996
rect 425789 684858 425855 684861
rect 569902 684858 569908 684860
rect 425789 684856 569908 684858
rect 425789 684800 425794 684856
rect 425850 684800 569908 684856
rect 425789 684798 569908 684800
rect 425789 684795 425855 684798
rect 569902 684796 569908 684798
rect 569972 684796 569978 684860
rect 361430 684660 361436 684724
rect 361500 684722 361506 684724
rect 545573 684722 545639 684725
rect 361500 684720 545639 684722
rect 361500 684664 545578 684720
rect 545634 684664 545639 684720
rect 361500 684662 545639 684664
rect 361500 684660 361506 684662
rect 545573 684659 545639 684662
rect 25446 684524 25452 684588
rect 25516 684586 25522 684588
rect 442533 684586 442599 684589
rect 25516 684584 442599 684586
rect 25516 684528 442538 684584
rect 442594 684528 442599 684584
rect 25516 684526 442599 684528
rect 25516 684524 25522 684526
rect 442533 684523 442599 684526
rect 453849 684586 453915 684589
rect 551502 684586 551508 684588
rect 453849 684584 551508 684586
rect 453849 684528 453854 684584
rect 453910 684528 551508 684584
rect 453849 684526 551508 684528
rect 453849 684523 453915 684526
rect 551502 684524 551508 684526
rect 551572 684524 551578 684588
rect -960 684164 480 684404
rect 409822 683844 409828 683908
rect 409892 683906 409898 683908
rect 583520 683906 584960 683996
rect 409892 683846 584960 683906
rect 409892 683844 409898 683846
rect 393078 683708 393084 683772
rect 393148 683770 393154 683772
rect 423857 683770 423923 683773
rect 393148 683768 423923 683770
rect 393148 683712 423862 683768
rect 423918 683712 423923 683768
rect 583520 683756 584960 683846
rect 393148 683710 423923 683712
rect 393148 683708 393154 683710
rect 423857 683707 423923 683710
rect 402094 683572 402100 683636
rect 402164 683634 402170 683636
rect 480529 683634 480595 683637
rect 402164 683632 480595 683634
rect 402164 683576 480534 683632
rect 480590 683576 480595 683632
rect 402164 683574 480595 683576
rect 402164 683572 402170 683574
rect 480529 683571 480595 683574
rect 375046 683436 375052 683500
rect 375116 683498 375122 683500
rect 413553 683498 413619 683501
rect 375116 683496 413619 683498
rect 375116 683440 413558 683496
rect 413614 683440 413619 683496
rect 375116 683438 413619 683440
rect 375116 683436 375122 683438
rect 413553 683435 413619 683438
rect 21357 683362 21423 683365
rect 502517 683362 502583 683365
rect 21357 683360 502583 683362
rect 21357 683304 21362 683360
rect 21418 683304 502522 683360
rect 502578 683304 502583 683360
rect 21357 683302 502583 683304
rect 21357 683299 21423 683302
rect 502517 683299 502583 683302
rect 26877 683226 26943 683229
rect 509509 683226 509575 683229
rect 26877 683224 509575 683226
rect 26877 683168 26882 683224
rect 26938 683168 509514 683224
rect 509570 683168 509575 683224
rect 26877 683166 509575 683168
rect 26877 683163 26943 683166
rect 509509 683163 509575 683166
rect 400806 682620 400812 682684
rect 400876 682682 400882 682684
rect 545113 682682 545179 682685
rect 400876 682680 545179 682682
rect 400876 682624 545118 682680
rect 545174 682624 545179 682680
rect 400876 682622 545179 682624
rect 400876 682620 400882 682622
rect 545113 682619 545179 682622
rect 371734 682484 371740 682548
rect 371804 682546 371810 682548
rect 530117 682546 530183 682549
rect 371804 682544 530183 682546
rect 371804 682488 530122 682544
rect 530178 682488 530183 682544
rect 371804 682486 530183 682488
rect 371804 682484 371810 682486
rect 530117 682483 530183 682486
rect 400990 682348 400996 682412
rect 401060 682410 401066 682412
rect 447685 682410 447751 682413
rect 401060 682408 447751 682410
rect 401060 682352 447690 682408
rect 447746 682352 447751 682408
rect 401060 682350 447751 682352
rect 401060 682348 401066 682350
rect 447685 682347 447751 682350
rect 526253 682410 526319 682413
rect 566958 682410 566964 682412
rect 526253 682408 566964 682410
rect 526253 682352 526258 682408
rect 526314 682352 566964 682408
rect 526253 682350 566964 682352
rect 526253 682347 526319 682350
rect 566958 682348 566964 682350
rect 567028 682348 567034 682412
rect 383510 682212 383516 682276
rect 383580 682274 383586 682276
rect 462497 682274 462563 682277
rect 383580 682272 462563 682274
rect 383580 682216 462502 682272
rect 462558 682216 462563 682272
rect 383580 682214 462563 682216
rect 383580 682212 383586 682214
rect 462497 682211 462563 682214
rect 528737 682274 528803 682277
rect 560518 682274 560524 682276
rect 528737 682272 560524 682274
rect 528737 682216 528742 682272
rect 528798 682216 560524 682272
rect 528737 682214 560524 682216
rect 528737 682211 528803 682214
rect 560518 682212 560524 682214
rect 560588 682212 560594 682276
rect 356646 682076 356652 682140
rect 356716 682138 356722 682140
rect 500493 682138 500559 682141
rect 356716 682136 500559 682138
rect 356716 682080 500498 682136
rect 500554 682080 500559 682136
rect 356716 682078 500559 682080
rect 356716 682076 356722 682078
rect 500493 682075 500559 682078
rect 531221 682138 531287 682141
rect 564617 682138 564683 682141
rect 531221 682136 564683 682138
rect 531221 682080 531226 682136
rect 531282 682080 564622 682136
rect 564678 682080 564683 682136
rect 531221 682078 564683 682080
rect 531221 682075 531287 682078
rect 564617 682075 564683 682078
rect 389766 681940 389772 682004
rect 389836 682002 389842 682004
rect 412909 682002 412975 682005
rect 389836 682000 412975 682002
rect 389836 681944 412914 682000
rect 412970 681944 412975 682000
rect 389836 681942 412975 681944
rect 389836 681940 389842 681942
rect 412909 681939 412975 681942
rect 546861 682002 546927 682005
rect 574134 682002 574140 682004
rect 546861 682000 574140 682002
rect 546861 681944 546866 682000
rect 546922 681944 574140 682000
rect 546861 681942 574140 681944
rect 546861 681939 546927 681942
rect 574134 681940 574140 681942
rect 574204 681940 574210 682004
rect 406510 681804 406516 681868
rect 406580 681866 406586 681868
rect 428365 681866 428431 681869
rect 406580 681864 428431 681866
rect 406580 681808 428370 681864
rect 428426 681808 428431 681864
rect 406580 681806 428431 681808
rect 406580 681804 406586 681806
rect 428365 681803 428431 681806
rect 548793 681866 548859 681869
rect 569401 681866 569467 681869
rect 548793 681864 569467 681866
rect 548793 681808 548798 681864
rect 548854 681808 569406 681864
rect 569462 681808 569467 681864
rect 548793 681806 569467 681808
rect 548793 681803 548859 681806
rect 569401 681803 569467 681806
rect 24669 681458 24735 681461
rect 532693 681458 532759 681461
rect 24669 681456 532759 681458
rect 24669 681400 24674 681456
rect 24730 681400 532698 681456
rect 532754 681400 532759 681456
rect 24669 681398 532759 681400
rect 24669 681395 24735 681398
rect 532693 681395 532759 681398
rect 171777 681322 171843 681325
rect 514753 681322 514819 681325
rect 171777 681320 514819 681322
rect 171777 681264 171782 681320
rect 171838 681264 514758 681320
rect 514814 681264 514819 681320
rect 171777 681262 514819 681264
rect 171777 681259 171843 681262
rect 514753 681259 514819 681262
rect 446857 681186 446923 681189
rect 570086 681186 570092 681188
rect 446857 681184 570092 681186
rect 446857 681128 446862 681184
rect 446918 681128 570092 681184
rect 446857 681126 570092 681128
rect 446857 681123 446923 681126
rect 570086 681124 570092 681126
rect 570156 681124 570162 681188
rect 363454 680988 363460 681052
rect 363524 681050 363530 681052
rect 488717 681050 488783 681053
rect 363524 681048 488783 681050
rect 363524 680992 488722 681048
rect 488778 680992 488783 681048
rect 363524 680990 488783 680992
rect 363524 680988 363530 680990
rect 488717 680987 488783 680990
rect 368974 680852 368980 680916
rect 369044 680914 369050 680916
rect 505093 680914 505159 680917
rect 369044 680912 505159 680914
rect 369044 680856 505098 680912
rect 505154 680856 505159 680912
rect 369044 680854 505159 680856
rect 369044 680852 369050 680854
rect 505093 680851 505159 680854
rect 511441 680914 511507 680917
rect 576945 680914 577011 680917
rect 511441 680912 577011 680914
rect 511441 680856 511446 680912
rect 511502 680856 576950 680912
rect 577006 680856 577011 680912
rect 511441 680854 577011 680856
rect 511441 680851 511507 680854
rect 576945 680851 577011 680854
rect 370630 680716 370636 680780
rect 370700 680778 370706 680780
rect 518985 680778 519051 680781
rect 370700 680776 519051 680778
rect 370700 680720 518990 680776
rect 519046 680720 519051 680776
rect 370700 680718 519051 680720
rect 370700 680716 370706 680718
rect 518985 680715 519051 680718
rect 410006 680580 410012 680644
rect 410076 680642 410082 680644
rect 580625 680642 580691 680645
rect 410076 680640 580691 680642
rect 410076 680584 580630 680640
rect 580686 680584 580691 680640
rect 410076 680582 580691 680584
rect 410076 680580 410082 680582
rect 580625 680579 580691 680582
rect 495157 680506 495223 680509
rect 578550 680506 578556 680508
rect 495157 680504 578556 680506
rect 495157 680448 495162 680504
rect 495218 680448 578556 680504
rect 495157 680446 578556 680448
rect 495157 680443 495223 680446
rect 578550 680444 578556 680446
rect 578620 680444 578626 680508
rect 403566 680308 403572 680372
rect 403636 680370 403642 680372
rect 411621 680370 411687 680373
rect 403636 680368 411687 680370
rect 403636 680312 411626 680368
rect 411682 680312 411687 680368
rect 403636 680310 411687 680312
rect 403636 680308 403642 680310
rect 411621 680307 411687 680310
rect 408861 680098 408927 680101
rect 408861 680096 425070 680098
rect 408861 680040 408866 680096
rect 408922 680040 425070 680096
rect 408861 680038 425070 680040
rect 408861 680035 408927 680038
rect 388294 679900 388300 679964
rect 388364 679962 388370 679964
rect 419993 679962 420059 679965
rect 388364 679960 420059 679962
rect 388364 679904 419998 679960
rect 420054 679904 420059 679960
rect 388364 679902 420059 679904
rect 425010 679962 425070 680038
rect 433517 679962 433583 679965
rect 425010 679960 433583 679962
rect 425010 679904 433522 679960
rect 433578 679904 433583 679960
rect 425010 679902 433583 679904
rect 388364 679900 388370 679902
rect 419993 679899 420059 679902
rect 433517 679899 433583 679902
rect 409638 679764 409644 679828
rect 409708 679826 409714 679828
rect 553117 679826 553183 679829
rect 409708 679824 553183 679826
rect 409708 679768 553122 679824
rect 553178 679768 553183 679824
rect 409708 679766 553183 679768
rect 409708 679764 409714 679766
rect 553117 679763 553183 679766
rect 406929 679690 406995 679693
rect 552422 679690 552428 679692
rect 406929 679688 552428 679690
rect 406929 679632 406934 679688
rect 406990 679632 552428 679688
rect 406929 679630 552428 679632
rect 406929 679627 406995 679630
rect 552422 679628 552428 679630
rect 552492 679628 552498 679692
rect 565118 679554 565124 679556
rect 410566 679494 565124 679554
rect 410566 679388 410626 679494
rect 565118 679492 565124 679494
rect 565188 679492 565194 679556
rect 552473 679418 552539 679421
rect 549884 679416 552539 679418
rect 549884 679360 552478 679416
rect 552534 679360 552539 679416
rect 549884 679358 552539 679360
rect 552473 679355 552539 679358
rect 552105 678738 552171 678741
rect 549884 678736 552171 678738
rect 549884 678680 552110 678736
rect 552166 678680 552171 678736
rect 549884 678678 552171 678680
rect 552105 678675 552171 678678
rect 408217 678330 408283 678333
rect 409822 678330 409828 678332
rect 408217 678328 409828 678330
rect 408217 678272 408222 678328
rect 408278 678272 409828 678328
rect 408217 678270 409828 678272
rect 408217 678267 408283 678270
rect 409822 678268 409828 678270
rect 409892 678268 409898 678332
rect 164918 678132 164924 678196
rect 164988 678194 164994 678196
rect 165521 678194 165587 678197
rect 164988 678192 165587 678194
rect 164988 678136 165526 678192
rect 165582 678136 165587 678192
rect 164988 678134 165587 678136
rect 164988 678132 164994 678134
rect 165521 678131 165587 678134
rect 407113 678058 407179 678061
rect 552013 678058 552079 678061
rect 407113 678056 410044 678058
rect 407113 678000 407118 678056
rect 407174 678000 410044 678056
rect 407113 677998 410044 678000
rect 549884 678056 552079 678058
rect 549884 678000 552018 678056
rect 552074 678000 552079 678056
rect 549884 677998 552079 678000
rect 407113 677995 407179 677998
rect 552013 677995 552079 677998
rect 153694 677724 153700 677788
rect 153764 677786 153770 677788
rect 346894 677786 346900 677788
rect 153764 677726 346900 677786
rect 153764 677724 153770 677726
rect 346894 677724 346900 677726
rect 346964 677724 346970 677788
rect 152406 677588 152412 677652
rect 152476 677650 152482 677652
rect 153101 677650 153167 677653
rect 152476 677648 153167 677650
rect 152476 677592 153106 677648
rect 153162 677592 153167 677648
rect 152476 677590 153167 677592
rect 152476 677588 152482 677590
rect 153101 677587 153167 677590
rect 324446 677588 324452 677652
rect 324516 677650 324522 677652
rect 325049 677650 325115 677653
rect 324516 677648 325115 677650
rect 324516 677592 325054 677648
rect 325110 677592 325115 677648
rect 324516 677590 325115 677592
rect 324516 677588 324522 677590
rect 325049 677587 325115 677590
rect 336774 677588 336780 677652
rect 336844 677650 336850 677652
rect 337561 677650 337627 677653
rect 336844 677648 337627 677650
rect 336844 677592 337566 677648
rect 337622 677592 337627 677648
rect 336844 677590 337627 677592
rect 336844 677588 336850 677590
rect 337561 677587 337627 677590
rect 407021 677650 407087 677653
rect 409822 677650 409828 677652
rect 407021 677648 409828 677650
rect 407021 677592 407026 677648
rect 407082 677592 409828 677648
rect 407021 677590 409828 677592
rect 407021 677587 407087 677590
rect 409822 677588 409828 677590
rect 409892 677588 409898 677652
rect 325785 677108 325851 677109
rect 325734 677044 325740 677108
rect 325804 677106 325851 677108
rect 325804 677104 325896 677106
rect 325846 677048 325896 677104
rect 325804 677046 325896 677048
rect 325804 677044 325851 677046
rect 325785 677043 325851 677044
rect 552013 676018 552079 676021
rect 549884 676016 552079 676018
rect 549884 675960 552018 676016
rect 552074 675960 552079 676016
rect 549884 675958 552079 675960
rect 552013 675955 552079 675958
rect 552473 674658 552539 674661
rect 549884 674656 552539 674658
rect 549884 674600 552478 674656
rect 552534 674600 552539 674656
rect 549884 674598 552539 674600
rect 552473 674595 552539 674598
rect 552054 673978 552060 673980
rect 549884 673918 552060 673978
rect 552054 673916 552060 673918
rect 552124 673916 552130 673980
rect 551502 673372 551508 673436
rect 551572 673434 551578 673436
rect 552238 673434 552244 673436
rect 551572 673374 552244 673434
rect 551572 673372 551578 673374
rect 552238 673372 552244 673374
rect 552308 673372 552314 673436
rect 549884 672490 550282 672550
rect 550222 672482 550282 672490
rect 552013 672482 552079 672485
rect 550222 672480 552079 672482
rect 550222 672424 552018 672480
rect 552074 672424 552079 672480
rect 550222 672422 552079 672424
rect 552013 672419 552079 672422
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect 171225 671258 171291 671261
rect 343633 671258 343699 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect 171090 671256 171291 671258
rect 171090 671220 171230 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 170568 671200 171230 671220
rect 171286 671200 171291 671256
rect 343222 671256 343699 671258
rect 343222 671220 343638 671256
rect 170568 671198 171291 671200
rect 170568 671160 171150 671198
rect 171225 671195 171291 671198
rect 342608 671200 343638 671220
rect 343694 671200 343699 671256
rect 342608 671198 343699 671200
rect 342608 671160 343282 671198
rect 343633 671195 343699 671198
rect 580901 670714 580967 670717
rect 583520 670714 584960 670804
rect 580901 670712 584960 670714
rect 580901 670656 580906 670712
rect 580962 670656 584960 670712
rect 580901 670654 584960 670656
rect 580901 670651 580967 670654
rect 407113 670578 407179 670581
rect 552749 670578 552815 670581
rect 407113 670576 410044 670578
rect 407113 670520 407118 670576
rect 407174 670520 410044 670576
rect 407113 670518 410044 670520
rect 549884 670576 552815 670578
rect 549884 670520 552754 670576
rect 552810 670520 552815 670576
rect 583520 670564 584960 670654
rect 549884 670518 552815 670520
rect 407113 670515 407179 670518
rect 552749 670515 552815 670518
rect 580942 669898 580948 669900
rect 549884 669838 580948 669898
rect 580942 669836 580948 669838
rect 581012 669836 581018 669900
rect 407113 669218 407179 669221
rect 407113 669216 410044 669218
rect 407113 669160 407118 669216
rect 407174 669160 410044 669216
rect 407113 669158 410044 669160
rect 407113 669155 407179 669158
rect 557574 668538 557580 668540
rect 549884 668478 557580 668538
rect 557574 668476 557580 668478
rect 557644 668476 557650 668540
rect 407113 667858 407179 667861
rect 563094 667858 563100 667860
rect 407113 667856 410044 667858
rect 407113 667800 407118 667856
rect 407174 667800 410044 667856
rect 407113 667798 410044 667800
rect 549884 667798 563100 667858
rect 407113 667795 407179 667798
rect 563094 667796 563100 667798
rect 563164 667796 563170 667860
rect 408401 667178 408467 667181
rect 408401 667176 410044 667178
rect 408401 667120 408406 667176
rect 408462 667120 410044 667176
rect 408401 667118 410044 667120
rect 408401 667115 408467 667118
rect 407113 666498 407179 666501
rect 570270 666498 570276 666500
rect 407113 666496 410044 666498
rect 407113 666440 407118 666496
rect 407174 666440 410044 666496
rect 407113 666438 410044 666440
rect 549884 666438 570276 666498
rect 407113 666435 407179 666438
rect 570270 666436 570276 666438
rect 570340 666436 570346 666500
rect 553117 665818 553183 665821
rect 549884 665816 553183 665818
rect 549884 665760 553122 665816
rect 553178 665760 553183 665816
rect 549884 665758 553183 665760
rect 553117 665755 553183 665758
rect 409873 665138 409939 665141
rect 409873 665136 410044 665138
rect 409873 665080 409878 665136
rect 409934 665080 410044 665136
rect 409873 665078 410044 665080
rect 409873 665075 409939 665078
rect 407113 663778 407179 663781
rect 565302 663778 565308 663780
rect 407113 663776 410044 663778
rect 407113 663720 407118 663776
rect 407174 663720 410044 663776
rect 407113 663718 410044 663720
rect 549884 663718 565308 663778
rect 407113 663715 407179 663718
rect 565302 663716 565308 663718
rect 565372 663716 565378 663780
rect 407205 662418 407271 662421
rect 407205 662416 410044 662418
rect 407205 662360 407210 662416
rect 407266 662360 410044 662416
rect 407205 662358 410044 662360
rect 407205 662355 407271 662358
rect 407113 661738 407179 661741
rect 552013 661738 552079 661741
rect 407113 661736 410044 661738
rect 407113 661680 407118 661736
rect 407174 661680 410044 661736
rect 407113 661678 410044 661680
rect 549884 661736 552079 661738
rect 549884 661680 552018 661736
rect 552074 661680 552079 661736
rect 549884 661678 552079 661680
rect 407113 661675 407179 661678
rect 552013 661675 552079 661678
rect 391054 660996 391060 661060
rect 391124 661058 391130 661060
rect 391124 660998 410044 661058
rect 391124 660996 391130 660998
rect 405590 658956 405596 659020
rect 405660 659018 405666 659020
rect 405660 658958 410044 659018
rect 405660 658956 405666 658958
rect -960 658202 480 658292
rect 3601 658202 3667 658205
rect -960 658200 3667 658202
rect -960 658144 3606 658200
rect 3662 658144 3667 658200
rect -960 658142 3667 658144
rect -960 658052 480 658142
rect 3601 658139 3667 658142
rect 377254 657596 377260 657660
rect 377324 657658 377330 657660
rect 377324 657598 410044 657658
rect 377324 657596 377330 657598
rect 583520 657236 584960 657476
rect 553301 656978 553367 656981
rect 549884 656976 553367 656978
rect 549884 656920 553306 656976
rect 553362 656920 553367 656976
rect 549884 656918 553367 656920
rect 553301 656915 553367 656918
rect 407113 654938 407179 654941
rect 407113 654936 410044 654938
rect 407113 654880 407118 654936
rect 407174 654880 410044 654936
rect 407113 654878 410044 654880
rect 407113 654875 407179 654878
rect 407113 654258 407179 654261
rect 552657 654258 552723 654261
rect 407113 654256 410044 654258
rect 407113 654200 407118 654256
rect 407174 654200 410044 654256
rect 407113 654198 410044 654200
rect 549884 654256 552723 654258
rect 549884 654200 552662 654256
rect 552718 654200 552723 654256
rect 549884 654198 552723 654200
rect 407113 654195 407179 654198
rect 552657 654195 552723 654198
rect 553301 653578 553367 653581
rect 549884 653576 553367 653578
rect 549884 653520 553306 653576
rect 553362 653520 553367 653576
rect 549884 653518 553367 653520
rect 553301 653515 553367 653518
rect 407113 652898 407179 652901
rect 407113 652896 410044 652898
rect 407113 652840 407118 652896
rect 407174 652840 410044 652896
rect 407113 652838 410044 652840
rect 407113 652835 407179 652838
rect 407113 652218 407179 652221
rect 407113 652216 410044 652218
rect 407113 652160 407118 652216
rect 407174 652160 410044 652216
rect 407113 652158 410044 652160
rect 407113 652155 407179 652158
rect 561622 650858 561628 650860
rect 549884 650798 561628 650858
rect 561622 650796 561628 650798
rect 561692 650796 561698 650860
rect 407297 650178 407363 650181
rect 407573 650178 407639 650181
rect 552657 650178 552723 650181
rect 407297 650176 410044 650178
rect 407297 650120 407302 650176
rect 407358 650120 407578 650176
rect 407634 650120 410044 650176
rect 407297 650118 410044 650120
rect 549884 650176 552723 650178
rect 549884 650120 552662 650176
rect 552718 650120 552723 650176
rect 549884 650118 552723 650120
rect 407297 650115 407363 650118
rect 407573 650115 407639 650118
rect 552657 650115 552723 650118
rect 407205 649498 407271 649501
rect 558862 649498 558868 649500
rect 407205 649496 410044 649498
rect 407205 649440 407210 649496
rect 407266 649440 410044 649496
rect 407205 649438 410044 649440
rect 549884 649438 558868 649498
rect 407205 649435 407271 649438
rect 558862 649436 558868 649438
rect 558932 649436 558938 649500
rect 407113 648818 407179 648821
rect 553301 648818 553367 648821
rect 407113 648816 410044 648818
rect 407113 648760 407118 648816
rect 407174 648760 410044 648816
rect 407113 648758 410044 648760
rect 549884 648816 553367 648818
rect 549884 648760 553306 648816
rect 553362 648760 553367 648816
rect 549884 648758 553367 648760
rect 407113 648755 407179 648758
rect 553301 648755 553367 648758
rect 408350 646716 408356 646780
rect 408420 646778 408426 646780
rect 552933 646778 552999 646781
rect 408420 646718 410044 646778
rect 549884 646776 552999 646778
rect 549884 646720 552938 646776
rect 552994 646720 552999 646776
rect 549884 646718 552999 646720
rect 408420 646716 408426 646718
rect 552933 646715 552999 646718
rect 578734 646098 578740 646100
rect 549884 646038 578740 646098
rect 578734 646036 578740 646038
rect 578804 646036 578810 646100
rect 407389 645418 407455 645421
rect 553301 645418 553367 645421
rect 407389 645416 410044 645418
rect 407389 645360 407394 645416
rect 407450 645360 410044 645416
rect 407389 645358 410044 645360
rect 549884 645416 553367 645418
rect 549884 645360 553306 645416
rect 553362 645360 553367 645416
rect 549884 645358 553367 645360
rect 407389 645355 407455 645358
rect 553301 645355 553367 645358
rect -960 644996 480 645236
rect 407113 644738 407179 644741
rect 552933 644738 552999 644741
rect 407113 644736 410044 644738
rect 407113 644680 407118 644736
rect 407174 644680 410044 644736
rect 407113 644678 410044 644680
rect 549884 644736 552999 644738
rect 549884 644680 552938 644736
rect 552994 644680 552999 644736
rect 549884 644678 552999 644680
rect 407113 644675 407179 644678
rect 552933 644675 552999 644678
rect 407205 644058 407271 644061
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 407205 644056 410044 644058
rect 407205 644000 407210 644056
rect 407266 644000 410044 644056
rect 407205 643998 410044 644000
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 407205 643995 407271 643998
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect 552565 642698 552631 642701
rect 550222 642696 552631 642698
rect 550222 642640 552570 642696
rect 552626 642640 552631 642696
rect 550222 642638 552631 642640
rect 550222 642630 550282 642638
rect 552565 642635 552631 642638
rect 407297 642154 407363 642157
rect 410014 642154 410074 642600
rect 549884 642570 550282 642630
rect 407297 642152 410074 642154
rect 407297 642096 407302 642152
rect 407358 642096 410074 642152
rect 407297 642094 410074 642096
rect 407297 642091 407363 642094
rect 407205 642018 407271 642021
rect 552013 642018 552079 642021
rect 407205 642016 410044 642018
rect 407205 641960 407210 642016
rect 407266 641960 410044 642016
rect 407205 641958 410044 641960
rect 549884 642016 552079 642018
rect 549884 641960 552018 642016
rect 552074 641960 552079 642016
rect 549884 641958 552079 641960
rect 407205 641955 407271 641958
rect 552013 641955 552079 641958
rect 407205 641338 407271 641341
rect 552054 641338 552060 641340
rect 407205 641336 410044 641338
rect 407205 641280 407210 641336
rect 407266 641280 410044 641336
rect 407205 641278 410044 641280
rect 549884 641278 552060 641338
rect 407205 641275 407271 641278
rect 552054 641276 552060 641278
rect 552124 641276 552130 641340
rect 407481 638074 407547 638077
rect 410014 638074 410074 638520
rect 549884 638490 550466 638550
rect 550406 638482 550466 638490
rect 552473 638482 552539 638485
rect 550406 638480 552539 638482
rect 550406 638424 552478 638480
rect 552534 638424 552539 638480
rect 550406 638422 552539 638424
rect 552473 638419 552539 638422
rect 407481 638072 410074 638074
rect 407481 638016 407486 638072
rect 407542 638016 410074 638072
rect 407481 638014 410074 638016
rect 407481 638011 407547 638014
rect 406326 637876 406332 637940
rect 406396 637938 406402 637940
rect 552013 637938 552079 637941
rect 406396 637878 410044 637938
rect 549884 637936 552079 637938
rect 549884 637880 552018 637936
rect 552074 637880 552079 637936
rect 549884 637878 552079 637880
rect 406396 637876 406402 637878
rect 552013 637875 552079 637878
rect 407205 637258 407271 637261
rect 407205 637256 410044 637258
rect 407205 637200 407210 637256
rect 407266 637200 410044 637256
rect 407205 637198 410044 637200
rect 407205 637195 407271 637198
rect 364926 635836 364932 635900
rect 364996 635898 365002 635900
rect 364996 635838 410044 635898
rect 364996 635836 365002 635838
rect 552565 634538 552631 634541
rect 549884 634536 552631 634538
rect 549884 634480 552570 634536
rect 552626 634480 552631 634536
rect 549884 634478 552631 634480
rect 552565 634475 552631 634478
rect 407205 633858 407271 633861
rect 557758 633858 557764 633860
rect 407205 633856 410044 633858
rect 407205 633800 407210 633856
rect 407266 633800 410044 633856
rect 407205 633798 410044 633800
rect 549884 633798 557764 633858
rect 407205 633795 407271 633798
rect 557758 633796 557764 633798
rect 557828 633796 557834 633860
rect 407205 632498 407271 632501
rect 407205 632496 410044 632498
rect 407205 632440 407210 632496
rect 407266 632440 410044 632496
rect 407205 632438 410044 632440
rect 407205 632435 407271 632438
rect -960 631940 480 632180
rect 407205 631818 407271 631821
rect 552013 631818 552079 631821
rect 407205 631816 410044 631818
rect 407205 631760 407210 631816
rect 407266 631760 410044 631816
rect 407205 631758 410044 631760
rect 549884 631816 552079 631818
rect 549884 631760 552018 631816
rect 552074 631760 552079 631816
rect 549884 631758 552079 631760
rect 407205 631755 407271 631758
rect 552013 631755 552079 631758
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 553301 630458 553367 630461
rect 549884 630456 553367 630458
rect 549884 630400 553306 630456
rect 553362 630400 553367 630456
rect 549884 630398 553367 630400
rect 553301 630395 553367 630398
rect 407205 629098 407271 629101
rect 407205 629096 410044 629098
rect 407205 629040 407210 629096
rect 407266 629040 410044 629096
rect 407205 629038 410044 629040
rect 407205 629035 407271 629038
rect 32857 628282 32923 628285
rect 34002 628282 34062 628894
rect 32857 628280 34062 628282
rect 32857 628224 32862 628280
rect 32918 628224 34062 628280
rect 32857 628222 34062 628224
rect 204161 628282 204227 628285
rect 206002 628282 206062 628894
rect 391790 628356 391796 628420
rect 391860 628418 391866 628420
rect 553342 628418 553348 628420
rect 391860 628358 410044 628418
rect 549884 628358 553348 628418
rect 391860 628356 391866 628358
rect 553342 628356 553348 628358
rect 553412 628356 553418 628420
rect 204161 628280 206062 628282
rect 204161 628224 204166 628280
rect 204222 628224 206062 628280
rect 204161 628222 206062 628224
rect 32857 628219 32923 628222
rect 204161 628219 204227 628222
rect 31569 628010 31635 628013
rect 203517 628010 203583 628013
rect 31569 628008 34062 628010
rect 31569 627952 31574 628008
rect 31630 627952 34062 628008
rect 31569 627950 34062 627952
rect 31569 627947 31635 627950
rect 34002 627942 34062 627950
rect 203517 628008 206062 628010
rect 203517 627952 203522 628008
rect 203578 627952 206062 628008
rect 203517 627950 206062 627952
rect 203517 627947 203583 627950
rect 206002 627942 206062 627950
rect 406142 627676 406148 627740
rect 406212 627738 406218 627740
rect 406212 627678 410044 627738
rect 406212 627676 406218 627678
rect 576894 627058 576900 627060
rect 549884 626998 576900 627058
rect 576894 626996 576900 626998
rect 576964 626996 576970 627060
rect 31385 625426 31451 625429
rect 34002 625426 34062 625766
rect 31385 625424 34062 625426
rect 31385 625368 31390 625424
rect 31446 625368 34062 625424
rect 31385 625366 34062 625368
rect 203609 625426 203675 625429
rect 206002 625426 206062 625766
rect 407389 625698 407455 625701
rect 407389 625696 410044 625698
rect 407389 625640 407394 625696
rect 407450 625640 410044 625696
rect 407389 625638 410044 625640
rect 407389 625635 407455 625638
rect 549884 625570 550466 625630
rect 550406 625562 550466 625570
rect 550406 625502 557550 625562
rect 203609 625424 206062 625426
rect 203609 625368 203614 625424
rect 203670 625368 206062 625424
rect 203609 625366 206062 625368
rect 31385 625363 31451 625366
rect 203609 625363 203675 625366
rect 557490 625290 557550 625502
rect 572662 625290 572668 625292
rect 557490 625230 572668 625290
rect 572662 625228 572668 625230
rect 572732 625228 572738 625292
rect 33041 624202 33107 624205
rect 34002 624202 34062 624814
rect 33041 624200 34062 624202
rect 33041 624144 33046 624200
rect 33102 624144 34062 624200
rect 33041 624142 34062 624144
rect 204069 624202 204135 624205
rect 206002 624202 206062 624814
rect 401358 624276 401364 624340
rect 401428 624338 401434 624340
rect 553301 624338 553367 624341
rect 401428 624278 410044 624338
rect 549884 624336 553367 624338
rect 549884 624280 553306 624336
rect 553362 624280 553367 624336
rect 549884 624278 553367 624280
rect 401428 624276 401434 624278
rect 553301 624275 553367 624278
rect 204069 624200 206062 624202
rect 204069 624144 204074 624200
rect 204130 624144 206062 624200
rect 204069 624142 206062 624144
rect 33041 624139 33107 624142
rect 204069 624139 204135 624142
rect 32765 622434 32831 622437
rect 34002 622434 34062 623046
rect 32765 622432 34062 622434
rect 32765 622376 32770 622432
rect 32826 622376 34062 622432
rect 32765 622374 34062 622376
rect 203977 622434 204043 622437
rect 206002 622434 206062 623046
rect 407205 622978 407271 622981
rect 551185 622978 551251 622981
rect 407205 622976 410044 622978
rect 407205 622920 407210 622976
rect 407266 622920 410044 622976
rect 407205 622918 410044 622920
rect 549884 622976 551251 622978
rect 549884 622920 551190 622976
rect 551246 622920 551251 622976
rect 549884 622918 551251 622920
rect 407205 622915 407271 622918
rect 551185 622915 551251 622918
rect 203977 622432 206062 622434
rect 203977 622376 203982 622432
rect 204038 622376 206062 622432
rect 203977 622374 206062 622376
rect 32765 622371 32831 622374
rect 203977 622371 204043 622374
rect 205541 621988 205607 621991
rect 205541 621986 206032 621988
rect 32949 621346 33015 621349
rect 34002 621346 34062 621958
rect 205541 621930 205546 621986
rect 205602 621930 206032 621986
rect 205541 621928 206032 621930
rect 205541 621925 205607 621928
rect 32949 621344 34062 621346
rect 32949 621288 32954 621344
rect 33010 621288 34062 621344
rect 32949 621286 34062 621288
rect 32949 621283 33015 621286
rect 553301 620258 553367 620261
rect 549884 620256 553367 620258
rect 549884 620200 553306 620256
rect 553362 620200 553367 620256
rect 549884 620198 553367 620200
rect 553301 620195 553367 620198
rect 31477 619714 31543 619717
rect 34002 619714 34062 620190
rect 31477 619712 34062 619714
rect 31477 619656 31482 619712
rect 31538 619656 34062 619712
rect 31477 619654 34062 619656
rect 203885 619714 203951 619717
rect 206002 619714 206062 620190
rect 203885 619712 206062 619714
rect 203885 619656 203890 619712
rect 203946 619656 206062 619712
rect 203885 619654 206062 619656
rect 31477 619651 31543 619654
rect 203885 619651 203951 619654
rect 395838 619516 395844 619580
rect 395908 619578 395914 619580
rect 395908 619518 410044 619578
rect 395908 619516 395914 619518
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 407205 618898 407271 618901
rect 407205 618896 410044 618898
rect 407205 618840 407210 618896
rect 407266 618840 410044 618896
rect 407205 618838 410044 618840
rect 407205 618835 407271 618838
rect 553301 617538 553367 617541
rect 549884 617536 553367 617538
rect 549884 617480 553306 617536
rect 553362 617480 553367 617536
rect 549884 617478 553367 617480
rect 553301 617475 553367 617478
rect 580809 617538 580875 617541
rect 583520 617538 584960 617628
rect 580809 617536 584960 617538
rect 580809 617480 580814 617536
rect 580870 617480 584960 617536
rect 580809 617478 584960 617480
rect 580809 617475 580875 617478
rect 583520 617388 584960 617478
rect 407297 616858 407363 616861
rect 407297 616856 410044 616858
rect 407297 616800 407302 616856
rect 407358 616800 410044 616856
rect 407297 616798 410044 616800
rect 407297 616795 407363 616798
rect 552749 616178 552815 616181
rect 549884 616176 552815 616178
rect 549884 616120 552754 616176
rect 552810 616120 552815 616176
rect 549884 616118 552815 616120
rect 552749 616115 552815 616118
rect 407297 614954 407363 614957
rect 410014 614954 410074 615468
rect 407297 614952 410074 614954
rect 407297 614896 407302 614952
rect 407358 614896 410074 614952
rect 407297 614894 410074 614896
rect 407297 614891 407363 614894
rect 407665 614818 407731 614821
rect 553301 614818 553367 614821
rect 407665 614816 410044 614818
rect 407665 614760 407670 614816
rect 407726 614760 410044 614816
rect 407665 614758 410044 614760
rect 549884 614816 553367 614818
rect 549884 614760 553306 614816
rect 553362 614760 553367 614816
rect 549884 614758 553367 614760
rect 407665 614755 407731 614758
rect 553301 614755 553367 614758
rect 553301 613458 553367 613461
rect 549884 613456 553367 613458
rect 549884 613400 553306 613456
rect 553362 613400 553367 613456
rect 549884 613398 553367 613400
rect 553301 613395 553367 613398
rect 407205 612778 407271 612781
rect 575606 612778 575612 612780
rect 407205 612776 410044 612778
rect 407205 612720 407210 612776
rect 407266 612720 410044 612776
rect 407205 612718 410044 612720
rect 549884 612718 575612 612778
rect 407205 612715 407271 612718
rect 575606 612716 575612 612718
rect 575676 612716 575682 612780
rect 559046 612098 559052 612100
rect 549884 612038 559052 612098
rect 559046 612036 559052 612038
rect 559116 612036 559122 612100
rect 172605 611418 172671 611421
rect 346301 611418 346367 611421
rect 171090 611416 172671 611418
rect 171090 611380 172610 611416
rect 170568 611360 172610 611380
rect 172666 611360 172671 611416
rect 343222 611416 346367 611418
rect 343222 611380 346306 611416
rect 170568 611358 172671 611360
rect 170568 611320 171150 611358
rect 172605 611355 172671 611358
rect 342608 611360 346306 611380
rect 346362 611360 346367 611416
rect 342608 611358 346367 611360
rect 342608 611320 343282 611358
rect 346301 611355 346367 611358
rect 388478 611356 388484 611420
rect 388548 611418 388554 611420
rect 553301 611418 553367 611421
rect 388548 611358 410044 611418
rect 549884 611416 553367 611418
rect 549884 611360 553306 611416
rect 553362 611360 553367 611416
rect 549884 611358 553367 611360
rect 388548 611356 388554 611358
rect 553301 611355 553367 611358
rect 553301 610738 553367 610741
rect 549884 610736 553367 610738
rect 549884 610680 553306 610736
rect 553362 610680 553367 610736
rect 549884 610678 553367 610680
rect 553301 610675 553367 610678
rect 173801 609786 173867 609789
rect 345013 609786 345079 609789
rect 171090 609784 173867 609786
rect 171090 609748 173806 609784
rect 170568 609728 173806 609748
rect 173862 609728 173867 609784
rect 343222 609784 345079 609786
rect 343222 609748 345018 609784
rect 170568 609726 173867 609728
rect 170568 609688 171150 609726
rect 173801 609723 173867 609726
rect 342608 609728 345018 609748
rect 345074 609728 345079 609784
rect 342608 609726 345079 609728
rect 342608 609688 343282 609726
rect 345013 609723 345079 609726
rect 407205 608698 407271 608701
rect 552473 608698 552539 608701
rect 407205 608696 410044 608698
rect 407205 608640 407210 608696
rect 407266 608640 410044 608696
rect 407205 608638 410044 608640
rect 550222 608696 552539 608698
rect 550222 608640 552478 608696
rect 552534 608640 552539 608696
rect 550222 608638 552539 608640
rect 407205 608635 407271 608638
rect 550222 608630 550282 608638
rect 552473 608635 552539 608638
rect 549884 608570 550282 608630
rect 173801 608426 173867 608429
rect 345105 608426 345171 608429
rect 171090 608424 173867 608426
rect 171090 608388 173806 608424
rect 170568 608368 173806 608388
rect 173862 608368 173867 608424
rect 343222 608424 345171 608426
rect 343222 608388 345110 608424
rect 170568 608366 173867 608368
rect 170568 608328 171150 608366
rect 173801 608363 173867 608366
rect 342608 608368 345110 608388
rect 345166 608368 345171 608424
rect 342608 608366 345171 608368
rect 342608 608328 343282 608366
rect 345105 608363 345171 608366
rect 556286 608018 556292 608020
rect 549884 607958 556292 608018
rect 556286 607956 556292 607958
rect 556356 607956 556362 608020
rect 407205 607338 407271 607341
rect 553301 607338 553367 607341
rect 407205 607336 410044 607338
rect 407205 607280 407210 607336
rect 407266 607280 410044 607336
rect 407205 607278 410044 607280
rect 549884 607336 553367 607338
rect 549884 607280 553306 607336
rect 553362 607280 553367 607336
rect 549884 607278 553367 607280
rect 407205 607275 407271 607278
rect 553301 607275 553367 607278
rect 172513 606930 172579 606933
rect 345565 606930 345631 606933
rect 171090 606928 172579 606930
rect 171090 606892 172518 606928
rect 170568 606872 172518 606892
rect 172574 606872 172579 606928
rect 343222 606928 345631 606930
rect 343222 606892 345570 606928
rect 170568 606870 172579 606872
rect 170568 606832 171150 606870
rect 172513 606867 172579 606870
rect 342608 606872 345570 606892
rect 345626 606872 345631 606928
rect 342608 606870 345631 606872
rect 342608 606832 343282 606870
rect 345565 606867 345631 606870
rect -960 606114 480 606204
rect 3693 606114 3759 606117
rect -960 606112 3759 606114
rect -960 606056 3698 606112
rect 3754 606056 3759 606112
rect -960 606054 3759 606056
rect -960 605964 480 606054
rect 3693 606051 3759 606054
rect 407941 605978 408007 605981
rect 550909 605978 550975 605981
rect 407941 605976 410044 605978
rect 407941 605920 407946 605976
rect 408002 605920 410044 605976
rect 407941 605918 410044 605920
rect 549884 605976 550975 605978
rect 549884 605920 550914 605976
rect 550970 605920 550975 605976
rect 549884 605918 550975 605920
rect 407941 605915 408007 605918
rect 550909 605915 550975 605918
rect 171317 605706 171383 605709
rect 345105 605706 345171 605709
rect 171090 605704 171383 605706
rect 171090 605668 171322 605704
rect 170568 605648 171322 605668
rect 171378 605648 171383 605704
rect 343222 605704 345171 605706
rect 343222 605668 345110 605704
rect 170568 605646 171383 605648
rect 170568 605608 171150 605646
rect 171317 605643 171383 605646
rect 342608 605648 345110 605668
rect 345166 605648 345171 605704
rect 342608 605646 345171 605648
rect 342608 605608 343282 605646
rect 345105 605643 345171 605646
rect 409462 604490 410044 604550
rect 387558 604420 387564 604484
rect 387628 604482 387634 604484
rect 409462 604482 409522 604490
rect 387628 604422 409522 604482
rect 387628 604420 387634 604422
rect 583520 604060 584960 604300
rect 552013 603938 552079 603941
rect 549884 603936 552079 603938
rect 549884 603880 552018 603936
rect 552074 603880 552079 603936
rect 549884 603878 552079 603880
rect 552013 603875 552079 603878
rect 553301 603258 553367 603261
rect 549884 603256 553367 603258
rect 549884 603200 553306 603256
rect 553362 603200 553367 603256
rect 549884 603198 553367 603200
rect 553301 603195 553367 603198
rect 407665 602578 407731 602581
rect 563278 602578 563284 602580
rect 407665 602576 410044 602578
rect 407665 602520 407670 602576
rect 407726 602520 410044 602576
rect 407665 602518 410044 602520
rect 549884 602518 563284 602578
rect 407665 602515 407731 602518
rect 563278 602516 563284 602518
rect 563348 602516 563354 602580
rect 31661 601762 31727 601765
rect 34002 601762 34062 601966
rect 31661 601760 34062 601762
rect 31661 601704 31666 601760
rect 31722 601704 34062 601760
rect 31661 601702 34062 601704
rect 203057 601762 203123 601765
rect 206002 601762 206062 601966
rect 407297 601898 407363 601901
rect 571374 601898 571380 601900
rect 407297 601896 410044 601898
rect 407297 601840 407302 601896
rect 407358 601840 410044 601896
rect 407297 601838 410044 601840
rect 549884 601838 571380 601898
rect 407297 601835 407363 601838
rect 571374 601836 571380 601838
rect 571444 601836 571450 601900
rect 203057 601760 206062 601762
rect 203057 601704 203062 601760
rect 203118 601704 206062 601760
rect 203057 601702 206062 601704
rect 31661 601699 31727 601702
rect 203057 601699 203123 601702
rect 407757 601218 407823 601221
rect 407757 601216 410044 601218
rect 407757 601160 407762 601216
rect 407818 601160 410044 601216
rect 407757 601158 410044 601160
rect 407757 601155 407823 601158
rect 550817 600538 550883 600541
rect 549884 600536 550883 600538
rect 549884 600480 550822 600536
rect 550878 600480 550883 600536
rect 549884 600478 550883 600480
rect 550817 600475 550883 600478
rect 32673 600402 32739 600405
rect 204897 600402 204963 600405
rect 32673 600400 34062 600402
rect 32673 600344 32678 600400
rect 32734 600344 34062 600400
rect 32673 600342 34062 600344
rect 32673 600339 32739 600342
rect 34002 600334 34062 600342
rect 204897 600400 206062 600402
rect 204897 600344 204902 600400
rect 204958 600344 206062 600400
rect 204897 600342 206062 600344
rect 204897 600339 204963 600342
rect 206002 600334 206062 600342
rect 31518 599388 31524 599452
rect 31588 599450 31594 599452
rect 34002 599450 34062 600062
rect 31588 599390 34062 599450
rect 203793 599450 203859 599453
rect 206002 599450 206062 600062
rect 560702 599858 560708 599860
rect 549884 599798 560708 599858
rect 560702 599796 560708 599798
rect 560772 599796 560778 599860
rect 203793 599448 206062 599450
rect 203793 599392 203798 599448
rect 203854 599392 206062 599448
rect 203793 599390 206062 599392
rect 31588 599388 31594 599390
rect 203793 599387 203859 599390
rect 407297 599178 407363 599181
rect 556102 599178 556108 599180
rect 407297 599176 410044 599178
rect 407297 599120 407302 599176
rect 407358 599120 410044 599176
rect 407297 599118 410044 599120
rect 549884 599118 556108 599178
rect 407297 599115 407363 599118
rect 556102 599116 556108 599118
rect 556172 599116 556178 599180
rect 378726 598436 378732 598500
rect 378796 598498 378802 598500
rect 552013 598498 552079 598501
rect 378796 598438 410044 598498
rect 549884 598496 552079 598498
rect 549884 598440 552018 598496
rect 552074 598440 552079 598496
rect 549884 598438 552079 598440
rect 378796 598436 378802 598438
rect 552013 598435 552079 598438
rect 552841 597818 552907 597821
rect 549884 597816 552907 597818
rect 549884 597760 552846 597816
rect 552902 597760 552907 597816
rect 549884 597758 552907 597760
rect 552841 597755 552907 597758
rect 407297 597138 407363 597141
rect 407297 597136 410044 597138
rect 407297 597080 407302 597136
rect 407358 597080 410044 597136
rect 407297 597078 410044 597080
rect 407297 597075 407363 597078
rect 550817 596458 550883 596461
rect 549884 596456 550883 596458
rect 549884 596400 550822 596456
rect 550878 596400 550883 596456
rect 549884 596398 550883 596400
rect 550817 596395 550883 596398
rect 407297 595098 407363 595101
rect 407297 595096 410044 595098
rect 407297 595040 407302 595096
rect 407358 595040 410044 595096
rect 407297 595038 410044 595040
rect 407297 595035 407363 595038
rect 407941 594418 408007 594421
rect 407941 594416 410044 594418
rect 407941 594360 407946 594416
rect 408002 594360 410044 594416
rect 407941 594358 410044 594360
rect 407941 594355 408007 594358
rect 371918 593676 371924 593740
rect 371988 593738 371994 593740
rect 371988 593678 410044 593738
rect 371988 593676 371994 593678
rect -960 592908 480 593148
rect 407297 593058 407363 593061
rect 407297 593056 410044 593058
rect 407297 593000 407302 593056
rect 407358 593000 410044 593056
rect 407297 592998 410044 593000
rect 407297 592995 407363 592998
rect 407297 591154 407363 591157
rect 410014 591154 410074 591600
rect 549884 591570 550282 591630
rect 550222 591562 550282 591570
rect 550222 591502 550650 591562
rect 550590 591426 550650 591502
rect 552473 591426 552539 591429
rect 550590 591424 552539 591426
rect 550590 591368 552478 591424
rect 552534 591368 552539 591424
rect 550590 591366 552539 591368
rect 552473 591363 552539 591366
rect 407297 591152 410074 591154
rect 407297 591096 407302 591152
rect 407358 591096 410074 591152
rect 407297 591094 410074 591096
rect 407297 591091 407363 591094
rect 397310 590956 397316 591020
rect 397380 591018 397386 591020
rect 552013 591018 552079 591021
rect 397380 590958 410044 591018
rect 549884 591016 552079 591018
rect 549884 590960 552018 591016
rect 552074 590960 552079 591016
rect 549884 590958 552079 590960
rect 397380 590956 397386 590958
rect 552013 590955 552079 590958
rect 580717 591018 580783 591021
rect 583520 591018 584960 591108
rect 580717 591016 584960 591018
rect 580717 590960 580722 591016
rect 580778 590960 584960 591016
rect 580717 590958 584960 590960
rect 580717 590955 580783 590958
rect 583520 590868 584960 590958
rect 50061 590612 50127 590613
rect 55857 590612 55923 590613
rect 50061 590608 50108 590612
rect 50172 590610 50178 590612
rect 55806 590610 55812 590612
rect 50061 590552 50066 590608
rect 50061 590548 50108 590552
rect 50172 590550 50218 590610
rect 55766 590550 55812 590610
rect 55876 590608 55923 590612
rect 55918 590552 55923 590608
rect 50172 590548 50178 590550
rect 55806 590548 55812 590550
rect 55876 590548 55923 590552
rect 50061 590547 50127 590548
rect 55857 590547 55923 590548
rect 60365 590612 60431 590613
rect 60365 590608 60412 590612
rect 60476 590610 60482 590612
rect 69013 590610 69079 590613
rect 74809 590612 74875 590613
rect 69790 590610 69796 590612
rect 60365 590552 60370 590608
rect 60365 590548 60412 590552
rect 60476 590550 60522 590610
rect 69013 590608 69796 590610
rect 69013 590552 69018 590608
rect 69074 590552 69796 590608
rect 69013 590550 69796 590552
rect 60476 590548 60482 590550
rect 60365 590547 60431 590548
rect 69013 590547 69079 590550
rect 69790 590548 69796 590550
rect 69860 590548 69866 590612
rect 74758 590610 74764 590612
rect 74718 590550 74764 590610
rect 74828 590608 74875 590612
rect 74870 590552 74875 590608
rect 74758 590548 74764 590550
rect 74828 590548 74875 590552
rect 77518 590548 77524 590612
rect 77588 590610 77594 590612
rect 77845 590610 77911 590613
rect 77588 590608 77911 590610
rect 77588 590552 77850 590608
rect 77906 590552 77911 590608
rect 77588 590550 77911 590552
rect 77588 590548 77594 590550
rect 74809 590547 74875 590548
rect 77845 590547 77911 590550
rect 99925 590612 99991 590613
rect 107561 590612 107627 590613
rect 99925 590608 99972 590612
rect 100036 590610 100042 590612
rect 107510 590610 107516 590612
rect 99925 590552 99930 590608
rect 99925 590548 99972 590552
rect 100036 590550 100082 590610
rect 107470 590550 107516 590610
rect 107580 590608 107627 590612
rect 107622 590552 107627 590608
rect 100036 590548 100042 590550
rect 107510 590548 107516 590550
rect 107580 590548 107627 590552
rect 99925 590547 99991 590548
rect 107561 590547 107627 590548
rect 127341 590612 127407 590613
rect 129733 590612 129799 590613
rect 127341 590608 127388 590612
rect 127452 590610 127458 590612
rect 127341 590552 127346 590608
rect 127341 590548 127388 590552
rect 127452 590550 127498 590610
rect 129733 590608 129780 590612
rect 129844 590610 129850 590612
rect 220813 590610 220879 590613
rect 223021 590612 223087 590613
rect 238385 590612 238451 590613
rect 221958 590610 221964 590612
rect 129733 590552 129738 590608
rect 127452 590548 127458 590550
rect 129733 590548 129780 590552
rect 129844 590550 129890 590610
rect 220813 590608 221964 590610
rect 220813 590552 220818 590608
rect 220874 590552 221964 590608
rect 220813 590550 221964 590552
rect 129844 590548 129850 590550
rect 127341 590547 127407 590548
rect 129733 590547 129799 590548
rect 220813 590547 220879 590550
rect 221958 590548 221964 590550
rect 222028 590548 222034 590612
rect 223021 590608 223068 590612
rect 223132 590610 223138 590612
rect 238334 590610 238340 590612
rect 223021 590552 223026 590608
rect 223021 590548 223068 590552
rect 223132 590550 223178 590610
rect 238294 590550 238340 590610
rect 238404 590608 238451 590612
rect 238446 590552 238451 590608
rect 223132 590548 223138 590550
rect 238334 590548 238340 590550
rect 238404 590548 238451 590552
rect 223021 590547 223087 590548
rect 238385 590547 238451 590548
rect 241513 590610 241579 590613
rect 246665 590612 246731 590613
rect 252369 590612 252435 590613
rect 241830 590610 241836 590612
rect 241513 590608 241836 590610
rect 241513 590552 241518 590608
rect 241574 590552 241836 590608
rect 241513 590550 241836 590552
rect 241513 590547 241579 590550
rect 241830 590548 241836 590550
rect 241900 590548 241906 590612
rect 246614 590610 246620 590612
rect 246574 590550 246620 590610
rect 246684 590608 246731 590612
rect 252318 590610 252324 590612
rect 246726 590552 246731 590608
rect 246614 590548 246620 590550
rect 246684 590548 246731 590552
rect 252278 590550 252324 590610
rect 252388 590608 252435 590612
rect 252430 590552 252435 590608
rect 252318 590548 252324 590550
rect 252388 590548 252435 590552
rect 246665 590547 246731 590548
rect 252369 590547 252435 590548
rect 273253 590610 273319 590613
rect 289537 590612 289603 590613
rect 292113 590612 292179 590613
rect 274214 590610 274220 590612
rect 273253 590608 274220 590610
rect 273253 590552 273258 590608
rect 273314 590552 274220 590608
rect 273253 590550 274220 590552
rect 273253 590547 273319 590550
rect 274214 590548 274220 590550
rect 274284 590548 274290 590612
rect 289486 590610 289492 590612
rect 289446 590550 289492 590610
rect 289556 590608 289603 590612
rect 292062 590610 292068 590612
rect 289598 590552 289603 590608
rect 289486 590548 289492 590550
rect 289556 590548 289603 590552
rect 292022 590550 292068 590610
rect 292132 590608 292179 590612
rect 292174 590552 292179 590608
rect 292062 590548 292068 590550
rect 292132 590548 292179 590552
rect 311934 590548 311940 590612
rect 312004 590610 312010 590612
rect 312077 590610 312143 590613
rect 312004 590608 312143 590610
rect 312004 590552 312082 590608
rect 312138 590552 312143 590608
rect 312004 590550 312143 590552
rect 312004 590548 312010 590550
rect 289537 590547 289603 590548
rect 292113 590547 292179 590548
rect 312077 590547 312143 590550
rect 48446 590412 48452 590476
rect 48516 590474 48522 590476
rect 75177 590474 75243 590477
rect 48516 590472 75243 590474
rect 48516 590416 75182 590472
rect 75238 590416 75243 590472
rect 48516 590414 75243 590416
rect 48516 590412 48522 590414
rect 75177 590411 75243 590414
rect 77293 590474 77359 590477
rect 77886 590474 77892 590476
rect 77293 590472 77892 590474
rect 77293 590416 77298 590472
rect 77354 590416 77892 590472
rect 77293 590414 77892 590416
rect 77293 590411 77359 590414
rect 77886 590412 77892 590414
rect 77956 590412 77962 590476
rect 78673 590474 78739 590477
rect 79910 590474 79916 590476
rect 78673 590472 79916 590474
rect 78673 590416 78678 590472
rect 78734 590416 79916 590472
rect 78673 590414 79916 590416
rect 78673 590411 78739 590414
rect 79910 590412 79916 590414
rect 79980 590412 79986 590476
rect 92473 590474 92539 590477
rect 93158 590474 93164 590476
rect 92473 590472 93164 590474
rect 92473 590416 92478 590472
rect 92534 590416 93164 590472
rect 92473 590414 93164 590416
rect 92473 590411 92539 590414
rect 93158 590412 93164 590414
rect 93228 590412 93234 590476
rect 97574 590412 97580 590476
rect 97644 590474 97650 590476
rect 351126 590474 351132 590476
rect 97644 590414 351132 590474
rect 97644 590412 97650 590414
rect 351126 590412 351132 590414
rect 351196 590412 351202 590476
rect 43478 590276 43484 590340
rect 43548 590338 43554 590340
rect 402421 590338 402487 590341
rect 43548 590336 402487 590338
rect 43548 590280 402426 590336
rect 402482 590280 402487 590336
rect 43548 590278 402487 590280
rect 43548 590276 43554 590278
rect 402421 590275 402487 590278
rect 43846 590140 43852 590204
rect 43916 590202 43922 590204
rect 405181 590202 405247 590205
rect 43916 590200 405247 590202
rect 43916 590144 405186 590200
rect 405242 590144 405247 590200
rect 43916 590142 405247 590144
rect 43916 590140 43922 590142
rect 405181 590139 405247 590142
rect 42517 590066 42583 590069
rect 405365 590066 405431 590069
rect 42517 590064 405431 590066
rect 42517 590008 42522 590064
rect 42578 590008 405370 590064
rect 405426 590008 405431 590064
rect 42517 590006 405431 590008
rect 42517 590003 42583 590006
rect 405365 590003 405431 590006
rect 35249 589930 35315 589933
rect 404905 589930 404971 589933
rect 35249 589928 404971 589930
rect 35249 589872 35254 589928
rect 35310 589872 404910 589928
rect 404966 589872 404971 589928
rect 35249 589870 404971 589872
rect 35249 589867 35315 589870
rect 404905 589867 404971 589870
rect 75177 589794 75243 589797
rect 122557 589796 122623 589797
rect 240593 589796 240659 589797
rect 85246 589794 85252 589796
rect 75177 589792 85252 589794
rect 75177 589736 75182 589792
rect 75238 589736 85252 589792
rect 75177 589734 85252 589736
rect 75177 589731 75243 589734
rect 85246 589732 85252 589734
rect 85316 589732 85322 589796
rect 122557 589792 122604 589796
rect 122668 589794 122674 589796
rect 240542 589794 240548 589796
rect 122557 589736 122562 589792
rect 122557 589732 122604 589736
rect 122668 589734 122714 589794
rect 240502 589734 240548 589794
rect 240612 589792 240659 589796
rect 240654 589736 240659 589792
rect 122668 589732 122674 589734
rect 240542 589732 240548 589734
rect 240612 589732 240659 589736
rect 255814 589732 255820 589796
rect 255884 589794 255890 589796
rect 256049 589794 256115 589797
rect 255884 589792 256115 589794
rect 255884 589736 256054 589792
rect 256110 589736 256115 589792
rect 255884 589734 256115 589736
rect 255884 589732 255890 589734
rect 122557 589731 122623 589732
rect 240593 589731 240659 589732
rect 256049 589731 256115 589734
rect 304574 589732 304580 589796
rect 304644 589794 304650 589796
rect 350574 589794 350580 589796
rect 304644 589734 350580 589794
rect 304644 589732 304650 589734
rect 350574 589732 350580 589734
rect 350644 589732 350650 589796
rect 67633 589658 67699 589661
rect 137277 589660 137343 589661
rect 68502 589658 68508 589660
rect 67633 589656 68508 589658
rect 67633 589600 67638 589656
rect 67694 589600 68508 589656
rect 67633 589598 68508 589600
rect 67633 589595 67699 589598
rect 68502 589596 68508 589598
rect 68572 589596 68578 589660
rect 137277 589656 137324 589660
rect 137388 589658 137394 589660
rect 278957 589658 279023 589661
rect 279366 589658 279372 589660
rect 137277 589600 137282 589656
rect 137277 589596 137324 589600
rect 137388 589598 137434 589658
rect 278957 589656 279372 589658
rect 278957 589600 278962 589656
rect 279018 589600 279372 589656
rect 278957 589598 279372 589600
rect 137388 589596 137394 589598
rect 137277 589595 137343 589596
rect 278957 589595 279023 589598
rect 279366 589596 279372 589598
rect 279436 589596 279442 589660
rect 329230 589596 329236 589660
rect 329300 589658 329306 589660
rect 329741 589658 329807 589661
rect 329300 589656 329807 589658
rect 329300 589600 329746 589656
rect 329802 589600 329807 589656
rect 329300 589598 329807 589600
rect 329300 589596 329306 589598
rect 329741 589595 329807 589598
rect 51073 589522 51139 589525
rect 52126 589522 52132 589524
rect 51073 589520 52132 589522
rect 51073 589464 51078 589520
rect 51134 589464 52132 589520
rect 51073 589462 52132 589464
rect 51073 589459 51139 589462
rect 52126 589460 52132 589462
rect 52196 589460 52202 589524
rect 53833 589522 53899 589525
rect 54518 589522 54524 589524
rect 53833 589520 54524 589522
rect 53833 589464 53838 589520
rect 53894 589464 54524 589520
rect 53833 589462 54524 589464
rect 53833 589459 53899 589462
rect 54518 589460 54524 589462
rect 54588 589460 54594 589524
rect 59486 589460 59492 589524
rect 59556 589522 59562 589524
rect 60641 589522 60707 589525
rect 59556 589520 60707 589522
rect 59556 589464 60646 589520
rect 60702 589464 60707 589520
rect 59556 589462 60707 589464
rect 59556 589460 59562 589462
rect 60641 589459 60707 589462
rect 62205 589522 62271 589525
rect 62614 589522 62620 589524
rect 62205 589520 62620 589522
rect 62205 589464 62210 589520
rect 62266 589464 62620 589520
rect 62205 589462 62620 589464
rect 62205 589459 62271 589462
rect 62614 589460 62620 589462
rect 62684 589460 62690 589524
rect 72182 589460 72188 589524
rect 72252 589522 72258 589524
rect 72417 589522 72483 589525
rect 72252 589520 72483 589522
rect 72252 589464 72422 589520
rect 72478 589464 72483 589520
rect 72252 589462 72483 589464
rect 72252 589460 72258 589462
rect 72417 589459 72483 589462
rect 74533 589522 74599 589525
rect 75678 589522 75684 589524
rect 74533 589520 75684 589522
rect 74533 589464 74538 589520
rect 74594 589464 75684 589520
rect 74533 589462 75684 589464
rect 74533 589459 74599 589462
rect 75678 589460 75684 589462
rect 75748 589460 75754 589524
rect 78673 589522 78739 589525
rect 79174 589522 79180 589524
rect 78673 589520 79180 589522
rect 78673 589464 78678 589520
rect 78734 589464 79180 589520
rect 78673 589462 79180 589464
rect 78673 589459 78739 589462
rect 79174 589460 79180 589462
rect 79244 589460 79250 589524
rect 80462 589460 80468 589524
rect 80532 589522 80538 589524
rect 81341 589522 81407 589525
rect 80532 589520 81407 589522
rect 80532 589464 81346 589520
rect 81402 589464 81407 589520
rect 80532 589462 81407 589464
rect 80532 589460 80538 589462
rect 81341 589459 81407 589462
rect 82302 589460 82308 589524
rect 82372 589522 82378 589524
rect 82721 589522 82787 589525
rect 82372 589520 82787 589522
rect 82372 589464 82726 589520
rect 82782 589464 82787 589520
rect 82372 589462 82787 589464
rect 82372 589460 82378 589462
rect 82721 589459 82787 589462
rect 84193 589522 84259 589525
rect 84878 589522 84884 589524
rect 84193 589520 84884 589522
rect 84193 589464 84198 589520
rect 84254 589464 84884 589520
rect 84193 589462 84884 589464
rect 84193 589459 84259 589462
rect 84878 589460 84884 589462
rect 84948 589460 84954 589524
rect 87270 589460 87276 589524
rect 87340 589522 87346 589524
rect 88241 589522 88307 589525
rect 87340 589520 88307 589522
rect 87340 589464 88246 589520
rect 88302 589464 88307 589520
rect 87340 589462 88307 589464
rect 87340 589460 87346 589462
rect 88241 589459 88307 589462
rect 88374 589460 88380 589524
rect 88444 589522 88450 589524
rect 89621 589522 89687 589525
rect 88444 589520 89687 589522
rect 88444 589464 89626 589520
rect 89682 589464 89687 589520
rect 88444 589462 89687 589464
rect 88444 589460 88450 589462
rect 89621 589459 89687 589462
rect 90030 589460 90036 589524
rect 90100 589522 90106 589524
rect 91001 589522 91067 589525
rect 90100 589520 91067 589522
rect 90100 589464 91006 589520
rect 91062 589464 91067 589520
rect 90100 589462 91067 589464
rect 90100 589460 90106 589462
rect 91001 589459 91067 589462
rect 104893 589524 104959 589525
rect 104893 589520 104940 589524
rect 105004 589522 105010 589524
rect 104893 589464 104898 589520
rect 104893 589460 104940 589464
rect 105004 589462 105050 589522
rect 105004 589460 105010 589462
rect 229134 589460 229140 589524
rect 229204 589522 229210 589524
rect 230197 589522 230263 589525
rect 229204 589520 230263 589522
rect 229204 589464 230202 589520
rect 230258 589464 230263 589520
rect 229204 589462 230263 589464
rect 229204 589460 229210 589462
rect 104893 589459 104959 589460
rect 230197 589459 230263 589462
rect 230473 589522 230539 589525
rect 231342 589522 231348 589524
rect 230473 589520 231348 589522
rect 230473 589464 230478 589520
rect 230534 589464 231348 589520
rect 230473 589462 231348 589464
rect 230473 589459 230539 589462
rect 231342 589460 231348 589462
rect 231412 589460 231418 589524
rect 234286 589460 234292 589524
rect 234356 589522 234362 589524
rect 234521 589522 234587 589525
rect 234356 589520 234587 589522
rect 234356 589464 234526 589520
rect 234582 589464 234587 589520
rect 234356 589462 234587 589464
rect 234356 589460 234362 589462
rect 234521 589459 234587 589462
rect 235993 589522 236059 589525
rect 237230 589522 237236 589524
rect 235993 589520 237236 589522
rect 235993 589464 235998 589520
rect 236054 589464 237236 589520
rect 235993 589462 237236 589464
rect 235993 589459 236059 589462
rect 237230 589460 237236 589462
rect 237300 589460 237306 589524
rect 239622 589460 239628 589524
rect 239692 589522 239698 589524
rect 239949 589522 240015 589525
rect 239692 589520 240015 589522
rect 239692 589464 239954 589520
rect 240010 589464 240015 589520
rect 239692 589462 240015 589464
rect 239692 589460 239698 589462
rect 239949 589459 240015 589462
rect 242198 589460 242204 589524
rect 242268 589522 242274 589524
rect 242801 589522 242867 589525
rect 242268 589520 242867 589522
rect 242268 589464 242806 589520
rect 242862 589464 242867 589520
rect 242268 589462 242867 589464
rect 242268 589460 242274 589462
rect 242801 589459 242867 589462
rect 244273 589522 244339 589525
rect 244406 589522 244412 589524
rect 244273 589520 244412 589522
rect 244273 589464 244278 589520
rect 244334 589464 244412 589520
rect 244273 589462 244412 589464
rect 244273 589459 244339 589462
rect 244406 589460 244412 589462
rect 244476 589460 244482 589524
rect 248413 589522 248479 589525
rect 251173 589524 251239 589525
rect 248822 589522 248828 589524
rect 248413 589520 248828 589522
rect 248413 589464 248418 589520
rect 248474 589464 248828 589520
rect 248413 589462 248828 589464
rect 248413 589459 248479 589462
rect 248822 589460 248828 589462
rect 248892 589460 248898 589524
rect 251173 589522 251220 589524
rect 251128 589520 251220 589522
rect 251128 589464 251178 589520
rect 251128 589462 251220 589464
rect 251173 589460 251220 589462
rect 251284 589460 251290 589524
rect 253933 589522 253999 589525
rect 254710 589522 254716 589524
rect 253933 589520 254716 589522
rect 253933 589464 253938 589520
rect 253994 589464 254716 589520
rect 253933 589462 254716 589464
rect 251173 589459 251239 589460
rect 253933 589459 253999 589462
rect 254710 589460 254716 589462
rect 254780 589460 254786 589524
rect 256918 589460 256924 589524
rect 256988 589522 256994 589524
rect 257981 589522 258047 589525
rect 256988 589520 258047 589522
rect 256988 589464 257986 589520
rect 258042 589464 258047 589520
rect 256988 589462 258047 589464
rect 256988 589460 256994 589462
rect 257981 589459 258047 589462
rect 259453 589522 259519 589525
rect 260414 589522 260420 589524
rect 259453 589520 260420 589522
rect 259453 589464 259458 589520
rect 259514 589464 260420 589520
rect 259453 589462 260420 589464
rect 259453 589459 259519 589462
rect 260414 589460 260420 589462
rect 260484 589460 260490 589524
rect 260833 589522 260899 589525
rect 262070 589522 262076 589524
rect 260833 589520 262076 589522
rect 260833 589464 260838 589520
rect 260894 589464 262076 589520
rect 260833 589462 262076 589464
rect 260833 589459 260899 589462
rect 262070 589460 262076 589462
rect 262140 589460 262146 589524
rect 264094 589460 264100 589524
rect 264164 589522 264170 589524
rect 264881 589522 264947 589525
rect 264164 589520 264947 589522
rect 264164 589464 264886 589520
rect 264942 589464 264947 589520
rect 264164 589462 264947 589464
rect 264164 589460 264170 589462
rect 264881 589459 264947 589462
rect 266353 589522 266419 589525
rect 266854 589522 266860 589524
rect 266353 589520 266860 589522
rect 266353 589464 266358 589520
rect 266414 589464 266860 589520
rect 266353 589462 266860 589464
rect 266353 589459 266419 589462
rect 266854 589460 266860 589462
rect 266924 589460 266930 589524
rect 293953 589522 294019 589525
rect 294454 589522 294460 589524
rect 293953 589520 294460 589522
rect 293953 589464 293958 589520
rect 294014 589464 294460 589520
rect 293953 589462 294460 589464
rect 293953 589459 294019 589462
rect 294454 589460 294460 589462
rect 294524 589460 294530 589524
rect 296713 589522 296779 589525
rect 299473 589524 299539 589525
rect 297030 589522 297036 589524
rect 296713 589520 297036 589522
rect 296713 589464 296718 589520
rect 296774 589464 297036 589520
rect 296713 589462 297036 589464
rect 296713 589459 296779 589462
rect 297030 589460 297036 589462
rect 297100 589460 297106 589524
rect 299422 589522 299428 589524
rect 299382 589462 299428 589522
rect 299492 589520 299539 589524
rect 299534 589464 299539 589520
rect 299422 589460 299428 589462
rect 299492 589460 299539 589464
rect 299473 589459 299539 589460
rect 300853 589522 300919 589525
rect 301814 589522 301820 589524
rect 300853 589520 301820 589522
rect 300853 589464 300858 589520
rect 300914 589464 301820 589520
rect 300853 589462 301820 589464
rect 300853 589459 300919 589462
rect 301814 589460 301820 589462
rect 301884 589460 301890 589524
rect 306373 589522 306439 589525
rect 306966 589522 306972 589524
rect 306373 589520 306972 589522
rect 306373 589464 306378 589520
rect 306434 589464 306972 589520
rect 306373 589462 306972 589464
rect 306373 589459 306439 589462
rect 306966 589460 306972 589462
rect 307036 589460 307042 589524
rect 309133 589522 309199 589525
rect 309358 589522 309364 589524
rect 309133 589520 309364 589522
rect 309133 589464 309138 589520
rect 309194 589464 309364 589520
rect 309133 589462 309364 589464
rect 309133 589459 309199 589462
rect 309358 589460 309364 589462
rect 309428 589460 309434 589524
rect 329414 589460 329420 589524
rect 329484 589522 329490 589524
rect 329649 589522 329715 589525
rect 329484 589520 329715 589522
rect 329484 589464 329654 589520
rect 329710 589464 329715 589520
rect 329484 589462 329715 589464
rect 329484 589460 329490 589462
rect 329649 589459 329715 589462
rect 51165 589388 51231 589389
rect 51165 589384 51212 589388
rect 51276 589386 51282 589388
rect 51165 589328 51170 589384
rect 51165 589324 51212 589328
rect 51276 589326 51322 589386
rect 51276 589324 51282 589326
rect 53598 589324 53604 589388
rect 53668 589386 53674 589388
rect 53741 589386 53807 589389
rect 53668 589384 53807 589386
rect 53668 589328 53746 589384
rect 53802 589328 53807 589384
rect 53668 589326 53807 589328
rect 53668 589324 53674 589326
rect 51165 589323 51231 589324
rect 53741 589323 53807 589326
rect 56685 589386 56751 589389
rect 57094 589386 57100 589388
rect 56685 589384 57100 589386
rect 56685 589328 56690 589384
rect 56746 589328 57100 589384
rect 56685 589326 57100 589328
rect 56685 589323 56751 589326
rect 57094 589324 57100 589326
rect 57164 589324 57170 589388
rect 57973 589386 58039 589389
rect 58198 589386 58204 589388
rect 57973 589384 58204 589386
rect 57973 589328 57978 589384
rect 58034 589328 58204 589384
rect 57973 589326 58204 589328
rect 57973 589323 58039 589326
rect 58198 589324 58204 589326
rect 58268 589324 58274 589388
rect 60733 589386 60799 589389
rect 61510 589386 61516 589388
rect 60733 589384 61516 589386
rect 60733 589328 60738 589384
rect 60794 589328 61516 589384
rect 60733 589326 61516 589328
rect 60733 589323 60799 589326
rect 61510 589324 61516 589326
rect 61580 589324 61586 589388
rect 62113 589386 62179 589389
rect 62246 589386 62252 589388
rect 62113 589384 62252 589386
rect 62113 589328 62118 589384
rect 62174 589328 62252 589384
rect 62113 589326 62252 589328
rect 62113 589323 62179 589326
rect 62246 589324 62252 589326
rect 62316 589324 62322 589388
rect 63493 589386 63559 589389
rect 64781 589388 64847 589389
rect 65425 589388 65491 589389
rect 64086 589386 64092 589388
rect 63493 589384 64092 589386
rect 63493 589328 63498 589384
rect 63554 589328 64092 589384
rect 63493 589326 64092 589328
rect 63493 589323 63559 589326
rect 64086 589324 64092 589326
rect 64156 589324 64162 589388
rect 64781 589384 64828 589388
rect 64892 589386 64898 589388
rect 65374 589386 65380 589388
rect 64781 589328 64786 589384
rect 64781 589324 64828 589328
rect 64892 589326 64938 589386
rect 65334 589326 65380 589386
rect 65444 589384 65491 589388
rect 66253 589388 66319 589389
rect 66253 589386 66300 589388
rect 65486 589328 65491 589384
rect 64892 589324 64898 589326
rect 65374 589324 65380 589326
rect 65444 589324 65491 589328
rect 66208 589384 66300 589386
rect 66208 589328 66258 589384
rect 66208 589326 66300 589328
rect 64781 589323 64847 589324
rect 65425 589323 65491 589324
rect 66253 589324 66300 589326
rect 66364 589324 66370 589388
rect 67398 589324 67404 589388
rect 67468 589386 67474 589388
rect 67541 589386 67607 589389
rect 67468 589384 67607 589386
rect 67468 589328 67546 589384
rect 67602 589328 67607 589384
rect 67468 589326 67607 589328
rect 67468 589324 67474 589326
rect 66253 589323 66319 589324
rect 67541 589323 67607 589326
rect 67725 589388 67791 589389
rect 67725 589384 67772 589388
rect 67836 589386 67842 589388
rect 67725 589328 67730 589384
rect 67725 589324 67772 589328
rect 67836 589326 67882 589386
rect 67836 589324 67842 589326
rect 70158 589324 70164 589388
rect 70228 589386 70234 589388
rect 70301 589386 70367 589389
rect 71129 589388 71195 589389
rect 71078 589386 71084 589388
rect 70228 589384 70367 589386
rect 70228 589328 70306 589384
rect 70362 589328 70367 589384
rect 70228 589326 70367 589328
rect 71038 589326 71084 589386
rect 71148 589384 71195 589388
rect 71190 589328 71195 589384
rect 70228 589324 70234 589326
rect 67725 589323 67791 589324
rect 70301 589323 70367 589326
rect 71078 589324 71084 589326
rect 71148 589324 71195 589328
rect 71129 589323 71195 589324
rect 71773 589386 71839 589389
rect 72366 589386 72372 589388
rect 71773 589384 72372 589386
rect 71773 589328 71778 589384
rect 71834 589328 72372 589384
rect 71773 589326 72372 589328
rect 71773 589323 71839 589326
rect 72366 589324 72372 589326
rect 72436 589324 72442 589388
rect 73153 589386 73219 589389
rect 73470 589386 73476 589388
rect 73153 589384 73476 589386
rect 73153 589328 73158 589384
rect 73214 589328 73476 589384
rect 73153 589326 73476 589328
rect 73153 589323 73219 589326
rect 73470 589324 73476 589326
rect 73540 589324 73546 589388
rect 75126 589324 75132 589388
rect 75196 589386 75202 589388
rect 75637 589386 75703 589389
rect 75196 589384 75703 589386
rect 75196 589328 75642 589384
rect 75698 589328 75703 589384
rect 75196 589326 75703 589328
rect 75196 589324 75202 589326
rect 75637 589323 75703 589326
rect 75913 589386 75979 589389
rect 76782 589386 76788 589388
rect 75913 589384 76788 589386
rect 75913 589328 75918 589384
rect 75974 589328 76788 589384
rect 75913 589326 76788 589328
rect 75913 589323 75979 589326
rect 76782 589324 76788 589326
rect 76852 589324 76858 589388
rect 81433 589386 81499 589389
rect 82629 589388 82695 589389
rect 81566 589386 81572 589388
rect 81433 589384 81572 589386
rect 81433 589328 81438 589384
rect 81494 589328 81572 589384
rect 81433 589326 81572 589328
rect 81433 589323 81499 589326
rect 81566 589324 81572 589326
rect 81636 589324 81642 589388
rect 82629 589386 82676 589388
rect 82584 589384 82676 589386
rect 82584 589328 82634 589384
rect 82584 589326 82676 589328
rect 82629 589324 82676 589326
rect 82740 589324 82746 589388
rect 83774 589324 83780 589388
rect 83844 589386 83850 589388
rect 84101 589386 84167 589389
rect 83844 589384 84167 589386
rect 83844 589328 84106 589384
rect 84162 589328 84167 589384
rect 83844 589326 84167 589328
rect 83844 589324 83850 589326
rect 82629 589323 82695 589324
rect 84101 589323 84167 589326
rect 85573 589386 85639 589389
rect 86166 589386 86172 589388
rect 85573 589384 86172 589386
rect 85573 589328 85578 589384
rect 85634 589328 86172 589384
rect 85573 589326 86172 589328
rect 85573 589323 85639 589326
rect 86166 589324 86172 589326
rect 86236 589324 86242 589388
rect 86953 589386 87019 589389
rect 87638 589386 87644 589388
rect 86953 589384 87644 589386
rect 86953 589328 86958 589384
rect 87014 589328 87644 589384
rect 86953 589326 87644 589328
rect 86953 589323 87019 589326
rect 87638 589324 87644 589326
rect 87708 589324 87714 589388
rect 89713 589386 89779 589389
rect 90909 589388 90975 589389
rect 89846 589386 89852 589388
rect 89713 589384 89852 589386
rect 89713 589328 89718 589384
rect 89774 589328 89852 589384
rect 89713 589326 89852 589328
rect 89713 589323 89779 589326
rect 89846 589324 89852 589326
rect 89916 589324 89922 589388
rect 90909 589386 90956 589388
rect 90864 589384 90956 589386
rect 90864 589328 90914 589384
rect 90864 589326 90956 589328
rect 90909 589324 90956 589326
rect 91020 589324 91026 589388
rect 91093 589386 91159 589389
rect 92054 589386 92060 589388
rect 91093 589384 92060 589386
rect 91093 589328 91098 589384
rect 91154 589328 92060 589384
rect 91093 589326 92060 589328
rect 90909 589323 90975 589324
rect 91093 589323 91159 589326
rect 92054 589324 92060 589326
rect 92124 589324 92130 589388
rect 92422 589324 92428 589388
rect 92492 589386 92498 589388
rect 93761 589386 93827 589389
rect 92492 589384 93827 589386
rect 92492 589328 93766 589384
rect 93822 589328 93827 589384
rect 92492 589326 93827 589328
rect 92492 589324 92498 589326
rect 93761 589323 93827 589326
rect 94998 589324 95004 589388
rect 95068 589386 95074 589388
rect 95141 589386 95207 589389
rect 95068 589384 95207 589386
rect 95068 589328 95146 589384
rect 95202 589328 95207 589384
rect 95068 589326 95207 589328
rect 95068 589324 95074 589326
rect 95141 589323 95207 589326
rect 102358 589324 102364 589388
rect 102428 589386 102434 589388
rect 103421 589386 103487 589389
rect 102428 589384 103487 589386
rect 102428 589328 103426 589384
rect 103482 589328 103487 589384
rect 102428 589326 103487 589328
rect 102428 589324 102434 589326
rect 103421 589323 103487 589326
rect 109902 589324 109908 589388
rect 109972 589386 109978 589388
rect 110321 589386 110387 589389
rect 109972 589384 110387 589386
rect 109972 589328 110326 589384
rect 110382 589328 110387 589384
rect 109972 589326 110387 589328
rect 109972 589324 109978 589326
rect 110321 589323 110387 589326
rect 112478 589324 112484 589388
rect 112548 589386 112554 589388
rect 113081 589386 113147 589389
rect 112548 589384 113147 589386
rect 112548 589328 113086 589384
rect 113142 589328 113147 589384
rect 112548 589326 113147 589328
rect 112548 589324 112554 589326
rect 113081 589323 113147 589326
rect 114870 589324 114876 589388
rect 114940 589386 114946 589388
rect 115841 589386 115907 589389
rect 114940 589384 115907 589386
rect 114940 589328 115846 589384
rect 115902 589328 115907 589384
rect 114940 589326 115907 589328
rect 114940 589324 114946 589326
rect 115841 589323 115907 589326
rect 117313 589386 117379 589389
rect 119981 589388 120047 589389
rect 117446 589386 117452 589388
rect 117313 589384 117452 589386
rect 117313 589328 117318 589384
rect 117374 589328 117452 589384
rect 117313 589326 117452 589328
rect 117313 589323 117379 589326
rect 117446 589324 117452 589326
rect 117516 589324 117522 589388
rect 119981 589384 120028 589388
rect 120092 589386 120098 589388
rect 119981 589328 119986 589384
rect 119981 589324 120028 589328
rect 120092 589326 120138 589386
rect 120092 589324 120098 589326
rect 124990 589324 124996 589388
rect 125060 589386 125066 589388
rect 125501 589386 125567 589389
rect 125060 589384 125567 589386
rect 125060 589328 125506 589384
rect 125562 589328 125567 589384
rect 125060 589326 125567 589328
rect 125060 589324 125066 589326
rect 119981 589323 120047 589324
rect 125501 589323 125567 589326
rect 132493 589388 132559 589389
rect 132493 589384 132540 589388
rect 132604 589386 132610 589388
rect 133873 589386 133939 589389
rect 134926 589386 134932 589388
rect 132493 589328 132498 589384
rect 132493 589324 132540 589328
rect 132604 589326 132650 589386
rect 133873 589384 134932 589386
rect 133873 589328 133878 589384
rect 133934 589328 134932 589384
rect 133873 589326 134932 589328
rect 132604 589324 132610 589326
rect 132493 589323 132559 589324
rect 133873 589323 133939 589326
rect 134926 589324 134932 589326
rect 134996 589324 135002 589388
rect 139894 589324 139900 589388
rect 139964 589386 139970 589388
rect 140681 589386 140747 589389
rect 157241 589388 157307 589389
rect 157190 589386 157196 589388
rect 139964 589384 140747 589386
rect 139964 589328 140686 589384
rect 140742 589328 140747 589384
rect 139964 589326 140747 589328
rect 157150 589326 157196 589386
rect 157260 589384 157307 589388
rect 157302 589328 157307 589384
rect 139964 589324 139970 589326
rect 140681 589323 140747 589326
rect 157190 589324 157196 589326
rect 157260 589324 157307 589328
rect 157374 589324 157380 589388
rect 157444 589386 157450 589388
rect 158621 589386 158687 589389
rect 157444 589384 158687 589386
rect 157444 589328 158626 589384
rect 158682 589328 158687 589384
rect 157444 589326 158687 589328
rect 157444 589324 157450 589326
rect 157241 589323 157307 589324
rect 158621 589323 158687 589326
rect 223573 589386 223639 589389
rect 224166 589386 224172 589388
rect 223573 589384 224172 589386
rect 223573 589328 223578 589384
rect 223634 589328 224172 589384
rect 223573 589326 224172 589328
rect 223573 589323 223639 589326
rect 224166 589324 224172 589326
rect 224236 589324 224242 589388
rect 225321 589386 225387 589389
rect 226609 589388 226675 589389
rect 225638 589386 225644 589388
rect 225321 589384 225644 589386
rect 225321 589328 225326 589384
rect 225382 589328 225644 589384
rect 225321 589326 225644 589328
rect 225321 589323 225387 589326
rect 225638 589324 225644 589326
rect 225708 589324 225714 589388
rect 226558 589386 226564 589388
rect 226518 589326 226564 589386
rect 226628 589384 226675 589388
rect 226670 589328 226675 589384
rect 226558 589324 226564 589326
rect 226628 589324 226675 589328
rect 227846 589324 227852 589388
rect 227916 589386 227922 589388
rect 229001 589386 229067 589389
rect 227916 589384 229067 589386
rect 227916 589328 229006 589384
rect 229062 589328 229067 589384
rect 227916 589326 229067 589328
rect 227916 589324 227922 589326
rect 226609 589323 226675 589324
rect 229001 589323 229067 589326
rect 230238 589324 230244 589388
rect 230308 589386 230314 589388
rect 230381 589386 230447 589389
rect 230308 589384 230447 589386
rect 230308 589328 230386 589384
rect 230442 589328 230447 589384
rect 230308 589326 230447 589328
rect 230308 589324 230314 589326
rect 230381 589323 230447 589326
rect 231853 589386 231919 589389
rect 232446 589386 232452 589388
rect 231853 589384 232452 589386
rect 231853 589328 231858 589384
rect 231914 589328 232452 589384
rect 231853 589326 232452 589328
rect 231853 589323 231919 589326
rect 232446 589324 232452 589326
rect 232516 589324 232522 589388
rect 233233 589386 233299 589389
rect 234613 589388 234679 589389
rect 236085 589388 236151 589389
rect 233550 589386 233556 589388
rect 233233 589384 233556 589386
rect 233233 589328 233238 589384
rect 233294 589328 233556 589384
rect 233233 589326 233556 589328
rect 233233 589323 233299 589326
rect 233550 589324 233556 589326
rect 233620 589324 233626 589388
rect 234613 589384 234660 589388
rect 234724 589386 234730 589388
rect 236085 589386 236132 589388
rect 234613 589328 234618 589384
rect 234613 589324 234660 589328
rect 234724 589326 234770 589386
rect 236040 589384 236132 589386
rect 236040 589328 236090 589384
rect 236040 589326 236132 589328
rect 234724 589324 234730 589326
rect 236085 589324 236132 589326
rect 236196 589324 236202 589388
rect 236678 589324 236684 589388
rect 236748 589386 236754 589388
rect 237281 589386 237347 589389
rect 236748 589384 237347 589386
rect 236748 589328 237286 589384
rect 237342 589328 237347 589384
rect 236748 589326 237347 589328
rect 236748 589324 236754 589326
rect 234613 589323 234679 589324
rect 236085 589323 236151 589324
rect 237281 589323 237347 589326
rect 239438 589324 239444 589388
rect 239508 589386 239514 589388
rect 240041 589386 240107 589389
rect 242893 589388 242959 589389
rect 242893 589386 242940 589388
rect 239508 589384 240107 589386
rect 239508 589328 240046 589384
rect 240102 589328 240107 589384
rect 239508 589326 240107 589328
rect 242848 589384 242940 589386
rect 242848 589328 242898 589384
rect 242848 589326 242940 589328
rect 239508 589324 239514 589326
rect 240041 589323 240107 589326
rect 242893 589324 242940 589326
rect 243004 589324 243010 589388
rect 244038 589324 244044 589388
rect 244108 589386 244114 589388
rect 244181 589386 244247 589389
rect 245561 589388 245627 589389
rect 247033 589388 247099 589389
rect 245510 589386 245516 589388
rect 244108 589384 244247 589386
rect 244108 589328 244186 589384
rect 244242 589328 244247 589384
rect 244108 589326 244247 589328
rect 245470 589326 245516 589386
rect 245580 589384 245627 589388
rect 245622 589328 245627 589384
rect 244108 589324 244114 589326
rect 242893 589323 242959 589324
rect 244181 589323 244247 589326
rect 245510 589324 245516 589326
rect 245580 589324 245627 589328
rect 246982 589324 246988 589388
rect 247052 589386 247099 589388
rect 247052 589384 247144 589386
rect 247094 589328 247144 589384
rect 247052 589326 247144 589328
rect 247052 589324 247099 589326
rect 247718 589324 247724 589388
rect 247788 589386 247794 589388
rect 248321 589386 248387 589389
rect 247788 589384 248387 589386
rect 247788 589328 248326 589384
rect 248382 589328 248387 589384
rect 247788 589326 248387 589328
rect 247788 589324 247794 589326
rect 245561 589323 245627 589324
rect 247033 589323 247099 589324
rect 248321 589323 248387 589326
rect 248505 589386 248571 589389
rect 249558 589386 249564 589388
rect 248505 589384 249564 589386
rect 248505 589328 248510 589384
rect 248566 589328 249564 589384
rect 248505 589326 249564 589328
rect 248505 589323 248571 589326
rect 249558 589324 249564 589326
rect 249628 589324 249634 589388
rect 249793 589386 249859 589389
rect 249926 589386 249932 589388
rect 249793 589384 249932 589386
rect 249793 589328 249798 589384
rect 249854 589328 249932 589384
rect 249793 589326 249932 589328
rect 249793 589323 249859 589326
rect 249926 589324 249932 589326
rect 249996 589324 250002 589388
rect 251265 589386 251331 589389
rect 251950 589386 251956 589388
rect 251265 589384 251956 589386
rect 251265 589328 251270 589384
rect 251326 589328 251956 589384
rect 251265 589326 251956 589328
rect 251265 589323 251331 589326
rect 251950 589324 251956 589326
rect 252020 589324 252026 589388
rect 253606 589324 253612 589388
rect 253676 589386 253682 589388
rect 253841 589386 253907 589389
rect 254117 589388 254183 589389
rect 254117 589386 254164 589388
rect 253676 589384 253907 589386
rect 253676 589328 253846 589384
rect 253902 589328 253907 589384
rect 253676 589326 253907 589328
rect 254072 589384 254164 589386
rect 254072 589328 254122 589384
rect 254072 589326 254164 589328
rect 253676 589324 253682 589326
rect 253841 589323 253907 589326
rect 254117 589324 254164 589326
rect 254228 589324 254234 589388
rect 257286 589324 257292 589388
rect 257356 589386 257362 589388
rect 257889 589386 257955 589389
rect 257356 589384 257955 589386
rect 257356 589328 257894 589384
rect 257950 589328 257955 589384
rect 257356 589326 257955 589328
rect 257356 589324 257362 589326
rect 254117 589323 254183 589324
rect 257889 589323 257955 589326
rect 258073 589386 258139 589389
rect 259269 589388 259335 589389
rect 258206 589386 258212 589388
rect 258073 589384 258212 589386
rect 258073 589328 258078 589384
rect 258134 589328 258212 589384
rect 258073 589326 258212 589328
rect 258073 589323 258139 589326
rect 258206 589324 258212 589326
rect 258276 589324 258282 589388
rect 259269 589386 259316 589388
rect 259224 589384 259316 589386
rect 259224 589328 259274 589384
rect 259224 589326 259316 589328
rect 259269 589324 259316 589326
rect 259380 589324 259386 589388
rect 259678 589324 259684 589388
rect 259748 589386 259754 589388
rect 260741 589386 260807 589389
rect 259748 589384 260807 589386
rect 259748 589328 260746 589384
rect 260802 589328 260807 589384
rect 259748 589326 260807 589328
rect 259748 589324 259754 589326
rect 259269 589323 259335 589324
rect 260741 589323 260807 589326
rect 261702 589324 261708 589388
rect 261772 589386 261778 589388
rect 262121 589386 262187 589389
rect 261772 589384 262187 589386
rect 261772 589328 262126 589384
rect 262182 589328 262187 589384
rect 261772 589326 262187 589328
rect 261772 589324 261778 589326
rect 262121 589323 262187 589326
rect 262990 589324 262996 589388
rect 263060 589386 263066 589388
rect 263501 589386 263567 589389
rect 263060 589384 263567 589386
rect 263060 589328 263506 589384
rect 263562 589328 263567 589384
rect 263060 589326 263567 589328
rect 263060 589324 263066 589326
rect 263501 589323 263567 589326
rect 264462 589324 264468 589388
rect 264532 589386 264538 589388
rect 264789 589386 264855 589389
rect 264532 589384 264855 589386
rect 264532 589328 264794 589384
rect 264850 589328 264855 589384
rect 264532 589326 264855 589328
rect 264532 589324 264538 589326
rect 264789 589323 264855 589326
rect 265198 589324 265204 589388
rect 265268 589386 265274 589388
rect 266261 589386 266327 589389
rect 265268 589384 266327 589386
rect 265268 589328 266266 589384
rect 266322 589328 266327 589384
rect 265268 589326 266327 589328
rect 265268 589324 265274 589326
rect 266261 589323 266327 589326
rect 269614 589324 269620 589388
rect 269684 589386 269690 589388
rect 270401 589386 270467 589389
rect 269684 589384 270467 589386
rect 269684 589328 270406 589384
rect 270462 589328 270467 589384
rect 269684 589326 270467 589328
rect 269684 589324 269690 589326
rect 270401 589323 270467 589326
rect 271873 589386 271939 589389
rect 272006 589386 272012 589388
rect 271873 589384 272012 589386
rect 271873 589328 271878 589384
rect 271934 589328 272012 589384
rect 271873 589326 272012 589328
rect 271873 589323 271939 589326
rect 272006 589324 272012 589326
rect 272076 589324 272082 589388
rect 276974 589324 276980 589388
rect 277044 589386 277050 589388
rect 277301 589386 277367 589389
rect 277044 589384 277367 589386
rect 277044 589328 277306 589384
rect 277362 589328 277367 589384
rect 277044 589326 277367 589328
rect 277044 589324 277050 589326
rect 277301 589323 277367 589326
rect 281942 589324 281948 589388
rect 282012 589386 282018 589388
rect 282821 589386 282887 589389
rect 282012 589384 282887 589386
rect 282012 589328 282826 589384
rect 282882 589328 282887 589384
rect 282012 589326 282887 589328
rect 282012 589324 282018 589326
rect 282821 589323 282887 589326
rect 284293 589386 284359 589389
rect 284518 589386 284524 589388
rect 284293 589384 284524 589386
rect 284293 589328 284298 589384
rect 284354 589328 284524 589384
rect 284293 589326 284524 589328
rect 284293 589323 284359 589326
rect 284518 589324 284524 589326
rect 284588 589324 284594 589388
rect 286910 589324 286916 589388
rect 286980 589386 286986 589388
rect 347078 589386 347084 589388
rect 286980 589326 347084 589386
rect 286980 589324 286986 589326
rect 347078 589324 347084 589326
rect 347148 589324 347154 589388
rect 407297 588978 407363 588981
rect 552013 588978 552079 588981
rect 407297 588976 410044 588978
rect 407297 588920 407302 588976
rect 407358 588920 410044 588976
rect 407297 588918 410044 588920
rect 549884 588976 552079 588978
rect 549884 588920 552018 588976
rect 552074 588920 552079 588976
rect 549884 588918 552079 588920
rect 407297 588915 407363 588918
rect 552013 588915 552079 588918
rect 77845 588570 77911 588573
rect 347998 588570 348004 588572
rect 77845 588568 348004 588570
rect 77845 588512 77850 588568
rect 77906 588512 348004 588568
rect 77845 588510 348004 588512
rect 77845 588507 77911 588510
rect 347998 588508 348004 588510
rect 348068 588508 348074 588572
rect 28901 587346 28967 587349
rect 402605 587346 402671 587349
rect 28901 587344 402671 587346
rect 28901 587288 28906 587344
rect 28962 587288 402610 587344
rect 402666 587288 402671 587344
rect 28901 587286 402671 587288
rect 28901 587283 28967 587286
rect 402605 587283 402671 587286
rect 23381 587210 23447 587213
rect 407757 587210 407823 587213
rect 23381 587208 407823 587210
rect 23381 587152 23386 587208
rect 23442 587152 407762 587208
rect 407818 587152 407823 587208
rect 23381 587150 407823 587152
rect 23381 587147 23447 587150
rect 407757 587147 407823 587150
rect 407297 586938 407363 586941
rect 552013 586938 552079 586941
rect 407297 586936 410044 586938
rect 407297 586880 407302 586936
rect 407358 586880 410044 586936
rect 407297 586878 410044 586880
rect 549884 586936 552079 586938
rect 549884 586880 552018 586936
rect 552074 586880 552079 586936
rect 549884 586878 552079 586880
rect 407297 586875 407363 586878
rect 552013 586875 552079 586878
rect 407941 586258 408007 586261
rect 567326 586258 567332 586260
rect 407941 586256 410044 586258
rect 407941 586200 407946 586256
rect 408002 586200 410044 586256
rect 407941 586198 410044 586200
rect 549884 586198 567332 586258
rect 407941 586195 408007 586198
rect 567326 586196 567332 586198
rect 567396 586196 567402 586260
rect 46790 585652 46796 585716
rect 46860 585714 46866 585716
rect 266353 585714 266419 585717
rect 46860 585712 266419 585714
rect 46860 585656 266358 585712
rect 266414 585656 266419 585712
rect 46860 585654 266419 585656
rect 46860 585652 46866 585654
rect 266353 585651 266419 585654
rect 407665 585578 407731 585581
rect 552013 585578 552079 585581
rect 407665 585576 410044 585578
rect 407665 585520 407670 585576
rect 407726 585520 410044 585576
rect 407665 585518 410044 585520
rect 549884 585576 552079 585578
rect 549884 585520 552018 585576
rect 552074 585520 552079 585576
rect 549884 585518 552079 585520
rect 407665 585515 407731 585518
rect 552013 585515 552079 585518
rect 381670 584836 381676 584900
rect 381740 584898 381746 584900
rect 553209 584898 553275 584901
rect 381740 584838 410044 584898
rect 549884 584896 553275 584898
rect 549884 584840 553214 584896
rect 553270 584840 553275 584896
rect 549884 584838 553275 584840
rect 381740 584836 381746 584838
rect 553209 584835 553275 584838
rect 72417 584490 72483 584493
rect 349470 584490 349476 584492
rect 72417 584488 349476 584490
rect 72417 584432 72422 584488
rect 72478 584432 349476 584488
rect 72417 584430 349476 584432
rect 72417 584427 72483 584430
rect 349470 584428 349476 584430
rect 349540 584428 349546 584492
rect 3693 584354 3759 584357
rect 399702 584354 399708 584356
rect 3693 584352 399708 584354
rect 3693 584296 3698 584352
rect 3754 584296 399708 584352
rect 3693 584294 399708 584296
rect 3693 584291 3759 584294
rect 399702 584292 399708 584294
rect 399772 584292 399778 584356
rect 71129 582994 71195 582997
rect 354438 582994 354444 582996
rect 71129 582992 354444 582994
rect 71129 582936 71134 582992
rect 71190 582936 354444 582992
rect 71129 582934 354444 582936
rect 71129 582931 71195 582934
rect 354438 582932 354444 582934
rect 354508 582932 354514 582996
rect 571558 582178 571564 582180
rect 549884 582118 571564 582178
rect 571558 582116 571564 582118
rect 571628 582116 571634 582180
rect 385534 581436 385540 581500
rect 385604 581498 385610 581500
rect 385604 581438 410044 581498
rect 385604 581436 385610 581438
rect 373390 580756 373396 580820
rect 373460 580818 373466 580820
rect 567510 580818 567516 580820
rect 373460 580758 410044 580818
rect 549884 580758 567516 580818
rect 373460 580756 373466 580758
rect 567510 580756 567516 580758
rect 567580 580756 567586 580820
rect 407297 580138 407363 580141
rect 407297 580136 410044 580138
rect -960 579852 480 580092
rect 407297 580080 407302 580136
rect 407358 580080 410044 580136
rect 407297 580078 410044 580080
rect 407297 580075 407363 580078
rect 552013 579458 552079 579461
rect 549884 579456 552079 579458
rect 549884 579400 552018 579456
rect 552074 579400 552079 579456
rect 549884 579398 552079 579400
rect 552013 579395 552079 579398
rect 359590 578716 359596 578780
rect 359660 578778 359666 578780
rect 359660 578718 410044 578778
rect 359660 578716 359666 578718
rect 408953 578098 409019 578101
rect 552013 578098 552079 578101
rect 408953 578096 410044 578098
rect 408953 578040 408958 578096
rect 409014 578040 410044 578096
rect 408953 578038 410044 578040
rect 549884 578096 552079 578098
rect 549884 578040 552018 578096
rect 552074 578040 552079 578096
rect 549884 578038 552079 578040
rect 408953 578035 409019 578038
rect 552013 578035 552079 578038
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect 407297 577418 407363 577421
rect 407297 577416 410044 577418
rect 407297 577360 407302 577416
rect 407358 577360 410044 577416
rect 407297 577358 410044 577360
rect 407297 577355 407363 577358
rect 407389 576738 407455 576741
rect 561806 576738 561812 576740
rect 407389 576736 410044 576738
rect 407389 576680 407394 576736
rect 407450 576680 410044 576736
rect 407389 576678 410044 576680
rect 549884 576678 561812 576738
rect 407389 576675 407455 576678
rect 561806 576676 561812 576678
rect 561876 576676 561882 576740
rect 45134 575996 45140 576060
rect 45204 576058 45210 576060
rect 273253 576058 273319 576061
rect 552013 576058 552079 576061
rect 45204 576056 273319 576058
rect 45204 576000 273258 576056
rect 273314 576000 273319 576056
rect 45204 575998 273319 576000
rect 549884 576056 552079 576058
rect 549884 576000 552018 576056
rect 552074 576000 552079 576056
rect 549884 575998 552079 576000
rect 45204 575996 45210 575998
rect 273253 575995 273319 575998
rect 552013 575995 552079 575998
rect 47158 574772 47164 574836
rect 47228 574834 47234 574836
rect 253933 574834 253999 574837
rect 47228 574832 253999 574834
rect 47228 574776 253938 574832
rect 253994 574776 253999 574832
rect 47228 574774 253999 574776
rect 47228 574772 47234 574774
rect 253933 574771 253999 574774
rect 46606 574636 46612 574700
rect 46676 574698 46682 574700
rect 300853 574698 300919 574701
rect 46676 574696 300919 574698
rect 46676 574640 300858 574696
rect 300914 574640 300919 574696
rect 46676 574638 300919 574640
rect 46676 574636 46682 574638
rect 300853 574635 300919 574638
rect 549884 574570 550282 574630
rect 550222 574562 550282 574570
rect 552013 574562 552079 574565
rect 550222 574560 552079 574562
rect 550222 574504 552018 574560
rect 552074 574504 552079 574560
rect 550222 574502 552079 574504
rect 552013 574499 552079 574502
rect 408033 574018 408099 574021
rect 552013 574018 552079 574021
rect 408033 574016 410044 574018
rect 408033 573960 408038 574016
rect 408094 573960 410044 574016
rect 408033 573958 410044 573960
rect 549884 574016 552079 574018
rect 549884 573960 552018 574016
rect 552074 573960 552079 574016
rect 549884 573958 552079 573960
rect 408033 573955 408099 573958
rect 552013 573955 552079 573958
rect 407665 573338 407731 573341
rect 407665 573336 410044 573338
rect 407665 573280 407670 573336
rect 407726 573280 410044 573336
rect 407665 573278 410044 573280
rect 407665 573275 407731 573278
rect 407297 572658 407363 572661
rect 407297 572656 410044 572658
rect 407297 572600 407302 572656
rect 407358 572600 410044 572656
rect 407297 572598 410044 572600
rect 407297 572595 407363 572598
rect 46974 572188 46980 572252
rect 47044 572250 47050 572252
rect 248413 572250 248479 572253
rect 47044 572248 248479 572250
rect 47044 572192 248418 572248
rect 248474 572192 248479 572248
rect 47044 572190 248479 572192
rect 47044 572188 47050 572190
rect 248413 572187 248479 572190
rect 90909 572114 90975 572117
rect 346342 572114 346348 572116
rect 90909 572112 346348 572114
rect 90909 572056 90914 572112
rect 90970 572056 346348 572112
rect 90909 572054 346348 572056
rect 90909 572051 90975 572054
rect 346342 572052 346348 572054
rect 346412 572052 346418 572116
rect 46422 571916 46428 571980
rect 46492 571978 46498 571980
rect 309133 571978 309199 571981
rect 46492 571976 309199 571978
rect 46492 571920 309138 571976
rect 309194 571920 309199 571976
rect 46492 571918 309199 571920
rect 46492 571916 46498 571918
rect 309133 571915 309199 571918
rect 409137 570618 409203 570621
rect 409137 570616 410044 570618
rect 409137 570560 409142 570616
rect 409198 570560 410044 570616
rect 409137 570558 410044 570560
rect 409137 570555 409203 570558
rect 407297 569938 407363 569941
rect 550766 569938 550772 569940
rect 407297 569936 410044 569938
rect 407297 569880 407302 569936
rect 407358 569880 410044 569936
rect 407297 569878 410044 569880
rect 549884 569878 550772 569938
rect 407297 569875 407363 569878
rect 550766 569876 550772 569878
rect 550836 569876 550842 569940
rect 130561 568850 130627 568853
rect 352046 568850 352052 568852
rect 130561 568848 352052 568850
rect 130561 568792 130566 568848
rect 130622 568792 352052 568848
rect 130561 568790 352052 568792
rect 130561 568787 130627 568790
rect 352046 568788 352052 568790
rect 352116 568788 352122 568852
rect 126053 568714 126119 568717
rect 376886 568714 376892 568716
rect 126053 568712 376892 568714
rect 126053 568656 126058 568712
rect 126114 568656 376892 568712
rect 126053 568654 376892 568656
rect 126053 568651 126119 568654
rect 376886 568652 376892 568654
rect 376956 568652 376962 568716
rect 553117 568578 553183 568581
rect 549884 568576 553183 568578
rect 549884 568520 553122 568576
rect 553178 568520 553183 568576
rect 549884 568518 553183 568520
rect 553117 568515 553183 568518
rect 347078 568244 347084 568308
rect 347148 568244 347154 568308
rect 347086 568036 347146 568244
rect 347078 567972 347084 568036
rect 347148 567972 347154 568036
rect 45318 567836 45324 567900
rect 45388 567898 45394 567900
rect 284293 567898 284359 567901
rect 45388 567896 284359 567898
rect 45388 567840 284298 567896
rect 284354 567840 284359 567896
rect 45388 567838 284359 567840
rect 45388 567836 45394 567838
rect 284293 567835 284359 567838
rect 407389 567898 407455 567901
rect 553301 567898 553367 567901
rect 407389 567896 410044 567898
rect 407389 567840 407394 567896
rect 407450 567840 410044 567896
rect 407389 567838 410044 567840
rect 549884 567896 553367 567898
rect 549884 567840 553306 567896
rect 553362 567840 553367 567896
rect 549884 567838 553367 567840
rect 407389 567835 407455 567838
rect 553301 567835 553367 567838
rect 308305 567354 308371 567357
rect 378910 567354 378916 567356
rect 308305 567352 378916 567354
rect 308305 567296 308310 567352
rect 308366 567296 378916 567352
rect 308305 567294 378916 567296
rect 308305 567291 308371 567294
rect 378910 567292 378916 567294
rect 378980 567292 378986 567356
rect 216857 567218 216923 567221
rect 381486 567218 381492 567220
rect 216857 567216 381492 567218
rect 216857 567160 216862 567216
rect 216918 567160 381492 567216
rect 216857 567158 381492 567160
rect 216857 567155 216923 567158
rect 381486 567156 381492 567158
rect 381556 567156 381562 567220
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 85481 566810 85547 566813
rect 369158 566810 369164 566812
rect 85481 566808 369164 566810
rect 85481 566752 85486 566808
rect 85542 566752 369164 566808
rect 85481 566750 369164 566752
rect 85481 566747 85547 566750
rect 369158 566748 369164 566750
rect 369228 566748 369234 566812
rect 190361 566674 190427 566677
rect 390134 566674 390140 566676
rect 190361 566672 390140 566674
rect 190361 566616 190366 566672
rect 190422 566616 390140 566672
rect 190361 566614 390140 566616
rect 190361 566611 190427 566614
rect 390134 566612 390140 566614
rect 390204 566612 390210 566676
rect 64781 566538 64847 566541
rect 347814 566538 347820 566540
rect 64781 566536 347820 566538
rect 64781 566480 64786 566536
rect 64842 566480 347820 566536
rect 64781 566478 347820 566480
rect 64781 566475 64847 566478
rect 347814 566476 347820 566478
rect 347884 566476 347890 566540
rect 568614 566538 568620 566540
rect 549884 566478 568620 566538
rect 568614 566476 568620 566478
rect 568684 566476 568690 566540
rect 53741 566402 53807 566405
rect 349102 566402 349108 566404
rect 53741 566400 349108 566402
rect 53741 566344 53746 566400
rect 53802 566344 349108 566400
rect 53741 566342 349108 566344
rect 53741 566339 53807 566342
rect 349102 566340 349108 566342
rect 349172 566340 349178 566404
rect 143441 566266 143507 566269
rect 360694 566266 360700 566268
rect 143441 566264 360700 566266
rect 143441 566208 143446 566264
rect 143502 566208 360700 566264
rect 143441 566206 360700 566208
rect 143441 566203 143507 566206
rect 360694 566204 360700 566206
rect 360764 566204 360770 566268
rect 109585 566130 109651 566133
rect 351862 566130 351868 566132
rect 109585 566128 351868 566130
rect 109585 566072 109590 566128
rect 109646 566072 351868 566128
rect 109585 566070 351868 566072
rect 109585 566067 109651 566070
rect 351862 566068 351868 566070
rect 351932 566068 351938 566132
rect 106181 565994 106247 565997
rect 373206 565994 373212 565996
rect 106181 565992 373212 565994
rect 106181 565936 106186 565992
rect 106242 565936 373212 565992
rect 106181 565934 373212 565936
rect 106181 565931 106247 565934
rect 373206 565932 373212 565934
rect 373276 565932 373282 565996
rect 365110 565796 365116 565860
rect 365180 565858 365186 565860
rect 365180 565798 410044 565858
rect 365180 565796 365186 565798
rect 346894 565116 346900 565180
rect 346964 565178 346970 565180
rect 347630 565178 347636 565180
rect 346964 565118 347636 565178
rect 346964 565116 346970 565118
rect 347630 565116 347636 565118
rect 347700 565116 347706 565180
rect 408309 565178 408375 565181
rect 553301 565178 553367 565181
rect 408309 565176 410044 565178
rect 408309 565120 408314 565176
rect 408370 565120 410044 565176
rect 408309 565118 410044 565120
rect 549884 565176 553367 565178
rect 549884 565120 553306 565176
rect 553362 565120 553367 565176
rect 549884 565118 553367 565120
rect 408309 565115 408375 565118
rect 553301 565115 553367 565118
rect 275001 564906 275067 564909
rect 395286 564906 395292 564908
rect 275001 564904 395292 564906
rect 275001 564848 275006 564904
rect 275062 564848 395292 564904
rect 275001 564846 395292 564848
rect 275001 564843 275067 564846
rect 395286 564844 395292 564846
rect 395356 564844 395362 564908
rect 195881 564770 195947 564773
rect 358261 564770 358327 564773
rect 195881 564768 358327 564770
rect 195881 564712 195886 564768
rect 195942 564712 358266 564768
rect 358322 564712 358327 564768
rect 195881 564710 358327 564712
rect 195881 564707 195947 564710
rect 358261 564707 358327 564710
rect 77937 564634 78003 564637
rect 398281 564634 398347 564637
rect 77937 564632 398347 564634
rect 77937 564576 77942 564632
rect 77998 564576 398286 564632
rect 398342 564576 398347 564632
rect 77937 564574 398347 564576
rect 77937 564571 78003 564574
rect 398281 564571 398347 564574
rect 59813 564498 59879 564501
rect 396574 564498 396580 564500
rect 59813 564496 396580 564498
rect 59813 564440 59818 564496
rect 59874 564440 396580 564496
rect 59813 564438 396580 564440
rect 59813 564435 59879 564438
rect 396574 564436 396580 564438
rect 396644 564436 396650 564500
rect 407389 564498 407455 564501
rect 550173 564498 550239 564501
rect 407389 564496 410044 564498
rect 407389 564440 407394 564496
rect 407450 564440 410044 564496
rect 407389 564438 410044 564440
rect 549884 564496 550239 564498
rect 549884 564440 550178 564496
rect 550234 564440 550239 564496
rect 549884 564438 550239 564440
rect 407389 564435 407455 564438
rect 550173 564435 550239 564438
rect 580533 564362 580599 564365
rect 583520 564362 584960 564452
rect 580533 564360 584960 564362
rect 580533 564304 580538 564360
rect 580594 564304 584960 564360
rect 580533 564302 584960 564304
rect 580533 564299 580599 564302
rect 583520 564212 584960 564302
rect 83089 563818 83155 563821
rect 376201 563818 376267 563821
rect 83089 563816 376267 563818
rect 83089 563760 83094 563816
rect 83150 563760 376206 563816
rect 376262 563760 376267 563816
rect 83089 563758 376267 563760
rect 83089 563755 83155 563758
rect 376201 563755 376267 563758
rect 277025 563682 277091 563685
rect 350942 563682 350948 563684
rect 277025 563680 350948 563682
rect 277025 563624 277030 563680
rect 277086 563624 350948 563680
rect 277025 563622 350948 563624
rect 277025 563619 277091 563622
rect 350942 563620 350948 563622
rect 351012 563620 351018 563684
rect 298921 563546 298987 563549
rect 380341 563546 380407 563549
rect 298921 563544 380407 563546
rect 298921 563488 298926 563544
rect 298982 563488 380346 563544
rect 380402 563488 380407 563544
rect 298921 563486 380407 563488
rect 298921 563483 298987 563486
rect 380341 563483 380407 563486
rect 180701 563410 180767 563413
rect 385769 563410 385835 563413
rect 180701 563408 385835 563410
rect 180701 563352 180706 563408
rect 180762 563352 385774 563408
rect 385830 563352 385835 563408
rect 180701 563350 385835 563352
rect 180701 563347 180767 563350
rect 385769 563347 385835 563350
rect 41270 563212 41276 563276
rect 41340 563274 41346 563276
rect 294321 563274 294387 563277
rect 41340 563272 294387 563274
rect 41340 563216 294326 563272
rect 294382 563216 294387 563272
rect 41340 563214 294387 563216
rect 41340 563212 41346 563214
rect 294321 563211 294387 563214
rect 297633 563274 297699 563277
rect 399518 563274 399524 563276
rect 297633 563272 399524 563274
rect 297633 563216 297638 563272
rect 297694 563216 399524 563272
rect 297633 563214 399524 563216
rect 297633 563211 297699 563214
rect 399518 563212 399524 563214
rect 399588 563212 399594 563276
rect 336181 563138 336247 563141
rect 360377 563138 360443 563141
rect 336181 563136 360443 563138
rect 336181 563080 336186 563136
rect 336242 563080 360382 563136
rect 360438 563080 360443 563136
rect 336181 563078 360443 563080
rect 336181 563075 336247 563078
rect 360377 563075 360443 563078
rect 48446 562668 48452 562732
rect 48516 562730 48522 562732
rect 121545 562730 121611 562733
rect 48516 562728 121611 562730
rect 48516 562672 121550 562728
rect 121606 562672 121611 562728
rect 48516 562670 121611 562672
rect 48516 562668 48522 562670
rect 121545 562667 121611 562670
rect 274449 562730 274515 562733
rect 388621 562730 388687 562733
rect 274449 562728 388687 562730
rect 274449 562672 274454 562728
rect 274510 562672 388626 562728
rect 388682 562672 388687 562728
rect 274449 562670 388687 562672
rect 274449 562667 274515 562670
rect 388621 562667 388687 562670
rect 27470 562532 27476 562596
rect 27540 562594 27546 562596
rect 48957 562594 49023 562597
rect 27540 562592 49023 562594
rect 27540 562536 48962 562592
rect 49018 562536 49023 562592
rect 27540 562534 49023 562536
rect 27540 562532 27546 562534
rect 48957 562531 49023 562534
rect 346342 562532 346348 562596
rect 346412 562594 346418 562596
rect 347446 562594 347452 562596
rect 346412 562534 347452 562594
rect 346412 562532 346418 562534
rect 347446 562532 347452 562534
rect 347516 562532 347522 562596
rect 41638 562396 41644 562460
rect 41708 562458 41714 562460
rect 89713 562458 89779 562461
rect 41708 562456 89779 562458
rect 41708 562400 89718 562456
rect 89774 562400 89779 562456
rect 41708 562398 89779 562400
rect 41708 562396 41714 562398
rect 89713 562395 89779 562398
rect 240041 562458 240107 562461
rect 356697 562458 356763 562461
rect 550909 562458 550975 562461
rect 240041 562456 356763 562458
rect 240041 562400 240046 562456
rect 240102 562400 356702 562456
rect 356758 562400 356763 562456
rect 240041 562398 356763 562400
rect 549884 562456 550975 562458
rect 549884 562400 550914 562456
rect 550970 562400 550975 562456
rect 549884 562398 550975 562400
rect 240041 562395 240107 562398
rect 356697 562395 356763 562398
rect 550909 562395 550975 562398
rect 47761 562322 47827 562325
rect 104341 562322 104407 562325
rect 47761 562320 104407 562322
rect 47761 562264 47766 562320
rect 47822 562264 104346 562320
rect 104402 562264 104407 562320
rect 47761 562262 104407 562264
rect 47761 562259 47827 562262
rect 104341 562259 104407 562262
rect 208761 562322 208827 562325
rect 365989 562322 366055 562325
rect 208761 562320 366055 562322
rect 208761 562264 208766 562320
rect 208822 562264 365994 562320
rect 366050 562264 366055 562320
rect 208761 562262 366055 562264
rect 208761 562259 208827 562262
rect 365989 562259 366055 562262
rect 27521 562186 27587 562189
rect 57973 562186 58039 562189
rect 27521 562184 58039 562186
rect 27521 562128 27526 562184
rect 27582 562128 57978 562184
rect 58034 562128 58039 562184
rect 27521 562126 58039 562128
rect 27521 562123 27587 562126
rect 57973 562123 58039 562126
rect 189441 562186 189507 562189
rect 359457 562186 359523 562189
rect 189441 562184 359523 562186
rect 189441 562128 189446 562184
rect 189502 562128 359462 562184
rect 359518 562128 359523 562184
rect 189441 562126 359523 562128
rect 189441 562123 189507 562126
rect 359457 562123 359523 562126
rect 25957 562050 26023 562053
rect 57421 562050 57487 562053
rect 25957 562048 57487 562050
rect 25957 561992 25962 562048
rect 26018 561992 57426 562048
rect 57482 561992 57487 562048
rect 25957 561990 57487 561992
rect 25957 561987 26023 561990
rect 57421 561987 57487 561990
rect 58525 562050 58591 562053
rect 170765 562050 170831 562053
rect 58525 562048 170831 562050
rect 58525 561992 58530 562048
rect 58586 561992 170770 562048
rect 170826 561992 170831 562048
rect 58525 561990 170831 561992
rect 58525 561987 58591 561990
rect 170765 561987 170831 561990
rect 201033 562050 201099 562053
rect 374494 562050 374500 562052
rect 201033 562048 374500 562050
rect 201033 561992 201038 562048
rect 201094 561992 374500 562048
rect 201033 561990 374500 561992
rect 201033 561987 201099 561990
rect 374494 561988 374500 561990
rect 374564 561988 374570 562052
rect 26141 561914 26207 561917
rect 59905 561914 59971 561917
rect 26141 561912 59971 561914
rect 26141 561856 26146 561912
rect 26202 561856 59910 561912
rect 59966 561856 59971 561912
rect 26141 561854 59971 561856
rect 26141 561851 26207 561854
rect 59905 561851 59971 561854
rect 60733 561914 60799 561917
rect 173893 561914 173959 561917
rect 60733 561912 173959 561914
rect 60733 561856 60738 561912
rect 60794 561856 173898 561912
rect 173954 561856 173959 561912
rect 60733 561854 173959 561856
rect 60733 561851 60799 561854
rect 173893 561851 173959 561854
rect 184841 561914 184907 561917
rect 365897 561914 365963 561917
rect 184841 561912 365963 561914
rect 184841 561856 184846 561912
rect 184902 561856 365902 561912
rect 365958 561856 365963 561912
rect 184841 561854 365963 561856
rect 184841 561851 184907 561854
rect 365897 561851 365963 561854
rect 30097 561778 30163 561781
rect 267917 561778 267983 561781
rect 30097 561776 267983 561778
rect 30097 561720 30102 561776
rect 30158 561720 267922 561776
rect 267978 561720 267983 561776
rect 30097 561718 267983 561720
rect 30097 561715 30163 561718
rect 267917 561715 267983 561718
rect 341977 561778 342043 561781
rect 367134 561778 367140 561780
rect 341977 561776 367140 561778
rect 341977 561720 341982 561776
rect 342038 561720 367140 561776
rect 341977 561718 367140 561720
rect 341977 561715 342043 561718
rect 367134 561716 367140 561718
rect 367204 561716 367210 561780
rect 348049 561642 348115 561645
rect 348366 561642 348372 561644
rect 348049 561640 348372 561642
rect 348049 561584 348054 561640
rect 348110 561584 348372 561640
rect 348049 561582 348372 561584
rect 348049 561579 348115 561582
rect 348366 561580 348372 561582
rect 348436 561580 348442 561644
rect 27337 561370 27403 561373
rect 330477 561370 330543 561373
rect 27337 561368 330543 561370
rect 27337 561312 27342 561368
rect 27398 561312 330482 561368
rect 330538 561312 330543 561368
rect 27337 561310 330543 561312
rect 27337 561307 27403 561310
rect 330477 561307 330543 561310
rect 43805 561234 43871 561237
rect 60733 561234 60799 561237
rect 43805 561232 60799 561234
rect 43805 561176 43810 561232
rect 43866 561176 60738 561232
rect 60794 561176 60799 561232
rect 43805 561174 60799 561176
rect 43805 561171 43871 561174
rect 60733 561171 60799 561174
rect 30005 561098 30071 561101
rect 63493 561098 63559 561101
rect 30005 561096 63559 561098
rect 30005 561040 30010 561096
rect 30066 561040 63498 561096
rect 63554 561040 63559 561096
rect 30005 561038 63559 561040
rect 30005 561035 30071 561038
rect 63493 561035 63559 561038
rect 340137 561098 340203 561101
rect 349286 561098 349292 561100
rect 340137 561096 349292 561098
rect 340137 561040 340142 561096
rect 340198 561040 349292 561096
rect 340137 561038 349292 561040
rect 340137 561035 340203 561038
rect 349286 561036 349292 561038
rect 349356 561036 349362 561100
rect 407389 561098 407455 561101
rect 553117 561098 553183 561101
rect 407389 561096 410044 561098
rect 407389 561040 407394 561096
rect 407450 561040 410044 561096
rect 407389 561038 410044 561040
rect 549884 561096 553183 561098
rect 549884 561040 553122 561096
rect 553178 561040 553183 561096
rect 549884 561038 553183 561040
rect 407389 561035 407455 561038
rect 553117 561035 553183 561038
rect 22645 560962 22711 560965
rect 56685 560962 56751 560965
rect 22645 560960 56751 560962
rect 22645 560904 22650 560960
rect 22706 560904 56690 560960
rect 56746 560904 56751 560960
rect 22645 560902 56751 560904
rect 22645 560899 22711 560902
rect 56685 560899 56751 560902
rect 207473 560962 207539 560965
rect 399334 560962 399340 560964
rect 207473 560960 399340 560962
rect 207473 560904 207478 560960
rect 207534 560904 399340 560960
rect 207473 560902 399340 560904
rect 207473 560899 207539 560902
rect 399334 560900 399340 560902
rect 399404 560900 399410 560964
rect 24577 560826 24643 560829
rect 311157 560826 311223 560829
rect 24577 560824 311223 560826
rect 24577 560768 24582 560824
rect 24638 560768 311162 560824
rect 311218 560768 311223 560824
rect 24577 560766 311223 560768
rect 24577 560763 24643 560766
rect 311157 560763 311223 560766
rect 328361 560690 328427 560693
rect 361757 560690 361823 560693
rect 328361 560688 361823 560690
rect 328361 560632 328366 560688
rect 328422 560632 361762 560688
rect 361818 560632 361823 560688
rect 328361 560630 361823 560632
rect 328361 560627 328427 560630
rect 361757 560627 361823 560630
rect 46238 560492 46244 560556
rect 46308 560554 46314 560556
rect 351361 560554 351427 560557
rect 46308 560552 351427 560554
rect 46308 560496 351366 560552
rect 351422 560496 351427 560552
rect 46308 560494 351427 560496
rect 46308 560492 46314 560494
rect 351361 560491 351427 560494
rect 63217 560418 63283 560421
rect 389950 560418 389956 560420
rect 63217 560416 389956 560418
rect 63217 560360 63222 560416
rect 63278 560360 389956 560416
rect 63217 560358 389956 560360
rect 63217 560355 63283 560358
rect 389950 560356 389956 560358
rect 390020 560356 390026 560420
rect 553301 560418 553367 560421
rect 549884 560416 553367 560418
rect 549884 560360 553306 560416
rect 553362 560360 553367 560416
rect 549884 560358 553367 560360
rect 553301 560355 553367 560358
rect 42241 560146 42307 560149
rect 58525 560146 58591 560149
rect 42241 560144 58591 560146
rect 42241 560088 42246 560144
rect 42302 560088 58530 560144
rect 58586 560088 58591 560144
rect 42241 560086 58591 560088
rect 42241 560083 42307 560086
rect 58525 560083 58591 560086
rect 32673 560010 32739 560013
rect 402421 560010 402487 560013
rect 32673 560008 402487 560010
rect 32673 559952 32678 560008
rect 32734 559952 402426 560008
rect 402482 559952 402487 560008
rect 32673 559950 402487 559952
rect 32673 559947 32739 559950
rect 402421 559947 402487 559950
rect 408033 559058 408099 559061
rect 408033 559056 410044 559058
rect 408033 559000 408038 559056
rect 408094 559000 410044 559056
rect 408033 558998 410044 559000
rect 408033 558995 408099 558998
rect 43345 558922 43411 558925
rect 47761 558922 47827 558925
rect 43345 558920 47827 558922
rect 43345 558864 43350 558920
rect 43406 558864 47766 558920
rect 47822 558864 47827 558920
rect 43345 558862 47827 558864
rect 43345 558859 43411 558862
rect 47761 558859 47827 558862
rect 347630 558860 347636 558924
rect 347700 558922 347706 558924
rect 349654 558922 349660 558924
rect 347700 558862 349660 558922
rect 347700 558860 347706 558862
rect 349654 558860 349660 558862
rect 349724 558860 349730 558924
rect 552933 558378 552999 558381
rect 549884 558376 552999 558378
rect 549884 558320 552938 558376
rect 552994 558320 552999 558376
rect 549884 558318 552999 558320
rect 552933 558315 552999 558318
rect 385718 557636 385724 557700
rect 385788 557698 385794 557700
rect 553301 557698 553367 557701
rect 385788 557638 410044 557698
rect 549884 557696 553367 557698
rect 549884 557640 553306 557696
rect 553362 557640 553367 557696
rect 549884 557638 553367 557640
rect 385788 557636 385794 557638
rect 553301 557635 553367 557638
rect 347630 557228 347636 557292
rect 347700 557228 347706 557292
rect 347638 557124 347698 557228
rect 46105 556610 46171 556613
rect 48086 556610 48146 557056
rect 407665 557018 407731 557021
rect 553301 557018 553367 557021
rect 407665 557016 410044 557018
rect 407665 556960 407670 557016
rect 407726 556960 410044 557016
rect 407665 556958 410044 556960
rect 549884 557016 553367 557018
rect 549884 556960 553306 557016
rect 553362 556960 553367 557016
rect 549884 556958 553367 556960
rect 407665 556955 407731 556958
rect 553301 556955 553367 556958
rect 46105 556608 48146 556610
rect 46105 556552 46110 556608
rect 46166 556552 48146 556608
rect 46105 556550 48146 556552
rect 46105 556547 46171 556550
rect 407389 556338 407455 556341
rect 553301 556338 553367 556341
rect 407389 556336 410044 556338
rect 407389 556280 407394 556336
rect 407450 556280 410044 556336
rect 407389 556278 410044 556280
rect 549884 556336 553367 556338
rect 549884 556280 553306 556336
rect 553362 556280 553367 556336
rect 549884 556278 553367 556280
rect 407389 556275 407455 556278
rect 553301 556275 553367 556278
rect 45921 556202 45987 556205
rect 48262 556202 48268 556204
rect 45921 556200 48268 556202
rect 45921 556144 45926 556200
rect 45982 556144 48268 556200
rect 45921 556142 48268 556144
rect 45921 556139 45987 556142
rect 48262 556140 48268 556142
rect 48332 556140 48338 556204
rect 407941 555658 408007 555661
rect 551093 555658 551159 555661
rect 407941 555656 410044 555658
rect 407941 555600 407946 555656
rect 408002 555600 410044 555656
rect 407941 555598 410044 555600
rect 549884 555656 551159 555658
rect 549884 555600 551098 555656
rect 551154 555600 551159 555656
rect 549884 555598 551159 555600
rect 407941 555595 408007 555598
rect 551093 555595 551159 555598
rect 350441 554434 350507 554437
rect 347852 554432 350507 554434
rect 347852 554376 350446 554432
rect 350502 554376 350507 554432
rect 347852 554374 350507 554376
rect 350441 554371 350507 554374
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 552013 553618 552079 553621
rect 550222 553616 552079 553618
rect 550222 553560 552018 553616
rect 552074 553560 552079 553616
rect 550222 553558 552079 553560
rect 550222 553550 550282 553558
rect 552013 553555 552079 553558
rect 549884 553490 550282 553550
rect 407481 552938 407547 552941
rect 561990 552938 561996 552940
rect 407481 552936 410044 552938
rect 407481 552880 407486 552936
rect 407542 552880 410044 552936
rect 407481 552878 410044 552880
rect 549884 552878 561996 552938
rect 407481 552875 407547 552878
rect 561990 552876 561996 552878
rect 562060 552876 562066 552940
rect 549884 552198 557550 552258
rect 557490 552122 557550 552198
rect 565854 552122 565860 552124
rect 557490 552062 565860 552122
rect 565854 552060 565860 552062
rect 565924 552060 565930 552124
rect 46105 551306 46171 551309
rect 48086 551306 48146 551616
rect 347822 551442 347882 551616
rect 407389 551578 407455 551581
rect 553301 551578 553367 551581
rect 407389 551576 410044 551578
rect 407389 551520 407394 551576
rect 407450 551520 410044 551576
rect 407389 551518 410044 551520
rect 549884 551576 553367 551578
rect 549884 551520 553306 551576
rect 553362 551520 553367 551576
rect 549884 551518 553367 551520
rect 407389 551515 407455 551518
rect 553301 551515 553367 551518
rect 350441 551442 350507 551445
rect 347822 551440 350507 551442
rect 347822 551384 350446 551440
rect 350502 551384 350507 551440
rect 347822 551382 350507 551384
rect 350441 551379 350507 551382
rect 46105 551304 48146 551306
rect 46105 551248 46110 551304
rect 46166 551248 48146 551304
rect 46105 551246 48146 551248
rect 46105 551243 46171 551246
rect 583520 551020 584960 551260
rect 46105 550898 46171 550901
rect 48086 550898 48146 550936
rect 46105 550896 48146 550898
rect 46105 550840 46110 550896
rect 46166 550840 48146 550896
rect 46105 550838 48146 550840
rect 407389 550898 407455 550901
rect 552013 550898 552079 550901
rect 407389 550896 410044 550898
rect 407389 550840 407394 550896
rect 407450 550840 410044 550896
rect 407389 550838 410044 550840
rect 549884 550896 552079 550898
rect 549884 550840 552018 550896
rect 552074 550840 552079 550896
rect 549884 550838 552079 550840
rect 46105 550835 46171 550838
rect 407389 550835 407455 550838
rect 552013 550835 552079 550838
rect 46105 549810 46171 549813
rect 48086 549810 48146 550256
rect 407389 550218 407455 550221
rect 407389 550216 410044 550218
rect 407389 550160 407394 550216
rect 407450 550160 410044 550216
rect 407389 550158 410044 550160
rect 407389 550155 407455 550158
rect 46105 549808 48146 549810
rect 46105 549752 46110 549808
rect 46166 549752 48146 549808
rect 46105 549750 48146 549752
rect 46105 549747 46171 549750
rect 553301 549538 553367 549541
rect 549884 549536 553367 549538
rect 549884 549480 553306 549536
rect 553362 549480 553367 549536
rect 549884 549478 553367 549480
rect 553301 549475 553367 549478
rect 350165 548994 350231 548997
rect 347852 548992 350231 548994
rect 347852 548936 350170 548992
rect 350226 548936 350231 548992
rect 347852 548934 350231 548936
rect 350165 548931 350231 548934
rect 46105 548314 46171 548317
rect 48086 548314 48146 548896
rect 407481 548858 407547 548861
rect 407481 548856 410044 548858
rect 407481 548800 407486 548856
rect 407542 548800 410044 548856
rect 407481 548798 410044 548800
rect 407481 548795 407547 548798
rect 46105 548312 48146 548314
rect 46105 548256 46110 548312
rect 46166 548256 48146 548312
rect 46105 548254 48146 548256
rect 46105 548251 46171 548254
rect 347822 547090 347882 547536
rect 407389 547498 407455 547501
rect 552105 547498 552171 547501
rect 407389 547496 410044 547498
rect 407389 547440 407394 547496
rect 407450 547440 410044 547496
rect 407389 547438 410044 547440
rect 549884 547496 552171 547498
rect 549884 547440 552110 547496
rect 552166 547440 552171 547496
rect 549884 547438 552171 547440
rect 407389 547435 407455 547438
rect 552105 547435 552171 547438
rect 350257 547090 350323 547093
rect 347822 547088 350323 547090
rect 347822 547032 350262 547088
rect 350318 547032 350323 547088
rect 347822 547030 350323 547032
rect 350257 547027 350323 547030
rect 37590 546484 37596 546548
rect 37660 546546 37666 546548
rect 48086 546546 48146 546856
rect 347822 546682 347882 546856
rect 560886 546818 560892 546820
rect 549884 546758 560892 546818
rect 560886 546756 560892 546758
rect 560956 546756 560962 546820
rect 350441 546682 350507 546685
rect 347822 546680 350507 546682
rect 347822 546624 350446 546680
rect 350502 546624 350507 546680
rect 347822 546622 350507 546624
rect 350441 546619 350507 546622
rect 37660 546486 48146 546546
rect 37660 546484 37666 546486
rect 46749 545730 46815 545733
rect 48086 545730 48146 546176
rect 408309 546138 408375 546141
rect 408309 546136 410044 546138
rect 408309 546080 408314 546136
rect 408370 546080 410044 546136
rect 408309 546078 410044 546080
rect 408309 546075 408375 546078
rect 46749 545728 48146 545730
rect 46749 545672 46754 545728
rect 46810 545672 48146 545728
rect 46749 545670 48146 545672
rect 46749 545667 46815 545670
rect 552105 545458 552171 545461
rect 549884 545456 552171 545458
rect 549884 545400 552110 545456
rect 552166 545400 552171 545456
rect 549884 545398 552171 545400
rect 552105 545395 552171 545398
rect 46749 544370 46815 544373
rect 48086 544370 48146 544816
rect 407389 544778 407455 544781
rect 574318 544778 574324 544780
rect 407389 544776 410044 544778
rect 407389 544720 407394 544776
rect 407450 544720 410044 544776
rect 407389 544718 410044 544720
rect 549884 544718 574324 544778
rect 407389 544715 407455 544718
rect 574318 544716 574324 544718
rect 574388 544716 574394 544780
rect 46749 544368 48146 544370
rect 46749 544312 46754 544368
rect 46810 544312 48146 544368
rect 46749 544310 48146 544312
rect 46749 544307 46815 544310
rect 46105 544234 46171 544237
rect 46105 544232 48116 544234
rect 46105 544176 46110 544232
rect 46166 544176 48116 544232
rect 46105 544174 48116 544176
rect 46105 544171 46171 544174
rect 407481 544098 407547 544101
rect 552565 544098 552631 544101
rect 407481 544096 410044 544098
rect 407481 544040 407486 544096
rect 407542 544040 410044 544096
rect 407481 544038 410044 544040
rect 549884 544096 552631 544098
rect 549884 544040 552570 544096
rect 552626 544040 552631 544096
rect 549884 544038 552631 544040
rect 407481 544035 407547 544038
rect 552565 544035 552631 544038
rect 347822 543010 347882 543456
rect 350441 543010 350507 543013
rect 347822 543008 350507 543010
rect 347822 542952 350446 543008
rect 350502 542952 350507 543008
rect 347822 542950 350507 542952
rect 350441 542947 350507 542950
rect 407389 542058 407455 542061
rect 407389 542056 410044 542058
rect 407389 542000 407394 542056
rect 407450 542000 410044 542056
rect 407389 541998 410044 542000
rect 407389 541995 407455 541998
rect 349153 541514 349219 541517
rect 347852 541512 349219 541514
rect 347852 541456 349158 541512
rect 349214 541456 349219 541512
rect 347852 541454 349219 541456
rect 349153 541451 349219 541454
rect 46749 541106 46815 541109
rect 48086 541106 48146 541416
rect 46749 541104 48146 541106
rect 46749 541048 46754 541104
rect 46810 541048 48146 541104
rect 46749 541046 48146 541048
rect 46749 541043 46815 541046
rect 349061 540970 349127 540973
rect 349286 540970 349292 540972
rect 349061 540968 349292 540970
rect -960 540684 480 540924
rect 349061 540912 349066 540968
rect 349122 540912 349292 540968
rect 349061 540910 349292 540912
rect 349061 540907 349127 540910
rect 349286 540908 349292 540910
rect 349356 540908 349362 540972
rect 553117 540698 553183 540701
rect 549884 540696 553183 540698
rect 549884 540640 553122 540696
rect 553178 540640 553183 540696
rect 549884 540638 553183 540640
rect 553117 540635 553183 540638
rect 553301 540018 553367 540021
rect 549884 540016 553367 540018
rect 549884 539960 553306 540016
rect 553362 539960 553367 540016
rect 549884 539958 553367 539960
rect 553301 539955 553367 539958
rect 551093 539338 551159 539341
rect 549884 539336 551159 539338
rect 549884 539280 551098 539336
rect 551154 539280 551159 539336
rect 549884 539278 551159 539280
rect 551093 539275 551159 539278
rect 347822 538386 347882 538696
rect 350441 538386 350507 538389
rect 347822 538384 350507 538386
rect 347822 538328 350446 538384
rect 350502 538328 350507 538384
rect 347822 538326 350507 538328
rect 350441 538323 350507 538326
rect 46749 538114 46815 538117
rect 46749 538112 48116 538114
rect 46749 538056 46754 538112
rect 46810 538056 48116 538112
rect 46749 538054 48116 538056
rect 46749 538051 46815 538054
rect 405406 537916 405412 537980
rect 405476 537978 405482 537980
rect 405476 537918 410044 537978
rect 405476 537916 405482 537918
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect 347822 537162 347882 537336
rect 350441 537162 350507 537165
rect 347822 537160 350507 537162
rect 347822 537104 350446 537160
rect 350502 537104 350507 537160
rect 347822 537102 350507 537104
rect 350441 537099 350507 537102
rect 552381 536618 552447 536621
rect 550222 536616 552447 536618
rect 550222 536560 552386 536616
rect 552442 536560 552447 536616
rect 550222 536558 552447 536560
rect 550222 536550 550282 536558
rect 552381 536555 552447 536558
rect 549884 536490 550282 536550
rect 553301 535938 553367 535941
rect 549884 535936 553367 535938
rect 549884 535880 553306 535936
rect 553362 535880 553367 535936
rect 549884 535878 553367 535880
rect 553301 535875 553367 535878
rect 347822 534714 347882 535296
rect 407297 535258 407363 535261
rect 553301 535258 553367 535261
rect 407297 535256 410044 535258
rect 407297 535200 407302 535256
rect 407358 535200 410044 535256
rect 407297 535198 410044 535200
rect 549884 535256 553367 535258
rect 549884 535200 553306 535256
rect 553362 535200 553367 535256
rect 549884 535198 553367 535200
rect 407297 535195 407363 535198
rect 553301 535195 553367 535198
rect 350441 534714 350507 534717
rect 347822 534712 350507 534714
rect 347822 534656 350446 534712
rect 350502 534656 350507 534712
rect 347822 534654 350507 534656
rect 350441 534651 350507 534654
rect 35750 534108 35756 534172
rect 35820 534170 35826 534172
rect 48086 534170 48146 534616
rect 556470 534578 556476 534580
rect 549884 534518 556476 534578
rect 556470 534516 556476 534518
rect 556540 534516 556546 534580
rect 35820 534110 48146 534170
rect 35820 534108 35826 534110
rect 46749 533354 46815 533357
rect 48086 533354 48146 533936
rect 347822 533490 347882 533936
rect 407297 533898 407363 533901
rect 552565 533898 552631 533901
rect 407297 533896 410044 533898
rect 407297 533840 407302 533896
rect 407358 533840 410044 533896
rect 407297 533838 410044 533840
rect 549884 533896 552631 533898
rect 549884 533840 552570 533896
rect 552626 533840 552631 533896
rect 549884 533838 552631 533840
rect 407297 533835 407363 533838
rect 552565 533835 552631 533838
rect 350257 533490 350323 533493
rect 347822 533488 350323 533490
rect 347822 533432 350262 533488
rect 350318 533432 350323 533488
rect 347822 533430 350323 533432
rect 350257 533427 350323 533430
rect 46749 533352 48146 533354
rect 46749 533296 46754 533352
rect 46810 533296 48146 533352
rect 46749 533294 48146 533296
rect 46749 533291 46815 533294
rect 347822 533082 347882 533256
rect 350441 533082 350507 533085
rect 347822 533080 350507 533082
rect 347822 533024 350446 533080
rect 350502 533024 350507 533080
rect 347822 533022 350507 533024
rect 350441 533019 350507 533022
rect 46749 532130 46815 532133
rect 48086 532130 48146 532576
rect 46749 532128 48146 532130
rect 46749 532072 46754 532128
rect 46810 532072 48146 532128
rect 46749 532070 48146 532072
rect 347822 532130 347882 532576
rect 552381 532538 552447 532541
rect 549884 532536 552447 532538
rect 549884 532480 552386 532536
rect 552442 532480 552447 532536
rect 549884 532478 552447 532480
rect 552381 532475 552447 532478
rect 350441 532130 350507 532133
rect 347822 532128 350507 532130
rect 347822 532072 350446 532128
rect 350502 532072 350507 532128
rect 347822 532070 350507 532072
rect 46749 532067 46815 532070
rect 350441 532067 350507 532070
rect 407297 531858 407363 531861
rect 557942 531858 557948 531860
rect 407297 531856 410044 531858
rect 407297 531800 407302 531856
rect 407358 531800 410044 531856
rect 407297 531798 410044 531800
rect 549884 531798 557948 531858
rect 407297 531795 407363 531798
rect 557942 531796 557948 531798
rect 558012 531796 558018 531860
rect 44030 530708 44036 530772
rect 44100 530770 44106 530772
rect 48086 530770 48146 531216
rect 44100 530710 48146 530770
rect 347822 530770 347882 531216
rect 553301 531178 553367 531181
rect 549884 531176 553367 531178
rect 549884 531120 553306 531176
rect 553362 531120 553367 531176
rect 549884 531118 553367 531120
rect 553301 531115 553367 531118
rect 350441 530770 350507 530773
rect 347822 530768 350507 530770
rect 347822 530712 350446 530768
rect 350502 530712 350507 530768
rect 347822 530710 350507 530712
rect 44100 530708 44106 530710
rect 350441 530707 350507 530710
rect 552381 530498 552447 530501
rect 549884 530496 552447 530498
rect 549884 530440 552386 530496
rect 552442 530440 552447 530496
rect 549884 530438 552447 530440
rect 552381 530435 552447 530438
rect 46749 529954 46815 529957
rect 46749 529952 48116 529954
rect 46749 529896 46754 529952
rect 46810 529896 48116 529952
rect 46749 529894 48116 529896
rect 46749 529891 46815 529894
rect 46105 529002 46171 529005
rect 48086 529002 48146 529176
rect 407614 529076 407620 529140
rect 407684 529138 407690 529140
rect 407684 529078 410044 529138
rect 407684 529076 407690 529078
rect 46105 529000 48146 529002
rect 46105 528944 46110 529000
rect 46166 528944 48146 529000
rect 46105 528942 48146 528944
rect 46105 528939 46171 528942
rect 553301 528458 553367 528461
rect 549884 528456 553367 528458
rect 549884 528400 553306 528456
rect 553362 528400 553367 528456
rect 549884 528398 553367 528400
rect 553301 528395 553367 528398
rect -960 527764 480 528004
rect 35566 527308 35572 527372
rect 35636 527370 35642 527372
rect 48086 527370 48146 527816
rect 35636 527310 48146 527370
rect 35636 527308 35642 527310
rect 39798 527172 39804 527236
rect 39868 527234 39874 527236
rect 350441 527234 350507 527237
rect 39868 527174 48116 527234
rect 347852 527232 350507 527234
rect 347852 527176 350446 527232
rect 350502 527176 350507 527232
rect 347852 527174 350507 527176
rect 39868 527172 39874 527174
rect 350441 527171 350507 527174
rect 358118 527036 358124 527100
rect 358188 527098 358194 527100
rect 358188 527038 410044 527098
rect 358188 527036 358194 527038
rect 46289 526554 46355 526557
rect 46289 526552 48116 526554
rect 46289 526496 46294 526552
rect 46350 526496 48116 526552
rect 46289 526494 48116 526496
rect 46289 526491 46355 526494
rect 347822 526282 347882 526456
rect 552381 526418 552447 526421
rect 549884 526416 552447 526418
rect 549884 526360 552386 526416
rect 552442 526360 552447 526416
rect 549884 526358 552447 526360
rect 552381 526355 552447 526358
rect 350441 526282 350507 526285
rect 347822 526280 350507 526282
rect 347822 526224 350446 526280
rect 350502 526224 350507 526280
rect 347822 526222 350507 526224
rect 350441 526219 350507 526222
rect 407113 525738 407179 525741
rect 552289 525738 552355 525741
rect 407113 525736 410044 525738
rect 407113 525680 407118 525736
rect 407174 525680 410044 525736
rect 407113 525678 410044 525680
rect 549884 525736 552355 525738
rect 549884 525680 552294 525736
rect 552350 525680 552355 525736
rect 549884 525678 552355 525680
rect 407113 525675 407179 525678
rect 552289 525675 552355 525678
rect 46749 525194 46815 525197
rect 46749 525192 48116 525194
rect 46749 525136 46754 525192
rect 46810 525136 48116 525192
rect 46749 525134 48116 525136
rect 46749 525131 46815 525134
rect 407297 525058 407363 525061
rect 407297 525056 410044 525058
rect 407297 525000 407302 525056
rect 407358 525000 410044 525056
rect 407297 524998 410044 525000
rect 407297 524995 407363 524998
rect 47393 524650 47459 524653
rect 47894 524650 47900 524652
rect 47393 524648 47900 524650
rect 47393 524592 47398 524648
rect 47454 524592 47900 524648
rect 47393 524590 47900 524592
rect 47393 524587 47459 524590
rect 47894 524588 47900 524590
rect 47964 524588 47970 524652
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 552473 524378 552539 524381
rect 549884 524376 552539 524378
rect 549884 524320 552478 524376
rect 552534 524320 552539 524376
rect 583520 524364 584960 524454
rect 549884 524318 552539 524320
rect 552473 524315 552539 524318
rect 347822 523290 347882 523736
rect 407297 523698 407363 523701
rect 407297 523696 410044 523698
rect 407297 523640 407302 523696
rect 407358 523640 410044 523696
rect 407297 523638 410044 523640
rect 407297 523635 407363 523638
rect 350441 523290 350507 523293
rect 347822 523288 350507 523290
rect 347822 523232 350446 523288
rect 350502 523232 350507 523288
rect 347822 523230 350507 523232
rect 350441 523227 350507 523230
rect 350257 523154 350323 523157
rect 347852 523152 350323 523154
rect 347852 523096 350262 523152
rect 350318 523096 350323 523152
rect 347852 523094 350323 523096
rect 350257 523091 350323 523094
rect 348417 523018 348483 523021
rect 350574 523018 350580 523020
rect 348417 523016 350580 523018
rect 348417 522960 348422 523016
rect 348478 522960 350580 523016
rect 348417 522958 350580 522960
rect 348417 522955 348483 522958
rect 350574 522956 350580 522958
rect 350644 522956 350650 523020
rect 407389 523018 407455 523021
rect 407389 523016 410044 523018
rect 407389 522960 407394 523016
rect 407450 522960 410044 523016
rect 407389 522958 410044 522960
rect 407389 522955 407455 522958
rect 407113 522338 407179 522341
rect 552013 522338 552079 522341
rect 407113 522336 410044 522338
rect 407113 522280 407118 522336
rect 407174 522280 410044 522336
rect 407113 522278 410044 522280
rect 549884 522336 552079 522338
rect 549884 522280 552018 522336
rect 552074 522280 552079 522336
rect 549884 522278 552079 522280
rect 407113 522275 407179 522278
rect 552013 522275 552079 522278
rect 45737 521794 45803 521797
rect 349889 521794 349955 521797
rect 45737 521792 48116 521794
rect 45737 521736 45742 521792
rect 45798 521736 48116 521792
rect 45737 521734 48116 521736
rect 347852 521792 349955 521794
rect 347852 521736 349894 521792
rect 349950 521736 349955 521792
rect 347852 521734 349955 521736
rect 45737 521731 45803 521734
rect 349889 521731 349955 521734
rect 391238 521596 391244 521660
rect 391308 521658 391314 521660
rect 552013 521658 552079 521661
rect 391308 521598 410044 521658
rect 549884 521656 552079 521658
rect 549884 521600 552018 521656
rect 552074 521600 552079 521656
rect 549884 521598 552079 521600
rect 391308 521596 391314 521598
rect 552013 521595 552079 521598
rect 45645 520706 45711 520709
rect 48086 520706 48146 521016
rect 552422 520978 552428 520980
rect 549884 520918 552428 520978
rect 552422 520916 552428 520918
rect 552492 520916 552498 520980
rect 45645 520704 48146 520706
rect 45645 520648 45650 520704
rect 45706 520648 48146 520704
rect 45645 520646 48146 520648
rect 45645 520643 45711 520646
rect 45553 520434 45619 520437
rect 350165 520434 350231 520437
rect 45553 520432 48116 520434
rect 45553 520376 45558 520432
rect 45614 520376 48116 520432
rect 45553 520374 48116 520376
rect 347852 520432 350231 520434
rect 347852 520376 350170 520432
rect 350226 520376 350231 520432
rect 347852 520374 350231 520376
rect 45553 520371 45619 520374
rect 350165 520371 350231 520374
rect 549884 519490 550282 519550
rect 550222 519482 550282 519490
rect 552013 519482 552079 519485
rect 550222 519480 552079 519482
rect 550222 519424 552018 519480
rect 552074 519424 552079 519480
rect 550222 519422 552079 519424
rect 552013 519419 552079 519422
rect 347822 518938 347882 518976
rect 353518 518938 353524 518940
rect 347822 518878 353524 518938
rect 353518 518876 353524 518878
rect 353588 518876 353594 518940
rect 552013 518938 552079 518941
rect 549884 518936 552079 518938
rect 549884 518880 552018 518936
rect 552074 518880 552079 518936
rect 549884 518878 552079 518880
rect 552013 518875 552079 518878
rect 407297 518258 407363 518261
rect 407297 518256 410044 518258
rect 407297 518200 407302 518256
rect 407358 518200 410044 518256
rect 407297 518198 410044 518200
rect 407297 518195 407363 518198
rect 350441 517714 350507 517717
rect 347852 517712 350507 517714
rect 347852 517656 350446 517712
rect 350502 517656 350507 517712
rect 347852 517654 350507 517656
rect 350441 517651 350507 517654
rect 407113 517578 407179 517581
rect 407113 517576 410044 517578
rect 407113 517520 407118 517576
rect 407174 517520 410044 517576
rect 407113 517518 410044 517520
rect 407113 517515 407179 517518
rect 45553 516626 45619 516629
rect 48086 516626 48146 516936
rect 45553 516624 48146 516626
rect 45553 516568 45558 516624
rect 45614 516568 48146 516624
rect 45553 516566 48146 516568
rect 347822 516626 347882 516936
rect 407297 516898 407363 516901
rect 552013 516898 552079 516901
rect 407297 516896 410044 516898
rect 407297 516840 407302 516896
rect 407358 516840 410044 516896
rect 407297 516838 410044 516840
rect 549884 516896 552079 516898
rect 549884 516840 552018 516896
rect 552074 516840 552079 516896
rect 549884 516838 552079 516840
rect 407297 516835 407363 516838
rect 552013 516835 552079 516838
rect 350257 516626 350323 516629
rect 347822 516624 350323 516626
rect 347822 516568 350262 516624
rect 350318 516568 350323 516624
rect 347822 516566 350323 516568
rect 45553 516563 45619 516566
rect 350257 516563 350323 516566
rect 347822 516218 347882 516256
rect 350441 516218 350507 516221
rect 347822 516216 350507 516218
rect 347822 516160 350446 516216
rect 350502 516160 350507 516216
rect 347822 516158 350507 516160
rect 350441 516155 350507 516158
rect 407113 516218 407179 516221
rect 407113 516216 410044 516218
rect 407113 516160 407118 516216
rect 407174 516160 410044 516216
rect 407113 516158 410044 516160
rect 407113 516155 407179 516158
rect 45553 515266 45619 515269
rect 48086 515266 48146 515576
rect 552381 515538 552447 515541
rect 549884 515536 552447 515538
rect 549884 515480 552386 515536
rect 552442 515480 552447 515536
rect 549884 515478 552447 515480
rect 552381 515475 552447 515478
rect 45553 515264 48146 515266
rect 45553 515208 45558 515264
rect 45614 515208 48146 515264
rect 45553 515206 48146 515208
rect 45553 515203 45619 515206
rect -960 514858 480 514948
rect 36670 514932 36676 514996
rect 36740 514994 36746 514996
rect 36740 514934 48116 514994
rect 36740 514932 36746 514934
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 407573 514858 407639 514861
rect 552013 514858 552079 514861
rect 407573 514856 410044 514858
rect 407573 514800 407578 514856
rect 407634 514800 410044 514856
rect 407573 514798 410044 514800
rect 549884 514856 552079 514858
rect 549884 514800 552018 514856
rect 552074 514800 552079 514856
rect 549884 514798 552079 514800
rect 407573 514795 407639 514798
rect 552013 514795 552079 514798
rect 46197 513906 46263 513909
rect 48086 513906 48146 514216
rect 46197 513904 48146 513906
rect 46197 513848 46202 513904
rect 46258 513848 48146 513904
rect 46197 513846 48146 513848
rect 46197 513843 46263 513846
rect 347822 513770 347882 514216
rect 350441 513770 350507 513773
rect 347822 513768 350507 513770
rect 347822 513712 350446 513768
rect 350502 513712 350507 513768
rect 347822 513710 350507 513712
rect 350441 513707 350507 513710
rect 347822 513498 347882 513536
rect 350257 513498 350323 513501
rect 347822 513496 350323 513498
rect 347822 513440 350262 513496
rect 350318 513440 350323 513496
rect 347822 513438 350323 513440
rect 350257 513435 350323 513438
rect 407113 512818 407179 512821
rect 407113 512816 410044 512818
rect 407113 512760 407118 512816
rect 407174 512760 410044 512816
rect 407113 512758 410044 512760
rect 407113 512755 407179 512758
rect 407113 512138 407179 512141
rect 407113 512136 410044 512138
rect 407113 512080 407118 512136
rect 407174 512080 410044 512136
rect 407113 512078 410044 512080
rect 407113 512075 407179 512078
rect 348049 512002 348115 512005
rect 348366 512002 348372 512004
rect 348049 512000 348372 512002
rect 348049 511944 348054 512000
rect 348110 511944 348372 512000
rect 348049 511942 348372 511944
rect 348049 511939 348115 511942
rect 348366 511940 348372 511942
rect 348436 511940 348442 512004
rect 348601 511594 348667 511597
rect 347852 511592 348667 511594
rect 347852 511536 348606 511592
rect 348662 511536 348667 511592
rect 347852 511534 348667 511536
rect 348601 511531 348667 511534
rect 583520 511172 584960 511412
rect 46013 510914 46079 510917
rect 46013 510912 48116 510914
rect 46013 510856 46018 510912
rect 46074 510856 48116 510912
rect 46013 510854 48116 510856
rect 46013 510851 46079 510854
rect 387006 510716 387012 510780
rect 387076 510778 387082 510780
rect 387076 510718 410044 510778
rect 387076 510716 387082 510718
rect 409045 510098 409111 510101
rect 553301 510098 553367 510101
rect 409045 510096 410044 510098
rect 409045 510040 409050 510096
rect 409106 510040 410044 510096
rect 409045 510038 410044 510040
rect 549884 510096 553367 510098
rect 549884 510040 553306 510096
rect 553362 510040 553367 510096
rect 549884 510038 553367 510040
rect 409045 510035 409111 510038
rect 553301 510035 553367 510038
rect 46749 509554 46815 509557
rect 46749 509552 48116 509554
rect 46749 509496 46754 509552
rect 46810 509496 48116 509552
rect 46749 509494 48116 509496
rect 46749 509491 46815 509494
rect 407113 509418 407179 509421
rect 407113 509416 410044 509418
rect 407113 509360 407118 509416
rect 407174 509360 410044 509416
rect 407113 509358 410044 509360
rect 407113 509355 407179 509358
rect 350441 508874 350507 508877
rect 347852 508872 350507 508874
rect 347852 508816 350446 508872
rect 350502 508816 350507 508872
rect 347852 508814 350507 508816
rect 350441 508811 350507 508814
rect 347822 507922 347882 508096
rect 407757 508058 407823 508061
rect 407757 508056 410044 508058
rect 407757 508000 407762 508056
rect 407818 508000 410044 508056
rect 407757 507998 410044 508000
rect 407757 507995 407823 507998
rect 350574 507922 350580 507924
rect 347822 507862 350580 507922
rect 350574 507860 350580 507862
rect 350644 507860 350650 507924
rect 41086 506908 41092 506972
rect 41156 506970 41162 506972
rect 48086 506970 48146 507416
rect 41156 506910 48146 506970
rect 347822 506970 347882 507416
rect 550633 507378 550699 507381
rect 549884 507376 550699 507378
rect 549884 507320 550638 507376
rect 550694 507320 550699 507376
rect 549884 507318 550699 507320
rect 550633 507315 550699 507318
rect 350441 506970 350507 506973
rect 347822 506968 350507 506970
rect 347822 506912 350446 506968
rect 350502 506912 350507 506968
rect 347822 506910 350507 506912
rect 41156 506908 41162 506910
rect 350441 506907 350507 506910
rect 356830 506636 356836 506700
rect 356900 506698 356906 506700
rect 356900 506638 410044 506698
rect 356900 506636 356906 506638
rect 347822 505610 347882 506056
rect 554814 506018 554820 506020
rect 549884 505958 554820 506018
rect 554814 505956 554820 505958
rect 554884 505956 554890 506020
rect 350441 505610 350507 505613
rect 347822 505608 350507 505610
rect 347822 505552 350446 505608
rect 350502 505552 350507 505608
rect 347822 505550 350507 505552
rect 350441 505547 350507 505550
rect 350257 505474 350323 505477
rect 347852 505472 350323 505474
rect 347852 505416 350262 505472
rect 350318 505416 350323 505472
rect 347852 505414 350323 505416
rect 350257 505411 350323 505414
rect 46749 505202 46815 505205
rect 48086 505202 48146 505376
rect 553301 505338 553367 505341
rect 549884 505336 553367 505338
rect 549884 505280 553306 505336
rect 553362 505280 553367 505336
rect 549884 505278 553367 505280
rect 553301 505275 553367 505278
rect 46749 505200 48146 505202
rect 46749 505144 46754 505200
rect 46810 505144 48146 505200
rect 46749 505142 48146 505144
rect 46749 505139 46815 505142
rect 553301 504658 553367 504661
rect 549884 504656 553367 504658
rect 549884 504600 553306 504656
rect 553362 504600 553367 504656
rect 549884 504598 553367 504600
rect 553301 504595 553367 504598
rect 47485 504114 47551 504117
rect 47485 504112 48116 504114
rect 47485 504056 47490 504112
rect 47546 504056 48116 504112
rect 47485 504054 48116 504056
rect 47485 504051 47551 504054
rect 347822 503842 347882 504016
rect 350441 503842 350507 503845
rect 347822 503840 350507 503842
rect 347822 503784 350446 503840
rect 350502 503784 350507 503840
rect 347822 503782 350507 503784
rect 350441 503779 350507 503782
rect 409462 502490 410044 502550
rect 549884 502490 550282 502550
rect 392526 502420 392532 502484
rect 392596 502482 392602 502484
rect 409462 502482 409522 502490
rect 392596 502422 409522 502482
rect 550222 502482 550282 502490
rect 553301 502482 553367 502485
rect 550222 502480 553367 502482
rect 550222 502424 553306 502480
rect 553362 502424 553367 502480
rect 550222 502422 553367 502424
rect 392596 502420 392602 502422
rect 553301 502419 553367 502422
rect 553301 501938 553367 501941
rect 549884 501936 553367 501938
rect -960 501802 480 501892
rect 549884 501880 553306 501936
rect 553362 501880 553367 501936
rect 549884 501878 553367 501880
rect 553301 501875 553367 501878
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 45829 501394 45895 501397
rect 45829 501392 48116 501394
rect 45829 501336 45834 501392
rect 45890 501336 48116 501392
rect 45829 501334 48116 501336
rect 45829 501331 45895 501334
rect 408309 501258 408375 501261
rect 553301 501258 553367 501261
rect 408309 501256 410044 501258
rect 408309 501200 408314 501256
rect 408370 501200 410044 501256
rect 408309 501198 410044 501200
rect 549884 501256 553367 501258
rect 549884 501200 553306 501256
rect 553362 501200 553367 501256
rect 549884 501198 553367 501200
rect 408309 501195 408375 501198
rect 553301 501195 553367 501198
rect 46749 500714 46815 500717
rect 46749 500712 48116 500714
rect 46749 500656 46754 500712
rect 46810 500656 48116 500712
rect 46749 500654 48116 500656
rect 46749 500651 46815 500654
rect 347822 500170 347882 500616
rect 407113 500578 407179 500581
rect 552289 500578 552355 500581
rect 407113 500576 410044 500578
rect 407113 500520 407118 500576
rect 407174 500520 410044 500576
rect 407113 500518 410044 500520
rect 549884 500576 552355 500578
rect 549884 500520 552294 500576
rect 552350 500520 552355 500576
rect 549884 500518 552355 500520
rect 407113 500515 407179 500518
rect 552289 500515 552355 500518
rect 350441 500170 350507 500173
rect 347822 500168 350507 500170
rect 347822 500112 350446 500168
rect 350502 500112 350507 500168
rect 347822 500110 350507 500112
rect 350441 500107 350507 500110
rect 349797 500034 349863 500037
rect 347852 500032 349863 500034
rect 347852 499976 349802 500032
rect 349858 499976 349863 500032
rect 347852 499974 349863 499976
rect 349797 499971 349863 499974
rect 38510 499700 38516 499764
rect 38580 499762 38586 499764
rect 48086 499762 48146 499936
rect 553301 499898 553367 499901
rect 549884 499896 553367 499898
rect 549884 499840 553306 499896
rect 553362 499840 553367 499896
rect 549884 499838 553367 499840
rect 553301 499835 553367 499838
rect 38580 499702 48146 499762
rect 38580 499700 38586 499702
rect 40718 498748 40724 498812
rect 40788 498810 40794 498812
rect 48086 498810 48146 499256
rect 40788 498750 48146 498810
rect 40788 498748 40794 498750
rect 347822 498266 347882 498576
rect 553301 498538 553367 498541
rect 549884 498536 553367 498538
rect 549884 498480 553306 498536
rect 553362 498480 553367 498536
rect 549884 498478 553367 498480
rect 553301 498475 553367 498478
rect 350441 498266 350507 498269
rect 347822 498264 350507 498266
rect 347822 498208 350446 498264
rect 350502 498208 350507 498264
rect 347822 498206 350507 498208
rect 350441 498203 350507 498206
rect 583520 497844 584960 498084
rect 45829 497314 45895 497317
rect 45829 497312 48116 497314
rect 45829 497256 45834 497312
rect 45890 497256 48116 497312
rect 45829 497254 48116 497256
rect 45829 497251 45895 497254
rect 407113 497178 407179 497181
rect 558126 497178 558132 497180
rect 407113 497176 410044 497178
rect 407113 497120 407118 497176
rect 407174 497120 410044 497176
rect 407113 497118 410044 497120
rect 549884 497118 558132 497178
rect 407113 497115 407179 497118
rect 558126 497116 558132 497118
rect 558196 497116 558202 497180
rect 46381 496090 46447 496093
rect 48086 496090 48146 496536
rect 553485 496498 553551 496501
rect 549884 496496 553551 496498
rect 549884 496440 553490 496496
rect 553546 496440 553551 496496
rect 549884 496438 553551 496440
rect 553485 496435 553551 496438
rect 46381 496088 48146 496090
rect 46381 496032 46386 496088
rect 46442 496032 48146 496088
rect 46381 496030 48146 496032
rect 46381 496027 46447 496030
rect 46749 495954 46815 495957
rect 46749 495952 48116 495954
rect 46749 495896 46754 495952
rect 46810 495896 48116 495952
rect 46749 495894 48116 495896
rect 46749 495891 46815 495894
rect 347822 495546 347882 495856
rect 407113 495818 407179 495821
rect 550357 495818 550423 495821
rect 407113 495816 410044 495818
rect 407113 495760 407118 495816
rect 407174 495760 410044 495816
rect 407113 495758 410044 495760
rect 549884 495816 550423 495818
rect 549884 495760 550362 495816
rect 550418 495760 550423 495816
rect 549884 495758 550423 495760
rect 407113 495755 407179 495758
rect 550357 495755 550423 495758
rect 350441 495546 350507 495549
rect 347822 495544 350507 495546
rect 347822 495488 350446 495544
rect 350502 495488 350507 495544
rect 347822 495486 350507 495488
rect 350441 495483 350507 495486
rect 46749 495274 46815 495277
rect 46749 495272 48116 495274
rect 46749 495216 46754 495272
rect 46810 495216 48116 495272
rect 46749 495214 48116 495216
rect 46749 495211 46815 495214
rect 46013 494594 46079 494597
rect 347822 494594 347882 495176
rect 350758 494594 350764 494596
rect 46013 494592 48116 494594
rect 46013 494536 46018 494592
rect 46074 494536 48116 494592
rect 46013 494534 48116 494536
rect 347822 494534 350764 494594
rect 46013 494531 46079 494534
rect 350758 494532 350764 494534
rect 350828 494532 350834 494596
rect 556654 494458 556660 494460
rect 549884 494398 556660 494458
rect 556654 494396 556660 494398
rect 556724 494396 556730 494460
rect 349429 493914 349495 493917
rect 347852 493912 349495 493914
rect 347852 493856 349434 493912
rect 349490 493856 349495 493912
rect 347852 493854 349495 493856
rect 349429 493851 349495 493854
rect 46749 493234 46815 493237
rect 48086 493234 48146 493816
rect 552657 493778 552723 493781
rect 549884 493776 552723 493778
rect 549884 493720 552662 493776
rect 552718 493720 552723 493776
rect 549884 493718 552723 493720
rect 552657 493715 552723 493718
rect 46749 493232 48146 493234
rect 46749 493176 46754 493232
rect 46810 493176 48146 493232
rect 46749 493174 48146 493176
rect 46749 493171 46815 493174
rect 407113 493098 407179 493101
rect 553117 493098 553183 493101
rect 407113 493096 410044 493098
rect 407113 493040 407118 493096
rect 407174 493040 410044 493096
rect 407113 493038 410044 493040
rect 549884 493096 553183 493098
rect 549884 493040 553122 493096
rect 553178 493040 553183 493096
rect 549884 493038 553183 493040
rect 407113 493035 407179 493038
rect 553117 493035 553183 493038
rect 347822 492010 347882 492456
rect 552565 492418 552631 492421
rect 549884 492416 552631 492418
rect 549884 492360 552570 492416
rect 552626 492360 552631 492416
rect 549884 492358 552631 492360
rect 552565 492355 552631 492358
rect 350257 492010 350323 492013
rect 347822 492008 350323 492010
rect 347822 491952 350262 492008
rect 350318 491952 350323 492008
rect 347822 491950 350323 491952
rect 350257 491947 350323 491950
rect 347822 491466 347882 491776
rect 553526 491738 553532 491740
rect 549884 491678 553532 491738
rect 553526 491676 553532 491678
rect 553596 491676 553602 491740
rect 350441 491466 350507 491469
rect 347822 491464 350507 491466
rect 347822 491408 350446 491464
rect 350502 491408 350507 491464
rect 347822 491406 350507 491408
rect 350441 491403 350507 491406
rect 46749 490650 46815 490653
rect 48086 490650 48146 491096
rect 46749 490648 48146 490650
rect 46749 490592 46754 490648
rect 46810 490592 48146 490648
rect 46749 490590 48146 490592
rect 347822 490650 347882 491096
rect 407113 491058 407179 491061
rect 407113 491056 410044 491058
rect 407113 491000 407118 491056
rect 407174 491000 410044 491056
rect 407113 490998 410044 491000
rect 407113 490995 407179 490998
rect 350441 490650 350507 490653
rect 347822 490648 350507 490650
rect 347822 490592 350446 490648
rect 350502 490592 350507 490648
rect 347822 490590 350507 490592
rect 46749 490587 46815 490590
rect 350441 490587 350507 490590
rect 46381 489970 46447 489973
rect 48086 489970 48146 490416
rect 347822 490242 347882 490416
rect 350257 490242 350323 490245
rect 347822 490240 350323 490242
rect 347822 490184 350262 490240
rect 350318 490184 350323 490240
rect 347822 490182 350323 490184
rect 350257 490179 350323 490182
rect 46381 489968 48146 489970
rect 46381 489912 46386 489968
rect 46442 489912 48146 489968
rect 46381 489910 48146 489912
rect 46381 489907 46447 489910
rect 46749 489834 46815 489837
rect 350165 489834 350231 489837
rect 46749 489832 48116 489834
rect 46749 489776 46754 489832
rect 46810 489776 48116 489832
rect 46749 489774 48116 489776
rect 347852 489832 350231 489834
rect 347852 489776 350170 489832
rect 350226 489776 350231 489832
rect 347852 489774 350231 489776
rect 46749 489771 46815 489774
rect 350165 489771 350231 489774
rect 407297 489698 407363 489701
rect 407297 489696 410044 489698
rect 407297 489640 407302 489696
rect 407358 489640 410044 489696
rect 407297 489638 410044 489640
rect 407297 489635 407363 489638
rect 407113 489018 407179 489021
rect 553301 489018 553367 489021
rect 407113 489016 410044 489018
rect 407113 488960 407118 489016
rect 407174 488960 410044 489016
rect 407113 488958 410044 488960
rect 549884 489016 553367 489018
rect 549884 488960 553306 489016
rect 553362 488960 553367 489016
rect 549884 488958 553367 488960
rect 407113 488955 407179 488958
rect 553301 488955 553367 488958
rect -960 488596 480 488836
rect 553301 488338 553367 488341
rect 549884 488336 553367 488338
rect 549884 488280 553306 488336
rect 553362 488280 553367 488336
rect 549884 488278 553367 488280
rect 553301 488275 553367 488278
rect 350257 487794 350323 487797
rect 347852 487792 350323 487794
rect 347852 487736 350262 487792
rect 350318 487736 350323 487792
rect 347852 487734 350323 487736
rect 350257 487731 350323 487734
rect 407113 487658 407179 487661
rect 407113 487656 410044 487658
rect 407113 487600 407118 487656
rect 407174 487600 410044 487656
rect 407113 487598 410044 487600
rect 407113 487595 407179 487598
rect 348366 487188 348372 487252
rect 348436 487250 348442 487252
rect 353937 487250 354003 487253
rect 348436 487248 354003 487250
rect 348436 487192 353942 487248
rect 353998 487192 354003 487248
rect 348436 487190 354003 487192
rect 348436 487188 348442 487190
rect 353937 487187 354003 487190
rect 44766 486508 44772 486572
rect 44836 486570 44842 486572
rect 48086 486570 48146 487016
rect 407113 486978 407179 486981
rect 407113 486976 410044 486978
rect 407113 486920 407118 486976
rect 407174 486920 410044 486976
rect 407113 486918 410044 486920
rect 407113 486915 407179 486918
rect 44836 486510 48146 486570
rect 44836 486508 44842 486510
rect 46749 485890 46815 485893
rect 48086 485890 48146 486336
rect 46749 485888 48146 485890
rect 46749 485832 46754 485888
rect 46810 485832 48146 485888
rect 46749 485830 48146 485832
rect 46749 485827 46815 485830
rect 41822 485148 41828 485212
rect 41892 485210 41898 485212
rect 48086 485210 48146 485656
rect 41892 485150 48146 485210
rect 347822 485210 347882 485656
rect 407021 485618 407087 485621
rect 407021 485616 410044 485618
rect 407021 485560 407026 485616
rect 407082 485560 410044 485616
rect 407021 485558 410044 485560
rect 407021 485555 407087 485558
rect 349981 485210 350047 485213
rect 347822 485208 350047 485210
rect 347822 485152 349986 485208
rect 350042 485152 350047 485208
rect 347822 485150 350047 485152
rect 41892 485148 41898 485150
rect 349981 485147 350047 485150
rect 46749 484802 46815 484805
rect 48086 484802 48146 484976
rect 407113 484938 407179 484941
rect 551553 484938 551619 484941
rect 407113 484936 410044 484938
rect 407113 484880 407118 484936
rect 407174 484880 410044 484936
rect 407113 484878 410044 484880
rect 549884 484936 551619 484938
rect 549884 484880 551558 484936
rect 551614 484880 551619 484936
rect 549884 484878 551619 484880
rect 407113 484875 407179 484878
rect 551553 484875 551619 484878
rect 46749 484800 48146 484802
rect 46749 484744 46754 484800
rect 46810 484744 48146 484800
rect 46749 484742 48146 484744
rect 46749 484739 46815 484742
rect 580349 484666 580415 484669
rect 583520 484666 584960 484756
rect 580349 484664 584960 484666
rect 580349 484608 580354 484664
rect 580410 484608 584960 484664
rect 580349 484606 584960 484608
rect 580349 484603 580415 484606
rect 583520 484516 584960 484606
rect 407113 484258 407179 484261
rect 552657 484258 552723 484261
rect 407113 484256 410044 484258
rect 407113 484200 407118 484256
rect 407174 484200 410044 484256
rect 407113 484198 410044 484200
rect 549884 484256 552723 484258
rect 549884 484200 552662 484256
rect 552718 484200 552723 484256
rect 549884 484198 552723 484200
rect 407113 484195 407179 484198
rect 552657 484195 552723 484198
rect 46749 483442 46815 483445
rect 48086 483442 48146 483616
rect 46749 483440 48146 483442
rect 46749 483384 46754 483440
rect 46810 483384 48146 483440
rect 46749 483382 48146 483384
rect 347822 483442 347882 483616
rect 407021 483578 407087 483581
rect 407021 483576 410044 483578
rect 407021 483520 407026 483576
rect 407082 483520 410044 483576
rect 407021 483518 410044 483520
rect 407021 483515 407087 483518
rect 350257 483442 350323 483445
rect 347822 483440 350323 483442
rect 347822 483384 350262 483440
rect 350318 483384 350323 483440
rect 347822 483382 350323 483384
rect 46749 483379 46815 483382
rect 350257 483379 350323 483382
rect 349102 483034 349108 483036
rect 347852 482974 349108 483034
rect 349102 482972 349108 482974
rect 349172 482972 349178 483036
rect 46473 482354 46539 482357
rect 46473 482352 48116 482354
rect 46473 482296 46478 482352
rect 46534 482296 48116 482352
rect 46473 482294 48116 482296
rect 46473 482291 46539 482294
rect 407113 482218 407179 482221
rect 407113 482216 410044 482218
rect 407113 482160 407118 482216
rect 407174 482160 410044 482216
rect 407113 482158 410044 482160
rect 407113 482155 407179 482158
rect 350441 481674 350507 481677
rect 347852 481672 350507 481674
rect 347852 481616 350446 481672
rect 350502 481616 350507 481672
rect 347852 481614 350507 481616
rect 350441 481611 350507 481614
rect 37038 480388 37044 480452
rect 37108 480450 37114 480452
rect 48086 480450 48146 480896
rect 347822 480722 347882 480896
rect 350257 480722 350323 480725
rect 347822 480720 350323 480722
rect 347822 480664 350262 480720
rect 350318 480664 350323 480720
rect 347822 480662 350323 480664
rect 350257 480659 350323 480662
rect 37108 480390 48146 480450
rect 37108 480388 37114 480390
rect 46657 480314 46723 480317
rect 350441 480314 350507 480317
rect 46657 480312 48116 480314
rect 46657 480256 46662 480312
rect 46718 480256 48116 480312
rect 46657 480254 48116 480256
rect 347852 480312 350507 480314
rect 347852 480256 350446 480312
rect 350502 480256 350507 480312
rect 347852 480254 350507 480256
rect 46657 480251 46723 480254
rect 350441 480251 350507 480254
rect 407113 480178 407179 480181
rect 552197 480178 552263 480181
rect 407113 480176 410044 480178
rect 407113 480120 407118 480176
rect 407174 480120 410044 480176
rect 407113 480118 410044 480120
rect 549884 480176 552263 480178
rect 549884 480120 552202 480176
rect 552258 480120 552263 480176
rect 549884 480118 552263 480120
rect 407113 480115 407179 480118
rect 552197 480115 552263 480118
rect 409229 479498 409295 479501
rect 559230 479498 559236 479500
rect 409229 479496 410044 479498
rect 409229 479440 409234 479496
rect 409290 479440 410044 479496
rect 409229 479438 410044 479440
rect 549884 479438 559236 479498
rect 409229 479435 409295 479438
rect 559230 479436 559236 479438
rect 559300 479436 559306 479500
rect 553301 478818 553367 478821
rect 549884 478816 553367 478818
rect 549884 478760 553306 478816
rect 553362 478760 553367 478816
rect 549884 478758 553367 478760
rect 553301 478755 553367 478758
rect 406929 478138 406995 478141
rect 406929 478136 410044 478138
rect 406929 478080 406934 478136
rect 406990 478080 410044 478136
rect 406929 478078 410044 478080
rect 406929 478075 406995 478078
rect 348325 477594 348391 477597
rect 347852 477592 348391 477594
rect 347852 477536 348330 477592
rect 348386 477536 348391 477592
rect 347852 477534 348391 477536
rect 348325 477531 348391 477534
rect 46749 476506 46815 476509
rect 48086 476506 48146 476816
rect 347822 476642 347882 476816
rect 409321 476778 409387 476781
rect 409321 476776 410044 476778
rect 409321 476720 409326 476776
rect 409382 476720 410044 476776
rect 409321 476718 410044 476720
rect 409321 476715 409387 476718
rect 350165 476642 350231 476645
rect 347822 476640 350231 476642
rect 347822 476584 350170 476640
rect 350226 476584 350231 476640
rect 347822 476582 350231 476584
rect 350165 476579 350231 476582
rect 46749 476504 48146 476506
rect 46749 476448 46754 476504
rect 46810 476448 48146 476504
rect 46749 476446 48146 476448
rect 46749 476443 46815 476446
rect 43846 476172 43852 476236
rect 43916 476234 43922 476236
rect 350257 476234 350323 476237
rect 43916 476174 48116 476234
rect 347852 476232 350323 476234
rect 347852 476176 350262 476232
rect 350318 476176 350323 476232
rect 347852 476174 350323 476176
rect 43916 476172 43922 476174
rect 350257 476171 350323 476174
rect 407297 476098 407363 476101
rect 552565 476098 552631 476101
rect 407297 476096 410044 476098
rect 407297 476040 407302 476096
rect 407358 476040 410044 476096
rect 407297 476038 410044 476040
rect 549884 476096 552631 476098
rect 549884 476040 552570 476096
rect 552626 476040 552631 476096
rect 549884 476038 552631 476040
rect 407297 476035 407363 476038
rect 552565 476035 552631 476038
rect -960 475540 480 475780
rect 46565 475554 46631 475557
rect 46565 475552 48116 475554
rect 46565 475496 46570 475552
rect 46626 475496 48116 475552
rect 46565 475494 48116 475496
rect 46565 475491 46631 475494
rect 347822 475010 347882 475456
rect 407113 475418 407179 475421
rect 553301 475418 553367 475421
rect 407113 475416 410044 475418
rect 407113 475360 407118 475416
rect 407174 475360 410044 475416
rect 407113 475358 410044 475360
rect 549884 475416 553367 475418
rect 549884 475360 553306 475416
rect 553362 475360 553367 475416
rect 549884 475358 553367 475360
rect 407113 475355 407179 475358
rect 553301 475355 553367 475358
rect 348693 475010 348759 475013
rect 347822 475008 348759 475010
rect 347822 474952 348698 475008
rect 348754 474952 348759 475008
rect 347822 474950 348759 474952
rect 348693 474947 348759 474950
rect 407297 474738 407363 474741
rect 407297 474736 410044 474738
rect 407297 474680 407302 474736
rect 407358 474680 410044 474736
rect 407297 474678 410044 474680
rect 407297 474675 407363 474678
rect 46105 474194 46171 474197
rect 46105 474192 48116 474194
rect 46105 474136 46110 474192
rect 46166 474136 48116 474192
rect 46105 474134 48116 474136
rect 46105 474131 46171 474134
rect 407113 474058 407179 474061
rect 407113 474056 410044 474058
rect 407113 474000 407118 474056
rect 407174 474000 410044 474056
rect 407113 473998 410044 474000
rect 407113 473995 407179 473998
rect 46565 473514 46631 473517
rect 350257 473514 350323 473517
rect 46565 473512 48116 473514
rect 46565 473456 46570 473512
rect 46626 473456 48116 473512
rect 46565 473454 48116 473456
rect 347852 473512 350323 473514
rect 347852 473456 350262 473512
rect 350318 473456 350323 473512
rect 347852 473454 350323 473456
rect 46565 473451 46631 473454
rect 350257 473451 350323 473454
rect 347822 472290 347882 472736
rect 565486 472698 565492 472700
rect 549884 472638 565492 472698
rect 565486 472636 565492 472638
rect 565556 472636 565562 472700
rect 350441 472290 350507 472293
rect 347822 472288 350507 472290
rect 347822 472232 350446 472288
rect 350502 472232 350507 472288
rect 347822 472230 350507 472232
rect 350441 472227 350507 472230
rect 409229 472018 409295 472021
rect 409229 472016 410044 472018
rect 409229 471960 409234 472016
rect 409290 471960 410044 472016
rect 409229 471958 410044 471960
rect 409229 471955 409295 471958
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 35382 470868 35388 470932
rect 35452 470930 35458 470932
rect 48086 470930 48146 471376
rect 583520 471324 584960 471414
rect 347773 471202 347839 471205
rect 347773 471200 347882 471202
rect 347773 471144 347778 471200
rect 347834 471144 347882 471200
rect 347773 471139 347882 471144
rect 35452 470870 48146 470930
rect 35452 470868 35458 470870
rect 347822 470764 347882 471139
rect 553301 470658 553367 470661
rect 549884 470656 553367 470658
rect 549884 470600 553306 470656
rect 553362 470600 553367 470656
rect 549884 470598 553367 470600
rect 553301 470595 553367 470598
rect 46749 469706 46815 469709
rect 48086 469706 48146 470016
rect 407113 469978 407179 469981
rect 553301 469978 553367 469981
rect 407113 469976 410044 469978
rect 407113 469920 407118 469976
rect 407174 469920 410044 469976
rect 407113 469918 410044 469920
rect 549884 469976 553367 469978
rect 549884 469920 553306 469976
rect 553362 469920 553367 469976
rect 549884 469918 553367 469920
rect 407113 469915 407179 469918
rect 553301 469915 553367 469918
rect 46749 469704 48146 469706
rect 46749 469648 46754 469704
rect 46810 469648 48146 469704
rect 46749 469646 48146 469648
rect 46749 469643 46815 469646
rect 349061 469298 349127 469301
rect 350942 469298 350948 469300
rect 349061 469296 350948 469298
rect 349061 469240 349066 469296
rect 349122 469240 350948 469296
rect 349061 469238 350948 469240
rect 349061 469235 349127 469238
rect 350942 469236 350948 469238
rect 351012 469236 351018 469300
rect 46565 468346 46631 468349
rect 48086 468346 48146 468656
rect 551001 468618 551067 468621
rect 550222 468616 551067 468618
rect 550222 468560 551006 468616
rect 551062 468560 551067 468616
rect 550222 468558 551067 468560
rect 550222 468550 550282 468558
rect 551001 468555 551067 468558
rect 46565 468344 48146 468346
rect 46565 468288 46570 468344
rect 46626 468288 48146 468344
rect 46565 468286 48146 468288
rect 46565 468283 46631 468286
rect 407113 468210 407179 468213
rect 410014 468210 410074 468520
rect 549884 468490 550282 468550
rect 407113 468208 410074 468210
rect 407113 468152 407118 468208
rect 407174 468152 410074 468208
rect 407113 468150 410074 468152
rect 407113 468147 407179 468150
rect 46749 468074 46815 468077
rect 46749 468072 48116 468074
rect 46749 468016 46754 468072
rect 46810 468016 48116 468072
rect 46749 468014 48116 468016
rect 46749 468011 46815 468014
rect 407297 467938 407363 467941
rect 407297 467936 410044 467938
rect 407297 467880 407302 467936
rect 407358 467880 410044 467936
rect 407297 467878 410044 467880
rect 407297 467875 407363 467878
rect 410014 466714 410074 467228
rect 407990 466654 410074 466714
rect 42006 466516 42012 466580
rect 42076 466578 42082 466580
rect 48086 466578 48146 466616
rect 42076 466518 48146 466578
rect 347822 466578 347882 466616
rect 350441 466578 350507 466581
rect 347822 466576 350507 466578
rect 347822 466520 350446 466576
rect 350502 466520 350507 466576
rect 347822 466518 350507 466520
rect 42076 466516 42082 466518
rect 350441 466515 350507 466518
rect 407990 466442 408050 466654
rect 408217 466578 408283 466581
rect 553301 466578 553367 466581
rect 408217 466576 410044 466578
rect 408217 466520 408222 466576
rect 408278 466520 410044 466576
rect 408217 466518 410044 466520
rect 549884 466576 553367 466578
rect 549884 466520 553306 466576
rect 553362 466520 553367 466576
rect 549884 466518 553367 466520
rect 408217 466515 408283 466518
rect 553301 466515 553367 466518
rect 408217 466442 408283 466445
rect 407990 466440 408283 466442
rect 407990 466384 408222 466440
rect 408278 466384 408283 466440
rect 407990 466382 408283 466384
rect 408217 466379 408283 466382
rect 350257 466034 350323 466037
rect 347852 466032 350323 466034
rect 347852 465976 350262 466032
rect 350318 465976 350323 466032
rect 347852 465974 350323 465976
rect 350257 465971 350323 465974
rect 407113 465898 407179 465901
rect 552013 465898 552079 465901
rect 407113 465896 410044 465898
rect 407113 465840 407118 465896
rect 407174 465840 410044 465896
rect 407113 465838 410044 465840
rect 549884 465896 552079 465898
rect 549884 465840 552018 465896
rect 552074 465840 552079 465896
rect 549884 465838 552079 465840
rect 407113 465835 407179 465838
rect 552013 465835 552079 465838
rect 36486 465156 36492 465220
rect 36556 465218 36562 465220
rect 48086 465218 48146 465256
rect 36556 465158 48146 465218
rect 347822 465218 347882 465256
rect 349429 465218 349495 465221
rect 347822 465216 349495 465218
rect 347822 465160 349434 465216
rect 349490 465160 349495 465216
rect 347822 465158 349495 465160
rect 36556 465156 36562 465158
rect 349429 465155 349495 465158
rect 46749 464266 46815 464269
rect 48086 464266 48146 464576
rect 46749 464264 48146 464266
rect 46749 464208 46754 464264
rect 46810 464208 48146 464264
rect 46749 464206 48146 464208
rect 46749 464203 46815 464206
rect 347822 463994 347882 464576
rect 549884 464410 550282 464470
rect 550222 464402 550282 464410
rect 552013 464402 552079 464405
rect 550222 464400 552079 464402
rect 550222 464344 552018 464400
rect 552074 464344 552079 464400
rect 550222 464342 552079 464344
rect 552013 464339 552079 464342
rect 350942 463994 350948 463996
rect 347822 463934 350948 463994
rect 350942 463932 350948 463934
rect 351012 463932 351018 463996
rect 45645 463858 45711 463861
rect 48086 463858 48146 463896
rect 45645 463856 48146 463858
rect 45645 463800 45650 463856
rect 45706 463800 48146 463856
rect 45645 463798 48146 463800
rect 407113 463858 407179 463861
rect 407113 463856 410044 463858
rect 407113 463800 407118 463856
rect 407174 463800 410044 463856
rect 407113 463798 410044 463800
rect 45645 463795 45711 463798
rect 407113 463795 407179 463798
rect 46749 463314 46815 463317
rect 46749 463312 48116 463314
rect 46749 463256 46754 463312
rect 46810 463256 48116 463312
rect 46749 463254 48116 463256
rect 46749 463251 46815 463254
rect 347822 462906 347882 463216
rect 407297 463178 407363 463181
rect 552013 463178 552079 463181
rect 407297 463176 410044 463178
rect 407297 463120 407302 463176
rect 407358 463120 410044 463176
rect 407297 463118 410044 463120
rect 549884 463176 552079 463178
rect 549884 463120 552018 463176
rect 552074 463120 552079 463176
rect 549884 463118 552079 463120
rect 407297 463115 407363 463118
rect 552013 463115 552079 463118
rect 350257 462906 350323 462909
rect 347822 462904 350323 462906
rect 347822 462848 350262 462904
rect 350318 462848 350323 462904
rect 347822 462846 350323 462848
rect 350257 462843 350323 462846
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect 350441 462634 350507 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect 347852 462632 350507 462634
rect 347852 462576 350446 462632
rect 350502 462576 350507 462632
rect 347852 462574 350507 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 350441 462571 350507 462574
rect 407113 462498 407179 462501
rect 407113 462496 410044 462498
rect 407113 462440 407118 462496
rect 407174 462440 410044 462496
rect 407113 462438 410044 462440
rect 407113 462435 407179 462438
rect 347822 461546 347882 461856
rect 407113 461818 407179 461821
rect 407113 461816 410044 461818
rect 407113 461760 407118 461816
rect 407174 461760 410044 461816
rect 407113 461758 410044 461760
rect 407113 461755 407179 461758
rect 350257 461546 350323 461549
rect 347822 461544 350323 461546
rect 347822 461488 350262 461544
rect 350318 461488 350323 461544
rect 347822 461486 350323 461488
rect 350257 461483 350323 461486
rect 46749 461002 46815 461005
rect 48086 461002 48146 461176
rect 347822 461138 347882 461176
rect 350441 461138 350507 461141
rect 347822 461136 350507 461138
rect 347822 461080 350446 461136
rect 350502 461080 350507 461136
rect 347822 461078 350507 461080
rect 350441 461075 350507 461078
rect 406653 461138 406719 461141
rect 406653 461136 410044 461138
rect 406653 461080 406658 461136
rect 406714 461080 410044 461136
rect 406653 461078 410044 461080
rect 406653 461075 406719 461078
rect 46749 461000 48146 461002
rect 46749 460944 46754 461000
rect 46810 460944 48146 461000
rect 46749 460942 48146 460944
rect 46749 460939 46815 460942
rect 552013 460458 552079 460461
rect 549884 460456 552079 460458
rect 549884 460400 552018 460456
rect 552074 460400 552079 460456
rect 549884 460398 552079 460400
rect 552013 460395 552079 460398
rect 46565 459914 46631 459917
rect 46565 459912 48116 459914
rect 46565 459856 46570 459912
rect 46626 459856 48116 459912
rect 46565 459854 48116 459856
rect 46565 459851 46631 459854
rect 347822 459642 347882 459816
rect 409597 459778 409663 459781
rect 550173 459778 550239 459781
rect 409597 459776 410044 459778
rect 409597 459720 409602 459776
rect 409658 459720 410044 459776
rect 409597 459718 410044 459720
rect 549884 459776 550239 459778
rect 549884 459720 550178 459776
rect 550234 459720 550239 459776
rect 549884 459718 550239 459720
rect 409597 459715 409663 459718
rect 550173 459715 550239 459718
rect 350441 459642 350507 459645
rect 347822 459640 350507 459642
rect 347822 459584 350446 459640
rect 350502 459584 350507 459640
rect 347822 459582 350507 459584
rect 350441 459579 350507 459582
rect 407113 459098 407179 459101
rect 552013 459098 552079 459101
rect 407113 459096 410044 459098
rect 407113 459040 407118 459096
rect 407174 459040 410044 459096
rect 407113 459038 410044 459040
rect 549884 459096 552079 459098
rect 549884 459040 552018 459096
rect 552074 459040 552079 459096
rect 549884 459038 552079 459040
rect 407113 459035 407179 459038
rect 552013 459035 552079 459038
rect 46749 458282 46815 458285
rect 48086 458282 48146 458456
rect 46749 458280 48146 458282
rect 46749 458224 46754 458280
rect 46810 458224 48146 458280
rect 46749 458222 48146 458224
rect 46749 458219 46815 458222
rect 583520 457996 584960 458236
rect 347822 457330 347882 457776
rect 408125 457738 408191 457741
rect 552013 457738 552079 457741
rect 408125 457736 410044 457738
rect 408125 457680 408130 457736
rect 408186 457680 410044 457736
rect 408125 457678 410044 457680
rect 549884 457736 552079 457738
rect 549884 457680 552018 457736
rect 552074 457680 552079 457736
rect 549884 457678 552079 457680
rect 408125 457675 408191 457678
rect 552013 457675 552079 457678
rect 350257 457330 350323 457333
rect 347822 457328 350323 457330
rect 347822 457272 350262 457328
rect 350318 457272 350323 457328
rect 347822 457270 350323 457272
rect 350257 457267 350323 457270
rect 43846 456860 43852 456924
rect 43916 456922 43922 456924
rect 48086 456922 48146 457096
rect 43916 456862 48146 456922
rect 347822 456922 347882 457096
rect 407113 457058 407179 457061
rect 407113 457056 410044 457058
rect 407113 457000 407118 457056
rect 407174 457000 410044 457056
rect 407113 456998 410044 457000
rect 407113 456995 407179 456998
rect 350441 456922 350507 456925
rect 347822 456920 350507 456922
rect 347822 456864 350446 456920
rect 350502 456864 350507 456920
rect 347822 456862 350507 456864
rect 43916 456860 43922 456862
rect 350441 456859 350507 456862
rect 46749 456514 46815 456517
rect 348233 456514 348299 456517
rect 46749 456512 48116 456514
rect 46749 456456 46754 456512
rect 46810 456456 48116 456512
rect 46749 456454 48116 456456
rect 347852 456512 348299 456514
rect 347852 456456 348238 456512
rect 348294 456456 348299 456512
rect 347852 456454 348299 456456
rect 46749 456451 46815 456454
rect 348233 456451 348299 456454
rect 552013 456378 552079 456381
rect 549884 456376 552079 456378
rect 549884 456320 552018 456376
rect 552074 456320 552079 456376
rect 549884 456318 552079 456320
rect 552013 456315 552079 456318
rect 46238 455772 46244 455836
rect 46308 455834 46314 455836
rect 349613 455834 349679 455837
rect 46308 455774 48116 455834
rect 347852 455832 349679 455834
rect 347852 455776 349618 455832
rect 349674 455776 349679 455832
rect 347852 455774 349679 455776
rect 46308 455772 46314 455774
rect 349613 455771 349679 455774
rect 407297 455698 407363 455701
rect 407297 455696 410044 455698
rect 407297 455640 407302 455696
rect 407358 455640 410044 455696
rect 407297 455638 410044 455640
rect 407297 455635 407363 455638
rect 407665 455018 407731 455021
rect 553301 455018 553367 455021
rect 407665 455016 410044 455018
rect 407665 454960 407670 455016
rect 407726 454960 410044 455016
rect 407665 454958 410044 454960
rect 549884 455016 553367 455018
rect 549884 454960 553306 455016
rect 553362 454960 553367 455016
rect 549884 454958 553367 454960
rect 407665 454955 407731 454958
rect 553301 454955 553367 454958
rect 347822 454202 347882 454376
rect 407113 454338 407179 454341
rect 552289 454338 552355 454341
rect 407113 454336 410044 454338
rect 407113 454280 407118 454336
rect 407174 454280 410044 454336
rect 407113 454278 410044 454280
rect 549884 454336 552355 454338
rect 549884 454280 552294 454336
rect 552350 454280 552355 454336
rect 549884 454278 552355 454280
rect 407113 454275 407179 454278
rect 552289 454275 552355 454278
rect 350441 454202 350507 454205
rect 347822 454200 350507 454202
rect 347822 454144 350446 454200
rect 350502 454144 350507 454200
rect 347822 454142 350507 454144
rect 350441 454139 350507 454142
rect 407113 453658 407179 453661
rect 552841 453658 552907 453661
rect 407113 453656 410044 453658
rect 407113 453600 407118 453656
rect 407174 453600 410044 453656
rect 407113 453598 410044 453600
rect 549884 453656 552907 453658
rect 549884 453600 552846 453656
rect 552902 453600 552907 453656
rect 549884 453598 552907 453600
rect 407113 453595 407179 453598
rect 552841 453595 552907 453598
rect 409597 452978 409663 452981
rect 409597 452976 410044 452978
rect 409597 452920 409602 452976
rect 409658 452920 410044 452976
rect 409597 452918 410044 452920
rect 409597 452915 409663 452918
rect 347822 451890 347882 452336
rect 350441 451890 350507 451893
rect 347822 451888 350507 451890
rect 347822 451832 350446 451888
rect 350502 451832 350507 451888
rect 347822 451830 350507 451832
rect 350441 451827 350507 451830
rect 347822 451485 347882 451656
rect 347822 451480 347931 451485
rect 347822 451424 347870 451480
rect 347926 451424 347931 451480
rect 347822 451422 347931 451424
rect 347865 451419 347931 451422
rect 407113 451346 407179 451349
rect 410014 451346 410074 451520
rect 549884 451490 550282 451550
rect 550222 451482 550282 451490
rect 552197 451482 552263 451485
rect 550222 451480 552263 451482
rect 550222 451424 552202 451480
rect 552258 451424 552263 451480
rect 550222 451422 552263 451424
rect 552197 451419 552263 451422
rect 407113 451344 410074 451346
rect 407113 451288 407118 451344
rect 407174 451288 410074 451344
rect 407113 451286 410074 451288
rect 407113 451283 407179 451286
rect 349705 451074 349771 451077
rect 347852 451072 349771 451074
rect 347852 451016 349710 451072
rect 349766 451016 349771 451072
rect 347852 451014 349771 451016
rect 349705 451011 349771 451014
rect 39614 450468 39620 450532
rect 39684 450530 39690 450532
rect 48086 450530 48146 450976
rect 39684 450470 48146 450530
rect 39684 450468 39690 450470
rect 46749 450394 46815 450397
rect 46749 450392 48116 450394
rect 46749 450336 46754 450392
rect 46810 450336 48116 450392
rect 46749 450334 48116 450336
rect 46749 450331 46815 450334
rect 347822 449986 347882 450296
rect 553301 450258 553367 450261
rect 549884 450256 553367 450258
rect 549884 450200 553306 450256
rect 553362 450200 553367 450256
rect 549884 450198 553367 450200
rect 553301 450195 553367 450198
rect 350441 449986 350507 449989
rect 347822 449984 350507 449986
rect 347822 449928 350446 449984
rect 350502 449928 350507 449984
rect 347822 449926 350507 449928
rect 350441 449923 350507 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 43662 449108 43668 449172
rect 43732 449170 43738 449172
rect 48086 449170 48146 449616
rect 407113 449578 407179 449581
rect 552565 449578 552631 449581
rect 407113 449576 410044 449578
rect 407113 449520 407118 449576
rect 407174 449520 410044 449576
rect 407113 449518 410044 449520
rect 549884 449576 552631 449578
rect 549884 449520 552570 449576
rect 552626 449520 552631 449576
rect 549884 449518 552631 449520
rect 407113 449515 407179 449518
rect 552565 449515 552631 449518
rect 43732 449110 48146 449170
rect 43732 449108 43738 449110
rect 552657 448898 552723 448901
rect 549884 448896 552723 448898
rect 549884 448840 552662 448896
rect 552718 448840 552723 448896
rect 549884 448838 552723 448840
rect 552657 448835 552723 448838
rect 347822 447810 347882 448256
rect 350441 447810 350507 447813
rect 347822 447808 350507 447810
rect 347822 447752 350446 447808
rect 350502 447752 350507 447808
rect 347822 447750 350507 447752
rect 350441 447747 350507 447750
rect 407297 447266 407363 447269
rect 410014 447266 410074 447440
rect 407297 447264 410074 447266
rect 407297 447208 407302 447264
rect 407358 447208 410074 447264
rect 407297 447206 410074 447208
rect 407297 447203 407363 447206
rect 347822 446450 347882 446896
rect 552565 446858 552631 446861
rect 549884 446856 552631 446858
rect 549884 446800 552570 446856
rect 552626 446800 552631 446856
rect 549884 446798 552631 446800
rect 552565 446795 552631 446798
rect 350257 446450 350323 446453
rect 347822 446448 350323 446450
rect 347822 446392 350262 446448
rect 350318 446392 350323 446448
rect 347822 446390 350323 446392
rect 350257 446387 350323 446390
rect 46749 445906 46815 445909
rect 48086 445906 48146 446216
rect 46749 445904 48146 445906
rect 46749 445848 46754 445904
rect 46810 445848 48146 445904
rect 46749 445846 48146 445848
rect 46749 445843 46815 445846
rect 347822 445773 347882 446216
rect 407113 446178 407179 446181
rect 407113 446176 410044 446178
rect 407113 446120 407118 446176
rect 407174 446120 410044 446176
rect 407113 446118 410044 446120
rect 407113 446115 407179 446118
rect 347822 445768 347931 445773
rect 347822 445712 347870 445768
rect 347926 445712 347931 445768
rect 347822 445710 347931 445712
rect 347865 445707 347931 445710
rect 350441 445634 350507 445637
rect 347852 445632 350507 445634
rect 347852 445576 350446 445632
rect 350502 445576 350507 445632
rect 347852 445574 350507 445576
rect 350441 445571 350507 445574
rect 46749 445090 46815 445093
rect 48086 445090 48146 445536
rect 552565 445498 552631 445501
rect 549884 445496 552631 445498
rect 549884 445440 552570 445496
rect 552626 445440 552631 445496
rect 549884 445438 552631 445440
rect 552565 445435 552631 445438
rect 46749 445088 48146 445090
rect 46749 445032 46754 445088
rect 46810 445032 48146 445088
rect 46749 445030 48146 445032
rect 46749 445027 46815 445030
rect 407113 444818 407179 444821
rect 407113 444816 410044 444818
rect 407113 444760 407118 444816
rect 407174 444760 410044 444816
rect 407113 444758 410044 444760
rect 407113 444755 407179 444758
rect 583520 444668 584960 444908
rect 46749 443322 46815 443325
rect 48086 443322 48146 443496
rect 553301 443458 553367 443461
rect 549884 443456 553367 443458
rect 549884 443400 553306 443456
rect 553362 443400 553367 443456
rect 549884 443398 553367 443400
rect 553301 443395 553367 443398
rect 46749 443320 48146 443322
rect 46749 443264 46754 443320
rect 46810 443264 48146 443320
rect 46749 443262 48146 443264
rect 46749 443259 46815 443262
rect 46657 442914 46723 442917
rect 46657 442912 48116 442914
rect 46657 442856 46662 442912
rect 46718 442856 48116 442912
rect 46657 442854 48116 442856
rect 46657 442851 46723 442854
rect 347822 441962 347882 442136
rect 407113 442098 407179 442101
rect 407113 442096 410044 442098
rect 407113 442040 407118 442096
rect 407174 442040 410044 442096
rect 407113 442038 410044 442040
rect 407113 442035 407179 442038
rect 349286 441962 349292 441964
rect 347822 441902 349292 441962
rect 349286 441900 349292 441902
rect 349356 441900 349362 441964
rect 407297 441418 407363 441421
rect 551502 441418 551508 441420
rect 407297 441416 410044 441418
rect 407297 441360 407302 441416
rect 407358 441360 410044 441416
rect 407297 441358 410044 441360
rect 549884 441358 551508 441418
rect 407297 441355 407363 441358
rect 551502 441356 551508 441358
rect 551572 441356 551578 441420
rect 347822 440602 347882 440776
rect 552289 440738 552355 440741
rect 549884 440736 552355 440738
rect 549884 440680 552294 440736
rect 552350 440680 552355 440736
rect 549884 440678 552355 440680
rect 552289 440675 552355 440678
rect 350441 440602 350507 440605
rect 347822 440600 350507 440602
rect 347822 440544 350446 440600
rect 350502 440544 350507 440600
rect 347822 440542 350507 440544
rect 350441 440539 350507 440542
rect 46013 439650 46079 439653
rect 48086 439650 48146 440096
rect 407113 440058 407179 440061
rect 407113 440056 410044 440058
rect 407113 440000 407118 440056
rect 407174 440000 410044 440056
rect 407113 439998 410044 440000
rect 407113 439995 407179 439998
rect 46013 439648 48146 439650
rect 46013 439592 46018 439648
rect 46074 439592 48146 439648
rect 46013 439590 48146 439592
rect 46013 439587 46079 439590
rect 46749 439106 46815 439109
rect 48086 439106 48146 439416
rect 46749 439104 48146 439106
rect 46749 439048 46754 439104
rect 46810 439048 48146 439104
rect 46749 439046 48146 439048
rect 46749 439043 46815 439046
rect 47025 438834 47091 438837
rect 47025 438832 48116 438834
rect 47025 438776 47030 438832
rect 47086 438776 48116 438832
rect 47025 438774 48116 438776
rect 47025 438771 47091 438774
rect 407481 438698 407547 438701
rect 553025 438698 553091 438701
rect 407481 438696 410044 438698
rect 407481 438640 407486 438696
rect 407542 438640 410044 438696
rect 407481 438638 410044 438640
rect 549884 438696 553091 438698
rect 549884 438640 553030 438696
rect 553086 438640 553091 438696
rect 549884 438638 553091 438640
rect 407481 438635 407547 438638
rect 553025 438635 553091 438638
rect 347822 437882 347882 438056
rect 406377 438018 406443 438021
rect 553301 438018 553367 438021
rect 406377 438016 410044 438018
rect 406377 437960 406382 438016
rect 406438 437960 410044 438016
rect 406377 437958 410044 437960
rect 549884 438016 553367 438018
rect 549884 437960 553306 438016
rect 553362 437960 553367 438016
rect 549884 437958 553367 437960
rect 406377 437955 406443 437958
rect 553301 437955 553367 437958
rect 350257 437882 350323 437885
rect 347822 437880 350323 437882
rect 347822 437824 350262 437880
rect 350318 437824 350323 437880
rect 347822 437822 350323 437824
rect 350257 437819 350323 437822
rect 407113 437338 407179 437341
rect 553025 437338 553091 437341
rect 407113 437336 410044 437338
rect 407113 437280 407118 437336
rect 407174 437280 410044 437336
rect 407113 437278 410044 437280
rect 549884 437336 553091 437338
rect 549884 437280 553030 437336
rect 553086 437280 553091 437336
rect 549884 437278 553091 437280
rect 407113 437275 407179 437278
rect 553025 437275 553091 437278
rect 350441 436794 350507 436797
rect 347852 436792 350507 436794
rect -960 436508 480 436748
rect 347852 436736 350446 436792
rect 350502 436736 350507 436792
rect 347852 436734 350507 436736
rect 350441 436731 350507 436734
rect 46749 436522 46815 436525
rect 48086 436522 48146 436696
rect 553301 436658 553367 436661
rect 549884 436656 553367 436658
rect 549884 436600 553306 436656
rect 553362 436600 553367 436656
rect 549884 436598 553367 436600
rect 553301 436595 553367 436598
rect 46749 436520 48146 436522
rect 46749 436464 46754 436520
rect 46810 436464 48146 436520
rect 46749 436462 48146 436464
rect 46749 436459 46815 436462
rect 407113 435978 407179 435981
rect 579838 435978 579844 435980
rect 407113 435976 410044 435978
rect 407113 435920 407118 435976
rect 407174 435920 410044 435976
rect 407113 435918 410044 435920
rect 549884 435918 579844 435978
rect 407113 435915 407179 435918
rect 579838 435916 579844 435918
rect 579908 435916 579914 435980
rect 347822 434890 347882 435336
rect 349102 434890 349108 434892
rect 347822 434830 349108 434890
rect 349102 434828 349108 434830
rect 349172 434828 349178 434892
rect 46749 434754 46815 434757
rect 350441 434754 350507 434757
rect 46749 434752 48116 434754
rect 46749 434696 46754 434752
rect 46810 434696 48116 434752
rect 46749 434694 48116 434696
rect 347852 434752 350507 434754
rect 347852 434696 350446 434752
rect 350502 434696 350507 434752
rect 347852 434694 350507 434696
rect 46749 434691 46815 434694
rect 350441 434691 350507 434694
rect 407205 434618 407271 434621
rect 407205 434616 410044 434618
rect 407205 434560 407210 434616
rect 407266 434560 410044 434616
rect 407205 434558 410044 434560
rect 407205 434555 407271 434558
rect 46749 433666 46815 433669
rect 48086 433666 48146 433976
rect 408125 433938 408191 433941
rect 408125 433936 410044 433938
rect 408125 433880 408130 433936
rect 408186 433880 410044 433936
rect 408125 433878 410044 433880
rect 408125 433875 408191 433878
rect 46749 433664 48146 433666
rect 46749 433608 46754 433664
rect 46810 433608 48146 433664
rect 46749 433606 48146 433608
rect 46749 433603 46815 433606
rect 349797 433394 349863 433397
rect 347852 433392 349863 433394
rect 347852 433336 349802 433392
rect 349858 433336 349863 433392
rect 347852 433334 349863 433336
rect 349797 433331 349863 433334
rect 406653 433258 406719 433261
rect 406653 433256 410044 433258
rect 406653 433200 406658 433256
rect 406714 433200 410044 433256
rect 406653 433198 410044 433200
rect 406653 433195 406719 433198
rect 46749 432034 46815 432037
rect 48086 432034 48146 432616
rect 552197 432578 552263 432581
rect 549884 432576 552263 432578
rect 549884 432520 552202 432576
rect 552258 432520 552263 432576
rect 549884 432518 552263 432520
rect 552197 432515 552263 432518
rect 46749 432032 48146 432034
rect 46749 431976 46754 432032
rect 46810 431976 48146 432032
rect 46749 431974 48146 431976
rect 46749 431971 46815 431974
rect 550265 431898 550331 431901
rect 549884 431896 550331 431898
rect 549884 431840 550270 431896
rect 550326 431840 550331 431896
rect 549884 431838 550331 431840
rect 550265 431835 550331 431838
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect 347822 430946 347882 431256
rect 350257 430946 350323 430949
rect 347822 430944 350323 430946
rect 347822 430888 350262 430944
rect 350318 430888 350323 430944
rect 347822 430886 350323 430888
rect 350257 430883 350323 430886
rect 350441 430674 350507 430677
rect 347852 430672 350507 430674
rect 347852 430616 350446 430672
rect 350502 430616 350507 430672
rect 347852 430614 350507 430616
rect 350441 430611 350507 430614
rect 409505 430538 409571 430541
rect 409505 430536 410044 430538
rect 409505 430480 409510 430536
rect 409566 430480 410044 430536
rect 409505 430478 410044 430480
rect 409505 430475 409571 430478
rect 45921 429994 45987 429997
rect 45921 429992 48116 429994
rect 45921 429936 45926 429992
rect 45982 429936 48116 429992
rect 45921 429934 48116 429936
rect 45921 429931 45987 429934
rect 407113 429858 407179 429861
rect 552197 429858 552263 429861
rect 407113 429856 410044 429858
rect 407113 429800 407118 429856
rect 407174 429800 410044 429856
rect 407113 429798 410044 429800
rect 549884 429856 552263 429858
rect 549884 429800 552202 429856
rect 552258 429800 552263 429856
rect 549884 429798 552263 429800
rect 407113 429795 407179 429798
rect 552197 429795 552263 429798
rect 44950 429252 44956 429316
rect 45020 429314 45026 429316
rect 45020 429254 48116 429314
rect 45020 429252 45026 429254
rect 407113 429178 407179 429181
rect 407113 429176 410044 429178
rect 407113 429120 407118 429176
rect 407174 429120 410044 429176
rect 407113 429118 410044 429120
rect 407113 429115 407179 429118
rect 46657 428362 46723 428365
rect 48086 428362 48146 428536
rect 409413 428498 409479 428501
rect 553025 428498 553091 428501
rect 409413 428496 410044 428498
rect 409413 428440 409418 428496
rect 409474 428440 410044 428496
rect 409413 428438 410044 428440
rect 549884 428496 553091 428498
rect 549884 428440 553030 428496
rect 553086 428440 553091 428496
rect 549884 428438 553091 428440
rect 409413 428435 409479 428438
rect 553025 428435 553091 428438
rect 46657 428360 48146 428362
rect 46657 428304 46662 428360
rect 46718 428304 48146 428360
rect 46657 428302 48146 428304
rect 46657 428299 46723 428302
rect 46749 427954 46815 427957
rect 350441 427954 350507 427957
rect 46749 427952 48116 427954
rect 46749 427896 46754 427952
rect 46810 427896 48116 427952
rect 46749 427894 48116 427896
rect 347852 427952 350507 427954
rect 347852 427896 350446 427952
rect 350502 427896 350507 427952
rect 347852 427894 350507 427896
rect 46749 427891 46815 427894
rect 350441 427891 350507 427894
rect 407205 427818 407271 427821
rect 407205 427816 410044 427818
rect 407205 427760 407210 427816
rect 407266 427760 410044 427816
rect 407205 427758 410044 427760
rect 407205 427755 407271 427758
rect 407113 427138 407179 427141
rect 407113 427136 410044 427138
rect 407113 427080 407118 427136
rect 407174 427080 410044 427136
rect 407113 427078 410044 427080
rect 407113 427075 407179 427078
rect 350441 426594 350507 426597
rect 347852 426592 350507 426594
rect 347852 426536 350446 426592
rect 350502 426536 350507 426592
rect 347852 426534 350507 426536
rect 350441 426531 350507 426534
rect 553025 426458 553091 426461
rect 549884 426456 553091 426458
rect 549884 426400 553030 426456
rect 553086 426400 553091 426456
rect 549884 426398 553091 426400
rect 553025 426395 553091 426398
rect 46657 425370 46723 425373
rect 48086 425370 48146 425816
rect 46657 425368 48146 425370
rect 46657 425312 46662 425368
rect 46718 425312 48146 425368
rect 46657 425310 48146 425312
rect 347822 425370 347882 425816
rect 407941 425778 408007 425781
rect 407941 425776 410044 425778
rect 407941 425720 407946 425776
rect 408002 425720 410044 425776
rect 407941 425718 410044 425720
rect 407941 425715 408007 425718
rect 350441 425370 350507 425373
rect 347822 425368 350507 425370
rect 347822 425312 350446 425368
rect 350502 425312 350507 425368
rect 347822 425310 350507 425312
rect 46657 425307 46723 425310
rect 350441 425307 350507 425310
rect 45645 425234 45711 425237
rect 45645 425232 48116 425234
rect 45645 425176 45650 425232
rect 45706 425176 48116 425232
rect 45645 425174 48116 425176
rect 45645 425171 45711 425174
rect 553025 425098 553091 425101
rect 549884 425096 553091 425098
rect 549884 425040 553030 425096
rect 553086 425040 553091 425096
rect 549884 425038 553091 425040
rect 553025 425035 553091 425038
rect 43478 424492 43484 424556
rect 43548 424554 43554 424556
rect 43548 424494 48116 424554
rect 43548 424492 43554 424494
rect 552933 424418 552999 424421
rect 549884 424416 552999 424418
rect 549884 424360 552938 424416
rect 552994 424360 552999 424416
rect 549884 424358 552999 424360
rect 552933 424355 552999 424358
rect 46749 423738 46815 423741
rect 48086 423738 48146 423776
rect 46749 423736 48146 423738
rect -960 423452 480 423692
rect 46749 423680 46754 423736
rect 46810 423680 48146 423736
rect 46749 423678 48146 423680
rect 407113 423738 407179 423741
rect 553025 423738 553091 423741
rect 407113 423736 410044 423738
rect 407113 423680 407118 423736
rect 407174 423680 410044 423736
rect 407113 423678 410044 423680
rect 549884 423736 553091 423738
rect 549884 423680 553030 423736
rect 553086 423680 553091 423736
rect 549884 423678 553091 423680
rect 46749 423675 46815 423678
rect 407113 423675 407179 423678
rect 553025 423675 553091 423678
rect 407113 423058 407179 423061
rect 407113 423056 410044 423058
rect 407113 423000 407118 423056
rect 407174 423000 410044 423056
rect 407113 422998 410044 423000
rect 407113 422995 407179 422998
rect 347822 422378 347882 422416
rect 350441 422378 350507 422381
rect 552013 422378 552079 422381
rect 347822 422376 350507 422378
rect 347822 422320 350446 422376
rect 350502 422320 350507 422376
rect 347822 422318 350507 422320
rect 549884 422376 552079 422378
rect 549884 422320 552018 422376
rect 552074 422320 552079 422376
rect 549884 422318 552079 422320
rect 350441 422315 350507 422318
rect 552013 422315 552079 422318
rect 46565 421290 46631 421293
rect 48086 421290 48146 421736
rect 46565 421288 48146 421290
rect 46565 421232 46570 421288
rect 46626 421232 48146 421288
rect 46565 421230 48146 421232
rect 347822 421290 347882 421736
rect 407849 421698 407915 421701
rect 552381 421698 552447 421701
rect 407849 421696 410044 421698
rect 407849 421640 407854 421696
rect 407910 421640 410044 421696
rect 407849 421638 410044 421640
rect 549884 421696 552447 421698
rect 549884 421640 552386 421696
rect 552442 421640 552447 421696
rect 549884 421638 552447 421640
rect 407849 421635 407915 421638
rect 552381 421635 552447 421638
rect 349981 421290 350047 421293
rect 347822 421288 350047 421290
rect 347822 421232 349986 421288
rect 350042 421232 350047 421288
rect 347822 421230 350047 421232
rect 46565 421227 46631 421230
rect 349981 421227 350047 421230
rect 45645 421018 45711 421021
rect 48086 421018 48146 421056
rect 45645 421016 48146 421018
rect 45645 420960 45650 421016
rect 45706 420960 48146 421016
rect 45645 420958 48146 420960
rect 347822 421018 347882 421056
rect 350441 421018 350507 421021
rect 552197 421018 552263 421021
rect 347822 421016 350507 421018
rect 347822 420960 350446 421016
rect 350502 420960 350507 421016
rect 347822 420958 350507 420960
rect 549884 421016 552263 421018
rect 549884 420960 552202 421016
rect 552258 420960 552263 421016
rect 549884 420958 552263 420960
rect 45645 420955 45711 420958
rect 350441 420955 350507 420958
rect 552197 420955 552263 420958
rect 45921 420066 45987 420069
rect 48086 420066 48146 420376
rect 407205 420338 407271 420341
rect 553025 420338 553091 420341
rect 407205 420336 410044 420338
rect 407205 420280 407210 420336
rect 407266 420280 410044 420336
rect 407205 420278 410044 420280
rect 549884 420336 553091 420338
rect 549884 420280 553030 420336
rect 553086 420280 553091 420336
rect 549884 420278 553091 420280
rect 407205 420275 407271 420278
rect 553025 420275 553091 420278
rect 45921 420064 48146 420066
rect 45921 420008 45926 420064
rect 45982 420008 48146 420064
rect 45921 420006 48146 420008
rect 45921 420003 45987 420006
rect 45645 419658 45711 419661
rect 48086 419658 48146 419696
rect 45645 419656 48146 419658
rect 45645 419600 45650 419656
rect 45706 419600 48146 419656
rect 45645 419598 48146 419600
rect 347822 419658 347882 419696
rect 350441 419658 350507 419661
rect 347822 419656 350507 419658
rect 347822 419600 350446 419656
rect 350502 419600 350507 419656
rect 347822 419598 350507 419600
rect 45645 419595 45711 419598
rect 350441 419595 350507 419598
rect 407113 419658 407179 419661
rect 407113 419656 410044 419658
rect 407113 419600 407118 419656
rect 407174 419600 410044 419656
rect 407113 419598 410044 419600
rect 407113 419595 407179 419598
rect 45921 418706 45987 418709
rect 48086 418706 48146 419016
rect 45921 418704 48146 418706
rect 45921 418648 45926 418704
rect 45982 418648 48146 418704
rect 45921 418646 48146 418648
rect 45921 418643 45987 418646
rect 35198 418372 35204 418436
rect 35268 418434 35274 418436
rect 347822 418434 347882 419016
rect 407113 418978 407179 418981
rect 407113 418976 410044 418978
rect 407113 418920 407118 418976
rect 407174 418920 410044 418976
rect 407113 418918 410044 418920
rect 407113 418915 407179 418918
rect 350441 418434 350507 418437
rect 35268 418374 48116 418434
rect 347822 418432 350507 418434
rect 347822 418376 350446 418432
rect 350502 418376 350507 418432
rect 347822 418374 350507 418376
rect 35268 418372 35274 418374
rect 350441 418371 350507 418374
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect 347822 416938 347882 416976
rect 350441 416938 350507 416941
rect 347822 416936 350507 416938
rect 347822 416880 350446 416936
rect 350502 416880 350507 416936
rect 347822 416878 350507 416880
rect 350441 416875 350507 416878
rect 45921 415986 45987 415989
rect 48086 415986 48146 416296
rect 407113 416258 407179 416261
rect 553025 416258 553091 416261
rect 407113 416256 410044 416258
rect 407113 416200 407118 416256
rect 407174 416200 410044 416256
rect 407113 416198 410044 416200
rect 549884 416256 553091 416258
rect 549884 416200 553030 416256
rect 553086 416200 553091 416256
rect 549884 416198 553091 416200
rect 407113 416195 407179 416198
rect 553025 416195 553091 416198
rect 45921 415984 48146 415986
rect 45921 415928 45926 415984
rect 45982 415928 48146 415984
rect 45921 415926 48146 415928
rect 45921 415923 45987 415926
rect 45645 415578 45711 415581
rect 48086 415578 48146 415616
rect 553025 415578 553091 415581
rect 45645 415576 48146 415578
rect 45645 415520 45650 415576
rect 45706 415520 48146 415576
rect 45645 415518 48146 415520
rect 549884 415576 553091 415578
rect 549884 415520 553030 415576
rect 553086 415520 553091 415576
rect 549884 415518 553091 415520
rect 45645 415515 45711 415518
rect 553025 415515 553091 415518
rect 347822 414490 347882 414936
rect 407113 414898 407179 414901
rect 407113 414896 410044 414898
rect 407113 414840 407118 414896
rect 407174 414840 410044 414896
rect 407113 414838 410044 414840
rect 407113 414835 407179 414838
rect 350257 414490 350323 414493
rect 347822 414488 350323 414490
rect 347822 414432 350262 414488
rect 350318 414432 350323 414488
rect 347822 414430 350323 414432
rect 350257 414427 350323 414430
rect 46749 414082 46815 414085
rect 48086 414082 48146 414256
rect 347822 414218 347882 414256
rect 350441 414218 350507 414221
rect 347822 414216 350507 414218
rect 347822 414160 350446 414216
rect 350502 414160 350507 414216
rect 347822 414158 350507 414160
rect 350441 414155 350507 414158
rect 46749 414080 48146 414082
rect 46749 414024 46754 414080
rect 46810 414024 48146 414080
rect 46749 414022 48146 414024
rect 46749 414019 46815 414022
rect 549884 413410 550282 413470
rect 550222 413402 550282 413410
rect 553025 413402 553091 413405
rect 550222 413400 553091 413402
rect 550222 413344 553030 413400
rect 553086 413344 553091 413400
rect 550222 413342 553091 413344
rect 553025 413339 553091 413342
rect 46422 412932 46428 412996
rect 46492 412994 46498 412996
rect 46492 412934 48116 412994
rect 46492 412932 46498 412934
rect 552381 412858 552447 412861
rect 549884 412856 552447 412858
rect 549884 412800 552386 412856
rect 552442 412800 552447 412856
rect 549884 412798 552447 412800
rect 552381 412795 552447 412798
rect 409505 412178 409571 412181
rect 409505 412176 410044 412178
rect 409505 412120 409510 412176
rect 409566 412120 410044 412176
rect 409505 412118 410044 412120
rect 409505 412115 409571 412118
rect 46749 411362 46815 411365
rect 48086 411362 48146 411536
rect 46749 411360 48146 411362
rect 46749 411304 46754 411360
rect 46810 411304 48146 411360
rect 46749 411302 48146 411304
rect 347822 411362 347882 411536
rect 407113 411498 407179 411501
rect 407113 411496 410044 411498
rect 407113 411440 407118 411496
rect 407174 411440 410044 411496
rect 407113 411438 410044 411440
rect 407113 411435 407179 411438
rect 350441 411362 350507 411365
rect 347822 411360 350507 411362
rect 347822 411304 350446 411360
rect 350502 411304 350507 411360
rect 347822 411302 350507 411304
rect 46749 411299 46815 411302
rect 350441 411299 350507 411302
rect 348141 410954 348207 410957
rect 347852 410952 348207 410954
rect 347852 410896 348146 410952
rect 348202 410896 348207 410952
rect 347852 410894 348207 410896
rect 348141 410891 348207 410894
rect 407113 410818 407179 410821
rect 553025 410818 553091 410821
rect 407113 410816 410044 410818
rect 407113 410760 407118 410816
rect 407174 410760 410044 410816
rect 407113 410758 410044 410760
rect 549884 410816 553091 410818
rect 549884 410760 553030 410816
rect 553086 410760 553091 410816
rect 549884 410758 553091 410760
rect 407113 410755 407179 410758
rect 553025 410755 553091 410758
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 349521 409594 349587 409597
rect 347852 409592 349587 409594
rect 347852 409536 349526 409592
rect 349582 409536 349587 409592
rect 347852 409534 349587 409536
rect 349521 409531 349587 409534
rect 407113 408778 407179 408781
rect 407113 408776 410044 408778
rect 407113 408720 407118 408776
rect 407174 408720 410044 408776
rect 407113 408718 410044 408720
rect 407113 408715 407179 408718
rect 46749 407690 46815 407693
rect 48086 407690 48146 408136
rect 46749 407688 48146 407690
rect 46749 407632 46754 407688
rect 46810 407632 48146 407688
rect 46749 407630 48146 407632
rect 46749 407627 46815 407630
rect 347822 407146 347882 407456
rect 367686 407356 367692 407420
rect 367756 407418 367762 407420
rect 552473 407418 552539 407421
rect 367756 407358 410044 407418
rect 549884 407416 552539 407418
rect 549884 407360 552478 407416
rect 552534 407360 552539 407416
rect 549884 407358 552539 407360
rect 367756 407356 367762 407358
rect 552473 407355 552539 407358
rect 353702 407146 353708 407148
rect 347822 407086 353708 407146
rect 353702 407084 353708 407086
rect 353772 407084 353778 407148
rect 407113 406058 407179 406061
rect 407113 406056 410044 406058
rect 407113 406000 407118 406056
rect 407174 406000 410044 406056
rect 407113 405998 410044 406000
rect 407113 405995 407179 405998
rect 347822 404970 347882 405416
rect 553025 405378 553091 405381
rect 549884 405376 553091 405378
rect 549884 405320 553030 405376
rect 553086 405320 553091 405376
rect 549884 405318 553091 405320
rect 553025 405315 553091 405318
rect 350257 404970 350323 404973
rect 347822 404968 350323 404970
rect 347822 404912 350262 404968
rect 350318 404912 350323 404968
rect 347822 404910 350323 404912
rect 350257 404907 350323 404910
rect 583520 404820 584960 405060
rect 347822 404426 347882 404736
rect 407205 404698 407271 404701
rect 554998 404698 555004 404700
rect 407205 404696 410044 404698
rect 407205 404640 407210 404696
rect 407266 404640 410044 404696
rect 407205 404638 410044 404640
rect 549884 404638 555004 404698
rect 407205 404635 407271 404638
rect 554998 404636 555004 404638
rect 555068 404636 555074 404700
rect 350441 404426 350507 404429
rect 347822 404424 350507 404426
rect 347822 404368 350446 404424
rect 350502 404368 350507 404424
rect 347822 404366 350507 404368
rect 350441 404363 350507 404366
rect 46749 403610 46815 403613
rect 48086 403610 48146 404056
rect 553025 404018 553091 404021
rect 549884 404016 553091 404018
rect 549884 403960 553030 404016
rect 553086 403960 553091 404016
rect 549884 403958 553091 403960
rect 553025 403955 553091 403958
rect 46749 403608 48146 403610
rect 46749 403552 46754 403608
rect 46810 403552 48146 403608
rect 46749 403550 48146 403552
rect 46749 403547 46815 403550
rect 553025 403338 553091 403341
rect 549884 403336 553091 403338
rect 549884 403280 553030 403336
rect 553086 403280 553091 403336
rect 549884 403278 553091 403280
rect 553025 403275 553091 403278
rect 39430 402052 39436 402116
rect 39500 402114 39506 402116
rect 48086 402114 48146 402696
rect 39500 402054 48146 402114
rect 39500 402052 39506 402054
rect 407757 401978 407823 401981
rect 407757 401976 410044 401978
rect 407757 401920 407762 401976
rect 407818 401920 410044 401976
rect 407757 401918 410044 401920
rect 407757 401915 407823 401918
rect 32990 400828 32996 400892
rect 33060 400890 33066 400892
rect 48086 400890 48146 401336
rect 33060 400830 48146 400890
rect 33060 400828 33066 400830
rect 46749 400346 46815 400349
rect 48086 400346 48146 400656
rect 46749 400344 48146 400346
rect 46749 400288 46754 400344
rect 46810 400288 48146 400344
rect 46749 400286 48146 400288
rect 347822 400346 347882 400656
rect 350441 400346 350507 400349
rect 347822 400344 350507 400346
rect 347822 400288 350446 400344
rect 350502 400288 350507 400344
rect 347822 400286 350507 400288
rect 46749 400283 46815 400286
rect 350441 400283 350507 400286
rect 407481 400346 407547 400349
rect 410014 400346 410074 400520
rect 549884 400490 550282 400550
rect 550222 400482 550282 400490
rect 553025 400482 553091 400485
rect 550222 400480 553091 400482
rect 550222 400424 553030 400480
rect 553086 400424 553091 400480
rect 550222 400422 553091 400424
rect 553025 400419 553091 400422
rect 407481 400344 410074 400346
rect 407481 400288 407486 400344
rect 407542 400288 410074 400344
rect 407481 400286 410074 400288
rect 407481 400283 407547 400286
rect 46749 399530 46815 399533
rect 48086 399530 48146 399976
rect 46749 399528 48146 399530
rect 46749 399472 46754 399528
rect 46810 399472 48146 399528
rect 46749 399470 48146 399472
rect 347822 399530 347882 399976
rect 350441 399530 350507 399533
rect 347822 399528 350507 399530
rect 347822 399472 350446 399528
rect 350502 399472 350507 399528
rect 347822 399470 350507 399472
rect 46749 399467 46815 399470
rect 350441 399467 350507 399470
rect 407113 399258 407179 399261
rect 407113 399256 410044 399258
rect 407113 399200 407118 399256
rect 407174 399200 410044 399256
rect 407113 399198 410044 399200
rect 407113 399195 407179 399198
rect 347822 397626 347882 397936
rect 407113 397898 407179 397901
rect 407113 397896 410044 397898
rect 407113 397840 407118 397896
rect 407174 397840 410044 397896
rect 407113 397838 410044 397840
rect 407113 397835 407179 397838
rect 350441 397626 350507 397629
rect 347822 397624 350507 397626
rect -960 397490 480 397580
rect 347822 397568 350446 397624
rect 350502 397568 350507 397624
rect 347822 397566 350507 397568
rect 350441 397563 350507 397566
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 40902 396612 40908 396676
rect 40972 396674 40978 396676
rect 48086 396674 48146 397256
rect 347822 396810 347882 397256
rect 350441 396810 350507 396813
rect 347822 396808 350507 396810
rect 347822 396752 350446 396808
rect 350502 396752 350507 396808
rect 347822 396750 350507 396752
rect 350441 396747 350507 396750
rect 349337 396674 349403 396677
rect 40972 396614 48146 396674
rect 347852 396672 349403 396674
rect 347852 396616 349342 396672
rect 349398 396616 349403 396672
rect 347852 396614 349403 396616
rect 40972 396612 40978 396614
rect 349337 396611 349403 396614
rect 348233 395926 348299 395929
rect 347852 395924 348299 395926
rect 347852 395868 348238 395924
rect 348294 395868 348299 395924
rect 347852 395866 348299 395868
rect 348233 395863 348299 395866
rect 407205 395858 407271 395861
rect 407205 395856 410044 395858
rect 407205 395800 407210 395856
rect 407266 395800 410044 395856
rect 407205 395798 410044 395800
rect 407205 395795 407271 395798
rect 46749 394770 46815 394773
rect 48086 394770 48146 395216
rect 46749 394768 48146 394770
rect 46749 394712 46754 394768
rect 46810 394712 48146 394768
rect 46749 394710 48146 394712
rect 347822 394770 347882 395216
rect 407113 395178 407179 395181
rect 553025 395178 553091 395181
rect 407113 395176 410044 395178
rect 407113 395120 407118 395176
rect 407174 395120 410044 395176
rect 407113 395118 410044 395120
rect 549884 395176 553091 395178
rect 549884 395120 553030 395176
rect 553086 395120 553091 395176
rect 549884 395118 553091 395120
rect 407113 395115 407179 395118
rect 553025 395115 553091 395118
rect 350257 394770 350323 394773
rect 347822 394768 350323 394770
rect 347822 394712 350262 394768
rect 350318 394712 350323 394768
rect 347822 394710 350323 394712
rect 46749 394707 46815 394710
rect 350257 394707 350323 394710
rect 350441 394634 350507 394637
rect 347852 394632 350507 394634
rect 347852 394576 350446 394632
rect 350502 394576 350507 394632
rect 347852 394574 350507 394576
rect 350441 394571 350507 394574
rect 46749 393546 46815 393549
rect 48086 393546 48146 393856
rect 407113 393818 407179 393821
rect 552197 393818 552263 393821
rect 407113 393816 410044 393818
rect 407113 393760 407118 393816
rect 407174 393760 410044 393816
rect 407113 393758 410044 393760
rect 549884 393816 552263 393818
rect 549884 393760 552202 393816
rect 552258 393760 552263 393816
rect 549884 393758 552263 393760
rect 407113 393755 407179 393758
rect 552197 393755 552263 393758
rect 46749 393544 48146 393546
rect 46749 393488 46754 393544
rect 46810 393488 48146 393544
rect 46749 393486 48146 393488
rect 46749 393483 46815 393486
rect 46105 392730 46171 392733
rect 48086 392730 48146 393176
rect 407573 393138 407639 393141
rect 407573 393136 410044 393138
rect 407573 393080 407578 393136
rect 407634 393080 410044 393136
rect 407573 393078 410044 393080
rect 407573 393075 407639 393078
rect 46105 392728 48146 392730
rect 46105 392672 46110 392728
rect 46166 392672 48146 392728
rect 46105 392670 48146 392672
rect 46105 392667 46171 392670
rect 46013 392186 46079 392189
rect 48086 392186 48146 392496
rect 347822 392322 347882 392496
rect 350441 392322 350507 392325
rect 347822 392320 350507 392322
rect 347822 392264 350446 392320
rect 350502 392264 350507 392320
rect 347822 392262 350507 392264
rect 350441 392259 350507 392262
rect 46013 392184 48146 392186
rect 46013 392128 46018 392184
rect 46074 392128 48146 392184
rect 46013 392126 48146 392128
rect 46013 392123 46079 392126
rect 347822 391370 347882 391816
rect 407205 391778 407271 391781
rect 553025 391778 553091 391781
rect 407205 391776 410044 391778
rect 407205 391720 407210 391776
rect 407266 391720 410044 391776
rect 407205 391718 410044 391720
rect 549884 391776 553091 391778
rect 549884 391720 553030 391776
rect 553086 391720 553091 391776
rect 549884 391718 553091 391720
rect 407205 391715 407271 391718
rect 553025 391715 553091 391718
rect 583520 391628 584960 391868
rect 349613 391370 349679 391373
rect 347822 391368 349679 391370
rect 347822 391312 349618 391368
rect 349674 391312 349679 391368
rect 347822 391310 349679 391312
rect 349613 391307 349679 391310
rect 348141 391166 348207 391169
rect 347852 391164 348207 391166
rect 36854 390628 36860 390692
rect 36924 390690 36930 390692
rect 48086 390690 48146 391136
rect 347852 391108 348146 391164
rect 348202 391108 348207 391164
rect 347852 391106 348207 391108
rect 348141 391103 348207 391106
rect 407113 391098 407179 391101
rect 553485 391098 553551 391101
rect 407113 391096 410044 391098
rect 407113 391040 407118 391096
rect 407174 391040 410044 391096
rect 407113 391038 410044 391040
rect 549884 391096 553551 391098
rect 549884 391040 553490 391096
rect 553546 391040 553551 391096
rect 549884 391038 553551 391040
rect 407113 391035 407179 391038
rect 553485 391035 553551 391038
rect 36924 390630 48146 390690
rect 36924 390628 36930 390630
rect 46473 390554 46539 390557
rect 46473 390552 48116 390554
rect 46473 390496 46478 390552
rect 46534 390496 48116 390552
rect 46473 390494 48116 390496
rect 46473 390491 46539 390494
rect 347822 390010 347882 390456
rect 553025 390418 553091 390421
rect 549884 390416 553091 390418
rect 549884 390360 553030 390416
rect 553086 390360 553091 390416
rect 549884 390358 553091 390360
rect 553025 390355 553091 390358
rect 350257 390010 350323 390013
rect 347822 390008 350323 390010
rect 347822 389952 350262 390008
rect 350318 389952 350323 390008
rect 347822 389950 350323 389952
rect 350257 389947 350323 389950
rect 350441 389874 350507 389877
rect 347852 389872 350507 389874
rect 347852 389816 350446 389872
rect 350502 389816 350507 389872
rect 347852 389814 350507 389816
rect 350441 389811 350507 389814
rect 46473 389330 46539 389333
rect 48086 389330 48146 389776
rect 407113 389738 407179 389741
rect 407113 389736 410044 389738
rect 407113 389680 407118 389736
rect 407174 389680 410044 389736
rect 407113 389678 410044 389680
rect 407113 389675 407179 389678
rect 46473 389328 48146 389330
rect 46473 389272 46478 389328
rect 46534 389272 48146 389328
rect 46473 389270 48146 389272
rect 46473 389267 46539 389270
rect 553025 388378 553091 388381
rect 549884 388376 553091 388378
rect 549884 388320 553030 388376
rect 553086 388320 553091 388376
rect 549884 388318 553091 388320
rect 553025 388315 553091 388318
rect 350441 387834 350507 387837
rect 347852 387832 350507 387834
rect 347852 387776 350446 387832
rect 350502 387776 350507 387832
rect 347852 387774 350507 387776
rect 350441 387771 350507 387774
rect 553025 387698 553091 387701
rect 549884 387696 553091 387698
rect 549884 387640 553030 387696
rect 553086 387640 553091 387696
rect 549884 387638 553091 387640
rect 553025 387635 553091 387638
rect 350257 387154 350323 387157
rect 347852 387152 350323 387154
rect 347852 387096 350262 387152
rect 350318 387096 350323 387152
rect 347852 387094 350323 387096
rect 350257 387091 350323 387094
rect 46473 386474 46539 386477
rect 46473 386472 48116 386474
rect 46473 386416 46478 386472
rect 46534 386416 48116 386472
rect 46473 386414 48116 386416
rect 46473 386411 46539 386414
rect 46105 385794 46171 385797
rect 349654 385794 349660 385796
rect 46105 385792 48116 385794
rect 46105 385736 46110 385792
rect 46166 385736 48116 385792
rect 46105 385734 48116 385736
rect 347852 385734 349660 385794
rect 46105 385731 46171 385734
rect 349654 385732 349660 385734
rect 349724 385732 349730 385796
rect 407113 385658 407179 385661
rect 553025 385658 553091 385661
rect 407113 385656 410044 385658
rect 407113 385600 407118 385656
rect 407174 385600 410044 385656
rect 407113 385598 410044 385600
rect 549884 385656 553091 385658
rect 549884 385600 553030 385656
rect 553086 385600 553091 385656
rect 549884 385598 553091 385600
rect 407113 385595 407179 385598
rect 553025 385595 553091 385598
rect 46473 385114 46539 385117
rect 350441 385114 350507 385117
rect 46473 385112 48116 385114
rect 46473 385056 46478 385112
rect 46534 385056 48116 385112
rect 46473 385054 48116 385056
rect 347852 385112 350507 385114
rect 347852 385056 350446 385112
rect 350502 385056 350507 385112
rect 347852 385054 350507 385056
rect 46473 385051 46539 385054
rect 350441 385051 350507 385054
rect 407113 384978 407179 384981
rect 407113 384976 410044 384978
rect 407113 384920 407118 384976
rect 407174 384920 410044 384976
rect 407113 384918 410044 384920
rect 407113 384915 407179 384918
rect -960 384284 480 384524
rect 349470 383754 349476 383756
rect 347852 383694 349476 383754
rect 349470 383692 349476 383694
rect 349540 383692 349546 383756
rect 46473 383074 46539 383077
rect 406469 383074 406535 383077
rect 410014 383074 410074 383520
rect 46473 383072 48116 383074
rect 46473 383016 46478 383072
rect 46534 383016 48116 383072
rect 46473 383014 48116 383016
rect 406469 383072 410074 383074
rect 406469 383016 406474 383072
rect 406530 383016 410074 383072
rect 406469 383014 410074 383016
rect 46473 383011 46539 383014
rect 406469 383011 406535 383014
rect 407113 382938 407179 382941
rect 407113 382936 410044 382938
rect 407113 382880 407118 382936
rect 407174 382880 410044 382936
rect 407113 382878 410044 382880
rect 407113 382875 407179 382878
rect 43478 382332 43484 382396
rect 43548 382394 43554 382396
rect 350257 382394 350323 382397
rect 43548 382334 48116 382394
rect 347852 382392 350323 382394
rect 347852 382336 350262 382392
rect 350318 382336 350323 382392
rect 347852 382334 350323 382336
rect 43548 382332 43554 382334
rect 350257 382331 350323 382334
rect 347822 381306 347882 381616
rect 407113 381578 407179 381581
rect 553025 381578 553091 381581
rect 407113 381576 410044 381578
rect 407113 381520 407118 381576
rect 407174 381520 410044 381576
rect 407113 381518 410044 381520
rect 549884 381576 553091 381578
rect 549884 381520 553030 381576
rect 553086 381520 553091 381576
rect 549884 381518 553091 381520
rect 407113 381515 407179 381518
rect 553025 381515 553091 381518
rect 350073 381306 350139 381309
rect 347822 381304 350139 381306
rect 347822 381248 350078 381304
rect 350134 381248 350139 381304
rect 347822 381246 350139 381248
rect 350073 381243 350139 381246
rect 46841 381034 46907 381037
rect 350257 381034 350323 381037
rect 46841 381032 48116 381034
rect 46841 380976 46846 381032
rect 46902 380976 48116 381032
rect 46841 380974 48116 380976
rect 347852 381032 350323 381034
rect 347852 380976 350262 381032
rect 350318 380976 350323 381032
rect 347852 380974 350323 380976
rect 46841 380971 46907 380974
rect 350257 380971 350323 380974
rect 46841 379810 46907 379813
rect 48086 379810 48146 380256
rect 46841 379808 48146 379810
rect 46841 379752 46846 379808
rect 46902 379752 48146 379808
rect 46841 379750 48146 379752
rect 347822 379810 347882 380256
rect 351177 379810 351243 379813
rect 347822 379808 351243 379810
rect 347822 379752 351182 379808
rect 351238 379752 351243 379808
rect 347822 379750 351243 379752
rect 46841 379747 46907 379750
rect 351177 379747 351243 379750
rect 349981 379538 350047 379541
rect 351126 379538 351132 379540
rect 349981 379536 351132 379538
rect 349981 379480 349986 379536
rect 350042 379480 351132 379536
rect 349981 379478 351132 379480
rect 349981 379475 350047 379478
rect 351126 379476 351132 379478
rect 351196 379476 351202 379540
rect 407113 378858 407179 378861
rect 550081 378858 550147 378861
rect 407113 378856 410044 378858
rect 407113 378800 407118 378856
rect 407174 378800 410044 378856
rect 407113 378798 410044 378800
rect 549884 378856 550147 378858
rect 549884 378800 550086 378856
rect 550142 378800 550147 378856
rect 549884 378798 550147 378800
rect 407113 378795 407179 378798
rect 550081 378795 550147 378798
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 47710 378184 47716 378248
rect 47780 378246 47786 378248
rect 47780 378186 48116 378246
rect 47780 378184 47786 378186
rect 407798 378116 407804 378180
rect 407868 378178 407874 378180
rect 553025 378178 553091 378181
rect 407868 378118 410044 378178
rect 549884 378176 553091 378178
rect 549884 378120 553030 378176
rect 553086 378120 553091 378176
rect 549884 378118 553091 378120
rect 407868 378116 407874 378118
rect 553025 378115 553091 378118
rect 347822 377226 347882 377536
rect 406745 377498 406811 377501
rect 553025 377498 553091 377501
rect 406745 377496 410044 377498
rect 406745 377440 406750 377496
rect 406806 377440 410044 377496
rect 406745 377438 410044 377440
rect 549884 377496 553091 377498
rect 549884 377440 553030 377496
rect 553086 377440 553091 377496
rect 549884 377438 553091 377440
rect 406745 377435 406811 377438
rect 553025 377435 553091 377438
rect 350257 377226 350323 377229
rect 347822 377224 350323 377226
rect 347822 377168 350262 377224
rect 350318 377168 350323 377224
rect 347822 377166 350323 377168
rect 350257 377163 350323 377166
rect 350073 376954 350139 376957
rect 347852 376952 350139 376954
rect 347852 376896 350078 376952
rect 350134 376896 350139 376952
rect 347852 376894 350139 376896
rect 350073 376891 350139 376894
rect 46473 376274 46539 376277
rect 46473 376272 48116 376274
rect 46473 376216 46478 376272
rect 46534 376216 48116 376272
rect 46473 376214 48116 376216
rect 46473 376211 46539 376214
rect 347822 375866 347882 376176
rect 350073 375866 350139 375869
rect 347822 375864 350139 375866
rect 347822 375808 350078 375864
rect 350134 375808 350139 375864
rect 347822 375806 350139 375808
rect 350073 375803 350139 375806
rect 350257 374914 350323 374917
rect 347852 374912 350323 374914
rect 347852 374856 350262 374912
rect 350318 374856 350323 374912
rect 347852 374854 350323 374856
rect 350257 374851 350323 374854
rect 32806 374036 32812 374100
rect 32876 374098 32882 374100
rect 48086 374098 48146 374136
rect 32876 374038 48146 374098
rect 408125 374098 408191 374101
rect 408125 374096 410044 374098
rect 408125 374040 408130 374096
rect 408186 374040 410044 374096
rect 408125 374038 410044 374040
rect 32876 374036 32882 374038
rect 408125 374035 408191 374038
rect 45001 373010 45067 373013
rect 48086 373010 48146 373456
rect 45001 373008 48146 373010
rect 45001 372952 45006 373008
rect 45062 372952 48146 373008
rect 45001 372950 48146 372952
rect 45001 372947 45067 372950
rect 347822 372874 347882 373456
rect 407113 373418 407179 373421
rect 407113 373416 410044 373418
rect 407113 373360 407118 373416
rect 407174 373360 410044 373416
rect 407113 373358 410044 373360
rect 407113 373355 407179 373358
rect 350257 372874 350323 372877
rect 347822 372872 350323 372874
rect 347822 372816 350262 372872
rect 350318 372816 350323 372872
rect 347822 372814 350323 372816
rect 350257 372811 350323 372814
rect 46841 372738 46907 372741
rect 48086 372738 48146 372776
rect 552197 372738 552263 372741
rect 46841 372736 48146 372738
rect 46841 372680 46846 372736
rect 46902 372680 48146 372736
rect 46841 372678 48146 372680
rect 549884 372736 552263 372738
rect 549884 372680 552202 372736
rect 552258 372680 552263 372736
rect 549884 372678 552263 372680
rect 46841 372675 46907 372678
rect 552197 372675 552263 372678
rect 46841 371514 46907 371517
rect 48086 371514 48146 372096
rect 406837 372058 406903 372061
rect 406837 372056 410044 372058
rect 406837 372000 406842 372056
rect 406898 372000 410044 372056
rect 406837 371998 410044 372000
rect 406837 371995 406903 371998
rect 46841 371512 48146 371514
rect -960 371228 480 371468
rect 46841 371456 46846 371512
rect 46902 371456 48146 371512
rect 46841 371454 48146 371456
rect 46841 371451 46907 371454
rect 347822 371378 347882 371416
rect 350257 371378 350323 371381
rect 552013 371378 552079 371381
rect 347822 371376 350323 371378
rect 347822 371320 350262 371376
rect 350318 371320 350323 371376
rect 347822 371318 350323 371320
rect 549884 371376 552079 371378
rect 549884 371320 552018 371376
rect 552074 371320 552079 371376
rect 549884 371318 552079 371320
rect 350257 371315 350323 371318
rect 552013 371315 552079 371318
rect 407113 370698 407179 370701
rect 553025 370698 553091 370701
rect 407113 370696 410044 370698
rect 407113 370640 407118 370696
rect 407174 370640 410044 370696
rect 407113 370638 410044 370640
rect 549884 370696 553091 370698
rect 549884 370640 553030 370696
rect 553086 370640 553091 370696
rect 549884 370638 553091 370640
rect 407113 370635 407179 370638
rect 553025 370635 553091 370638
rect 350073 370154 350139 370157
rect 347852 370152 350139 370154
rect 347852 370096 350078 370152
rect 350134 370096 350139 370152
rect 347852 370094 350139 370096
rect 350073 370091 350139 370094
rect 46841 368930 46907 368933
rect 48086 368930 48146 369376
rect 403750 369276 403756 369340
rect 403820 369338 403826 369340
rect 552197 369338 552263 369341
rect 403820 369278 410044 369338
rect 549884 369336 552263 369338
rect 549884 369280 552202 369336
rect 552258 369280 552263 369336
rect 549884 369278 552263 369280
rect 403820 369276 403826 369278
rect 552197 369275 552263 369278
rect 46841 368928 48146 368930
rect 46841 368872 46846 368928
rect 46902 368872 48146 368928
rect 46841 368870 48146 368872
rect 46841 368867 46907 368870
rect 348325 368726 348391 368729
rect 347852 368724 348391 368726
rect 347852 368668 348330 368724
rect 348386 368668 348391 368724
rect 347852 368666 348391 368668
rect 348325 368663 348391 368666
rect 553025 368658 553091 368661
rect 549884 368656 553091 368658
rect 549884 368600 553030 368656
rect 553086 368600 553091 368656
rect 549884 368598 553091 368600
rect 553025 368595 553091 368598
rect 46841 367570 46907 367573
rect 48086 367570 48146 368016
rect 552013 367978 552079 367981
rect 549884 367976 552079 367978
rect 549884 367920 552018 367976
rect 552074 367920 552079 367976
rect 549884 367918 552079 367920
rect 552013 367915 552079 367918
rect 46841 367568 48146 367570
rect 46841 367512 46846 367568
rect 46902 367512 48146 367568
rect 46841 367510 48146 367512
rect 46841 367507 46907 367510
rect 549884 366490 550282 366550
rect 550222 366482 550282 366490
rect 552933 366482 552999 366485
rect 550222 366480 552999 366482
rect 550222 366424 552938 366480
rect 552994 366424 552999 366480
rect 550222 366422 552999 366424
rect 552933 366419 552999 366422
rect 46013 366074 46079 366077
rect 46013 366072 48116 366074
rect 46013 366016 46018 366072
rect 46074 366016 48116 366072
rect 46013 366014 48116 366016
rect 46013 366011 46079 366014
rect 553025 365938 553091 365941
rect 549884 365936 553091 365938
rect 549884 365880 553030 365936
rect 553086 365880 553091 365936
rect 549884 365878 553091 365880
rect 553025 365875 553091 365878
rect 351085 365394 351151 365397
rect 347852 365392 351151 365394
rect 347852 365336 351090 365392
rect 351146 365336 351151 365392
rect 347852 365334 351151 365336
rect 351085 365331 351151 365334
rect 552013 365258 552079 365261
rect 549884 365256 552079 365258
rect 549884 365200 552018 365256
rect 552074 365200 552079 365256
rect 549884 365198 552079 365200
rect 552013 365195 552079 365198
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect 347822 364578 347882 364616
rect 351085 364578 351151 364581
rect 347822 364576 351151 364578
rect 347822 364520 351090 364576
rect 351146 364520 351151 364576
rect 347822 364518 351151 364520
rect 351085 364515 351151 364518
rect 409689 364578 409755 364581
rect 409689 364576 410044 364578
rect 409689 364520 409694 364576
rect 409750 364520 410044 364576
rect 409689 364518 410044 364520
rect 409689 364515 409755 364518
rect 46841 363490 46907 363493
rect 48086 363490 48146 363936
rect 46841 363488 48146 363490
rect 46841 363432 46846 363488
rect 46902 363432 48146 363488
rect 46841 363430 48146 363432
rect 46841 363427 46907 363430
rect 347822 363354 347882 363936
rect 553577 363898 553643 363901
rect 549884 363896 553643 363898
rect 549884 363840 553582 363896
rect 553638 363840 553643 363896
rect 549884 363838 553643 363840
rect 553577 363835 553643 363838
rect 350073 363354 350139 363357
rect 347822 363352 350139 363354
rect 347822 363296 350078 363352
rect 350134 363296 350139 363352
rect 347822 363294 350139 363296
rect 350073 363291 350139 363294
rect 408033 362538 408099 362541
rect 408033 362536 410044 362538
rect 408033 362480 408038 362536
rect 408094 362480 410044 362536
rect 408033 362478 410044 362480
rect 408033 362475 408099 362478
rect 407113 361178 407179 361181
rect 552933 361178 552999 361181
rect 407113 361176 410044 361178
rect 407113 361120 407118 361176
rect 407174 361120 410044 361176
rect 407113 361118 410044 361120
rect 549884 361176 552999 361178
rect 549884 361120 552938 361176
rect 552994 361120 552999 361176
rect 549884 361118 552999 361120
rect 407113 361115 407179 361118
rect 552933 361115 552999 361118
rect 407113 360498 407179 360501
rect 553025 360498 553091 360501
rect 407113 360496 410044 360498
rect 407113 360440 407118 360496
rect 407174 360440 410044 360496
rect 407113 360438 410044 360440
rect 549884 360496 553091 360498
rect 549884 360440 553030 360496
rect 553086 360440 553091 360496
rect 549884 360438 553091 360440
rect 407113 360435 407179 360438
rect 553025 360435 553091 360438
rect 45093 359410 45159 359413
rect 48086 359410 48146 359856
rect 45093 359408 48146 359410
rect 45093 359352 45098 359408
rect 45154 359352 48146 359408
rect 45093 359350 48146 359352
rect 45093 359347 45159 359350
rect 347822 358866 347882 359176
rect 350257 358866 350323 358869
rect 347822 358864 350323 358866
rect 347822 358808 350262 358864
rect 350318 358808 350323 358864
rect 347822 358806 350323 358808
rect 350257 358803 350323 358806
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 347822 358322 347882 358496
rect 552933 358458 552999 358461
rect 549884 358456 552999 358458
rect 549884 358400 552938 358456
rect 552994 358400 552999 358456
rect 549884 358398 552999 358400
rect 552933 358395 552999 358398
rect 350257 358322 350323 358325
rect 347822 358320 350323 358322
rect 347822 358264 350262 358320
rect 350318 358264 350323 358320
rect 347822 358262 350323 358264
rect 350257 358259 350323 358262
rect 46841 357914 46907 357917
rect 46841 357912 48116 357914
rect 46841 357856 46846 357912
rect 46902 357856 48116 357912
rect 46841 357854 48116 357856
rect 46841 357851 46907 357854
rect 409454 357716 409460 357780
rect 409524 357778 409530 357780
rect 553025 357778 553091 357781
rect 409524 357718 410044 357778
rect 549884 357776 553091 357778
rect 549884 357720 553030 357776
rect 553086 357720 553091 357776
rect 549884 357718 553091 357720
rect 409524 357716 409530 357718
rect 553025 357715 553091 357718
rect 347822 356690 347882 357136
rect 407113 357098 407179 357101
rect 407113 357096 410044 357098
rect 407113 357040 407118 357096
rect 407174 357040 410044 357096
rect 407113 357038 410044 357040
rect 407113 357035 407179 357038
rect 350257 356690 350323 356693
rect 347822 356688 350323 356690
rect 347822 356632 350262 356688
rect 350318 356632 350323 356688
rect 347822 356630 350323 356632
rect 350257 356627 350323 356630
rect 406837 356418 406903 356421
rect 406837 356416 410044 356418
rect 406837 356360 406842 356416
rect 406898 356360 410044 356416
rect 406837 356358 410044 356360
rect 406837 356355 406903 356358
rect 350257 355874 350323 355877
rect 347852 355872 350323 355874
rect 347852 355816 350262 355872
rect 350318 355816 350323 355872
rect 347852 355814 350323 355816
rect 350257 355811 350323 355814
rect 553025 355738 553091 355741
rect 549884 355736 553091 355738
rect 549884 355680 553030 355736
rect 553086 355680 553091 355736
rect 549884 355678 553091 355680
rect 553025 355675 553091 355678
rect 46473 354786 46539 354789
rect 48086 354786 48146 355096
rect 46473 354784 48146 354786
rect 46473 354728 46478 354784
rect 46534 354728 48146 354784
rect 46473 354726 48146 354728
rect 347822 354786 347882 355096
rect 350257 354786 350323 354789
rect 347822 354784 350323 354786
rect 347822 354728 350262 354784
rect 350318 354728 350323 354784
rect 347822 354726 350323 354728
rect 46473 354723 46539 354726
rect 350257 354723 350323 354726
rect 552381 354378 552447 354381
rect 549884 354376 552447 354378
rect 549884 354320 552386 354376
rect 552442 354320 552447 354376
rect 549884 354318 552447 354320
rect 552381 354315 552447 354318
rect 407113 353698 407179 353701
rect 553025 353698 553091 353701
rect 407113 353696 410044 353698
rect 407113 353640 407118 353696
rect 407174 353640 410044 353696
rect 407113 353638 410044 353640
rect 549884 353696 553091 353698
rect 549884 353640 553030 353696
rect 553086 353640 553091 353696
rect 549884 353638 553091 353640
rect 407113 353635 407179 353638
rect 553025 353635 553091 353638
rect 46473 353154 46539 353157
rect 46473 353152 48116 353154
rect 46473 353096 46478 353152
rect 46534 353096 48116 353152
rect 46473 353094 48116 353096
rect 46473 353091 46539 353094
rect 407205 353018 407271 353021
rect 407205 353016 410044 353018
rect 407205 352960 407210 353016
rect 407266 352960 410044 353016
rect 407205 352958 410044 352960
rect 407205 352955 407271 352958
rect 407113 352338 407179 352341
rect 407113 352336 410044 352338
rect 407113 352280 407118 352336
rect 407174 352280 410044 352336
rect 407113 352278 410044 352280
rect 407113 352275 407179 352278
rect 583520 351780 584960 352020
rect 407113 351658 407179 351661
rect 552841 351658 552907 351661
rect 407113 351656 410044 351658
rect 407113 351600 407118 351656
rect 407174 351600 410044 351656
rect 407113 351598 410044 351600
rect 549884 351656 552907 351658
rect 549884 351600 552846 351656
rect 552902 351600 552907 351656
rect 549884 351598 552907 351600
rect 407113 351595 407179 351598
rect 552841 351595 552907 351598
rect 347822 350706 347882 351016
rect 553117 350978 553183 350981
rect 549884 350976 553183 350978
rect 549884 350920 553122 350976
rect 553178 350920 553183 350976
rect 549884 350918 553183 350920
rect 553117 350915 553183 350918
rect 350257 350706 350323 350709
rect 347822 350704 350323 350706
rect 347822 350648 350262 350704
rect 350318 350648 350323 350704
rect 347822 350646 350323 350648
rect 350257 350643 350323 350646
rect 347822 349890 347882 350336
rect 350073 349890 350139 349893
rect 347822 349888 350139 349890
rect 347822 349832 350078 349888
rect 350134 349832 350139 349888
rect 347822 349830 350139 349832
rect 350073 349827 350139 349830
rect 46473 349210 46539 349213
rect 48086 349210 48146 349656
rect 347822 349482 347882 349656
rect 350257 349482 350323 349485
rect 347822 349480 350323 349482
rect 347822 349424 350262 349480
rect 350318 349424 350323 349480
rect 347822 349422 350323 349424
rect 350257 349419 350323 349422
rect 46473 349208 48146 349210
rect 46473 349152 46478 349208
rect 46534 349152 48146 349208
rect 46473 349150 48146 349152
rect 407113 349210 407179 349213
rect 410014 349210 410074 349520
rect 549884 349490 550282 349550
rect 550222 349482 550282 349490
rect 553117 349482 553183 349485
rect 550222 349480 553183 349482
rect 550222 349424 553122 349480
rect 553178 349424 553183 349480
rect 550222 349422 553183 349424
rect 553117 349419 553183 349422
rect 407113 349208 410074 349210
rect 407113 349152 407118 349208
rect 407174 349152 410074 349208
rect 407113 349150 410074 349152
rect 46473 349147 46539 349150
rect 407113 349147 407179 349150
rect 46473 347170 46539 347173
rect 48086 347170 48146 347616
rect 553025 347578 553091 347581
rect 549884 347576 553091 347578
rect 549884 347520 553030 347576
rect 553086 347520 553091 347576
rect 549884 347518 553091 347520
rect 553025 347515 553091 347518
rect 46473 347168 48146 347170
rect 46473 347112 46478 347168
rect 46534 347112 48146 347168
rect 46473 347110 48146 347112
rect 46473 347107 46539 347110
rect 349245 347034 349311 347037
rect 347852 347032 349311 347034
rect 347852 346976 349250 347032
rect 349306 346976 349311 347032
rect 347852 346974 349311 346976
rect 349245 346971 349311 346974
rect 407113 346898 407179 346901
rect 553117 346898 553183 346901
rect 407113 346896 410044 346898
rect 407113 346840 407118 346896
rect 407174 346840 410044 346896
rect 407113 346838 410044 346840
rect 549884 346896 553183 346898
rect 549884 346840 553122 346896
rect 553178 346840 553183 346896
rect 549884 346838 553183 346840
rect 407113 346835 407179 346838
rect 553117 346835 553183 346838
rect 347822 345810 347882 346256
rect 350257 345810 350323 345813
rect 347822 345808 350323 345810
rect 347822 345752 350262 345808
rect 350318 345752 350323 345808
rect 347822 345750 350323 345752
rect 350257 345747 350323 345750
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 46473 345130 46539 345133
rect 48086 345130 48146 345576
rect 406745 345266 406811 345269
rect 410014 345266 410074 345440
rect 406745 345264 410074 345266
rect 406745 345208 406750 345264
rect 406806 345208 410074 345264
rect 406745 345206 410074 345208
rect 406745 345203 406811 345206
rect 46473 345128 48146 345130
rect 46473 345072 46478 345128
rect 46534 345072 48146 345128
rect 46473 345070 48146 345072
rect 46473 345067 46539 345070
rect 347822 344450 347882 344896
rect 407113 344858 407179 344861
rect 407113 344856 410044 344858
rect 407113 344800 407118 344856
rect 407174 344800 410044 344856
rect 407113 344798 410044 344800
rect 407113 344795 407179 344798
rect 350073 344450 350139 344453
rect 347822 344448 350139 344450
rect 347822 344392 350078 344448
rect 350134 344392 350139 344448
rect 347822 344390 350139 344392
rect 350073 344387 350139 344390
rect 347822 344042 347882 344216
rect 350257 344042 350323 344045
rect 347822 344040 350323 344042
rect 347822 343984 350262 344040
rect 350318 343984 350323 344040
rect 347822 343982 350323 343984
rect 350257 343979 350323 343982
rect 407113 343498 407179 343501
rect 553025 343498 553091 343501
rect 407113 343496 410044 343498
rect 407113 343440 407118 343496
rect 407174 343440 410044 343496
rect 407113 343438 410044 343440
rect 549884 343496 553091 343498
rect 549884 343440 553030 343496
rect 553086 343440 553091 343496
rect 549884 343438 553091 343440
rect 407113 343435 407179 343438
rect 553025 343435 553091 343438
rect 409689 342818 409755 342821
rect 552013 342818 552079 342821
rect 409689 342816 410044 342818
rect 409689 342760 409694 342816
rect 409750 342760 410044 342816
rect 409689 342758 410044 342760
rect 549884 342816 552079 342818
rect 549884 342760 552018 342816
rect 552074 342760 552079 342816
rect 549884 342758 552079 342760
rect 409689 342755 409755 342758
rect 552013 342755 552079 342758
rect 350993 342274 351059 342277
rect 347852 342272 351059 342274
rect 347852 342216 350998 342272
rect 351054 342216 351059 342272
rect 347852 342214 351059 342216
rect 350993 342211 351059 342214
rect 407113 340778 407179 340781
rect 553577 340778 553643 340781
rect 407113 340776 410044 340778
rect 407113 340720 407118 340776
rect 407174 340720 410044 340776
rect 407113 340718 410044 340720
rect 549884 340776 553643 340778
rect 549884 340720 553582 340776
rect 553638 340720 553643 340776
rect 549884 340718 553643 340720
rect 407113 340715 407179 340718
rect 553577 340715 553643 340718
rect 552933 340098 552999 340101
rect 549884 340096 552999 340098
rect 549884 340040 552938 340096
rect 552994 340040 552999 340096
rect 549884 340038 552999 340040
rect 552933 340035 552999 340038
rect 45277 339554 45343 339557
rect 45277 339552 48116 339554
rect 45277 339496 45282 339552
rect 45338 339496 48116 339552
rect 45277 339494 48116 339496
rect 45277 339491 45343 339494
rect 407113 339418 407179 339421
rect 407113 339416 410044 339418
rect 407113 339360 407118 339416
rect 407174 339360 410044 339416
rect 407113 339358 410044 339360
rect 407113 339355 407179 339358
rect 553117 338738 553183 338741
rect 549884 338736 553183 338738
rect 549884 338680 553122 338736
rect 553178 338680 553183 338736
rect 549884 338678 553183 338680
rect 553117 338675 553183 338678
rect 583520 338452 584960 338692
rect 350993 338194 351059 338197
rect 347852 338192 351059 338194
rect 347852 338136 350998 338192
rect 351054 338136 351059 338192
rect 347852 338134 351059 338136
rect 350993 338131 351059 338134
rect 46473 336834 46539 336837
rect 46473 336832 48116 336834
rect 46473 336776 46478 336832
rect 46534 336776 48116 336832
rect 46473 336774 48116 336776
rect 46473 336771 46539 336774
rect 407113 336698 407179 336701
rect 550214 336698 550220 336700
rect 407113 336696 410044 336698
rect 407113 336640 407118 336696
rect 407174 336640 410044 336696
rect 407113 336638 410044 336640
rect 549884 336638 550220 336698
rect 407113 336635 407179 336638
rect 550214 336636 550220 336638
rect 550284 336636 550290 336700
rect 347957 336562 348023 336565
rect 347822 336560 348023 336562
rect 347822 336504 347962 336560
rect 348018 336504 348023 336560
rect 347822 336502 348023 336504
rect 347822 336124 347882 336502
rect 347957 336499 348023 336502
rect 553025 336018 553091 336021
rect 549884 336016 553091 336018
rect 549884 335960 553030 336016
rect 553086 335960 553091 336016
rect 549884 335958 553091 335960
rect 553025 335955 553091 335958
rect 47025 335474 47091 335477
rect 47025 335472 48116 335474
rect 47025 335416 47030 335472
rect 47086 335416 48116 335472
rect 47025 335414 48116 335416
rect 47025 335411 47091 335414
rect 408125 335338 408191 335341
rect 553117 335338 553183 335341
rect 408125 335336 410044 335338
rect 408125 335280 408130 335336
rect 408186 335280 410044 335336
rect 408125 335278 410044 335280
rect 549884 335336 553183 335338
rect 549884 335280 553122 335336
rect 553178 335280 553183 335336
rect 549884 335278 553183 335280
rect 408125 335275 408191 335278
rect 553117 335275 553183 335278
rect 409781 334658 409847 334661
rect 552841 334658 552907 334661
rect 409781 334656 410044 334658
rect 409781 334600 409786 334656
rect 409842 334600 410044 334656
rect 409781 334598 410044 334600
rect 549884 334656 552907 334658
rect 549884 334600 552846 334656
rect 552902 334600 552907 334656
rect 549884 334598 552907 334600
rect 409781 334595 409847 334598
rect 552841 334595 552907 334598
rect 350349 334114 350415 334117
rect 347852 334112 350415 334114
rect 347852 334056 350354 334112
rect 350410 334056 350415 334112
rect 347852 334054 350415 334056
rect 350349 334051 350415 334054
rect 551185 333978 551251 333981
rect 549884 333976 551251 333978
rect 549884 333920 551190 333976
rect 551246 333920 551251 333976
rect 549884 333918 551251 333920
rect 551185 333915 551251 333918
rect 347822 332754 347882 333336
rect 350349 332754 350415 332757
rect 347822 332752 350415 332754
rect 347822 332696 350354 332752
rect 350410 332696 350415 332752
rect 347822 332694 350415 332696
rect 350349 332691 350415 332694
rect 407389 332618 407455 332621
rect 407389 332616 410044 332618
rect 407389 332560 407394 332616
rect 407450 332560 410044 332616
rect 407389 332558 410044 332560
rect 407389 332555 407455 332558
rect -960 332196 480 332436
rect 347822 331122 347882 331296
rect 395470 331196 395476 331260
rect 395540 331258 395546 331260
rect 552565 331258 552631 331261
rect 395540 331198 410044 331258
rect 549884 331256 552631 331258
rect 549884 331200 552570 331256
rect 552626 331200 552631 331256
rect 549884 331198 552631 331200
rect 395540 331196 395546 331198
rect 552565 331195 552631 331198
rect 347957 331122 348023 331125
rect 347822 331120 348023 331122
rect 347822 331064 347962 331120
rect 348018 331064 348023 331120
rect 347822 331062 348023 331064
rect 347957 331059 348023 331062
rect 46473 330714 46539 330717
rect 348182 330714 348188 330716
rect 46473 330712 48116 330714
rect 46473 330656 46478 330712
rect 46534 330656 48116 330712
rect 46473 330654 48116 330656
rect 347852 330654 348188 330714
rect 46473 330651 46539 330654
rect 348182 330652 348188 330654
rect 348252 330652 348258 330716
rect 407113 330578 407179 330581
rect 407113 330576 410044 330578
rect 407113 330520 407118 330576
rect 407174 330520 410044 330576
rect 407113 330518 410044 330520
rect 407113 330515 407179 330518
rect 47485 329898 47551 329901
rect 48086 329898 48146 329936
rect 47485 329896 48146 329898
rect 47485 329840 47490 329896
rect 47546 329840 48146 329896
rect 47485 329838 48146 329840
rect 347822 329898 347882 329936
rect 350349 329898 350415 329901
rect 347822 329896 350415 329898
rect 347822 329840 350354 329896
rect 350410 329840 350415 329896
rect 347822 329838 350415 329840
rect 47485 329835 47551 329838
rect 350349 329835 350415 329838
rect 46473 328946 46539 328949
rect 48086 328946 48146 329256
rect 46473 328944 48146 328946
rect 46473 328888 46478 328944
rect 46534 328888 48146 328944
rect 46473 328886 48146 328888
rect 347822 328946 347882 329256
rect 350349 328946 350415 328949
rect 347822 328944 350415 328946
rect 347822 328888 350354 328944
rect 350410 328888 350415 328944
rect 347822 328886 350415 328888
rect 46473 328883 46539 328886
rect 350349 328883 350415 328886
rect 407113 328538 407179 328541
rect 407113 328536 410044 328538
rect 407113 328480 407118 328536
rect 407174 328480 410044 328536
rect 407113 328478 410044 328480
rect 407113 328475 407179 328478
rect 47301 327994 47367 327997
rect 47301 327992 48116 327994
rect 47301 327936 47306 327992
rect 47362 327936 48116 327992
rect 47301 327934 48116 327936
rect 47301 327931 47367 327934
rect 407113 327858 407179 327861
rect 553025 327858 553091 327861
rect 407113 327856 410044 327858
rect 407113 327800 407118 327856
rect 407174 327800 410044 327856
rect 407113 327798 410044 327800
rect 549884 327856 553091 327858
rect 549884 327800 553030 327856
rect 553086 327800 553091 327856
rect 549884 327798 553091 327800
rect 407113 327795 407179 327798
rect 553025 327795 553091 327798
rect 553117 327178 553183 327181
rect 549884 327176 553183 327178
rect 549884 327120 553122 327176
rect 553178 327120 553183 327176
rect 549884 327118 553183 327120
rect 553117 327115 553183 327118
rect 553025 326498 553091 326501
rect 549884 326496 553091 326498
rect 549884 326440 553030 326496
rect 553086 326440 553091 326496
rect 549884 326438 553091 326440
rect 553025 326435 553091 326438
rect 347822 325818 347882 325856
rect 350349 325818 350415 325821
rect 347822 325816 350415 325818
rect 347822 325760 350354 325816
rect 350410 325760 350415 325816
rect 347822 325758 350415 325760
rect 350349 325755 350415 325758
rect 407113 325818 407179 325821
rect 553117 325818 553183 325821
rect 407113 325816 410044 325818
rect 407113 325760 407118 325816
rect 407174 325760 410044 325816
rect 407113 325758 410044 325760
rect 549884 325816 553183 325818
rect 549884 325760 553122 325816
rect 553178 325760 553183 325816
rect 549884 325758 553183 325760
rect 407113 325755 407179 325758
rect 553117 325755 553183 325758
rect 46473 325274 46539 325277
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 46473 325272 48116 325274
rect 46473 325216 46478 325272
rect 46534 325216 48116 325272
rect 46473 325214 48116 325216
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 46473 325211 46539 325214
rect 580165 325211 580231 325214
rect 407205 325138 407271 325141
rect 407205 325136 410044 325138
rect 407205 325080 407210 325136
rect 407266 325080 410044 325136
rect 583520 325124 584960 325214
rect 407205 325078 410044 325080
rect 407205 325075 407271 325078
rect 350257 324594 350323 324597
rect 347852 324592 350323 324594
rect 347852 324536 350262 324592
rect 350318 324536 350323 324592
rect 347852 324534 350323 324536
rect 350257 324531 350323 324534
rect 407205 323778 407271 323781
rect 551001 323778 551067 323781
rect 407205 323776 410044 323778
rect 407205 323720 407210 323776
rect 407266 323720 410044 323776
rect 407205 323718 410044 323720
rect 549884 323776 551067 323778
rect 549884 323720 551006 323776
rect 551062 323720 551067 323776
rect 549884 323718 551067 323720
rect 407205 323715 407271 323718
rect 551001 323715 551067 323718
rect 46841 323098 46907 323101
rect 48086 323098 48146 323136
rect 46841 323096 48146 323098
rect 46841 323040 46846 323096
rect 46902 323040 48146 323096
rect 46841 323038 48146 323040
rect 407113 323098 407179 323101
rect 407113 323096 410044 323098
rect 407113 323040 407118 323096
rect 407174 323040 410044 323096
rect 407113 323038 410044 323040
rect 46841 323035 46907 323038
rect 407113 323035 407179 323038
rect 407205 322418 407271 322421
rect 552013 322418 552079 322421
rect 407205 322416 410044 322418
rect 407205 322360 407210 322416
rect 407266 322360 410044 322416
rect 407205 322358 410044 322360
rect 549884 322416 552079 322418
rect 549884 322360 552018 322416
rect 552074 322360 552079 322416
rect 549884 322358 552079 322360
rect 407205 322355 407271 322358
rect 552013 322355 552079 322358
rect 46841 321738 46907 321741
rect 48086 321738 48146 321776
rect 46841 321736 48146 321738
rect 46841 321680 46846 321736
rect 46902 321680 48146 321736
rect 46841 321678 48146 321680
rect 347822 321738 347882 321776
rect 350349 321738 350415 321741
rect 347822 321736 350415 321738
rect 347822 321680 350354 321736
rect 350410 321680 350415 321736
rect 347822 321678 350415 321680
rect 46841 321675 46907 321678
rect 350349 321675 350415 321678
rect 407113 321738 407179 321741
rect 407113 321736 410044 321738
rect 407113 321680 407118 321736
rect 407174 321680 410044 321736
rect 407113 321678 410044 321680
rect 407113 321675 407179 321678
rect 44725 321604 44791 321605
rect 44725 321602 44772 321604
rect 44680 321600 44772 321602
rect 44680 321544 44730 321600
rect 44680 321542 44772 321544
rect 44725 321540 44772 321542
rect 44836 321540 44842 321604
rect 44725 321539 44791 321540
rect 347822 320650 347882 321096
rect 407297 321058 407363 321061
rect 407297 321056 410044 321058
rect 407297 321000 407302 321056
rect 407358 321000 410044 321056
rect 407297 320998 410044 321000
rect 407297 320995 407363 320998
rect 350349 320650 350415 320653
rect 347822 320648 350415 320650
rect 347822 320592 350354 320648
rect 350410 320592 350415 320648
rect 347822 320590 350415 320592
rect 350349 320587 350415 320590
rect 46841 320242 46907 320245
rect 48086 320242 48146 320416
rect 46841 320240 48146 320242
rect 46841 320184 46846 320240
rect 46902 320184 48146 320240
rect 46841 320182 48146 320184
rect 46841 320179 46907 320182
rect -960 319140 480 319380
rect 347822 319290 347882 319736
rect 409873 319698 409939 319701
rect 409873 319696 410044 319698
rect 409873 319640 409878 319696
rect 409934 319640 410044 319696
rect 409873 319638 410044 319640
rect 409873 319635 409939 319638
rect 350349 319290 350415 319293
rect 347822 319288 350415 319290
rect 347822 319232 350354 319288
rect 350410 319232 350415 319288
rect 347822 319230 350415 319232
rect 350349 319227 350415 319230
rect 350257 319154 350323 319157
rect 347852 319152 350323 319154
rect 347852 319096 350262 319152
rect 350318 319096 350323 319152
rect 347852 319094 350323 319096
rect 350257 319091 350323 319094
rect 46841 319018 46907 319021
rect 48086 319018 48146 319056
rect 46841 319016 48146 319018
rect 46841 318960 46846 319016
rect 46902 318960 48146 319016
rect 46841 318958 48146 318960
rect 408401 319018 408467 319021
rect 408401 319016 410044 319018
rect 408401 318960 408406 319016
rect 408462 318960 410044 319016
rect 408401 318958 410044 318960
rect 46841 318955 46907 318958
rect 408401 318955 408467 318958
rect 46289 318474 46355 318477
rect 46289 318472 48116 318474
rect 46289 318416 46294 318472
rect 46350 318416 48116 318472
rect 46289 318414 48116 318416
rect 46289 318411 46355 318414
rect 347822 317794 347882 318376
rect 409413 318338 409479 318341
rect 553025 318338 553091 318341
rect 409413 318336 410044 318338
rect 409413 318280 409418 318336
rect 409474 318280 410044 318336
rect 409413 318278 410044 318280
rect 549884 318336 553091 318338
rect 549884 318280 553030 318336
rect 553086 318280 553091 318336
rect 549884 318278 553091 318280
rect 409413 318275 409479 318278
rect 553025 318275 553091 318278
rect 350349 317794 350415 317797
rect 347822 317792 350415 317794
rect 347822 317736 350354 317792
rect 350410 317736 350415 317792
rect 347822 317734 350415 317736
rect 350349 317731 350415 317734
rect 553117 317658 553183 317661
rect 549884 317656 553183 317658
rect 549884 317600 553122 317656
rect 553178 317600 553183 317656
rect 549884 317598 553183 317600
rect 553117 317595 553183 317598
rect 409781 316978 409847 316981
rect 409781 316976 410044 316978
rect 409781 316920 409786 316976
rect 409842 316920 410044 316976
rect 409781 316918 410044 316920
rect 409781 316915 409847 316918
rect 553117 316298 553183 316301
rect 549884 316296 553183 316298
rect 549884 316240 553122 316296
rect 553178 316240 553183 316296
rect 549884 316238 553183 316240
rect 553117 316235 553183 316238
rect 347822 315210 347882 315656
rect 407113 315618 407179 315621
rect 553710 315618 553716 315620
rect 407113 315616 410044 315618
rect 407113 315560 407118 315616
rect 407174 315560 410044 315616
rect 407113 315558 410044 315560
rect 549884 315558 553716 315618
rect 407113 315555 407179 315558
rect 553710 315556 553716 315558
rect 553780 315556 553786 315620
rect 350257 315210 350323 315213
rect 347822 315208 350323 315210
rect 347822 315152 350262 315208
rect 350318 315152 350323 315208
rect 347822 315150 350323 315152
rect 350257 315147 350323 315150
rect 350349 315074 350415 315077
rect 347852 315072 350415 315074
rect 347852 315016 350354 315072
rect 350410 315016 350415 315072
rect 347852 315014 350415 315016
rect 350349 315011 350415 315014
rect 46289 314802 46355 314805
rect 48086 314802 48146 314976
rect 553117 314938 553183 314941
rect 549884 314936 553183 314938
rect 549884 314880 553122 314936
rect 553178 314880 553183 314936
rect 549884 314878 553183 314880
rect 553117 314875 553183 314878
rect 46289 314800 48146 314802
rect 46289 314744 46294 314800
rect 46350 314744 48146 314800
rect 46289 314742 48146 314744
rect 46289 314739 46355 314742
rect 553025 314258 553091 314261
rect 549884 314256 553091 314258
rect 549884 314200 553030 314256
rect 553086 314200 553091 314256
rect 549884 314198 553091 314200
rect 553025 314195 553091 314198
rect 347822 312354 347882 312936
rect 408033 312898 408099 312901
rect 553117 312898 553183 312901
rect 408033 312896 410044 312898
rect 408033 312840 408038 312896
rect 408094 312840 410044 312896
rect 408033 312838 410044 312840
rect 549884 312896 553183 312898
rect 549884 312840 553122 312896
rect 553178 312840 553183 312896
rect 549884 312838 553183 312840
rect 408033 312835 408099 312838
rect 553117 312835 553183 312838
rect 350349 312354 350415 312357
rect 347822 312352 350415 312354
rect 347822 312296 350354 312352
rect 350410 312296 350415 312352
rect 347822 312294 350415 312296
rect 350349 312291 350415 312294
rect 580441 312082 580507 312085
rect 583520 312082 584960 312172
rect 580441 312080 584960 312082
rect 580441 312024 580446 312080
rect 580502 312024 584960 312080
rect 580441 312022 584960 312024
rect 580441 312019 580507 312022
rect 583520 311932 584960 312022
rect 46105 310994 46171 310997
rect 48086 310994 48146 311576
rect 347822 311130 347882 311576
rect 350073 311130 350139 311133
rect 347822 311128 350139 311130
rect 347822 311072 350078 311128
rect 350134 311072 350139 311128
rect 347822 311070 350139 311072
rect 350073 311067 350139 311070
rect 407205 311130 407271 311133
rect 410014 311130 410074 311440
rect 549884 311410 550282 311470
rect 550222 311402 550282 311410
rect 553025 311402 553091 311405
rect 550222 311400 553091 311402
rect 550222 311344 553030 311400
rect 553086 311344 553091 311400
rect 550222 311342 553091 311344
rect 553025 311339 553091 311342
rect 407205 311128 410074 311130
rect 407205 311072 407210 311128
rect 407266 311072 410074 311128
rect 407205 311070 410074 311072
rect 407205 311067 407271 311070
rect 46105 310992 48146 310994
rect 46105 310936 46110 310992
rect 46166 310936 48146 310992
rect 46105 310934 48146 310936
rect 46105 310931 46171 310934
rect 407113 310858 407179 310861
rect 553117 310858 553183 310861
rect 407113 310856 410044 310858
rect 407113 310800 407118 310856
rect 407174 310800 410044 310856
rect 407113 310798 410044 310800
rect 549884 310856 553183 310858
rect 549884 310800 553122 310856
rect 553178 310800 553183 310856
rect 549884 310798 553183 310800
rect 407113 310795 407179 310798
rect 553117 310795 553183 310798
rect 46289 310314 46355 310317
rect 46289 310312 48116 310314
rect 46289 310256 46294 310312
rect 46350 310256 48116 310312
rect 46289 310254 48116 310256
rect 46289 310251 46355 310254
rect 407113 310178 407179 310181
rect 553117 310178 553183 310181
rect 407113 310176 410044 310178
rect 407113 310120 407118 310176
rect 407174 310120 410044 310176
rect 407113 310118 410044 310120
rect 549884 310176 553183 310178
rect 549884 310120 553122 310176
rect 553178 310120 553183 310176
rect 549884 310118 553183 310120
rect 407113 310115 407179 310118
rect 553117 310115 553183 310118
rect 46105 309226 46171 309229
rect 48086 309226 48146 309536
rect 46105 309224 48146 309226
rect 46105 309168 46110 309224
rect 46166 309168 48146 309224
rect 46105 309166 48146 309168
rect 46105 309163 46171 309166
rect 347822 308410 347882 308856
rect 553117 308818 553183 308821
rect 549884 308816 553183 308818
rect 549884 308760 553122 308816
rect 553178 308760 553183 308816
rect 549884 308758 553183 308760
rect 553117 308755 553183 308758
rect 350349 308410 350415 308413
rect 347822 308408 350415 308410
rect 347822 308352 350354 308408
rect 350410 308352 350415 308408
rect 347822 308350 350415 308352
rect 350349 308347 350415 308350
rect 407113 308138 407179 308141
rect 407113 308136 410044 308138
rect 407113 308080 407118 308136
rect 407174 308080 410044 308136
rect 407113 308078 410044 308080
rect 407113 308075 407179 308078
rect 552013 307458 552079 307461
rect 549884 307456 552079 307458
rect 549884 307400 552018 307456
rect 552074 307400 552079 307456
rect 549884 307398 552079 307400
rect 552013 307395 552079 307398
rect 407113 306778 407179 306781
rect 407113 306776 410044 306778
rect 407113 306720 407118 306776
rect 407174 306720 410044 306776
rect 407113 306718 410044 306720
rect 407113 306715 407179 306718
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 409270 306036 409276 306100
rect 409340 306098 409346 306100
rect 552197 306098 552263 306101
rect 409340 306038 410044 306098
rect 549884 306096 552263 306098
rect 549884 306040 552202 306096
rect 552258 306040 552263 306096
rect 549884 306038 552263 306040
rect 409340 306036 409346 306038
rect 552197 306035 552263 306038
rect 407113 305418 407179 305421
rect 553117 305418 553183 305421
rect 407113 305416 410044 305418
rect 407113 305360 407118 305416
rect 407174 305360 410044 305416
rect 407113 305358 410044 305360
rect 549884 305416 553183 305418
rect 549884 305360 553122 305416
rect 553178 305360 553183 305416
rect 549884 305358 553183 305360
rect 407113 305355 407179 305358
rect 553117 305355 553183 305358
rect 41638 304948 41644 305012
rect 41708 305010 41714 305012
rect 47301 305010 47367 305013
rect 41708 305008 47367 305010
rect 41708 304952 47306 305008
rect 47362 304952 47367 305008
rect 41708 304950 47367 304952
rect 41708 304948 41714 304950
rect 47301 304947 47367 304950
rect 347822 304330 347882 304776
rect 350441 304330 350507 304333
rect 347822 304328 350507 304330
rect 347822 304272 350446 304328
rect 350502 304272 350507 304328
rect 347822 304270 350507 304272
rect 350441 304267 350507 304270
rect 41638 303588 41644 303652
rect 41708 303650 41714 303652
rect 48086 303650 48146 304096
rect 407113 304058 407179 304061
rect 407113 304056 410044 304058
rect 407113 304000 407118 304056
rect 407174 304000 410044 304056
rect 407113 303998 410044 304000
rect 407113 303995 407179 303998
rect 41708 303590 48146 303650
rect 41708 303588 41714 303590
rect 46381 302970 46447 302973
rect 48086 302970 48146 303416
rect 46381 302968 48146 302970
rect 46381 302912 46386 302968
rect 46442 302912 48146 302968
rect 46381 302910 48146 302912
rect 347822 302970 347882 303416
rect 350441 302970 350507 302973
rect 347822 302968 350507 302970
rect 347822 302912 350446 302968
rect 350502 302912 350507 302968
rect 347822 302910 350507 302912
rect 46381 302907 46447 302910
rect 350441 302907 350507 302910
rect 46289 302290 46355 302293
rect 46246 302288 46355 302290
rect 46246 302232 46294 302288
rect 46350 302232 46355 302288
rect 46246 302227 46355 302232
rect 347822 302290 347882 302736
rect 407941 302698 408007 302701
rect 407941 302696 410044 302698
rect 407941 302640 407946 302696
rect 408002 302640 410044 302696
rect 407941 302638 410044 302640
rect 407941 302635 408007 302638
rect 349153 302290 349219 302293
rect 347822 302288 349219 302290
rect 347822 302232 349158 302288
rect 349214 302232 349219 302288
rect 347822 302230 349219 302232
rect 349153 302227 349219 302230
rect 46246 302154 46306 302227
rect 46246 302094 48116 302154
rect 407205 302018 407271 302021
rect 553025 302018 553091 302021
rect 407205 302016 410044 302018
rect 407205 301960 407210 302016
rect 407266 301960 410044 302016
rect 407205 301958 410044 301960
rect 549884 302016 553091 302018
rect 549884 301960 553030 302016
rect 553086 301960 553091 302016
rect 549884 301958 553091 301960
rect 407205 301955 407271 301958
rect 553025 301955 553091 301958
rect 46381 300930 46447 300933
rect 48086 300930 48146 301376
rect 347822 301066 347882 301376
rect 407113 301338 407179 301341
rect 553117 301338 553183 301341
rect 407113 301336 410044 301338
rect 407113 301280 407118 301336
rect 407174 301280 410044 301336
rect 407113 301278 410044 301280
rect 549884 301336 553183 301338
rect 549884 301280 553122 301336
rect 553178 301280 553183 301336
rect 549884 301278 553183 301280
rect 407113 301275 407179 301278
rect 553117 301275 553183 301278
rect 350441 301066 350507 301069
rect 347822 301064 350507 301066
rect 347822 301008 350446 301064
rect 350502 301008 350507 301064
rect 347822 301006 350507 301008
rect 350441 301003 350507 301006
rect 46381 300928 48146 300930
rect 46381 300872 46386 300928
rect 46442 300872 48146 300928
rect 46381 300870 48146 300872
rect 46381 300867 46447 300870
rect 347822 300250 347882 300696
rect 407481 300658 407547 300661
rect 553117 300658 553183 300661
rect 407481 300656 410044 300658
rect 407481 300600 407486 300656
rect 407542 300600 410044 300656
rect 407481 300598 410044 300600
rect 549884 300656 553183 300658
rect 549884 300600 553122 300656
rect 553178 300600 553183 300656
rect 549884 300598 553183 300600
rect 407481 300595 407547 300598
rect 553117 300595 553183 300598
rect 350441 300250 350507 300253
rect 347822 300248 350507 300250
rect 347822 300192 350446 300248
rect 350502 300192 350507 300248
rect 347822 300190 350507 300192
rect 350441 300187 350507 300190
rect 407113 299978 407179 299981
rect 407113 299976 410044 299978
rect 407113 299920 407118 299976
rect 407174 299920 410044 299976
rect 407113 299918 410044 299920
rect 407113 299915 407179 299918
rect 347822 298890 347882 299336
rect 350441 298890 350507 298893
rect 347822 298888 350507 298890
rect 347822 298832 350446 298888
rect 350502 298832 350507 298888
rect 347822 298830 350507 298832
rect 350441 298827 350507 298830
rect 46381 298210 46447 298213
rect 48086 298210 48146 298656
rect 407573 298618 407639 298621
rect 407573 298616 410044 298618
rect 407573 298560 407578 298616
rect 407634 298560 410044 298616
rect 583520 298604 584960 298844
rect 407573 298558 410044 298560
rect 407573 298555 407639 298558
rect 46381 298208 48146 298210
rect 46381 298152 46386 298208
rect 46442 298152 48146 298208
rect 46381 298150 48146 298152
rect 46381 298147 46447 298150
rect 47209 298074 47275 298077
rect 47209 298072 48116 298074
rect 47209 298016 47214 298072
rect 47270 298016 48116 298072
rect 47209 298014 48116 298016
rect 47209 298011 47275 298014
rect 550081 297938 550147 297941
rect 549884 297936 550147 297938
rect 549884 297880 550086 297936
rect 550142 297880 550147 297936
rect 549884 297878 550147 297880
rect 550081 297875 550147 297878
rect 46381 297122 46447 297125
rect 48086 297122 48146 297296
rect 553117 297258 553183 297261
rect 549884 297256 553183 297258
rect 549884 297200 553122 297256
rect 553178 297200 553183 297256
rect 549884 297198 553183 297200
rect 553117 297195 553183 297198
rect 46381 297120 48146 297122
rect 46381 297064 46386 297120
rect 46442 297064 48146 297120
rect 46381 297062 48146 297064
rect 46381 297059 46447 297062
rect 350441 296714 350507 296717
rect 347852 296712 350507 296714
rect 347852 296656 350446 296712
rect 350502 296656 350507 296712
rect 347852 296654 350507 296656
rect 350441 296651 350507 296654
rect 348049 296442 348115 296445
rect 347822 296440 348115 296442
rect 347822 296384 348054 296440
rect 348110 296384 348115 296440
rect 347822 296382 348115 296384
rect 347822 296004 347882 296382
rect 348049 296379 348115 296382
rect 407113 295898 407179 295901
rect 407113 295896 410044 295898
rect 407113 295840 407118 295896
rect 407174 295840 410044 295896
rect 407113 295838 410044 295840
rect 407113 295835 407179 295838
rect 349429 295492 349495 295493
rect 349429 295490 349476 295492
rect 349384 295488 349476 295490
rect 349384 295432 349434 295488
rect 349384 295430 349476 295432
rect 349429 295428 349476 295430
rect 349540 295428 349546 295492
rect 349429 295427 349495 295428
rect 350441 295354 350507 295357
rect 347852 295352 350507 295354
rect 347852 295296 350446 295352
rect 350502 295296 350507 295352
rect 347852 295294 350507 295296
rect 350441 295291 350507 295294
rect 350441 293994 350507 293997
rect 347852 293992 350507 293994
rect 347852 293936 350446 293992
rect 350502 293936 350507 293992
rect 347852 293934 350507 293936
rect 350441 293931 350507 293934
rect 408401 293994 408467 293997
rect 410014 293994 410074 294440
rect 408401 293992 410074 293994
rect 408401 293936 408406 293992
rect 408462 293936 410074 293992
rect 408401 293934 410074 293936
rect 408401 293931 408467 293934
rect 407205 293858 407271 293861
rect 407205 293856 410044 293858
rect 407205 293800 407210 293856
rect 407266 293800 410044 293856
rect 407205 293798 410044 293800
rect 407205 293795 407271 293798
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 46381 292906 46447 292909
rect 48086 292906 48146 293216
rect 404854 293116 404860 293180
rect 404924 293178 404930 293180
rect 552013 293178 552079 293181
rect 404924 293118 410044 293178
rect 549884 293176 552079 293178
rect 549884 293120 552018 293176
rect 552074 293120 552079 293176
rect 549884 293118 552079 293120
rect 404924 293116 404930 293118
rect 552013 293115 552079 293118
rect 554037 293178 554103 293181
rect 566222 293178 566228 293180
rect 554037 293176 566228 293178
rect 554037 293120 554042 293176
rect 554098 293120 566228 293176
rect 554037 293118 566228 293120
rect 554037 293115 554103 293118
rect 566222 293116 566228 293118
rect 566292 293116 566298 293180
rect 46381 292904 48146 292906
rect 46381 292848 46386 292904
rect 46442 292848 48146 292904
rect 46381 292846 48146 292848
rect 46381 292843 46447 292846
rect 43621 292634 43687 292637
rect 44766 292634 44772 292636
rect 43621 292632 44772 292634
rect 43621 292576 43626 292632
rect 43682 292576 44772 292632
rect 43621 292574 44772 292576
rect 43621 292571 43687 292574
rect 44766 292572 44772 292574
rect 44836 292572 44842 292636
rect 46105 292634 46171 292637
rect 46105 292632 48116 292634
rect 46105 292576 46110 292632
rect 46166 292576 48116 292632
rect 46105 292574 48116 292576
rect 46105 292571 46171 292574
rect 407113 292498 407179 292501
rect 553117 292498 553183 292501
rect 407113 292496 410044 292498
rect 407113 292440 407118 292496
rect 407174 292440 410044 292496
rect 407113 292438 410044 292440
rect 549884 292496 553183 292498
rect 549884 292440 553122 292496
rect 553178 292440 553183 292496
rect 549884 292438 553183 292440
rect 407113 292435 407179 292438
rect 553117 292435 553183 292438
rect 46381 291546 46447 291549
rect 48086 291546 48146 291856
rect 407205 291818 407271 291821
rect 552013 291818 552079 291821
rect 407205 291816 410044 291818
rect 407205 291760 407210 291816
rect 407266 291760 410044 291816
rect 407205 291758 410044 291760
rect 549884 291816 552079 291818
rect 549884 291760 552018 291816
rect 552074 291760 552079 291816
rect 549884 291758 552079 291760
rect 407205 291755 407271 291758
rect 552013 291755 552079 291758
rect 46381 291544 48146 291546
rect 46381 291488 46386 291544
rect 46442 291488 48146 291544
rect 46381 291486 48146 291488
rect 46381 291483 46447 291486
rect 553117 290458 553183 290461
rect 549884 290456 553183 290458
rect 549884 290400 553122 290456
rect 553178 290400 553183 290456
rect 549884 290398 553183 290400
rect 553117 290395 553183 290398
rect 407113 289778 407179 289781
rect 553025 289778 553091 289781
rect 407113 289776 410044 289778
rect 407113 289720 407118 289776
rect 407174 289720 410044 289776
rect 407113 289718 410044 289720
rect 549884 289776 553091 289778
rect 549884 289720 553030 289776
rect 553086 289720 553091 289776
rect 549884 289718 553091 289720
rect 407113 289715 407179 289718
rect 553025 289715 553091 289718
rect 347822 288826 347882 289136
rect 407297 289098 407363 289101
rect 553117 289098 553183 289101
rect 407297 289096 410044 289098
rect 407297 289040 407302 289096
rect 407358 289040 410044 289096
rect 407297 289038 410044 289040
rect 549884 289096 553183 289098
rect 549884 289040 553122 289096
rect 553178 289040 553183 289096
rect 549884 289038 553183 289040
rect 407297 289035 407363 289038
rect 553117 289035 553183 289038
rect 350441 288826 350507 288829
rect 347822 288824 350507 288826
rect 347822 288768 350446 288824
rect 350502 288768 350507 288824
rect 347822 288766 350507 288768
rect 350441 288763 350507 288766
rect 349245 288554 349311 288557
rect 347852 288552 349311 288554
rect 347852 288496 349250 288552
rect 349306 288496 349311 288552
rect 347852 288494 349311 288496
rect 349245 288491 349311 288494
rect 47526 288424 47532 288488
rect 47596 288486 47602 288488
rect 47596 288426 48116 288486
rect 47596 288424 47602 288426
rect 407205 288418 407271 288421
rect 407205 288416 410044 288418
rect 407205 288360 407210 288416
rect 407266 288360 410044 288416
rect 407205 288358 410044 288360
rect 407205 288355 407271 288358
rect 347822 287194 347882 287776
rect 407113 287738 407179 287741
rect 553117 287738 553183 287741
rect 407113 287736 410044 287738
rect 407113 287680 407118 287736
rect 407174 287680 410044 287736
rect 407113 287678 410044 287680
rect 549884 287736 553183 287738
rect 549884 287680 553122 287736
rect 553178 287680 553183 287736
rect 549884 287678 553183 287680
rect 407113 287675 407179 287678
rect 553117 287675 553183 287678
rect 350441 287194 350507 287197
rect 347822 287192 350507 287194
rect 347822 287136 350446 287192
rect 350502 287136 350507 287192
rect 347822 287134 350507 287136
rect 350441 287131 350507 287134
rect 407113 287058 407179 287061
rect 407113 287056 410044 287058
rect 407113 287000 407118 287056
rect 407174 287000 410044 287056
rect 407113 286998 410044 287000
rect 407113 286995 407179 286998
rect 347998 286786 348004 286788
rect 347822 286726 348004 286786
rect 347822 286484 347882 286726
rect 347998 286724 348004 286726
rect 348068 286724 348074 286788
rect 46381 285834 46447 285837
rect 48086 285834 48146 286416
rect 567694 286378 567700 286380
rect 549884 286318 567700 286378
rect 567694 286316 567700 286318
rect 567764 286316 567770 286380
rect 350441 285834 350507 285837
rect 46381 285832 48146 285834
rect 46381 285776 46386 285832
rect 46442 285776 48146 285832
rect 46381 285774 48146 285776
rect 347852 285832 350507 285834
rect 347852 285776 350446 285832
rect 350502 285776 350507 285832
rect 347852 285774 350507 285776
rect 46381 285771 46447 285774
rect 350441 285771 350507 285774
rect 583520 285276 584960 285516
rect 350349 285154 350415 285157
rect 347852 285152 350415 285154
rect 347852 285096 350354 285152
rect 350410 285096 350415 285152
rect 347852 285094 350415 285096
rect 350349 285091 350415 285094
rect 409137 285018 409203 285021
rect 409137 285016 410044 285018
rect 409137 284960 409142 285016
rect 409198 284960 410044 285016
rect 409137 284958 410044 284960
rect 409137 284955 409203 284958
rect 46238 284276 46244 284340
rect 46308 284338 46314 284340
rect 48086 284338 48146 284376
rect 46308 284278 48146 284338
rect 347822 284338 347882 284376
rect 349429 284338 349495 284341
rect 347822 284336 349495 284338
rect 347822 284280 349434 284336
rect 349490 284280 349495 284336
rect 347822 284278 349495 284280
rect 46308 284276 46314 284278
rect 349429 284275 349495 284278
rect 407113 284338 407179 284341
rect 407113 284336 410044 284338
rect 407113 284280 407118 284336
rect 407174 284280 410044 284336
rect 407113 284278 410044 284280
rect 407113 284275 407179 284278
rect 44909 283250 44975 283253
rect 48086 283250 48146 283696
rect 407205 283658 407271 283661
rect 553117 283658 553183 283661
rect 407205 283656 410044 283658
rect 407205 283600 407210 283656
rect 407266 283600 410044 283656
rect 407205 283598 410044 283600
rect 549884 283656 553183 283658
rect 549884 283600 553122 283656
rect 553178 283600 553183 283656
rect 549884 283598 553183 283600
rect 407205 283595 407271 283598
rect 553117 283595 553183 283598
rect 44909 283248 48146 283250
rect 44909 283192 44914 283248
rect 44970 283192 48146 283248
rect 44909 283190 48146 283192
rect 44909 283187 44975 283190
rect 46422 282916 46428 282980
rect 46492 282978 46498 282980
rect 47393 282978 47459 282981
rect 46492 282976 47459 282978
rect 46492 282920 47398 282976
rect 47454 282920 47459 282976
rect 46492 282918 47459 282920
rect 46492 282916 46498 282918
rect 47393 282915 47459 282918
rect 407113 282978 407179 282981
rect 407113 282976 410044 282978
rect 407113 282920 407118 282976
rect 407174 282920 410044 282976
rect 407113 282918 410044 282920
rect 407113 282915 407179 282918
rect 46841 281890 46907 281893
rect 48086 281890 48146 282336
rect 551369 282298 551435 282301
rect 549884 282296 551435 282298
rect 549884 282240 551374 282296
rect 551430 282240 551435 282296
rect 549884 282238 551435 282240
rect 551369 282235 551435 282238
rect 46841 281888 48146 281890
rect 46841 281832 46846 281888
rect 46902 281832 48146 281888
rect 46841 281830 48146 281832
rect 46841 281827 46907 281830
rect 45645 281618 45711 281621
rect 48086 281618 48146 281656
rect 553117 281618 553183 281621
rect 45645 281616 48146 281618
rect 45645 281560 45650 281616
rect 45706 281560 48146 281616
rect 45645 281558 48146 281560
rect 549884 281616 553183 281618
rect 549884 281560 553122 281616
rect 553178 281560 553183 281616
rect 549884 281558 553183 281560
rect 45645 281555 45711 281558
rect 553117 281555 553183 281558
rect 347822 280530 347882 280976
rect 553025 280938 553091 280941
rect 549884 280936 553091 280938
rect 549884 280880 553030 280936
rect 553086 280880 553091 280936
rect 549884 280878 553091 280880
rect 553025 280875 553091 280878
rect 349245 280530 349311 280533
rect 347822 280528 349311 280530
rect 347822 280472 349250 280528
rect 349306 280472 349311 280528
rect 347822 280470 349311 280472
rect 349245 280467 349311 280470
rect 553117 280258 553183 280261
rect 549884 280256 553183 280258
rect -960 279972 480 280212
rect 549884 280200 553122 280256
rect 553178 280200 553183 280256
rect 549884 280198 553183 280200
rect 553117 280195 553183 280198
rect 350717 279714 350783 279717
rect 347852 279712 350783 279714
rect 347852 279656 350722 279712
rect 350778 279656 350783 279712
rect 347852 279654 350783 279656
rect 350717 279651 350783 279654
rect 407205 279578 407271 279581
rect 553117 279578 553183 279581
rect 407205 279576 410044 279578
rect 407205 279520 407210 279576
rect 407266 279520 410044 279576
rect 407205 279518 410044 279520
rect 549884 279576 553183 279578
rect 549884 279520 553122 279576
rect 553178 279520 553183 279576
rect 549884 279518 553183 279520
rect 407205 279515 407271 279518
rect 553117 279515 553183 279518
rect 407113 278898 407179 278901
rect 553117 278898 553183 278901
rect 407113 278896 410044 278898
rect 407113 278840 407118 278896
rect 407174 278840 410044 278896
rect 407113 278838 410044 278840
rect 549884 278896 553183 278898
rect 549884 278840 553122 278896
rect 553178 278840 553183 278896
rect 549884 278838 553183 278840
rect 407113 278835 407179 278838
rect 553117 278835 553183 278838
rect 354438 278762 354444 278764
rect 347822 278702 354444 278762
rect 347822 278324 347882 278702
rect 354438 278700 354444 278702
rect 354508 278700 354514 278764
rect 46841 277810 46907 277813
rect 48086 277810 48146 278256
rect 46841 277808 48146 277810
rect 46841 277752 46846 277808
rect 46902 277752 48146 277808
rect 46841 277750 48146 277752
rect 46841 277747 46907 277750
rect 347822 277538 347882 277576
rect 350441 277538 350507 277541
rect 347822 277536 350507 277538
rect 347822 277480 350446 277536
rect 350502 277480 350507 277536
rect 347822 277478 350507 277480
rect 350441 277475 350507 277478
rect 409638 277476 409644 277540
rect 409708 277538 409714 277540
rect 553117 277538 553183 277541
rect 409708 277478 410044 277538
rect 550222 277536 553183 277538
rect 550222 277480 553122 277536
rect 553178 277480 553183 277536
rect 550222 277478 553183 277480
rect 409708 277476 409714 277478
rect 550222 277470 550282 277478
rect 553117 277475 553183 277478
rect 549884 277410 550282 277470
rect 407849 276858 407915 276861
rect 407849 276856 410044 276858
rect 407849 276800 407854 276856
rect 407910 276800 410044 276856
rect 407849 276798 410044 276800
rect 407849 276795 407915 276798
rect 347822 276042 347882 276216
rect 407113 276178 407179 276181
rect 553025 276178 553091 276181
rect 407113 276176 410044 276178
rect 407113 276120 407118 276176
rect 407174 276120 410044 276176
rect 407113 276118 410044 276120
rect 549884 276176 553091 276178
rect 549884 276120 553030 276176
rect 553086 276120 553091 276176
rect 549884 276118 553091 276120
rect 407113 276115 407179 276118
rect 553025 276115 553091 276118
rect 350717 276042 350783 276045
rect 347822 276040 350783 276042
rect 347822 275984 350722 276040
rect 350778 275984 350783 276040
rect 347822 275982 350783 275984
rect 350717 275979 350783 275982
rect 350441 275634 350507 275637
rect 347852 275632 350507 275634
rect 347852 275576 350446 275632
rect 350502 275576 350507 275632
rect 347852 275574 350507 275576
rect 350441 275571 350507 275574
rect 407113 275498 407179 275501
rect 407113 275496 410044 275498
rect 407113 275440 407118 275496
rect 407174 275440 410044 275496
rect 407113 275438 410044 275440
rect 407113 275435 407179 275438
rect 553117 274818 553183 274821
rect 549884 274816 553183 274818
rect 549884 274760 553122 274816
rect 553178 274760 553183 274816
rect 549884 274758 553183 274760
rect 553117 274755 553183 274758
rect 46841 273730 46907 273733
rect 48086 273730 48146 274176
rect 347822 273866 347882 274176
rect 350349 273866 350415 273869
rect 347822 273864 350415 273866
rect 347822 273808 350354 273864
rect 350410 273808 350415 273864
rect 347822 273806 350415 273808
rect 350349 273803 350415 273806
rect 46841 273728 48146 273730
rect 46841 273672 46846 273728
rect 46902 273672 48146 273728
rect 46841 273670 48146 273672
rect 46841 273667 46907 273670
rect 47209 273322 47275 273325
rect 48086 273322 48146 273496
rect 347822 273458 347882 273496
rect 350441 273458 350507 273461
rect 553117 273458 553183 273461
rect 347822 273456 350507 273458
rect 347822 273400 350446 273456
rect 350502 273400 350507 273456
rect 347822 273398 350507 273400
rect 549884 273456 553183 273458
rect 549884 273400 553122 273456
rect 553178 273400 553183 273456
rect 549884 273398 553183 273400
rect 350441 273395 350507 273398
rect 553117 273395 553183 273398
rect 47209 273320 48146 273322
rect 47209 273264 47214 273320
rect 47270 273264 48146 273320
rect 47209 273262 48146 273264
rect 47209 273259 47275 273262
rect 347822 272234 347882 272816
rect 403934 272716 403940 272780
rect 404004 272778 404010 272780
rect 404004 272718 410044 272778
rect 404004 272716 404010 272718
rect 350809 272234 350875 272237
rect 347822 272232 350875 272234
rect 347822 272176 350814 272232
rect 350870 272176 350875 272232
rect 347822 272174 350875 272176
rect 350809 272171 350875 272174
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 407113 271418 407179 271421
rect 550725 271418 550791 271421
rect 407113 271416 410044 271418
rect 407113 271360 407118 271416
rect 407174 271360 410044 271416
rect 407113 271358 410044 271360
rect 549884 271416 550791 271418
rect 549884 271360 550730 271416
rect 550786 271360 550791 271416
rect 549884 271358 550791 271360
rect 407113 271355 407179 271358
rect 550725 271355 550791 271358
rect 553117 270738 553183 270741
rect 549884 270736 553183 270738
rect 549884 270680 553122 270736
rect 553178 270680 553183 270736
rect 549884 270678 553183 270680
rect 553117 270675 553183 270678
rect 47117 270194 47183 270197
rect 350441 270194 350507 270197
rect 47117 270192 48116 270194
rect 47117 270136 47122 270192
rect 47178 270136 48116 270192
rect 47117 270134 48116 270136
rect 347852 270192 350507 270194
rect 347852 270136 350446 270192
rect 350502 270136 350507 270192
rect 347852 270134 350507 270136
rect 47117 270131 47183 270134
rect 350441 270131 350507 270134
rect 407113 270058 407179 270061
rect 407113 270056 410044 270058
rect 407113 270000 407118 270056
rect 407174 270000 410044 270056
rect 407113 269998 410044 270000
rect 407113 269995 407179 269998
rect 349981 268834 350047 268837
rect 347852 268832 350047 268834
rect 347852 268776 349986 268832
rect 350042 268776 350047 268832
rect 347852 268774 350047 268776
rect 349981 268771 350047 268774
rect 46473 268290 46539 268293
rect 48086 268290 48146 268736
rect 550725 268698 550791 268701
rect 549884 268696 550791 268698
rect 549884 268640 550730 268696
rect 550786 268640 550791 268696
rect 549884 268638 550791 268640
rect 550725 268635 550791 268638
rect 46473 268288 48146 268290
rect 46473 268232 46478 268288
rect 46534 268232 48146 268288
rect 46473 268230 48146 268232
rect 46473 268227 46539 268230
rect 350441 268154 350507 268157
rect 347852 268152 350507 268154
rect 347852 268096 350446 268152
rect 350502 268096 350507 268152
rect 347852 268094 350507 268096
rect 350441 268091 350507 268094
rect 46381 267882 46447 267885
rect 48086 267882 48146 268056
rect 407113 268018 407179 268021
rect 407113 268016 410044 268018
rect 407113 267960 407118 268016
rect 407174 267960 410044 268016
rect 407113 267958 410044 267960
rect 407113 267955 407179 267958
rect 46381 267880 48146 267882
rect 46381 267824 46386 267880
rect 46442 267824 48146 267880
rect 46381 267822 48146 267824
rect 46381 267819 46447 267822
rect -960 267052 480 267292
rect 347822 266794 347882 267376
rect 407757 267338 407823 267341
rect 407757 267336 410044 267338
rect 407757 267280 407762 267336
rect 407818 267280 410044 267336
rect 407757 267278 410044 267280
rect 407757 267275 407823 267278
rect 350441 266794 350507 266797
rect 347822 266792 350507 266794
rect 347822 266736 350446 266792
rect 350502 266736 350507 266792
rect 347822 266734 350507 266736
rect 350441 266731 350507 266734
rect 553117 266658 553183 266661
rect 549884 266656 553183 266658
rect 549884 266600 553122 266656
rect 553178 266600 553183 266656
rect 549884 266598 553183 266600
rect 553117 266595 553183 266598
rect 552013 265298 552079 265301
rect 549884 265296 552079 265298
rect 549884 265240 552018 265296
rect 552074 265240 552079 265296
rect 549884 265238 552079 265240
rect 552013 265235 552079 265238
rect 355358 264964 355364 265028
rect 355428 265026 355434 265028
rect 360377 265026 360443 265029
rect 355428 265024 360443 265026
rect 355428 264968 360382 265024
rect 360438 264968 360443 265024
rect 355428 264966 360443 264968
rect 355428 264964 355434 264966
rect 360377 264963 360443 264966
rect 45185 264754 45251 264757
rect 45185 264752 48116 264754
rect 45185 264696 45190 264752
rect 45246 264696 48116 264752
rect 45185 264694 48116 264696
rect 45185 264691 45251 264694
rect 552841 264618 552907 264621
rect 549884 264616 552907 264618
rect 549884 264560 552846 264616
rect 552902 264560 552907 264616
rect 549884 264558 552907 264560
rect 552841 264555 552907 264558
rect 347822 263938 347882 263976
rect 350441 263938 350507 263941
rect 347822 263936 350507 263938
rect 347822 263880 350446 263936
rect 350502 263880 350507 263936
rect 347822 263878 350507 263880
rect 350441 263875 350507 263878
rect 407113 263938 407179 263941
rect 553117 263938 553183 263941
rect 407113 263936 410044 263938
rect 407113 263880 407118 263936
rect 407174 263880 410044 263936
rect 407113 263878 410044 263880
rect 549884 263936 553183 263938
rect 549884 263880 553122 263936
rect 553178 263880 553183 263936
rect 549884 263878 553183 263880
rect 407113 263875 407179 263878
rect 553117 263875 553183 263878
rect 347822 262850 347882 263296
rect 552013 263258 552079 263261
rect 549884 263256 552079 263258
rect 549884 263200 552018 263256
rect 552074 263200 552079 263256
rect 549884 263198 552079 263200
rect 552013 263195 552079 263198
rect 362902 262924 362908 262988
rect 362972 262986 362978 262988
rect 364241 262986 364307 262989
rect 362972 262984 364307 262986
rect 362972 262928 364246 262984
rect 364302 262928 364307 262984
rect 362972 262926 364307 262928
rect 362972 262924 362978 262926
rect 364241 262923 364307 262926
rect 348049 262850 348115 262853
rect 347822 262848 348115 262850
rect 347822 262792 348054 262848
rect 348110 262792 348115 262848
rect 347822 262790 348115 262792
rect 348049 262787 348115 262790
rect 350625 262714 350691 262717
rect 347852 262712 350691 262714
rect 347852 262656 350630 262712
rect 350686 262656 350691 262712
rect 347852 262654 350691 262656
rect 350625 262651 350691 262654
rect 31334 262244 31340 262308
rect 31404 262306 31410 262308
rect 48086 262306 48146 262616
rect 407113 262578 407179 262581
rect 550398 262578 550404 262580
rect 407113 262576 410044 262578
rect 407113 262520 407118 262576
rect 407174 262520 410044 262576
rect 407113 262518 410044 262520
rect 549884 262518 550404 262578
rect 407113 262515 407179 262518
rect 550398 262516 550404 262518
rect 550468 262516 550474 262580
rect 31404 262246 48146 262306
rect 31404 262244 31410 262246
rect 407113 261898 407179 261901
rect 552013 261898 552079 261901
rect 407113 261896 410044 261898
rect 407113 261840 407118 261896
rect 407174 261840 410044 261896
rect 407113 261838 410044 261840
rect 549884 261896 552079 261898
rect 549884 261840 552018 261896
rect 552074 261840 552079 261896
rect 549884 261838 552079 261840
rect 407113 261835 407179 261838
rect 552013 261835 552079 261838
rect 350441 261354 350507 261357
rect 347852 261352 350507 261354
rect 347852 261296 350446 261352
rect 350502 261296 350507 261352
rect 347852 261294 350507 261296
rect 350441 261291 350507 261294
rect 408401 259994 408467 259997
rect 410014 259994 410074 260440
rect 549884 260410 550466 260470
rect 550406 260402 550466 260410
rect 552105 260402 552171 260405
rect 550406 260400 552171 260402
rect 550406 260344 552110 260400
rect 552166 260344 552171 260400
rect 550406 260342 552171 260344
rect 552105 260339 552171 260342
rect 408401 259992 410074 259994
rect 408401 259936 408406 259992
rect 408462 259936 410074 259992
rect 408401 259934 410074 259936
rect 408401 259931 408467 259934
rect 407113 259858 407179 259861
rect 552013 259858 552079 259861
rect 407113 259856 410044 259858
rect 407113 259800 407118 259856
rect 407174 259800 410044 259856
rect 407113 259798 410044 259800
rect 549884 259856 552079 259858
rect 549884 259800 552018 259856
rect 552074 259800 552079 259856
rect 549884 259798 552079 259800
rect 407113 259795 407179 259798
rect 552013 259795 552079 259798
rect 347822 258770 347882 259216
rect 552105 259178 552171 259181
rect 549884 259176 552171 259178
rect 549884 259120 552110 259176
rect 552166 259120 552171 259176
rect 549884 259118 552171 259120
rect 552105 259115 552171 259118
rect 579061 258906 579127 258909
rect 583520 258906 584960 258996
rect 579061 258904 584960 258906
rect 579061 258848 579066 258904
rect 579122 258848 584960 258904
rect 579061 258846 584960 258848
rect 579061 258843 579127 258846
rect 350441 258770 350507 258773
rect 347822 258768 350507 258770
rect 347822 258712 350446 258768
rect 350502 258712 350507 258768
rect 583520 258756 584960 258846
rect 347822 258710 350507 258712
rect 350441 258707 350507 258710
rect 46013 258362 46079 258365
rect 48086 258362 48146 258536
rect 552013 258498 552079 258501
rect 549884 258496 552079 258498
rect 549884 258440 552018 258496
rect 552074 258440 552079 258496
rect 549884 258438 552079 258440
rect 552013 258435 552079 258438
rect 46013 258360 48146 258362
rect 46013 258304 46018 258360
rect 46074 258304 48146 258360
rect 46013 258302 48146 258304
rect 46013 258299 46079 258302
rect 47669 257954 47735 257957
rect 349889 257954 349955 257957
rect 47669 257952 48116 257954
rect 47669 257896 47674 257952
rect 47730 257896 48116 257952
rect 47669 257894 48116 257896
rect 347852 257952 349955 257954
rect 347852 257896 349894 257952
rect 349950 257896 349955 257952
rect 347852 257894 349955 257896
rect 47669 257891 47735 257894
rect 349889 257891 349955 257894
rect 407205 257818 407271 257821
rect 552013 257818 552079 257821
rect 407205 257816 410044 257818
rect 407205 257760 407210 257816
rect 407266 257760 410044 257816
rect 407205 257758 410044 257760
rect 549884 257816 552079 257818
rect 549884 257760 552018 257816
rect 552074 257760 552079 257816
rect 549884 257758 552079 257760
rect 407205 257755 407271 257758
rect 552013 257755 552079 257758
rect 46473 256730 46539 256733
rect 48086 256730 48146 257176
rect 407113 257138 407179 257141
rect 407113 257136 410044 257138
rect 407113 257080 407118 257136
rect 407174 257080 410044 257136
rect 407113 257078 410044 257080
rect 407113 257075 407179 257078
rect 46473 256728 48146 256730
rect 46473 256672 46478 256728
rect 46534 256672 48146 256728
rect 46473 256670 48146 256672
rect 46473 256667 46539 256670
rect 347822 256050 347882 256496
rect 350349 256050 350415 256053
rect 347822 256048 350415 256050
rect 347822 255992 350354 256048
rect 350410 255992 350415 256048
rect 347822 255990 350415 255992
rect 350349 255987 350415 255990
rect 347822 255370 347882 255816
rect 350441 255370 350507 255373
rect 347822 255368 350507 255370
rect 347822 255312 350446 255368
rect 350502 255312 350507 255368
rect 347822 255310 350507 255312
rect 350441 255307 350507 255310
rect 407113 255098 407179 255101
rect 552105 255098 552171 255101
rect 407113 255096 410044 255098
rect 407113 255040 407118 255096
rect 407174 255040 410044 255096
rect 407113 255038 410044 255040
rect 549884 255096 552171 255098
rect 549884 255040 552110 255096
rect 552166 255040 552171 255096
rect 549884 255038 552171 255040
rect 407113 255035 407179 255038
rect 552105 255035 552171 255038
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 26877 254010 26943 254013
rect 27470 254010 27476 254012
rect 26877 254008 27476 254010
rect 26877 253952 26882 254008
rect 26938 253952 27476 254008
rect 26877 253950 27476 253952
rect 26877 253947 26943 253950
rect 27470 253948 27476 253950
rect 27540 253948 27546 254012
rect 46841 254010 46907 254013
rect 48086 254010 48146 254456
rect 46841 254008 48146 254010
rect 46841 253952 46846 254008
rect 46902 253952 48146 254008
rect 46841 253950 48146 253952
rect 347822 254010 347882 254456
rect 407481 254418 407547 254421
rect 552013 254418 552079 254421
rect 407481 254416 410044 254418
rect 407481 254360 407486 254416
rect 407542 254360 410044 254416
rect 407481 254358 410044 254360
rect 549884 254416 552079 254418
rect 549884 254360 552018 254416
rect 552074 254360 552079 254416
rect 549884 254358 552079 254360
rect 407481 254355 407547 254358
rect 552013 254355 552079 254358
rect 350441 254010 350507 254013
rect 347822 254008 350507 254010
rect 347822 253952 350446 254008
rect 350502 253952 350507 254008
rect 347822 253950 350507 253952
rect 46841 253947 46907 253950
rect 350441 253947 350507 253950
rect 553117 253738 553183 253741
rect 549884 253736 553183 253738
rect 549884 253680 553122 253736
rect 553178 253680 553183 253736
rect 549884 253678 553183 253680
rect 553117 253675 553183 253678
rect 553117 252378 553183 252381
rect 549884 252376 553183 252378
rect 549884 252320 553122 252376
rect 553178 252320 553183 252376
rect 549884 252318 553183 252320
rect 553117 252315 553183 252318
rect 45369 251834 45435 251837
rect 45369 251832 48116 251834
rect 45369 251776 45374 251832
rect 45430 251776 48116 251832
rect 45369 251774 48116 251776
rect 45369 251771 45435 251774
rect 407113 251698 407179 251701
rect 407113 251696 410044 251698
rect 407113 251640 407118 251696
rect 407174 251640 410044 251696
rect 407113 251638 410044 251640
rect 407113 251635 407179 251638
rect 407113 251018 407179 251021
rect 407113 251016 410044 251018
rect 407113 250960 407118 251016
rect 407174 250960 410044 251016
rect 407113 250958 410044 250960
rect 407113 250955 407179 250958
rect 347822 250202 347882 250376
rect 407205 250338 407271 250341
rect 552013 250338 552079 250341
rect 407205 250336 410044 250338
rect 407205 250280 407210 250336
rect 407266 250280 410044 250336
rect 407205 250278 410044 250280
rect 549884 250336 552079 250338
rect 549884 250280 552018 250336
rect 552074 250280 552079 250336
rect 549884 250278 552079 250280
rect 407205 250275 407271 250278
rect 552013 250275 552079 250278
rect 350441 250202 350507 250205
rect 347822 250200 350507 250202
rect 347822 250144 350446 250200
rect 350502 250144 350507 250200
rect 347822 250142 350507 250144
rect 350441 250139 350507 250142
rect 407757 249658 407823 249661
rect 566038 249658 566044 249660
rect 407757 249656 410044 249658
rect 407757 249600 407762 249656
rect 407818 249600 410044 249656
rect 407757 249598 410044 249600
rect 549884 249598 566044 249658
rect 407757 249595 407823 249598
rect 566038 249596 566044 249598
rect 566108 249596 566114 249660
rect 347822 248842 347882 249016
rect 350441 248842 350507 248845
rect 347822 248840 350507 248842
rect 347822 248784 350446 248840
rect 350502 248784 350507 248840
rect 347822 248782 350507 248784
rect 350441 248779 350507 248782
rect 553117 248298 553183 248301
rect 549884 248296 553183 248298
rect 549884 248240 553122 248296
rect 553178 248240 553183 248296
rect 549884 248238 553183 248240
rect 553117 248235 553183 248238
rect 349521 247754 349587 247757
rect 347852 247752 349587 247754
rect 347852 247696 349526 247752
rect 349582 247696 349587 247752
rect 347852 247694 349587 247696
rect 349521 247691 349587 247694
rect 46841 247482 46907 247485
rect 48086 247482 48146 247656
rect 550633 247618 550699 247621
rect 549884 247616 550699 247618
rect 549884 247560 550638 247616
rect 550694 247560 550699 247616
rect 549884 247558 550699 247560
rect 550633 247555 550699 247558
rect 46841 247480 48146 247482
rect 46841 247424 46846 247480
rect 46902 247424 48146 247480
rect 46841 247422 48146 247424
rect 46841 247419 46907 247422
rect 46606 247284 46612 247348
rect 46676 247346 46682 247348
rect 46676 247286 48146 247346
rect 46676 247284 46682 247286
rect 46054 247012 46060 247076
rect 46124 247074 46130 247076
rect 46657 247074 46723 247077
rect 46124 247072 46723 247074
rect 46124 247016 46662 247072
rect 46718 247016 46723 247072
rect 48086 247044 48146 247286
rect 46124 247014 46723 247016
rect 46124 247012 46130 247014
rect 46657 247011 46723 247014
rect 407205 246938 407271 246941
rect 553117 246938 553183 246941
rect 407205 246936 410044 246938
rect 407205 246880 407210 246936
rect 407266 246880 410044 246936
rect 407205 246878 410044 246880
rect 549884 246936 553183 246938
rect 549884 246880 553122 246936
rect 553178 246880 553183 246936
rect 549884 246878 553183 246880
rect 407205 246875 407271 246878
rect 553117 246875 553183 246878
rect 46841 245850 46907 245853
rect 48086 245850 48146 246296
rect 347822 245986 347882 246296
rect 407113 246258 407179 246261
rect 552197 246258 552263 246261
rect 407113 246256 410044 246258
rect 407113 246200 407118 246256
rect 407174 246200 410044 246256
rect 407113 246198 410044 246200
rect 549884 246256 552263 246258
rect 549884 246200 552202 246256
rect 552258 246200 552263 246256
rect 549884 246198 552263 246200
rect 407113 246195 407179 246198
rect 552197 246195 552263 246198
rect 350441 245986 350507 245989
rect 347822 245984 350507 245986
rect 347822 245928 350446 245984
rect 350502 245928 350507 245984
rect 347822 245926 350507 245928
rect 350441 245923 350507 245926
rect 46841 245848 48146 245850
rect 46841 245792 46846 245848
rect 46902 245792 48146 245848
rect 46841 245790 48146 245792
rect 46841 245787 46907 245790
rect 349613 245714 349679 245717
rect 347852 245712 349679 245714
rect 347852 245656 349618 245712
rect 349674 245656 349679 245712
rect 347852 245654 349679 245656
rect 349613 245651 349679 245654
rect 408953 245578 409019 245581
rect 408953 245576 410044 245578
rect 408953 245520 408958 245576
rect 409014 245520 410044 245576
rect 408953 245518 410044 245520
rect 408953 245515 409019 245518
rect 583520 245428 584960 245668
rect 347822 244490 347882 244936
rect 407113 244898 407179 244901
rect 553117 244898 553183 244901
rect 407113 244896 410044 244898
rect 407113 244840 407118 244896
rect 407174 244840 410044 244896
rect 407113 244838 410044 244840
rect 549884 244896 553183 244898
rect 549884 244840 553122 244896
rect 553178 244840 553183 244896
rect 549884 244838 553183 244840
rect 407113 244835 407179 244838
rect 553117 244835 553183 244838
rect 350533 244490 350599 244493
rect 347822 244488 350599 244490
rect 347822 244432 350538 244488
rect 350594 244432 350599 244488
rect 347822 244430 350599 244432
rect 350533 244427 350599 244430
rect 46565 244356 46631 244357
rect 46565 244354 46612 244356
rect 46520 244352 46612 244354
rect 46520 244296 46570 244352
rect 46520 244294 46612 244296
rect 46565 244292 46612 244294
rect 46676 244292 46682 244356
rect 46790 244292 46796 244356
rect 46860 244354 46866 244356
rect 350441 244354 350507 244357
rect 46860 244294 48116 244354
rect 347852 244352 350507 244354
rect 347852 244296 350446 244352
rect 350502 244296 350507 244352
rect 347852 244294 350507 244296
rect 46860 244292 46866 244294
rect 46565 244291 46631 244292
rect 350441 244291 350507 244294
rect 347822 243266 347882 243576
rect 350441 243266 350507 243269
rect 347822 243264 350507 243266
rect 347822 243208 350446 243264
rect 350502 243208 350507 243264
rect 347822 243206 350507 243208
rect 350441 243203 350507 243206
rect 44817 242994 44883 242997
rect 349981 242994 350047 242997
rect 44817 242992 48116 242994
rect 44817 242936 44822 242992
rect 44878 242936 48116 242992
rect 44817 242934 48116 242936
rect 347852 242992 350047 242994
rect 347852 242936 349986 242992
rect 350042 242936 350047 242992
rect 347852 242934 350047 242936
rect 44817 242931 44883 242934
rect 349981 242931 350047 242934
rect 407573 242994 407639 242997
rect 410014 242994 410074 243440
rect 549884 243410 550466 243470
rect 550406 243402 550466 243410
rect 552197 243402 552263 243405
rect 550406 243400 552263 243402
rect 550406 243344 552202 243400
rect 552258 243344 552263 243400
rect 550406 243342 552263 243344
rect 552197 243339 552263 243342
rect 407573 242992 410074 242994
rect 407573 242936 407578 242992
rect 407634 242936 410074 242992
rect 407573 242934 410074 242936
rect 407573 242931 407639 242934
rect 409822 242796 409828 242860
rect 409892 242858 409898 242860
rect 552013 242858 552079 242861
rect 409892 242798 410044 242858
rect 549884 242856 552079 242858
rect 549884 242800 552018 242856
rect 552074 242800 552079 242856
rect 549884 242798 552079 242800
rect 409892 242796 409898 242798
rect 552013 242795 552079 242798
rect 406101 242450 406167 242453
rect 410006 242450 410012 242452
rect 406101 242448 410012 242450
rect 406101 242392 406106 242448
rect 406162 242392 410012 242448
rect 406101 242390 410012 242392
rect 406101 242387 406167 242390
rect 410006 242388 410012 242390
rect 410076 242388 410082 242452
rect 393129 242314 393195 242317
rect 410006 242314 410012 242316
rect 393129 242312 410012 242314
rect 393129 242256 393134 242312
rect 393190 242256 410012 242312
rect 393129 242254 410012 242256
rect 393129 242251 393195 242254
rect 410006 242252 410012 242254
rect 410076 242252 410082 242316
rect 407113 242178 407179 242181
rect 407113 242176 410044 242178
rect 407113 242120 407118 242176
rect 407174 242120 410044 242176
rect 407113 242118 410044 242120
rect 407113 242115 407179 242118
rect 44398 241436 44404 241500
rect 44468 241498 44474 241500
rect 44725 241498 44791 241501
rect 44468 241496 44791 241498
rect 44468 241440 44730 241496
rect 44786 241440 44791 241496
rect 44468 241438 44791 241440
rect 44468 241436 44474 241438
rect 44725 241435 44791 241438
rect 409505 241226 409571 241229
rect 410014 241226 410074 241468
rect 409505 241224 410074 241226
rect -960 241090 480 241180
rect 409505 241168 409510 241224
rect 409566 241168 410074 241224
rect 409505 241166 410074 241168
rect 409505 241163 409571 241166
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 45134 240892 45140 240956
rect 45204 240954 45210 240956
rect 45204 240894 48116 240954
rect 45204 240892 45210 240894
rect 409505 240818 409571 240821
rect 550265 240818 550331 240821
rect 409505 240816 410044 240818
rect 409505 240760 409510 240816
rect 409566 240760 410044 240816
rect 409505 240758 410044 240760
rect 549884 240816 550331 240818
rect 549884 240760 550270 240816
rect 550326 240760 550331 240816
rect 549884 240758 550331 240760
rect 409505 240755 409571 240758
rect 550265 240755 550331 240758
rect 376201 240546 376267 240549
rect 564985 240546 565051 240549
rect 376201 240544 565051 240546
rect 376201 240488 376206 240544
rect 376262 240488 564990 240544
rect 565046 240488 565051 240544
rect 376201 240486 565051 240488
rect 376201 240483 376267 240486
rect 564985 240483 565051 240486
rect 409454 240348 409460 240412
rect 409524 240410 409530 240412
rect 410333 240410 410399 240413
rect 409524 240408 410399 240410
rect 409524 240352 410338 240408
rect 410394 240352 410399 240408
rect 409524 240350 410399 240352
rect 409524 240348 409530 240350
rect 410333 240347 410399 240350
rect 363873 240138 363939 240141
rect 572069 240138 572135 240141
rect 363873 240136 572135 240138
rect 363873 240080 363878 240136
rect 363934 240080 572074 240136
rect 572130 240080 572135 240136
rect 363873 240078 572135 240080
rect 363873 240075 363939 240078
rect 572069 240075 572135 240078
rect 375281 240002 375347 240005
rect 578785 240002 578851 240005
rect 375281 240000 578851 240002
rect 375281 239944 375286 240000
rect 375342 239944 578790 240000
rect 578846 239944 578851 240000
rect 375281 239942 578851 239944
rect 375281 239939 375347 239942
rect 578785 239939 578851 239942
rect 386454 239804 386460 239868
rect 386524 239866 386530 239868
rect 387701 239866 387767 239869
rect 386524 239864 387767 239866
rect 386524 239808 387706 239864
rect 387762 239808 387767 239864
rect 386524 239806 387767 239808
rect 386524 239804 386530 239806
rect 387701 239803 387767 239806
rect 408401 239866 408467 239869
rect 560385 239866 560451 239869
rect 408401 239864 560451 239866
rect 408401 239808 408406 239864
rect 408462 239808 560390 239864
rect 560446 239808 560451 239864
rect 408401 239806 560451 239808
rect 408401 239803 408467 239806
rect 560385 239803 560451 239806
rect 548374 239668 548380 239732
rect 548444 239730 548450 239732
rect 565813 239730 565879 239733
rect 548444 239728 565879 239730
rect 548444 239672 565818 239728
rect 565874 239672 565879 239728
rect 548444 239670 565879 239672
rect 548444 239668 548450 239670
rect 565813 239667 565879 239670
rect 547086 239532 547092 239596
rect 547156 239594 547162 239596
rect 565077 239594 565143 239597
rect 547156 239592 565143 239594
rect 547156 239536 565082 239592
rect 565138 239536 565143 239592
rect 547156 239534 565143 239536
rect 547156 239532 547162 239534
rect 565077 239531 565143 239534
rect 347822 239322 347882 239496
rect 537477 239458 537543 239461
rect 571609 239458 571675 239461
rect 537477 239456 571675 239458
rect 537477 239400 537482 239456
rect 537538 239400 571614 239456
rect 571670 239400 571675 239456
rect 537477 239398 571675 239400
rect 537477 239395 537543 239398
rect 571609 239395 571675 239398
rect 350441 239322 350507 239325
rect 347822 239320 350507 239322
rect 347822 239264 350446 239320
rect 350502 239264 350507 239320
rect 347822 239262 350507 239264
rect 350441 239259 350507 239262
rect 544469 239322 544535 239325
rect 561765 239322 561831 239325
rect 544469 239320 561831 239322
rect 544469 239264 544474 239320
rect 544530 239264 561770 239320
rect 561826 239264 561831 239320
rect 544469 239262 561831 239264
rect 544469 239259 544535 239262
rect 561765 239259 561831 239262
rect 350441 238914 350507 238917
rect 347852 238912 350507 238914
rect 347852 238856 350446 238912
rect 350502 238856 350507 238912
rect 347852 238854 350507 238856
rect 350441 238851 350507 238854
rect 399477 238778 399543 238781
rect 509233 238778 509299 238781
rect 399477 238776 509299 238778
rect 399477 238720 399482 238776
rect 399538 238720 509238 238776
rect 509294 238720 509299 238776
rect 399477 238718 509299 238720
rect 399477 238715 399543 238718
rect 509233 238715 509299 238718
rect 387241 238642 387307 238645
rect 548149 238642 548215 238645
rect 387241 238640 548215 238642
rect 387241 238584 387246 238640
rect 387302 238584 548154 238640
rect 548210 238584 548215 238640
rect 387241 238582 548215 238584
rect 387241 238579 387307 238582
rect 548149 238579 548215 238582
rect 551093 238642 551159 238645
rect 551502 238642 551508 238644
rect 551093 238640 551508 238642
rect 551093 238584 551098 238640
rect 551154 238584 551508 238640
rect 551093 238582 551508 238584
rect 551093 238579 551159 238582
rect 551502 238580 551508 238582
rect 551572 238580 551578 238644
rect 399702 238444 399708 238508
rect 399772 238506 399778 238508
rect 458173 238506 458239 238509
rect 399772 238504 458239 238506
rect 399772 238448 458178 238504
rect 458234 238448 458239 238504
rect 399772 238446 458239 238448
rect 399772 238444 399778 238446
rect 458173 238443 458239 238446
rect 525609 238506 525675 238509
rect 546217 238506 546283 238509
rect 525609 238504 546283 238506
rect 525609 238448 525614 238504
rect 525670 238448 546222 238504
rect 546278 238448 546283 238504
rect 525609 238446 546283 238448
rect 525609 238443 525675 238446
rect 546217 238443 546283 238446
rect 520181 238370 520247 238373
rect 549478 238370 549484 238372
rect 520181 238368 549484 238370
rect 520181 238312 520186 238368
rect 520242 238312 549484 238368
rect 520181 238310 549484 238312
rect 520181 238307 520247 238310
rect 549478 238308 549484 238310
rect 549548 238308 549554 238372
rect 46657 238234 46723 238237
rect 393221 238234 393287 238237
rect 545062 238234 545068 238236
rect 46657 238232 48116 238234
rect 46657 238176 46662 238232
rect 46718 238176 48116 238232
rect 46657 238174 48116 238176
rect 393221 238232 545068 238234
rect 393221 238176 393226 238232
rect 393282 238176 545068 238232
rect 393221 238174 545068 238176
rect 46657 238171 46723 238174
rect 393221 238171 393287 238174
rect 545062 238172 545068 238174
rect 545132 238172 545138 238236
rect 388897 238098 388963 238101
rect 544009 238098 544075 238101
rect 388897 238096 544075 238098
rect 388897 238040 388902 238096
rect 388958 238040 544014 238096
rect 544070 238040 544075 238096
rect 388897 238038 544075 238040
rect 388897 238035 388963 238038
rect 544009 238035 544075 238038
rect 358537 237962 358603 237965
rect 537569 237962 537635 237965
rect 358537 237960 537635 237962
rect 358537 237904 358542 237960
rect 358598 237904 537574 237960
rect 537630 237904 537635 237960
rect 358537 237902 537635 237904
rect 358537 237899 358603 237902
rect 537569 237899 537635 237902
rect 45185 237418 45251 237421
rect 48086 237418 48146 237456
rect 549253 237418 549319 237421
rect 45185 237416 48146 237418
rect 45185 237360 45190 237416
rect 45246 237360 48146 237416
rect 45185 237358 48146 237360
rect 548750 237416 549319 237418
rect 548750 237360 549258 237416
rect 549314 237360 549319 237416
rect 548750 237358 549319 237360
rect 45185 237355 45251 237358
rect 379053 237282 379119 237285
rect 545481 237282 545547 237285
rect 548750 237282 548810 237358
rect 549253 237355 549319 237358
rect 379053 237280 545547 237282
rect 379053 237224 379058 237280
rect 379114 237224 545486 237280
rect 545542 237224 545547 237280
rect 379053 237222 545547 237224
rect 379053 237219 379119 237222
rect 545481 237219 545547 237222
rect 545622 237222 548810 237282
rect 548977 237282 549043 237285
rect 552238 237282 552244 237284
rect 548977 237280 552244 237282
rect 548977 237224 548982 237280
rect 549038 237224 552244 237280
rect 548977 237222 552244 237224
rect 381813 237146 381879 237149
rect 545622 237146 545682 237222
rect 548977 237219 549043 237222
rect 552238 237220 552244 237222
rect 552308 237220 552314 237284
rect 381813 237144 545682 237146
rect 381813 237088 381818 237144
rect 381874 237088 545682 237144
rect 381813 237086 545682 237088
rect 545757 237146 545823 237149
rect 551686 237146 551692 237148
rect 545757 237144 551692 237146
rect 545757 237088 545762 237144
rect 545818 237088 551692 237144
rect 545757 237086 551692 237088
rect 381813 237083 381879 237086
rect 545757 237083 545823 237086
rect 551686 237084 551692 237086
rect 551756 237084 551762 237148
rect 409638 236948 409644 237012
rect 409708 237010 409714 237012
rect 574829 237010 574895 237013
rect 409708 237008 574895 237010
rect 409708 236952 574834 237008
rect 574890 236952 574895 237008
rect 409708 236950 574895 236952
rect 409708 236948 409714 236950
rect 574829 236947 574895 236950
rect 545481 236874 545547 236877
rect 553025 236874 553091 236877
rect 545481 236872 553091 236874
rect 545481 236816 545486 236872
rect 545542 236816 553030 236872
rect 553086 236816 553091 236872
rect 545481 236814 553091 236816
rect 545481 236811 545547 236814
rect 553025 236811 553091 236814
rect 386321 236602 386387 236605
rect 538806 236602 538812 236604
rect 386321 236600 538812 236602
rect 386321 236544 386326 236600
rect 386382 236544 538812 236600
rect 386321 236542 538812 236544
rect 386321 236539 386387 236542
rect 538806 236540 538812 236542
rect 538876 236540 538882 236604
rect 350441 236194 350507 236197
rect 347852 236192 350507 236194
rect 347852 236136 350446 236192
rect 350502 236136 350507 236192
rect 347852 236134 350507 236136
rect 350441 236131 350507 236134
rect 46381 236058 46447 236061
rect 48086 236058 48146 236096
rect 46381 236056 48146 236058
rect 46381 236000 46386 236056
rect 46442 236000 48146 236056
rect 46381 235998 48146 236000
rect 46381 235995 46447 235998
rect 393078 235452 393084 235516
rect 393148 235514 393154 235516
rect 541249 235514 541315 235517
rect 393148 235512 541315 235514
rect 393148 235456 541254 235512
rect 541310 235456 541315 235512
rect 393148 235454 541315 235456
rect 393148 235452 393154 235454
rect 541249 235451 541315 235454
rect 347822 235106 347882 235416
rect 402094 235316 402100 235380
rect 402164 235378 402170 235380
rect 556889 235378 556955 235381
rect 402164 235376 556955 235378
rect 402164 235320 556894 235376
rect 556950 235320 556955 235376
rect 402164 235318 556955 235320
rect 402164 235316 402170 235318
rect 556889 235315 556955 235318
rect 388253 235242 388319 235245
rect 561070 235242 561076 235244
rect 388253 235240 561076 235242
rect 388253 235184 388258 235240
rect 388314 235184 561076 235240
rect 388253 235182 561076 235184
rect 388253 235179 388319 235182
rect 561070 235180 561076 235182
rect 561140 235180 561146 235244
rect 350441 235106 350507 235109
rect 347822 235104 350507 235106
rect 347822 235048 350446 235104
rect 350502 235048 350507 235104
rect 347822 235046 350507 235048
rect 350441 235043 350507 235046
rect 46657 234698 46723 234701
rect 48086 234698 48146 234736
rect 46657 234696 48146 234698
rect 46657 234640 46662 234696
rect 46718 234640 48146 234696
rect 46657 234638 48146 234640
rect 46657 234635 46723 234638
rect 402789 234290 402855 234293
rect 540237 234290 540303 234293
rect 402789 234288 540303 234290
rect 402789 234232 402794 234288
rect 402850 234232 540242 234288
rect 540298 234232 540303 234288
rect 402789 234230 540303 234232
rect 402789 234227 402855 234230
rect 540237 234227 540303 234230
rect 401358 234092 401364 234156
rect 401428 234154 401434 234156
rect 538990 234154 538996 234156
rect 401428 234094 538996 234154
rect 401428 234092 401434 234094
rect 538990 234092 538996 234094
rect 539060 234092 539066 234156
rect 396625 234018 396691 234021
rect 546953 234018 547019 234021
rect 396625 234016 547019 234018
rect 396625 233960 396630 234016
rect 396686 233960 546958 234016
rect 547014 233960 547019 234016
rect 396625 233958 547019 233960
rect 396625 233955 396691 233958
rect 546953 233955 547019 233958
rect 397177 233882 397243 233885
rect 573081 233882 573147 233885
rect 397177 233880 573147 233882
rect 397177 233824 397182 233880
rect 397238 233824 573086 233880
rect 573142 233824 573147 233880
rect 397177 233822 573147 233824
rect 397177 233819 397243 233822
rect 573081 233819 573147 233822
rect 45921 233474 45987 233477
rect 45921 233472 48116 233474
rect 45921 233416 45926 233472
rect 45982 233416 48116 233472
rect 45921 233414 48116 233416
rect 45921 233411 45987 233414
rect 390461 232930 390527 232933
rect 545246 232930 545252 232932
rect 390461 232928 545252 232930
rect 390461 232872 390466 232928
rect 390522 232872 545252 232928
rect 390461 232870 545252 232872
rect 390461 232867 390527 232870
rect 545246 232868 545252 232870
rect 545316 232868 545322 232932
rect 387558 232732 387564 232796
rect 387628 232794 387634 232796
rect 550817 232794 550883 232797
rect 387628 232792 550883 232794
rect 387628 232736 550822 232792
rect 550878 232736 550883 232792
rect 387628 232734 550883 232736
rect 387628 232732 387634 232734
rect 550817 232731 550883 232734
rect 45553 232250 45619 232253
rect 48086 232250 48146 232696
rect 45553 232248 48146 232250
rect 45553 232192 45558 232248
rect 45614 232192 48146 232248
rect 45553 232190 48146 232192
rect 347822 232250 347882 232696
rect 384941 232658 385007 232661
rect 562174 232658 562180 232660
rect 384941 232656 562180 232658
rect 384941 232600 384946 232656
rect 385002 232600 562180 232656
rect 384941 232598 562180 232600
rect 384941 232595 385007 232598
rect 562174 232596 562180 232598
rect 562244 232596 562250 232660
rect 357014 232460 357020 232524
rect 357084 232522 357090 232524
rect 553209 232522 553275 232525
rect 357084 232520 553275 232522
rect 357084 232464 553214 232520
rect 553270 232464 553275 232520
rect 357084 232462 553275 232464
rect 357084 232460 357090 232462
rect 553209 232459 553275 232462
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 350441 232250 350507 232253
rect 347822 232248 350507 232250
rect 347822 232192 350446 232248
rect 350502 232192 350507 232248
rect 583520 232236 584960 232326
rect 347822 232190 350507 232192
rect 45553 232187 45619 232190
rect 350441 232187 350507 232190
rect 46013 230890 46079 230893
rect 48086 230890 48146 231336
rect 46013 230888 48146 230890
rect 46013 230832 46018 230888
rect 46074 230832 48146 230888
rect 46013 230830 48146 230832
rect 46013 230827 46079 230830
rect 45553 230618 45619 230621
rect 48086 230618 48146 230656
rect 45553 230616 48146 230618
rect 45553 230560 45558 230616
rect 45614 230560 48146 230616
rect 45553 230558 48146 230560
rect 347822 230618 347882 230656
rect 350441 230618 350507 230621
rect 347822 230616 350507 230618
rect 347822 230560 350446 230616
rect 350502 230560 350507 230616
rect 347822 230558 350507 230560
rect 45553 230555 45619 230558
rect 350441 230555 350507 230558
rect 410241 230346 410307 230349
rect 539174 230346 539180 230348
rect 410241 230344 539180 230346
rect 410241 230288 410246 230344
rect 410302 230288 539180 230344
rect 410241 230286 539180 230288
rect 410241 230283 410307 230286
rect 539174 230284 539180 230286
rect 539244 230284 539250 230348
rect 386137 230210 386203 230213
rect 546033 230210 546099 230213
rect 386137 230208 546099 230210
rect 386137 230152 386142 230208
rect 386198 230152 546038 230208
rect 546094 230152 546099 230208
rect 386137 230150 546099 230152
rect 386137 230147 386203 230150
rect 546033 230147 546099 230150
rect 385953 230074 386019 230077
rect 549437 230074 549503 230077
rect 385953 230072 549503 230074
rect 385953 230016 385958 230072
rect 386014 230016 549442 230072
rect 549498 230016 549503 230072
rect 385953 230014 549503 230016
rect 385953 230011 386019 230014
rect 549437 230011 549503 230014
rect 383101 229938 383167 229941
rect 547965 229938 548031 229941
rect 383101 229936 548031 229938
rect 383101 229880 383106 229936
rect 383162 229880 547970 229936
rect 548026 229880 548031 229936
rect 383101 229878 548031 229880
rect 383101 229875 383167 229878
rect 547965 229875 548031 229878
rect 47577 229802 47643 229805
rect 47894 229802 47900 229804
rect 47577 229800 47900 229802
rect 47577 229744 47582 229800
rect 47638 229744 47900 229800
rect 47577 229742 47900 229744
rect 47577 229739 47643 229742
rect 47894 229740 47900 229742
rect 47964 229740 47970 229804
rect 391790 229740 391796 229804
rect 391860 229802 391866 229804
rect 581545 229802 581611 229805
rect 391860 229800 581611 229802
rect 391860 229744 581550 229800
rect 581606 229744 581611 229800
rect 391860 229742 581611 229744
rect 391860 229740 391866 229742
rect 581545 229739 581611 229742
rect 47158 229332 47164 229396
rect 47228 229394 47234 229396
rect 47228 229334 48116 229394
rect 47228 229332 47234 229334
rect 347822 229258 347882 229296
rect 350441 229258 350507 229261
rect 347822 229256 350507 229258
rect 347822 229200 350446 229256
rect 350502 229200 350507 229256
rect 347822 229198 350507 229200
rect 350441 229195 350507 229198
rect -960 227884 480 228124
rect 45553 227898 45619 227901
rect 48086 227898 48146 227936
rect 45553 227896 48146 227898
rect 45553 227840 45558 227896
rect 45614 227840 48146 227896
rect 45553 227838 48146 227840
rect 45553 227835 45619 227838
rect 46289 226674 46355 226677
rect 46289 226672 48116 226674
rect 46289 226616 46294 226672
rect 46350 226616 48116 226672
rect 46289 226614 48116 226616
rect 46289 226611 46355 226614
rect 347822 225042 347882 225216
rect 349521 225042 349587 225045
rect 347822 225040 349587 225042
rect 347822 224984 349526 225040
rect 349582 224984 349587 225040
rect 347822 224982 349587 224984
rect 349521 224979 349587 224982
rect 44766 224844 44772 224908
rect 44836 224906 44842 224908
rect 46381 224906 46447 224909
rect 44836 224904 46447 224906
rect 44836 224848 46386 224904
rect 46442 224848 46447 224904
rect 44836 224846 46447 224848
rect 44836 224844 44842 224846
rect 46381 224843 46447 224846
rect 35065 224226 35131 224229
rect 44582 224226 44588 224228
rect 35065 224224 44588 224226
rect 35065 224168 35070 224224
rect 35126 224168 44588 224224
rect 35065 224166 44588 224168
rect 35065 224163 35131 224166
rect 44582 224164 44588 224166
rect 44652 224164 44658 224228
rect 46657 224090 46723 224093
rect 48086 224090 48146 224536
rect 46657 224088 48146 224090
rect 46657 224032 46662 224088
rect 46718 224032 48146 224088
rect 46657 224030 48146 224032
rect 46657 224027 46723 224030
rect 350441 222594 350507 222597
rect 347852 222592 350507 222594
rect 347852 222536 350446 222592
rect 350502 222536 350507 222592
rect 347852 222534 350507 222536
rect 350441 222531 350507 222534
rect 46657 222458 46723 222461
rect 48086 222458 48146 222496
rect 46657 222456 48146 222458
rect 46657 222400 46662 222456
rect 46718 222400 48146 222456
rect 46657 222398 48146 222400
rect 46657 222395 46723 222398
rect 46565 221370 46631 221373
rect 48086 221370 48146 221816
rect 46565 221368 48146 221370
rect 46565 221312 46570 221368
rect 46626 221312 48146 221368
rect 46565 221310 48146 221312
rect 46565 221307 46631 221310
rect 347822 221234 347882 221816
rect 350441 221234 350507 221237
rect 347822 221232 350507 221234
rect 347822 221176 350446 221232
rect 350502 221176 350507 221232
rect 347822 221174 350507 221176
rect 350441 221171 350507 221174
rect 46657 221098 46723 221101
rect 48086 221098 48146 221136
rect 46657 221096 48146 221098
rect 46657 221040 46662 221096
rect 46718 221040 48146 221096
rect 46657 221038 48146 221040
rect 46657 221035 46723 221038
rect 47158 220764 47164 220828
rect 47228 220826 47234 220828
rect 47393 220826 47459 220829
rect 47228 220824 47459 220826
rect 47228 220768 47398 220824
rect 47454 220768 47459 220824
rect 47228 220766 47459 220768
rect 47228 220764 47234 220766
rect 47393 220763 47459 220766
rect 46974 220492 46980 220556
rect 47044 220554 47050 220556
rect 47044 220494 48116 220554
rect 47044 220492 47050 220494
rect 347822 220010 347882 220456
rect 349981 220010 350047 220013
rect 347822 220008 350047 220010
rect 347822 219952 349986 220008
rect 350042 219952 350047 220008
rect 347822 219950 350047 219952
rect 349981 219947 350047 219950
rect 46105 218650 46171 218653
rect 48086 218650 48146 219096
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 46105 218648 48146 218650
rect 46105 218592 46110 218648
rect 46166 218592 48146 218648
rect 46105 218590 48146 218592
rect 46105 218587 46171 218590
rect 46657 218378 46723 218381
rect 48086 218378 48146 218416
rect 46657 218376 48146 218378
rect 46657 218320 46662 218376
rect 46718 218320 48146 218376
rect 46657 218318 48146 218320
rect 46657 218315 46723 218318
rect 347822 218106 347882 218416
rect 350441 218106 350507 218109
rect 347822 218104 350507 218106
rect 347822 218048 350446 218104
rect 350502 218048 350507 218104
rect 347822 218046 350507 218048
rect 350441 218043 350507 218046
rect 46289 217290 46355 217293
rect 48086 217290 48146 217736
rect 347822 217562 347882 217736
rect 350441 217562 350507 217565
rect 347822 217560 350507 217562
rect 347822 217504 350446 217560
rect 350502 217504 350507 217560
rect 347822 217502 350507 217504
rect 350441 217499 350507 217502
rect 46289 217288 48146 217290
rect 46289 217232 46294 217288
rect 46350 217232 48146 217288
rect 46289 217230 48146 217232
rect 46289 217227 46355 217230
rect 350349 217154 350415 217157
rect 347852 217152 350415 217154
rect 347852 217096 350354 217152
rect 350410 217096 350415 217152
rect 347852 217094 350415 217096
rect 350349 217091 350415 217094
rect 46657 216746 46723 216749
rect 48086 216746 48146 217056
rect 46657 216744 48146 216746
rect 46657 216688 46662 216744
rect 46718 216688 48146 216744
rect 46657 216686 48146 216688
rect 46657 216683 46723 216686
rect 46657 215386 46723 215389
rect 48086 215386 48146 215696
rect 46657 215384 48146 215386
rect 46657 215328 46662 215384
rect 46718 215328 48146 215384
rect 46657 215326 48146 215328
rect 347822 215386 347882 215696
rect 350441 215386 350507 215389
rect 347822 215384 350507 215386
rect 347822 215328 350446 215384
rect 350502 215328 350507 215384
rect 347822 215326 350507 215328
rect 46657 215323 46723 215326
rect 350441 215323 350507 215326
rect -960 214828 480 215068
rect 348550 214508 348556 214572
rect 348620 214570 348626 214572
rect 352649 214570 352715 214573
rect 348620 214568 352715 214570
rect 348620 214512 352654 214568
rect 352710 214512 352715 214568
rect 348620 214510 352715 214512
rect 348620 214508 348626 214510
rect 352649 214507 352715 214510
rect 45461 214026 45527 214029
rect 48086 214026 48146 214336
rect 45461 214024 48146 214026
rect 45461 213968 45466 214024
rect 45522 213968 48146 214024
rect 45461 213966 48146 213968
rect 45461 213963 45527 213966
rect 347822 213210 347882 213656
rect 350441 213210 350507 213213
rect 347822 213208 350507 213210
rect 347822 213152 350446 213208
rect 350502 213152 350507 213208
rect 347822 213150 350507 213152
rect 350441 213147 350507 213150
rect 44582 212604 44588 212668
rect 44652 212666 44658 212668
rect 45829 212666 45895 212669
rect 44652 212664 45895 212666
rect 44652 212608 45834 212664
rect 45890 212608 45895 212664
rect 44652 212606 45895 212608
rect 44652 212604 44658 212606
rect 45829 212603 45895 212606
rect 34973 211850 35039 211853
rect 44766 211850 44772 211852
rect 34973 211848 44772 211850
rect 34973 211792 34978 211848
rect 35034 211792 44772 211848
rect 34973 211790 44772 211792
rect 34973 211787 35039 211790
rect 44766 211788 44772 211790
rect 44836 211788 44842 211852
rect 45553 211306 45619 211309
rect 48086 211306 48146 211616
rect 45553 211304 48146 211306
rect 45553 211248 45558 211304
rect 45614 211248 48146 211304
rect 45553 211246 48146 211248
rect 45553 211243 45619 211246
rect 44582 210428 44588 210492
rect 44652 210490 44658 210492
rect 46933 210490 46999 210493
rect 44652 210488 46999 210490
rect 44652 210432 46938 210488
rect 46994 210432 46999 210488
rect 44652 210430 46999 210432
rect 44652 210428 44658 210430
rect 46933 210427 46999 210430
rect 45318 210292 45324 210356
rect 45388 210354 45394 210356
rect 45388 210294 48116 210354
rect 45388 210292 45394 210294
rect 347822 209946 347882 210256
rect 350441 209946 350507 209949
rect 347822 209944 350507 209946
rect 347822 209888 350446 209944
rect 350502 209888 350507 209944
rect 347822 209886 350507 209888
rect 350441 209883 350507 209886
rect 47117 209674 47183 209677
rect 48078 209674 48084 209676
rect 47117 209672 48084 209674
rect 47117 209616 47122 209672
rect 47178 209616 48084 209672
rect 47117 209614 48084 209616
rect 47117 209611 47183 209614
rect 48078 209612 48084 209614
rect 48148 209612 48154 209676
rect 42057 209538 42123 209541
rect 47158 209538 47164 209540
rect 42057 209536 47164 209538
rect 42057 209480 42062 209536
rect 42118 209480 47164 209536
rect 42057 209478 47164 209480
rect 42057 209475 42123 209478
rect 47158 209476 47164 209478
rect 47228 209476 47234 209540
rect 347822 209130 347882 209576
rect 350441 209130 350507 209133
rect 347822 209128 350507 209130
rect 347822 209072 350446 209128
rect 350502 209072 350507 209128
rect 347822 209070 350507 209072
rect 350441 209067 350507 209070
rect 347822 207770 347882 208216
rect 350441 207770 350507 207773
rect 347822 207768 350507 207770
rect 347822 207712 350446 207768
rect 350502 207712 350507 207768
rect 347822 207710 350507 207712
rect 350441 207707 350507 207710
rect 45553 207634 45619 207637
rect 45553 207632 48116 207634
rect 45553 207576 45558 207632
rect 45614 207576 48116 207632
rect 45553 207574 48116 207576
rect 45553 207571 45619 207574
rect 347822 207362 347882 207536
rect 350349 207362 350415 207365
rect 347822 207360 350415 207362
rect 347822 207304 350354 207360
rect 350410 207304 350415 207360
rect 347822 207302 350415 207304
rect 350349 207299 350415 207302
rect 45645 206954 45711 206957
rect 350441 206954 350507 206957
rect 45645 206952 48116 206954
rect 45645 206896 45650 206952
rect 45706 206896 48116 206952
rect 45645 206894 48116 206896
rect 347852 206952 350507 206954
rect 347852 206896 350446 206952
rect 350502 206896 350507 206952
rect 347852 206894 350507 206896
rect 45645 206891 45711 206894
rect 350441 206891 350507 206894
rect 406142 206212 406148 206276
rect 406212 206274 406218 206276
rect 523033 206274 523099 206277
rect 406212 206272 523099 206274
rect 406212 206216 523038 206272
rect 523094 206216 523099 206272
rect 406212 206214 523099 206216
rect 406212 206212 406218 206214
rect 523033 206211 523099 206214
rect 45645 206002 45711 206005
rect 48086 206002 48146 206176
rect 45645 206000 48146 206002
rect 45645 205944 45650 206000
rect 45706 205944 48146 206000
rect 45645 205942 48146 205944
rect 45645 205939 45711 205942
rect 583520 205580 584960 205820
rect 347822 205050 347882 205496
rect 350349 205050 350415 205053
rect 347822 205048 350415 205050
rect 347822 204992 350354 205048
rect 350410 204992 350415 205048
rect 347822 204990 350415 204992
rect 350349 204987 350415 204990
rect 356697 204914 356763 204917
rect 542670 204914 542676 204916
rect 356697 204912 542676 204914
rect 356697 204856 356702 204912
rect 356758 204856 542676 204912
rect 356697 204854 542676 204856
rect 356697 204851 356763 204854
rect 542670 204852 542676 204854
rect 542740 204852 542746 204916
rect 350441 204234 350507 204237
rect 347852 204232 350507 204234
rect 347852 204176 350446 204232
rect 350502 204176 350507 204232
rect 347852 204174 350507 204176
rect 350441 204171 350507 204174
rect 46657 203690 46723 203693
rect 48086 203690 48146 204136
rect 46657 203688 48146 203690
rect 46657 203632 46662 203688
rect 46718 203632 48146 203688
rect 46657 203630 48146 203632
rect 46657 203627 46723 203630
rect 347822 203282 347882 203456
rect 350441 203282 350507 203285
rect 347822 203280 350507 203282
rect 347822 203224 350446 203280
rect 350502 203224 350507 203280
rect 347822 203222 350507 203224
rect 350441 203219 350507 203222
rect 46381 202874 46447 202877
rect 46381 202872 48116 202874
rect 46381 202816 46386 202872
rect 46442 202816 48116 202872
rect 46381 202814 48116 202816
rect 46381 202811 46447 202814
rect 347822 202330 347882 202776
rect 349337 202330 349403 202333
rect 347822 202328 349403 202330
rect 347822 202272 349342 202328
rect 349398 202272 349403 202328
rect 347822 202270 349403 202272
rect 349337 202267 349403 202270
rect -960 201922 480 202012
rect 2957 201922 3023 201925
rect -960 201920 3023 201922
rect -960 201864 2962 201920
rect 3018 201864 3023 201920
rect -960 201862 3023 201864
rect -960 201772 480 201862
rect 2957 201859 3023 201862
rect 46381 201650 46447 201653
rect 48086 201650 48146 202096
rect 347822 201922 347882 202096
rect 350441 201922 350507 201925
rect 347822 201920 350507 201922
rect 347822 201864 350446 201920
rect 350502 201864 350507 201920
rect 347822 201862 350507 201864
rect 350441 201859 350507 201862
rect 46381 201648 48146 201650
rect 46381 201592 46386 201648
rect 46442 201592 48146 201648
rect 46381 201590 48146 201592
rect 46381 201587 46447 201590
rect 37641 201380 37707 201381
rect 37590 201378 37596 201380
rect 37550 201318 37596 201378
rect 37660 201376 37707 201380
rect 37702 201320 37707 201376
rect 37590 201316 37596 201318
rect 37660 201316 37707 201320
rect 347630 201316 347636 201380
rect 347700 201378 347706 201380
rect 352046 201378 352052 201380
rect 347700 201318 352052 201378
rect 347700 201316 347706 201318
rect 352046 201316 352052 201318
rect 352116 201316 352122 201380
rect 37641 201315 37707 201316
rect 47301 201242 47367 201245
rect 47894 201242 47900 201244
rect 47301 201240 47900 201242
rect 47301 201184 47306 201240
rect 47362 201184 47900 201240
rect 47301 201182 47900 201184
rect 47301 201179 47367 201182
rect 47894 201180 47900 201182
rect 47964 201180 47970 201244
rect 37549 201106 37615 201109
rect 37549 201104 45570 201106
rect 37549 201048 37554 201104
rect 37610 201048 45570 201104
rect 37549 201046 45570 201048
rect 37549 201043 37615 201046
rect 45510 200562 45570 201046
rect 47761 200970 47827 200973
rect 48262 200970 48268 200972
rect 47761 200968 48268 200970
rect 47761 200912 47766 200968
rect 47822 200912 48268 200968
rect 47761 200910 48268 200912
rect 47761 200907 47827 200910
rect 48262 200908 48268 200910
rect 48332 200908 48338 200972
rect 347630 200908 347636 200972
rect 347700 200970 347706 200972
rect 552749 200970 552815 200973
rect 347700 200968 552815 200970
rect 347700 200912 552754 200968
rect 552810 200912 552815 200968
rect 347700 200910 552815 200912
rect 347700 200908 347706 200910
rect 552749 200907 552815 200910
rect 48262 200562 48268 200564
rect 45510 200502 48268 200562
rect 48262 200500 48268 200502
rect 48332 200500 48338 200564
rect 347681 200426 347747 200429
rect 351361 200426 351427 200429
rect 347681 200424 351427 200426
rect 347681 200368 347686 200424
rect 347742 200368 351366 200424
rect 351422 200368 351427 200424
rect 347681 200366 351427 200368
rect 347681 200363 347747 200366
rect 351361 200363 351427 200366
rect 347773 200292 347839 200293
rect 347773 200290 347820 200292
rect 347728 200288 347820 200290
rect 347728 200232 347778 200288
rect 347728 200230 347820 200232
rect 347773 200228 347820 200230
rect 347884 200228 347890 200292
rect 347773 200227 347839 200228
rect 46749 200154 46815 200157
rect 48262 200154 48268 200156
rect 46749 200152 48268 200154
rect 46749 200096 46754 200152
rect 46810 200096 48268 200152
rect 46749 200094 48268 200096
rect 46749 200091 46815 200094
rect 48262 200092 48268 200094
rect 48332 200092 48338 200156
rect 37181 199882 37247 199885
rect 356973 199882 357039 199885
rect 37181 199880 357039 199882
rect 37181 199824 37186 199880
rect 37242 199824 356978 199880
rect 357034 199824 357039 199880
rect 37181 199822 357039 199824
rect 37181 199819 37247 199822
rect 356973 199819 357039 199822
rect 36537 199746 36603 199749
rect 347630 199746 347636 199748
rect 36537 199744 347636 199746
rect 36537 199688 36542 199744
rect 36598 199688 347636 199744
rect 36537 199686 347636 199688
rect 36537 199683 36603 199686
rect 347630 199684 347636 199686
rect 347700 199684 347706 199748
rect 257981 199610 258047 199613
rect 356646 199610 356652 199612
rect 257981 199608 356652 199610
rect 257981 199552 257986 199608
rect 258042 199552 356652 199608
rect 257981 199550 356652 199552
rect 257981 199547 258047 199550
rect 356646 199548 356652 199550
rect 356716 199548 356722 199612
rect 296069 199474 296135 199477
rect 359406 199474 359412 199476
rect 296069 199472 359412 199474
rect 296069 199416 296074 199472
rect 296130 199416 359412 199472
rect 296069 199414 359412 199416
rect 296069 199411 296135 199414
rect 359406 199412 359412 199414
rect 359476 199412 359482 199476
rect 346894 199276 346900 199340
rect 346964 199338 346970 199340
rect 347681 199338 347747 199341
rect 346964 199336 347747 199338
rect 346964 199280 347686 199336
rect 347742 199280 347747 199336
rect 346964 199278 347747 199280
rect 346964 199276 346970 199278
rect 347681 199275 347747 199278
rect 34145 199202 34211 199205
rect 257889 199202 257955 199205
rect 34145 199200 257955 199202
rect 34145 199144 34150 199200
rect 34206 199144 257894 199200
rect 257950 199144 257955 199200
rect 34145 199142 257955 199144
rect 34145 199139 34211 199142
rect 257889 199139 257955 199142
rect 347630 199140 347636 199204
rect 347700 199202 347706 199204
rect 347773 199202 347839 199205
rect 347700 199200 347839 199202
rect 347700 199144 347778 199200
rect 347834 199144 347839 199200
rect 347700 199142 347839 199144
rect 347700 199140 347706 199142
rect 347773 199139 347839 199142
rect 47393 199066 47459 199069
rect 295333 199066 295399 199069
rect 47393 199064 295399 199066
rect 47393 199008 47398 199064
rect 47454 199008 295338 199064
rect 295394 199008 295399 199064
rect 47393 199006 295399 199008
rect 47393 199003 47459 199006
rect 295333 199003 295399 199006
rect 84101 198930 84167 198933
rect 369301 198930 369367 198933
rect 84101 198928 369367 198930
rect 84101 198872 84106 198928
rect 84162 198872 369306 198928
rect 369362 198872 369367 198928
rect 84101 198870 369367 198872
rect 84101 198867 84167 198870
rect 369301 198867 369367 198870
rect 33041 198794 33107 198797
rect 153653 198794 153719 198797
rect 33041 198792 153719 198794
rect 33041 198736 33046 198792
rect 33102 198736 153658 198792
rect 153714 198736 153719 198792
rect 33041 198734 153719 198736
rect 33041 198731 33107 198734
rect 153653 198731 153719 198734
rect 247033 198794 247099 198797
rect 560753 198794 560819 198797
rect 247033 198792 560819 198794
rect 247033 198736 247038 198792
rect 247094 198736 560758 198792
rect 560814 198736 560819 198792
rect 247033 198734 560819 198736
rect 247033 198731 247099 198734
rect 560753 198731 560819 198734
rect 34881 198658 34947 198661
rect 53833 198658 53899 198661
rect 34881 198656 53899 198658
rect 34881 198600 34886 198656
rect 34942 198600 53838 198656
rect 53894 198600 53899 198656
rect 34881 198598 53899 198600
rect 34881 198595 34947 198598
rect 53833 198595 53899 198598
rect 58985 198658 59051 198661
rect 560702 198658 560708 198660
rect 58985 198656 560708 198658
rect 58985 198600 58990 198656
rect 59046 198600 560708 198656
rect 58985 198598 560708 198600
rect 58985 198595 59051 198598
rect 560702 198596 560708 198598
rect 560772 198596 560778 198660
rect 28073 198522 28139 198525
rect 422293 198522 422359 198525
rect 28073 198520 422359 198522
rect 28073 198464 28078 198520
rect 28134 198464 422298 198520
rect 422354 198464 422359 198520
rect 28073 198462 422359 198464
rect 28073 198459 28139 198462
rect 422293 198459 422359 198462
rect 29453 198386 29519 198389
rect 412725 198386 412791 198389
rect 29453 198384 412791 198386
rect 29453 198328 29458 198384
rect 29514 198328 412730 198384
rect 412786 198328 412791 198384
rect 29453 198326 412791 198328
rect 29453 198323 29519 198326
rect 412725 198323 412791 198326
rect 49969 198250 50035 198253
rect 403566 198250 403572 198252
rect 49969 198248 403572 198250
rect 49969 198192 49974 198248
rect 50030 198192 403572 198248
rect 49969 198190 403572 198192
rect 49969 198187 50035 198190
rect 403566 198188 403572 198190
rect 403636 198188 403642 198252
rect 46197 198114 46263 198117
rect 93117 198114 93183 198117
rect 46197 198112 93183 198114
rect 46197 198056 46202 198112
rect 46258 198056 93122 198112
rect 93178 198056 93183 198112
rect 46197 198054 93183 198056
rect 46197 198051 46263 198054
rect 93117 198051 93183 198054
rect 94405 198114 94471 198117
rect 364926 198114 364932 198116
rect 94405 198112 364932 198114
rect 94405 198056 94410 198112
rect 94466 198056 364932 198112
rect 94405 198054 364932 198056
rect 94405 198051 94471 198054
rect 364926 198052 364932 198054
rect 364996 198052 365002 198116
rect 122741 197978 122807 197981
rect 368974 197978 368980 197980
rect 122741 197976 368980 197978
rect 122741 197920 122746 197976
rect 122802 197920 368980 197976
rect 122741 197918 368980 197920
rect 122741 197915 122807 197918
rect 368974 197916 368980 197918
rect 369044 197916 369050 197980
rect 38377 197842 38443 197845
rect 82813 197842 82879 197845
rect 38377 197840 82879 197842
rect 38377 197784 38382 197840
rect 38438 197784 82818 197840
rect 82874 197784 82879 197840
rect 38377 197782 82879 197784
rect 38377 197779 38443 197782
rect 82813 197779 82879 197782
rect 53189 197434 53255 197437
rect 54477 197434 54543 197437
rect 53189 197432 54543 197434
rect 53189 197376 53194 197432
rect 53250 197376 54482 197432
rect 54538 197376 54543 197432
rect 53189 197374 54543 197376
rect 53189 197371 53255 197374
rect 54477 197371 54543 197374
rect 561438 197372 561444 197436
rect 561508 197434 561514 197436
rect 564617 197434 564683 197437
rect 561508 197432 564683 197434
rect 561508 197376 564622 197432
rect 564678 197376 564683 197432
rect 561508 197374 564683 197376
rect 561508 197372 561514 197374
rect 564617 197371 564683 197374
rect 83457 197298 83523 197301
rect 560886 197298 560892 197300
rect 83457 197296 560892 197298
rect 83457 197240 83462 197296
rect 83518 197240 560892 197296
rect 83457 197238 560892 197240
rect 83457 197235 83523 197238
rect 560886 197236 560892 197238
rect 560956 197236 560962 197300
rect 60273 197162 60339 197165
rect 400990 197162 400996 197164
rect 60273 197160 400996 197162
rect 60273 197104 60278 197160
rect 60334 197104 400996 197160
rect 60273 197102 400996 197104
rect 60273 197099 60339 197102
rect 400990 197100 400996 197102
rect 401060 197100 401066 197164
rect 31518 196964 31524 197028
rect 31588 197026 31594 197028
rect 342345 197026 342411 197029
rect 31588 197024 342411 197026
rect 31588 196968 342350 197024
rect 342406 196968 342411 197024
rect 31588 196966 342411 196968
rect 31588 196964 31594 196966
rect 342345 196963 342411 196966
rect 227713 196890 227779 196893
rect 348366 196890 348372 196892
rect 227713 196888 348372 196890
rect 227713 196832 227718 196888
rect 227774 196832 348372 196888
rect 227713 196830 348372 196832
rect 227713 196827 227779 196830
rect 348366 196828 348372 196830
rect 348436 196828 348442 196892
rect 59118 196556 59124 196620
rect 59188 196618 59194 196620
rect 407798 196618 407804 196620
rect 59188 196558 407804 196618
rect 59188 196556 59194 196558
rect 407798 196556 407804 196558
rect 407868 196556 407874 196620
rect 158161 195938 158227 195941
rect 347630 195938 347636 195940
rect 158161 195936 347636 195938
rect 158161 195880 158166 195936
rect 158222 195880 347636 195936
rect 158161 195878 347636 195880
rect 158161 195875 158227 195878
rect 347630 195876 347636 195878
rect 347700 195876 347706 195940
rect 38193 195802 38259 195805
rect 228357 195802 228423 195805
rect 38193 195800 228423 195802
rect 38193 195744 38198 195800
rect 38254 195744 228362 195800
rect 228418 195744 228423 195800
rect 38193 195742 228423 195744
rect 38193 195739 38259 195742
rect 228357 195739 228423 195742
rect 41045 195666 41111 195669
rect 87689 195666 87755 195669
rect 41045 195664 87755 195666
rect 41045 195608 41050 195664
rect 41106 195608 87694 195664
rect 87750 195608 87755 195664
rect 41045 195606 87755 195608
rect 41045 195603 41111 195606
rect 87689 195603 87755 195606
rect 200021 195666 200087 195669
rect 363454 195666 363460 195668
rect 200021 195664 363460 195666
rect 200021 195608 200026 195664
rect 200082 195608 363460 195664
rect 200021 195606 363460 195608
rect 200021 195603 200087 195606
rect 363454 195604 363460 195606
rect 363524 195604 363530 195668
rect 39757 195530 39823 195533
rect 48078 195530 48084 195532
rect 39757 195528 48084 195530
rect 39757 195472 39762 195528
rect 39818 195472 48084 195528
rect 39757 195470 48084 195472
rect 39757 195467 39823 195470
rect 48078 195468 48084 195470
rect 48148 195468 48154 195532
rect 58341 195530 58407 195533
rect 349981 195530 350047 195533
rect 58341 195528 350047 195530
rect 58341 195472 58346 195528
rect 58402 195472 349986 195528
rect 350042 195472 350047 195528
rect 58341 195470 350047 195472
rect 58341 195467 58407 195470
rect 349981 195467 350047 195470
rect 43713 195394 43779 195397
rect 412725 195394 412791 195397
rect 43713 195392 412791 195394
rect 43713 195336 43718 195392
rect 43774 195336 412730 195392
rect 412786 195336 412791 195392
rect 43713 195334 412791 195336
rect 43713 195331 43779 195334
rect 412725 195331 412791 195334
rect 46841 195258 46907 195261
rect 452837 195258 452903 195261
rect 46841 195256 452903 195258
rect 46841 195200 46846 195256
rect 46902 195200 452842 195256
rect 452898 195200 452903 195256
rect 46841 195198 452903 195200
rect 46841 195195 46907 195198
rect 452837 195195 452903 195198
rect 2957 194578 3023 194581
rect 387006 194578 387012 194580
rect 2957 194576 387012 194578
rect 2957 194520 2962 194576
rect 3018 194520 387012 194576
rect 2957 194518 387012 194520
rect 2957 194515 3023 194518
rect 387006 194516 387012 194518
rect 387076 194516 387082 194580
rect 57646 193972 57652 194036
rect 57716 194034 57722 194036
rect 563605 194034 563671 194037
rect 57716 194032 563671 194034
rect 57716 193976 563610 194032
rect 563666 193976 563671 194032
rect 57716 193974 563671 193976
rect 57716 193972 57722 193974
rect 563605 193971 563671 193974
rect 53046 193836 53052 193900
rect 53116 193898 53122 193900
rect 566825 193898 566891 193901
rect 53116 193896 566891 193898
rect 53116 193840 566830 193896
rect 566886 193840 566891 193896
rect 53116 193838 566891 193840
rect 53116 193836 53122 193838
rect 566825 193835 566891 193838
rect 31385 193218 31451 193221
rect 531313 193218 531379 193221
rect 31385 193216 531379 193218
rect 31385 193160 31390 193216
rect 31446 193160 531318 193216
rect 531374 193160 531379 193216
rect 31385 193158 531379 193160
rect 31385 193155 31451 193158
rect 531313 193155 531379 193158
rect 49182 192884 49188 192948
rect 49252 192946 49258 192948
rect 139393 192946 139459 192949
rect 49252 192944 139459 192946
rect 49252 192888 139398 192944
rect 139454 192888 139459 192944
rect 49252 192886 139459 192888
rect 49252 192884 49258 192886
rect 139393 192883 139459 192886
rect 53414 192748 53420 192812
rect 53484 192810 53490 192812
rect 373390 192810 373396 192812
rect 53484 192750 373396 192810
rect 53484 192748 53490 192750
rect 373390 192748 373396 192750
rect 373460 192748 373466 192812
rect 44398 192612 44404 192676
rect 44468 192674 44474 192676
rect 453481 192674 453547 192677
rect 44468 192672 453547 192674
rect 44468 192616 453486 192672
rect 453542 192616 453547 192672
rect 44468 192614 453547 192616
rect 44468 192612 44474 192614
rect 453481 192611 453547 192614
rect 2773 192538 2839 192541
rect 551093 192538 551159 192541
rect 2773 192536 551159 192538
rect 2773 192480 2778 192536
rect 2834 192480 551098 192536
rect 551154 192480 551159 192536
rect 2773 192478 551159 192480
rect 2773 192475 2839 192478
rect 551093 192475 551159 192478
rect 580257 192538 580323 192541
rect 583520 192538 584960 192628
rect 580257 192536 584960 192538
rect 580257 192480 580262 192536
rect 580318 192480 584960 192536
rect 580257 192478 584960 192480
rect 580257 192475 580323 192478
rect 583520 192388 584960 192478
rect 54886 190980 54892 191044
rect 54956 191042 54962 191044
rect 366541 191042 366607 191045
rect 54956 191040 366607 191042
rect 54956 190984 366546 191040
rect 366602 190984 366607 191040
rect 54956 190982 366607 190984
rect 54956 190980 54962 190982
rect 366541 190979 366607 190982
rect 85665 190362 85731 190365
rect 377397 190362 377463 190365
rect 85665 190360 377463 190362
rect 85665 190304 85670 190360
rect 85726 190304 377402 190360
rect 377458 190304 377463 190360
rect 85665 190302 377463 190304
rect 85665 190299 85731 190302
rect 377397 190299 377463 190302
rect 270585 190090 270651 190093
rect 562041 190090 562107 190093
rect 270585 190088 562107 190090
rect 270585 190032 270590 190088
rect 270646 190032 562046 190088
rect 562102 190032 562107 190088
rect 270585 190030 562107 190032
rect 270585 190027 270651 190030
rect 562041 190027 562107 190030
rect 56777 189954 56843 189957
rect 350942 189954 350948 189956
rect 56777 189952 350948 189954
rect 56777 189896 56782 189952
rect 56838 189896 350948 189952
rect 56777 189894 350948 189896
rect 56777 189891 56843 189894
rect 350942 189892 350948 189894
rect 351012 189892 351018 189956
rect 54518 189756 54524 189820
rect 54588 189818 54594 189820
rect 395470 189818 395476 189820
rect 54588 189758 395476 189818
rect 54588 189756 54594 189758
rect 395470 189756 395476 189758
rect 395540 189756 395546 189820
rect 157885 189682 157951 189685
rect 563697 189682 563763 189685
rect 157885 189680 563763 189682
rect 157885 189624 157890 189680
rect 157946 189624 563702 189680
rect 563758 189624 563763 189680
rect 157885 189622 563763 189624
rect 157885 189619 157951 189622
rect 563697 189619 563763 189622
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 172053 188866 172119 188869
rect 350574 188866 350580 188868
rect 172053 188864 350580 188866
rect 172053 188808 172058 188864
rect 172114 188808 350580 188864
rect 172053 188806 350580 188808
rect 172053 188803 172119 188806
rect 350574 188804 350580 188806
rect 350644 188804 350650 188868
rect 41822 188668 41828 188732
rect 41892 188730 41898 188732
rect 275737 188730 275803 188733
rect 41892 188728 275803 188730
rect 41892 188672 275742 188728
rect 275798 188672 275803 188728
rect 41892 188670 275803 188672
rect 41892 188668 41898 188670
rect 275737 188667 275803 188670
rect 81249 188594 81315 188597
rect 381670 188594 381676 188596
rect 81249 188592 381676 188594
rect 81249 188536 81254 188592
rect 81310 188536 381676 188592
rect 81249 188534 381676 188536
rect 81249 188531 81315 188534
rect 381670 188532 381676 188534
rect 381740 188532 381746 188596
rect 54702 188396 54708 188460
rect 54772 188458 54778 188460
rect 371918 188458 371924 188460
rect 54772 188398 371924 188458
rect 54772 188396 54778 188398
rect 371918 188396 371924 188398
rect 371988 188396 371994 188460
rect 48773 188322 48839 188325
rect 378726 188322 378732 188324
rect 48773 188320 378732 188322
rect 48773 188264 48778 188320
rect 48834 188264 378732 188320
rect 48773 188262 378732 188264
rect 48773 188259 48839 188262
rect 378726 188260 378732 188262
rect 378796 188260 378802 188324
rect 55070 187308 55076 187372
rect 55140 187370 55146 187372
rect 367686 187370 367692 187372
rect 55140 187310 367692 187370
rect 55140 187308 55146 187310
rect 367686 187308 367692 187310
rect 367756 187308 367762 187372
rect 31753 187234 31819 187237
rect 385718 187234 385724 187236
rect 31753 187232 385724 187234
rect 31753 187176 31758 187232
rect 31814 187176 385724 187232
rect 31753 187174 385724 187176
rect 31753 187171 31819 187174
rect 385718 187172 385724 187174
rect 385788 187172 385794 187236
rect 43662 187036 43668 187100
rect 43732 187098 43738 187100
rect 427077 187098 427143 187101
rect 43732 187096 427143 187098
rect 43732 187040 427082 187096
rect 427138 187040 427143 187096
rect 43732 187038 427143 187040
rect 43732 187036 43738 187038
rect 427077 187035 427143 187038
rect 32397 186962 32463 186965
rect 547505 186962 547571 186965
rect 32397 186960 547571 186962
rect 32397 186904 32402 186960
rect 32458 186904 547510 186960
rect 547566 186904 547571 186960
rect 32397 186902 547571 186904
rect 32397 186899 32463 186902
rect 547505 186899 547571 186902
rect 61326 185812 61332 185876
rect 61396 185874 61402 185876
rect 368565 185874 368631 185877
rect 61396 185872 368631 185874
rect 61396 185816 368570 185872
rect 368626 185816 368631 185872
rect 61396 185814 368631 185816
rect 61396 185812 61402 185814
rect 368565 185811 368631 185814
rect 36670 185676 36676 185740
rect 36740 185738 36746 185740
rect 458173 185738 458239 185741
rect 36740 185736 458239 185738
rect 36740 185680 458178 185736
rect 458234 185680 458239 185736
rect 36740 185678 458239 185680
rect 36740 185676 36746 185678
rect 458173 185675 458239 185678
rect 46238 185540 46244 185604
rect 46308 185602 46314 185604
rect 539542 185602 539548 185604
rect 46308 185542 539548 185602
rect 46308 185540 46314 185542
rect 539542 185540 539548 185542
rect 539612 185540 539618 185604
rect 61510 184860 61516 184924
rect 61580 184922 61586 184924
rect 364701 184922 364767 184925
rect 61580 184920 364767 184922
rect 61580 184864 364706 184920
rect 364762 184864 364767 184920
rect 61580 184862 364767 184864
rect 61580 184860 61586 184862
rect 364701 184859 364767 184862
rect 33685 184786 33751 184789
rect 349470 184786 349476 184788
rect 33685 184784 349476 184786
rect 33685 184728 33690 184784
rect 33746 184728 349476 184784
rect 33685 184726 349476 184728
rect 33685 184723 33751 184726
rect 349470 184724 349476 184726
rect 349540 184724 349546 184788
rect 58566 184588 58572 184652
rect 58636 184650 58642 184652
rect 407614 184650 407620 184652
rect 58636 184590 407620 184650
rect 58636 184588 58642 184590
rect 407614 184588 407620 184590
rect 407684 184588 407690 184652
rect 27613 184514 27679 184517
rect 392526 184514 392532 184516
rect 27613 184512 392532 184514
rect 27613 184456 27618 184512
rect 27674 184456 392532 184512
rect 27613 184454 392532 184456
rect 27613 184451 27679 184454
rect 392526 184452 392532 184454
rect 392596 184452 392602 184516
rect 43478 184316 43484 184380
rect 43548 184378 43554 184380
rect 460565 184378 460631 184381
rect 43548 184376 460631 184378
rect 43548 184320 460570 184376
rect 460626 184320 460631 184376
rect 43548 184318 460631 184320
rect 43548 184316 43554 184318
rect 460565 184315 460631 184318
rect 50838 184180 50844 184244
rect 50908 184242 50914 184244
rect 566549 184242 566615 184245
rect 50908 184240 566615 184242
rect 50908 184184 566554 184240
rect 566610 184184 566615 184240
rect 50908 184182 566615 184184
rect 50908 184180 50914 184182
rect 566549 184179 566615 184182
rect 147673 184106 147739 184109
rect 350758 184106 350764 184108
rect 147673 184104 350764 184106
rect 147673 184048 147678 184104
rect 147734 184048 350764 184104
rect 147673 184046 350764 184048
rect 147673 184043 147739 184046
rect 350758 184044 350764 184046
rect 350828 184044 350834 184108
rect 382273 183698 382339 183701
rect 383510 183698 383516 183700
rect 382273 183696 383516 183698
rect 382273 183640 382278 183696
rect 382334 183640 383516 183696
rect 382273 183638 383516 183640
rect 382273 183635 382339 183638
rect 383510 183636 383516 183638
rect 383580 183636 383586 183700
rect 40309 183290 40375 183293
rect 349286 183290 349292 183292
rect 40309 183288 349292 183290
rect 40309 183232 40314 183288
rect 40370 183232 349292 183288
rect 40309 183230 349292 183232
rect 40309 183227 40375 183230
rect 349286 183228 349292 183230
rect 349356 183228 349362 183292
rect 49550 183092 49556 183156
rect 49620 183154 49626 183156
rect 382774 183154 382780 183156
rect 49620 183094 382780 183154
rect 49620 183092 49626 183094
rect 382774 183092 382780 183094
rect 382844 183092 382850 183156
rect 54293 183018 54359 183021
rect 404854 183018 404860 183020
rect 54293 183016 404860 183018
rect 54293 182960 54298 183016
rect 54354 182960 404860 183016
rect 54293 182958 404860 182960
rect 54293 182955 54359 182958
rect 404854 182956 404860 182958
rect 404924 182956 404930 183020
rect 35566 182820 35572 182884
rect 35636 182882 35642 182884
rect 497273 182882 497339 182885
rect 35636 182880 497339 182882
rect 35636 182824 497278 182880
rect 497334 182824 497339 182880
rect 35636 182822 497339 182824
rect 35636 182820 35642 182822
rect 497273 182819 497339 182822
rect 237741 182066 237807 182069
rect 371734 182066 371740 182068
rect 237741 182064 371740 182066
rect 237741 182008 237746 182064
rect 237802 182008 371740 182064
rect 237741 182006 371740 182008
rect 237741 182003 237807 182006
rect 371734 182004 371740 182006
rect 371804 182004 371810 182068
rect 159173 181930 159239 181933
rect 348550 181930 348556 181932
rect 159173 181928 348556 181930
rect 159173 181872 159178 181928
rect 159234 181872 348556 181928
rect 159173 181870 348556 181872
rect 159173 181867 159239 181870
rect 348550 181868 348556 181870
rect 348620 181868 348626 181932
rect 57830 181732 57836 181796
rect 57900 181794 57906 181796
rect 365110 181794 365116 181796
rect 57900 181734 365116 181794
rect 57900 181732 57906 181734
rect 365110 181732 365116 181734
rect 365180 181732 365186 181796
rect 52310 181596 52316 181660
rect 52380 181658 52386 181660
rect 369485 181658 369551 181661
rect 52380 181656 369551 181658
rect 52380 181600 369490 181656
rect 369546 181600 369551 181656
rect 52380 181598 369551 181600
rect 52380 181596 52386 181598
rect 369485 181595 369551 181598
rect 47710 181460 47716 181524
rect 47780 181522 47786 181524
rect 377029 181522 377095 181525
rect 47780 181520 377095 181522
rect 47780 181464 377034 181520
rect 377090 181464 377095 181520
rect 47780 181462 377095 181464
rect 47780 181460 47786 181462
rect 377029 181459 377095 181462
rect 55857 181386 55923 181389
rect 385534 181386 385540 181388
rect 55857 181384 385540 181386
rect 55857 181328 55862 181384
rect 55918 181328 385540 181384
rect 55857 181326 385540 181328
rect 55857 181323 55923 181326
rect 385534 181324 385540 181326
rect 385604 181324 385610 181388
rect 59854 180508 59860 180572
rect 59924 180570 59930 180572
rect 366081 180570 366147 180573
rect 59924 180568 366147 180570
rect 59924 180512 366086 180568
rect 366142 180512 366147 180568
rect 59924 180510 366147 180512
rect 59924 180508 59930 180510
rect 366081 180507 366147 180510
rect 50654 180372 50660 180436
rect 50724 180434 50730 180436
rect 358118 180434 358124 180436
rect 50724 180374 358124 180434
rect 50724 180372 50730 180374
rect 358118 180372 358124 180374
rect 358188 180372 358194 180436
rect 39798 180236 39804 180300
rect 39868 180298 39874 180300
rect 492765 180298 492831 180301
rect 39868 180296 492831 180298
rect 39868 180240 492770 180296
rect 492826 180240 492831 180296
rect 39868 180238 492831 180240
rect 39868 180236 39874 180238
rect 492765 180235 492831 180238
rect 67633 180162 67699 180165
rect 539726 180162 539732 180164
rect 67633 180160 539732 180162
rect 67633 180104 67638 180160
rect 67694 180104 539732 180160
rect 67633 180102 539732 180104
rect 67633 180099 67699 180102
rect 539726 180100 539732 180102
rect 539796 180100 539802 180164
rect 46238 179964 46244 180028
rect 46308 180026 46314 180028
rect 552054 180026 552060 180028
rect 46308 179966 552060 180026
rect 46308 179964 46314 179966
rect 552054 179964 552060 179966
rect 552124 179964 552130 180028
rect 49325 179210 49391 179213
rect 353518 179210 353524 179212
rect 49325 179208 353524 179210
rect 49325 179152 49330 179208
rect 49386 179152 353524 179208
rect 49325 179150 353524 179152
rect 49325 179147 49391 179150
rect 353518 179148 353524 179150
rect 353588 179148 353594 179212
rect 580073 179210 580139 179213
rect 583520 179210 584960 179300
rect 580073 179208 584960 179210
rect 580073 179152 580078 179208
rect 580134 179152 584960 179208
rect 580073 179150 584960 179152
rect 580073 179147 580139 179150
rect 49366 179012 49372 179076
rect 49436 179074 49442 179076
rect 386454 179074 386460 179076
rect 49436 179014 386460 179074
rect 49436 179012 49442 179014
rect 386454 179012 386460 179014
rect 386524 179012 386530 179076
rect 583520 179060 584960 179150
rect 39665 178938 39731 178941
rect 388478 178938 388484 178940
rect 39665 178936 388484 178938
rect 39665 178880 39670 178936
rect 39726 178880 388484 178936
rect 39665 178878 388484 178880
rect 39665 178875 39731 178878
rect 388478 178876 388484 178878
rect 388548 178876 388554 178940
rect 51625 178802 51691 178805
rect 403750 178802 403756 178804
rect 51625 178800 403756 178802
rect 51625 178744 51630 178800
rect 51686 178744 403756 178800
rect 51625 178742 403756 178744
rect 51625 178739 51691 178742
rect 403750 178740 403756 178742
rect 403820 178740 403826 178804
rect 39246 178604 39252 178668
rect 39316 178666 39322 178668
rect 394141 178666 394207 178669
rect 39316 178664 394207 178666
rect 39316 178608 394146 178664
rect 394202 178608 394207 178664
rect 39316 178606 394207 178608
rect 39316 178604 39322 178606
rect 394141 178603 394207 178606
rect 60406 177652 60412 177716
rect 60476 177714 60482 177716
rect 386413 177714 386479 177717
rect 60476 177712 386479 177714
rect 60476 177656 386418 177712
rect 386474 177656 386479 177712
rect 60476 177654 386479 177656
rect 60476 177652 60482 177654
rect 386413 177651 386479 177654
rect 52126 177516 52132 177580
rect 52196 177578 52202 177580
rect 391054 177578 391060 177580
rect 52196 177518 391060 177578
rect 52196 177516 52202 177518
rect 391054 177516 391060 177518
rect 391124 177516 391130 177580
rect 44950 177380 44956 177444
rect 45020 177442 45026 177444
rect 396165 177442 396231 177445
rect 45020 177440 396231 177442
rect 45020 177384 396170 177440
rect 396226 177384 396231 177440
rect 45020 177382 396231 177384
rect 45020 177380 45026 177382
rect 396165 177379 396231 177382
rect 45134 177244 45140 177308
rect 45204 177306 45210 177308
rect 577221 177306 577287 177309
rect 45204 177304 577287 177306
rect 45204 177248 577226 177304
rect 577282 177248 577287 177304
rect 45204 177246 577287 177248
rect 45204 177244 45210 177246
rect 577221 177243 577287 177246
rect 50889 176626 50955 176629
rect 353702 176626 353708 176628
rect 50889 176624 353708 176626
rect 50889 176568 50894 176624
rect 50950 176568 353708 176624
rect 50889 176566 353708 176568
rect 50889 176563 50955 176566
rect 353702 176564 353708 176566
rect 353772 176564 353778 176628
rect 48078 176428 48084 176492
rect 48148 176490 48154 176492
rect 367134 176490 367140 176492
rect 48148 176430 367140 176490
rect 48148 176428 48154 176430
rect 367134 176428 367140 176430
rect 367204 176428 367210 176492
rect 53230 176292 53236 176356
rect 53300 176354 53306 176356
rect 380157 176354 380223 176357
rect 53300 176352 380223 176354
rect 53300 176296 380162 176352
rect 380218 176296 380223 176352
rect 53300 176294 380223 176296
rect 53300 176292 53306 176294
rect 380157 176291 380223 176294
rect 39798 176156 39804 176220
rect 39868 176218 39874 176220
rect 373349 176218 373415 176221
rect 39868 176216 373415 176218
rect 39868 176160 373354 176216
rect 373410 176160 373415 176216
rect 39868 176158 373415 176160
rect 39868 176156 39874 176158
rect 373349 176155 373415 176158
rect 38285 176082 38351 176085
rect 391238 176082 391244 176084
rect 38285 176080 391244 176082
rect -960 175796 480 176036
rect 38285 176024 38290 176080
rect 38346 176024 391244 176080
rect 38285 176022 391244 176024
rect 38285 176019 38351 176022
rect 391238 176020 391244 176022
rect 391308 176020 391314 176084
rect 73337 175946 73403 175949
rect 541198 175946 541204 175948
rect 73337 175944 541204 175946
rect 73337 175888 73342 175944
rect 73398 175888 541204 175944
rect 73337 175886 541204 175888
rect 73337 175883 73403 175886
rect 541198 175884 541204 175886
rect 541268 175884 541274 175948
rect 313089 175810 313155 175813
rect 400806 175810 400812 175812
rect 313089 175808 400812 175810
rect 313089 175752 313094 175808
rect 313150 175752 400812 175808
rect 313089 175750 400812 175752
rect 313089 175747 313155 175750
rect 400806 175748 400812 175750
rect 400876 175748 400882 175812
rect 53598 174796 53604 174860
rect 53668 174858 53674 174860
rect 389817 174858 389883 174861
rect 53668 174856 389883 174858
rect 53668 174800 389822 174856
rect 389878 174800 389883 174856
rect 53668 174798 389883 174800
rect 53668 174796 53674 174798
rect 389817 174795 389883 174798
rect 43662 174660 43668 174724
rect 43732 174722 43738 174724
rect 383009 174722 383075 174725
rect 43732 174720 383075 174722
rect 43732 174664 383014 174720
rect 383070 174664 383075 174720
rect 43732 174662 383075 174664
rect 43732 174660 43738 174662
rect 383009 174659 383075 174662
rect 55622 174524 55628 174588
rect 55692 174586 55698 174588
rect 397085 174586 397151 174589
rect 55692 174584 397151 174586
rect 55692 174528 397090 174584
rect 397146 174528 397151 174584
rect 55692 174526 397151 174528
rect 55692 174524 55698 174526
rect 397085 174523 397151 174526
rect 39430 173164 39436 173228
rect 39500 173226 39506 173228
rect 539777 173226 539843 173229
rect 39500 173224 539843 173226
rect 39500 173168 539782 173224
rect 539838 173168 539843 173224
rect 39500 173166 539843 173168
rect 39500 173164 39506 173166
rect 539777 173163 539843 173166
rect 52453 171730 52519 171733
rect 403934 171730 403940 171732
rect 52453 171728 403940 171730
rect 52453 171672 52458 171728
rect 52514 171672 403940 171728
rect 52453 171670 403940 171672
rect 52453 171667 52519 171670
rect 403934 171668 403940 171670
rect 404004 171668 404010 171732
rect 50470 170308 50476 170372
rect 50540 170370 50546 170372
rect 389766 170370 389772 170372
rect 50540 170310 389772 170370
rect 50540 170308 50546 170310
rect 389766 170308 389772 170310
rect 389836 170308 389842 170372
rect 57789 169010 57855 169013
rect 356830 169010 356836 169012
rect 57789 169008 356836 169010
rect 57789 168952 57794 169008
rect 57850 168952 356836 169008
rect 57789 168950 356836 168952
rect 57789 168947 57855 168950
rect 356830 168948 356836 168950
rect 356900 168948 356906 169012
rect 58750 167860 58756 167924
rect 58820 167922 58826 167924
rect 349102 167922 349108 167924
rect 58820 167862 349108 167922
rect 58820 167860 58826 167862
rect 349102 167860 349108 167862
rect 349172 167860 349178 167924
rect 40718 167724 40724 167788
rect 40788 167786 40794 167788
rect 372337 167786 372403 167789
rect 40788 167784 372403 167786
rect 40788 167728 372342 167784
rect 372398 167728 372403 167784
rect 40788 167726 372403 167728
rect 40788 167724 40794 167726
rect 372337 167723 372403 167726
rect 387149 167786 387215 167789
rect 542670 167786 542676 167788
rect 387149 167784 542676 167786
rect 387149 167728 387154 167784
rect 387210 167728 542676 167784
rect 387149 167726 542676 167728
rect 387149 167723 387215 167726
rect 542670 167724 542676 167726
rect 542740 167724 542746 167788
rect 42006 167588 42012 167652
rect 42076 167650 42082 167652
rect 488901 167650 488967 167653
rect 42076 167648 488967 167650
rect 42076 167592 488906 167648
rect 488962 167592 488967 167648
rect 42076 167590 488967 167592
rect 42076 167588 42082 167590
rect 488901 167587 488967 167590
rect 405406 166364 405412 166428
rect 405476 166426 405482 166428
rect 547638 166426 547644 166428
rect 405476 166366 547644 166426
rect 405476 166364 405482 166366
rect 547638 166364 547644 166366
rect 547708 166364 547714 166428
rect 405590 166228 405596 166292
rect 405660 166290 405666 166292
rect 560702 166290 560708 166292
rect 405660 166230 560708 166290
rect 405660 166228 405666 166230
rect 560702 166228 560708 166230
rect 560772 166228 560778 166292
rect 583520 165732 584960 165972
rect 404169 165202 404235 165205
rect 543958 165202 543964 165204
rect 404169 165200 543964 165202
rect 404169 165144 404174 165200
rect 404230 165144 543964 165200
rect 404169 165142 543964 165144
rect 404169 165139 404235 165142
rect 543958 165140 543964 165142
rect 544028 165140 544034 165204
rect 397310 165004 397316 165068
rect 397380 165066 397386 165068
rect 566365 165066 566431 165069
rect 397380 165064 566431 165066
rect 397380 165008 566370 165064
rect 566426 165008 566431 165064
rect 397380 165006 566431 165008
rect 397380 165004 397386 165006
rect 566365 165003 566431 165006
rect 35198 164868 35204 164932
rect 35268 164930 35274 164932
rect 490189 164930 490255 164933
rect 35268 164928 490255 164930
rect 35268 164872 490194 164928
rect 490250 164872 490255 164928
rect 35268 164870 490255 164872
rect 35268 164868 35274 164870
rect 490189 164867 490255 164870
rect 390134 163508 390140 163572
rect 390204 163570 390210 163572
rect 552054 163570 552060 163572
rect 390204 163510 552060 163570
rect 390204 163508 390210 163510
rect 552054 163508 552060 163510
rect 552124 163508 552130 163572
rect 369158 163372 369164 163436
rect 369228 163434 369234 163436
rect 551502 163434 551508 163436
rect 369228 163374 551508 163434
rect 369228 163372 369234 163374
rect 551502 163372 551508 163374
rect 551572 163372 551578 163436
rect -960 162740 480 162980
rect 409638 162420 409644 162484
rect 409708 162482 409714 162484
rect 555233 162482 555299 162485
rect 409708 162480 555299 162482
rect 409708 162424 555238 162480
rect 555294 162424 555299 162480
rect 409708 162422 555299 162424
rect 409708 162420 409714 162422
rect 555233 162419 555299 162422
rect 388621 162346 388687 162349
rect 551645 162346 551711 162349
rect 388621 162344 551711 162346
rect 388621 162288 388626 162344
rect 388682 162288 551650 162344
rect 551706 162288 551711 162344
rect 388621 162286 551711 162288
rect 388621 162283 388687 162286
rect 551645 162283 551711 162286
rect 388437 162210 388503 162213
rect 577221 162210 577287 162213
rect 388437 162208 577287 162210
rect 388437 162152 388442 162208
rect 388498 162152 577226 162208
rect 577282 162152 577287 162208
rect 388437 162150 577287 162152
rect 388437 162147 388503 162150
rect 577221 162147 577287 162150
rect 39614 162012 39620 162076
rect 39684 162074 39690 162076
rect 502425 162074 502491 162077
rect 39684 162072 502491 162074
rect 39684 162016 502430 162072
rect 502486 162016 502491 162072
rect 39684 162014 502491 162016
rect 39684 162012 39690 162014
rect 502425 162011 502491 162014
rect 399518 160924 399524 160988
rect 399588 160986 399594 160988
rect 552606 160986 552612 160988
rect 399588 160926 552612 160986
rect 399588 160924 399594 160926
rect 552606 160924 552612 160926
rect 552676 160924 552682 160988
rect 378910 160788 378916 160852
rect 378980 160850 378986 160852
rect 551185 160850 551251 160853
rect 378980 160848 551251 160850
rect 378980 160792 551190 160848
rect 551246 160792 551251 160848
rect 378980 160790 551251 160792
rect 378980 160788 378986 160790
rect 551185 160787 551251 160790
rect 373206 160652 373212 160716
rect 373276 160714 373282 160716
rect 552238 160714 552244 160716
rect 373276 160654 552244 160714
rect 373276 160652 373282 160654
rect 552238 160652 552244 160654
rect 552308 160652 552314 160716
rect 410006 159700 410012 159764
rect 410076 159762 410082 159764
rect 563462 159762 563468 159764
rect 410076 159702 563468 159762
rect 410076 159700 410082 159702
rect 563462 159700 563468 159702
rect 563532 159700 563538 159764
rect 363597 159626 363663 159629
rect 540094 159626 540100 159628
rect 363597 159624 540100 159626
rect 363597 159568 363602 159624
rect 363658 159568 540100 159624
rect 363597 159566 540100 159568
rect 363597 159563 363663 159566
rect 540094 159564 540100 159566
rect 540164 159564 540170 159628
rect 57462 159428 57468 159492
rect 57532 159490 57538 159492
rect 362902 159490 362908 159492
rect 57532 159430 362908 159490
rect 57532 159428 57538 159430
rect 362902 159428 362908 159430
rect 362972 159428 362978 159492
rect 395286 159428 395292 159492
rect 395356 159490 395362 159492
rect 573357 159490 573423 159493
rect 395356 159488 573423 159490
rect 395356 159432 573362 159488
rect 573418 159432 573423 159488
rect 395356 159430 573423 159432
rect 395356 159428 395362 159430
rect 573357 159427 573423 159430
rect 64505 159354 64571 159357
rect 553301 159354 553367 159357
rect 64505 159352 553367 159354
rect 64505 159296 64510 159352
rect 64566 159296 553306 159352
rect 553362 159296 553367 159352
rect 64505 159294 553367 159296
rect 64505 159291 64571 159294
rect 553301 159291 553367 159294
rect 395838 158612 395844 158676
rect 395908 158674 395914 158676
rect 537937 158674 538003 158677
rect 395908 158672 538003 158674
rect 395908 158616 537942 158672
rect 537998 158616 538003 158672
rect 395908 158614 538003 158616
rect 395908 158612 395914 158614
rect 537937 158611 538003 158614
rect 385493 158538 385559 158541
rect 541014 158538 541020 158540
rect 385493 158536 541020 158538
rect 385493 158480 385498 158536
rect 385554 158480 541020 158536
rect 385493 158478 541020 158480
rect 385493 158475 385559 158478
rect 541014 158476 541020 158478
rect 541084 158476 541090 158540
rect 358261 158402 358327 158405
rect 545430 158402 545436 158404
rect 358261 158400 545436 158402
rect 358261 158344 358266 158400
rect 358322 158344 545436 158400
rect 358261 158342 545436 158344
rect 358261 158339 358327 158342
rect 545430 158340 545436 158342
rect 545500 158340 545506 158404
rect 60038 158204 60044 158268
rect 60108 158266 60114 158268
rect 376845 158266 376911 158269
rect 60108 158264 376911 158266
rect 60108 158208 376850 158264
rect 376906 158208 376911 158264
rect 60108 158206 376911 158208
rect 60108 158204 60114 158206
rect 376845 158203 376911 158206
rect 377489 158266 377555 158269
rect 553894 158266 553900 158268
rect 377489 158264 553900 158266
rect 377489 158208 377494 158264
rect 377550 158208 553900 158264
rect 377489 158206 553900 158208
rect 377489 158203 377555 158206
rect 553894 158204 553900 158206
rect 553964 158204 553970 158268
rect 46054 158068 46060 158132
rect 46124 158130 46130 158132
rect 539910 158130 539916 158132
rect 46124 158070 539916 158130
rect 46124 158068 46130 158070
rect 539910 158068 539916 158070
rect 539980 158068 539986 158132
rect 32806 157932 32812 157996
rect 32876 157994 32882 157996
rect 547270 157994 547276 157996
rect 32876 157934 547276 157994
rect 32876 157932 32882 157934
rect 547270 157932 547276 157934
rect 547340 157932 547346 157996
rect 375046 156980 375052 157044
rect 375116 157042 375122 157044
rect 548006 157042 548012 157044
rect 375116 156982 548012 157042
rect 375116 156980 375122 156982
rect 548006 156980 548012 156982
rect 548076 156980 548082 157044
rect 359457 156906 359523 156909
rect 542854 156906 542860 156908
rect 359457 156904 542860 156906
rect 359457 156848 359462 156904
rect 359518 156848 542860 156904
rect 359457 156846 542860 156848
rect 359457 156843 359523 156846
rect 542854 156844 542860 156846
rect 542924 156844 542930 156908
rect 366357 156770 366423 156773
rect 571977 156770 572043 156773
rect 366357 156768 572043 156770
rect 366357 156712 366362 156768
rect 366418 156712 571982 156768
rect 572038 156712 572043 156768
rect 366357 156710 572043 156712
rect 366357 156707 366423 156710
rect 571977 156707 572043 156710
rect 36486 156572 36492 156636
rect 36556 156634 36562 156636
rect 384573 156634 384639 156637
rect 36556 156632 384639 156634
rect 36556 156576 384578 156632
rect 384634 156576 384639 156632
rect 36556 156574 384639 156576
rect 36556 156572 36562 156574
rect 384573 156571 384639 156574
rect 406326 156572 406332 156636
rect 406396 156634 406402 156636
rect 563605 156634 563671 156637
rect 406396 156632 563671 156634
rect 406396 156576 563610 156632
rect 563666 156576 563671 156632
rect 406396 156574 563671 156576
rect 406396 156572 406402 156574
rect 563605 156571 563671 156574
rect 46473 155954 46539 155957
rect 355358 155954 355364 155956
rect 46473 155952 355364 155954
rect 46473 155896 46478 155952
rect 46534 155896 355364 155952
rect 46473 155894 355364 155896
rect 46473 155891 46539 155894
rect 355358 155892 355364 155894
rect 355428 155892 355434 155956
rect 366449 155954 366515 155957
rect 544326 155954 544332 155956
rect 366449 155952 544332 155954
rect 366449 155896 366454 155952
rect 366510 155896 544332 155952
rect 366449 155894 544332 155896
rect 366449 155891 366515 155894
rect 544326 155892 544332 155894
rect 544396 155892 544402 155956
rect 50286 155756 50292 155820
rect 50356 155818 50362 155820
rect 376886 155818 376892 155820
rect 50356 155758 376892 155818
rect 50356 155756 50362 155758
rect 376886 155756 376892 155758
rect 376956 155756 376962 155820
rect 377581 155818 377647 155821
rect 543038 155818 543044 155820
rect 377581 155816 543044 155818
rect 377581 155760 377586 155816
rect 377642 155760 543044 155816
rect 377581 155758 543044 155760
rect 377581 155755 377647 155758
rect 543038 155756 543044 155758
rect 543108 155756 543114 155820
rect 35382 155620 35388 155684
rect 35452 155682 35458 155684
rect 440601 155682 440667 155685
rect 35452 155680 440667 155682
rect 35452 155624 440606 155680
rect 440662 155624 440667 155680
rect 35452 155622 440667 155624
rect 35452 155620 35458 155622
rect 440601 155619 440667 155622
rect 59302 155484 59308 155548
rect 59372 155546 59378 155548
rect 488533 155546 488599 155549
rect 59372 155544 488599 155546
rect 59372 155488 488538 155544
rect 488594 155488 488599 155544
rect 59372 155486 488599 155488
rect 59372 155484 59378 155486
rect 488533 155483 488599 155486
rect 46606 155348 46612 155412
rect 46676 155410 46682 155412
rect 543774 155410 543780 155412
rect 46676 155350 543780 155410
rect 46676 155348 46682 155350
rect 543774 155348 543780 155350
rect 543844 155348 543850 155412
rect 28441 155274 28507 155277
rect 566038 155274 566044 155276
rect 28441 155272 566044 155274
rect 28441 155216 28446 155272
rect 28502 155216 566044 155272
rect 28441 155214 566044 155216
rect 28441 155211 28507 155214
rect 566038 155212 566044 155214
rect 566108 155212 566114 155276
rect 410190 155076 410196 155140
rect 410260 155138 410266 155140
rect 573265 155138 573331 155141
rect 410260 155136 573331 155138
rect 410260 155080 573270 155136
rect 573326 155080 573331 155136
rect 410260 155078 573331 155080
rect 410260 155076 410266 155078
rect 573265 155075 573331 155078
rect 406510 153988 406516 154052
rect 406580 154050 406586 154052
rect 547873 154050 547939 154053
rect 406580 154048 547939 154050
rect 406580 153992 547878 154048
rect 547934 153992 547939 154048
rect 406580 153990 547939 153992
rect 406580 153988 406586 153990
rect 547873 153987 547939 153990
rect 381486 153852 381492 153916
rect 381556 153914 381562 153916
rect 541382 153914 541388 153916
rect 381556 153854 541388 153914
rect 381556 153852 381562 153854
rect 541382 153852 541388 153854
rect 541452 153852 541458 153916
rect 57278 153716 57284 153780
rect 57348 153778 57354 153780
rect 359590 153778 359596 153780
rect 57348 153718 359596 153778
rect 57348 153716 57354 153718
rect 359590 153716 359596 153718
rect 359660 153716 359666 153780
rect 360694 153716 360700 153780
rect 360764 153778 360770 153780
rect 552422 153778 552428 153780
rect 360764 153718 552428 153778
rect 360764 153716 360770 153718
rect 552422 153716 552428 153718
rect 552492 153716 552498 153780
rect 35801 153098 35867 153101
rect 129549 153098 129615 153101
rect 35801 153096 129615 153098
rect 35801 153040 35806 153096
rect 35862 153040 129554 153096
rect 129610 153040 129615 153096
rect 35801 153038 129615 153040
rect 35801 153035 35867 153038
rect 129549 153035 129615 153038
rect 292481 153098 292547 153101
rect 370589 153100 370655 153101
rect 347078 153098 347084 153100
rect 292481 153096 347084 153098
rect 292481 153040 292486 153096
rect 292542 153040 347084 153096
rect 292481 153038 347084 153040
rect 292481 153035 292547 153038
rect 347078 153036 347084 153038
rect 347148 153036 347154 153100
rect 370589 153096 370636 153100
rect 370700 153098 370706 153100
rect 370589 153040 370594 153096
rect 370589 153036 370636 153040
rect 370700 153038 370746 153098
rect 370700 153036 370706 153038
rect 396574 153036 396580 153100
rect 396644 153098 396650 153100
rect 447685 153098 447751 153101
rect 396644 153096 447751 153098
rect 396644 153040 447690 153096
rect 447746 153040 447751 153096
rect 396644 153038 447751 153040
rect 396644 153036 396650 153038
rect 370589 153035 370655 153036
rect 447685 153035 447751 153038
rect 34237 152962 34303 152965
rect 145649 152962 145715 152965
rect 34237 152960 145715 152962
rect 34237 152904 34242 152960
rect 34298 152904 145654 152960
rect 145710 152904 145715 152960
rect 34237 152902 145715 152904
rect 34237 152899 34303 152902
rect 145649 152899 145715 152902
rect 213913 152962 213979 152965
rect 355174 152962 355180 152964
rect 213913 152960 355180 152962
rect 213913 152904 213918 152960
rect 213974 152904 355180 152960
rect 213913 152902 355180 152904
rect 213913 152899 213979 152902
rect 355174 152900 355180 152902
rect 355244 152900 355250 152964
rect 398281 152962 398347 152965
rect 463785 152962 463851 152965
rect 398281 152960 463851 152962
rect 398281 152904 398286 152960
rect 398342 152904 463790 152960
rect 463846 152904 463851 152960
rect 398281 152902 463851 152904
rect 398281 152899 398347 152902
rect 463785 152899 463851 152902
rect 44725 152826 44791 152829
rect 170121 152826 170187 152829
rect 44725 152824 170187 152826
rect 44725 152768 44730 152824
rect 44786 152768 170126 152824
rect 170182 152768 170187 152824
rect 44725 152766 170187 152768
rect 44725 152763 44791 152766
rect 170121 152763 170187 152766
rect 197169 152826 197235 152829
rect 357014 152826 357020 152828
rect 197169 152824 357020 152826
rect 197169 152768 197174 152824
rect 197230 152768 357020 152824
rect 197169 152766 357020 152768
rect 197169 152763 197235 152766
rect 357014 152764 357020 152766
rect 357084 152764 357090 152828
rect 389950 152764 389956 152828
rect 390020 152826 390026 152828
rect 482461 152826 482527 152829
rect 390020 152824 482527 152826
rect 390020 152768 482466 152824
rect 482522 152768 482527 152824
rect 390020 152766 482527 152768
rect 390020 152764 390026 152766
rect 482461 152763 482527 152766
rect 20621 152690 20687 152693
rect 153377 152690 153443 152693
rect 20621 152688 153443 152690
rect 20621 152632 20626 152688
rect 20682 152632 153382 152688
rect 153438 152632 153443 152688
rect 20621 152630 153443 152632
rect 20621 152627 20687 152630
rect 153377 152627 153443 152630
rect 179137 152690 179203 152693
rect 388294 152690 388300 152692
rect 179137 152688 388300 152690
rect 179137 152632 179142 152688
rect 179198 152632 388300 152688
rect 179137 152630 388300 152632
rect 179137 152627 179203 152630
rect 388294 152628 388300 152630
rect 388364 152628 388370 152692
rect 399334 152628 399340 152692
rect 399404 152690 399410 152692
rect 498561 152690 498627 152693
rect 399404 152688 498627 152690
rect 399404 152632 498566 152688
rect 498622 152632 498627 152688
rect 399404 152630 498627 152632
rect 399404 152628 399410 152630
rect 498561 152627 498627 152630
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 61929 152554 61995 152557
rect 287697 152554 287763 152557
rect 61929 152552 287763 152554
rect 61929 152496 61934 152552
rect 61990 152496 287702 152552
rect 287758 152496 287763 152552
rect 61929 152494 287763 152496
rect 61929 152491 61995 152494
rect 287697 152491 287763 152494
rect 291193 152554 291259 152557
rect 346894 152554 346900 152556
rect 291193 152552 346900 152554
rect 291193 152496 291198 152552
rect 291254 152496 346900 152552
rect 291193 152494 346900 152496
rect 291193 152491 291259 152494
rect 346894 152492 346900 152494
rect 346964 152492 346970 152556
rect 374494 152492 374500 152556
rect 374564 152554 374570 152556
rect 563646 152554 563652 152556
rect 374564 152494 563652 152554
rect 374564 152492 374570 152494
rect 563646 152492 563652 152494
rect 563716 152492 563722 152556
rect 583520 152540 584960 152630
rect 72877 152418 72943 152421
rect 377254 152418 377260 152420
rect 72877 152416 377260 152418
rect 72877 152360 72882 152416
rect 72938 152360 377260 152416
rect 72877 152358 377260 152360
rect 72877 152355 72943 152358
rect 377254 152356 377260 152358
rect 377324 152356 377330 152420
rect 408534 152356 408540 152420
rect 408604 152418 408610 152420
rect 409045 152418 409111 152421
rect 408604 152416 409111 152418
rect 408604 152360 409050 152416
rect 409106 152360 409111 152416
rect 408604 152358 409111 152360
rect 408604 152356 408610 152358
rect 409045 152355 409111 152358
rect 409822 152356 409828 152420
rect 409892 152418 409898 152420
rect 546677 152418 546743 152421
rect 409892 152416 546743 152418
rect 409892 152360 546682 152416
rect 546738 152360 546743 152416
rect 409892 152358 546743 152360
rect 409892 152356 409898 152358
rect 546677 152355 546743 152358
rect 317597 152282 317663 152285
rect 351862 152282 351868 152284
rect 317597 152280 351868 152282
rect 317597 152224 317602 152280
rect 317658 152224 351868 152280
rect 317597 152222 351868 152224
rect 317597 152219 317663 152222
rect 351862 152220 351868 152222
rect 351932 152220 351938 152284
rect 360193 152282 360259 152285
rect 361430 152282 361436 152284
rect 360193 152280 361436 152282
rect 360193 152224 360198 152280
rect 360254 152224 361436 152280
rect 360193 152222 361436 152224
rect 360193 152219 360259 152222
rect 361430 152220 361436 152222
rect 361500 152220 361506 152284
rect 541249 151738 541315 151741
rect 541566 151738 541572 151740
rect 541249 151736 541572 151738
rect 541249 151680 541254 151736
rect 541310 151680 541572 151736
rect 541249 151678 541572 151680
rect 541249 151675 541315 151678
rect 541566 151676 541572 151678
rect 541636 151676 541642 151740
rect 60958 151540 60964 151604
rect 61028 151602 61034 151604
rect 117313 151602 117379 151605
rect 61028 151600 117379 151602
rect 61028 151544 117318 151600
rect 117374 151544 117379 151600
rect 61028 151542 117379 151544
rect 61028 151540 61034 151542
rect 117313 151539 117379 151542
rect 47669 151466 47735 151469
rect 365713 151466 365779 151469
rect 47669 151464 365779 151466
rect 47669 151408 47674 151464
rect 47730 151408 365718 151464
rect 365774 151408 365779 151464
rect 47669 151406 365779 151408
rect 47669 151403 47735 151406
rect 365713 151403 365779 151406
rect 391841 151466 391907 151469
rect 566406 151466 566412 151468
rect 391841 151464 566412 151466
rect 391841 151408 391846 151464
rect 391902 151408 566412 151464
rect 391841 151406 566412 151408
rect 391841 151403 391907 151406
rect 566406 151404 566412 151406
rect 566476 151404 566482 151468
rect 28257 151330 28323 151333
rect 548190 151330 548196 151332
rect 28257 151328 548196 151330
rect 28257 151272 28262 151328
rect 28318 151272 548196 151328
rect 28257 151270 548196 151272
rect 28257 151267 28323 151270
rect 548190 151268 548196 151270
rect 548260 151268 548266 151332
rect 21633 151194 21699 151197
rect 544142 151194 544148 151196
rect 21633 151192 544148 151194
rect 21633 151136 21638 151192
rect 21694 151136 544148 151192
rect 21633 151134 544148 151136
rect 21633 151131 21699 151134
rect 544142 151132 544148 151134
rect 544212 151132 544218 151196
rect 27061 151058 27127 151061
rect 549713 151058 549779 151061
rect 27061 151056 549779 151058
rect 27061 151000 27066 151056
rect 27122 151000 549718 151056
rect 549774 151000 549779 151056
rect 27061 150998 549779 151000
rect 27061 150995 27127 150998
rect 549713 150995 549779 150998
rect 46013 150514 46079 150517
rect 46606 150514 46612 150516
rect 46013 150512 46612 150514
rect 46013 150456 46018 150512
rect 46074 150456 46612 150512
rect 46013 150454 46612 150456
rect 46013 150451 46079 150454
rect 46606 150452 46612 150454
rect 46676 150452 46682 150516
rect 538857 150378 538923 150381
rect 569493 150378 569559 150381
rect 538857 150376 569559 150378
rect 538857 150320 538862 150376
rect 538918 150320 569498 150376
rect 569554 150320 569559 150376
rect 538857 150318 569559 150320
rect 538857 150315 538923 150318
rect 569493 150315 569559 150318
rect 539225 150242 539291 150245
rect 540973 150242 541039 150245
rect 563789 150242 563855 150245
rect 539225 150240 540898 150242
rect 539225 150184 539230 150240
rect 539286 150184 540898 150240
rect 539225 150182 540898 150184
rect 539225 150179 539291 150182
rect 388989 150106 389055 150109
rect 399937 150106 400003 150109
rect 540605 150106 540671 150109
rect 388989 150104 393330 150106
rect 388989 150048 388994 150104
rect 389050 150048 393330 150104
rect 388989 150046 393330 150048
rect 388989 150043 389055 150046
rect 393270 149970 393330 150046
rect 399937 150104 540671 150106
rect 399937 150048 399942 150104
rect 399998 150048 540610 150104
rect 540666 150048 540671 150104
rect 399937 150046 540671 150048
rect 540838 150106 540898 150182
rect 540973 150240 563855 150242
rect 540973 150184 540978 150240
rect 541034 150184 563794 150240
rect 563850 150184 563855 150240
rect 540973 150182 563855 150184
rect 540973 150179 541039 150182
rect 563789 150179 563855 150182
rect 545614 150106 545620 150108
rect 540838 150046 545620 150106
rect 399937 150043 400003 150046
rect 540605 150043 540671 150046
rect 545614 150044 545620 150046
rect 545684 150044 545690 150108
rect 548701 149970 548767 149973
rect 393270 149968 548767 149970
rect -960 149834 480 149924
rect 393270 149912 548706 149968
rect 548762 149912 548767 149968
rect 393270 149910 548767 149912
rect 548701 149907 548767 149910
rect 3509 149834 3575 149837
rect 540145 149834 540211 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect 539948 149832 540211 149834
rect 539948 149776 540150 149832
rect 540206 149776 540211 149832
rect 539948 149774 540211 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 540145 149771 540211 149774
rect 540421 149290 540487 149293
rect 554221 149290 554287 149293
rect 540421 149288 554287 149290
rect 540421 149232 540426 149288
rect 540482 149232 554226 149288
rect 554282 149232 554287 149288
rect 540421 149230 554287 149232
rect 540421 149227 540487 149230
rect 554221 149227 554287 149230
rect 540237 149154 540303 149157
rect 540237 149152 540346 149154
rect 540237 149096 540242 149152
rect 540298 149096 540346 149152
rect 540237 149091 540346 149096
rect 549662 149092 549668 149156
rect 549732 149154 549738 149156
rect 550173 149154 550239 149157
rect 549732 149152 550239 149154
rect 549732 149096 550178 149152
rect 550234 149096 550239 149152
rect 549732 149094 550239 149096
rect 549732 149092 549738 149094
rect 550173 149091 550239 149094
rect 540286 149018 540346 149091
rect 542118 149018 542124 149020
rect 540286 148958 542124 149018
rect 542118 148956 542124 148958
rect 542188 148956 542194 149020
rect 539358 148820 539364 148884
rect 539428 148882 539434 148884
rect 544469 148882 544535 148885
rect 539428 148880 544535 148882
rect 539428 148824 544474 148880
rect 544530 148824 544535 148880
rect 539428 148822 544535 148824
rect 539428 148820 539434 148822
rect 544469 148819 544535 148822
rect 539358 147868 539364 147932
rect 539428 147868 539434 147932
rect 541382 147868 541388 147932
rect 541452 147930 541458 147932
rect 541525 147930 541591 147933
rect 541452 147928 541591 147930
rect 541452 147872 541530 147928
rect 541586 147872 541591 147928
rect 541452 147870 541591 147872
rect 541452 147868 541458 147870
rect 55489 147522 55555 147525
rect 60590 147522 60596 147524
rect 55489 147520 60596 147522
rect 55489 147464 55494 147520
rect 55550 147464 60596 147520
rect 55489 147462 60596 147464
rect 55489 147459 55555 147462
rect 60590 147460 60596 147462
rect 60660 147460 60666 147524
rect 539366 147522 539426 147868
rect 541525 147867 541591 147870
rect 543089 147794 543155 147797
rect 540470 147792 543155 147794
rect 540470 147736 543094 147792
rect 543150 147736 543155 147792
rect 540470 147734 543155 147736
rect 540470 147661 540530 147734
rect 543089 147731 543155 147734
rect 540421 147656 540530 147661
rect 540421 147600 540426 147656
rect 540482 147600 540530 147656
rect 540421 147598 540530 147600
rect 540421 147595 540487 147598
rect 541934 147596 541940 147660
rect 542004 147658 542010 147660
rect 549437 147658 549503 147661
rect 542004 147656 549503 147658
rect 542004 147600 549442 147656
rect 549498 147600 549503 147656
rect 542004 147598 549503 147600
rect 542004 147596 542010 147598
rect 549437 147595 549503 147598
rect 551461 147522 551527 147525
rect 539366 147520 551527 147522
rect 539366 147464 551466 147520
rect 551522 147464 551527 147520
rect 539366 147462 551527 147464
rect 551461 147459 551527 147462
rect 539358 147324 539364 147388
rect 539428 147386 539434 147388
rect 540145 147386 540211 147389
rect 539428 147384 540211 147386
rect 539428 147328 540150 147384
rect 540206 147328 540211 147384
rect 539428 147326 540211 147328
rect 539428 147324 539434 147326
rect 540145 147323 540211 147326
rect 59670 147188 59676 147252
rect 59740 147250 59746 147252
rect 60590 147250 60596 147252
rect 59740 147190 60596 147250
rect 59740 147188 59746 147190
rect 60590 147188 60596 147190
rect 60660 147188 60666 147252
rect 539358 147188 539364 147252
rect 539428 147250 539434 147252
rect 540329 147250 540395 147253
rect 539428 147248 540395 147250
rect 539428 147192 540334 147248
rect 540390 147192 540395 147248
rect 539428 147190 540395 147192
rect 539428 147188 539434 147190
rect 540329 147187 540395 147190
rect 547965 147114 548031 147117
rect 547965 147112 548074 147114
rect 547965 147056 547970 147112
rect 548026 147056 548074 147112
rect 547965 147051 548074 147056
rect 540329 146978 540395 146981
rect 541014 146978 541020 146980
rect 540329 146976 541020 146978
rect 540329 146920 540334 146976
rect 540390 146920 541020 146976
rect 540329 146918 541020 146920
rect 540329 146915 540395 146918
rect 541014 146916 541020 146918
rect 541084 146916 541090 146980
rect 548014 146845 548074 147051
rect 58934 146780 58940 146844
rect 59004 146842 59010 146844
rect 60038 146842 60044 146844
rect 59004 146782 60044 146842
rect 59004 146780 59010 146782
rect 60038 146780 60044 146782
rect 60108 146780 60114 146844
rect 548014 146840 548123 146845
rect 548014 146784 548062 146840
rect 548118 146784 548123 146840
rect 548014 146782 548123 146784
rect 548057 146779 548123 146782
rect 59077 146570 59143 146573
rect 60590 146570 60596 146572
rect 59077 146568 60596 146570
rect 59077 146512 59082 146568
rect 59138 146512 60596 146568
rect 59077 146510 60596 146512
rect 59077 146507 59143 146510
rect 60590 146508 60596 146510
rect 60660 146508 60666 146572
rect 543549 146434 543615 146437
rect 539948 146432 543615 146434
rect 539948 146376 543554 146432
rect 543610 146376 543615 146432
rect 539948 146374 543615 146376
rect 543549 146371 543615 146374
rect 57881 145754 57947 145757
rect 542997 145754 543063 145757
rect 57881 145752 60076 145754
rect 57881 145696 57886 145752
rect 57942 145696 60076 145752
rect 57881 145694 60076 145696
rect 539948 145752 543063 145754
rect 539948 145696 543002 145752
rect 543058 145696 543063 145752
rect 539948 145694 543063 145696
rect 57881 145691 57947 145694
rect 542997 145691 543063 145694
rect 542537 144802 542603 144805
rect 542854 144802 542860 144804
rect 542537 144800 542860 144802
rect 542537 144744 542542 144800
rect 542598 144744 542860 144800
rect 542537 144742 542860 144744
rect 542537 144739 542603 144742
rect 542854 144740 542860 144742
rect 542924 144740 542930 144804
rect 543590 144740 543596 144804
rect 543660 144802 543666 144804
rect 543917 144802 543983 144805
rect 543660 144800 543983 144802
rect 543660 144744 543922 144800
rect 543978 144744 543983 144800
rect 543660 144742 543983 144744
rect 543660 144740 543666 144742
rect 543917 144739 543983 144742
rect 57646 142972 57652 143036
rect 57716 143034 57722 143036
rect 543089 143034 543155 143037
rect 57716 142974 60076 143034
rect 539948 143032 543155 143034
rect 539948 142976 543094 143032
rect 543150 142976 543155 143032
rect 539948 142974 543155 142976
rect 57716 142972 57722 142974
rect 543089 142971 543155 142974
rect 543181 142354 543247 142357
rect 539948 142352 543247 142354
rect 539948 142296 543186 142352
rect 543242 142296 543247 142352
rect 539948 142294 543247 142296
rect 543181 142291 543247 142294
rect 57881 141674 57947 141677
rect 543181 141674 543247 141677
rect 57881 141672 60076 141674
rect 57881 141616 57886 141672
rect 57942 141616 60076 141672
rect 57881 141614 60076 141616
rect 539948 141672 543247 141674
rect 539948 141616 543186 141672
rect 543242 141616 543247 141672
rect 539948 141614 543247 141616
rect 57881 141611 57947 141614
rect 543181 141611 543247 141614
rect 49601 141402 49667 141405
rect 59486 141402 59492 141404
rect 49601 141400 59492 141402
rect 49601 141344 49606 141400
rect 49662 141344 59492 141400
rect 49601 141342 59492 141344
rect 49601 141339 49667 141342
rect 59486 141340 59492 141342
rect 59556 141340 59562 141404
rect 542118 141204 542124 141268
rect 542188 141266 542194 141268
rect 546585 141266 546651 141269
rect 542188 141264 546651 141266
rect 542188 141208 546590 141264
rect 546646 141208 546651 141264
rect 542188 141206 546651 141208
rect 542188 141204 542194 141206
rect 546585 141203 546651 141206
rect 541382 141068 541388 141132
rect 541452 141130 541458 141132
rect 543038 141130 543044 141132
rect 541452 141070 543044 141130
rect 541452 141068 541458 141070
rect 543038 141068 543044 141070
rect 543108 141068 543114 141132
rect 59353 140994 59419 140997
rect 60406 140994 60412 140996
rect 59353 140992 60412 140994
rect 59353 140936 59358 140992
rect 59414 140936 60412 140992
rect 59353 140934 60412 140936
rect 59353 140931 59419 140934
rect 60406 140932 60412 140934
rect 60476 140932 60482 140996
rect 543641 140994 543707 140997
rect 539948 140992 543707 140994
rect 539948 140936 543646 140992
rect 543702 140936 543707 140992
rect 539948 140934 543707 140936
rect 543641 140931 543707 140934
rect 542302 140796 542308 140860
rect 542372 140858 542378 140860
rect 542537 140858 542603 140861
rect 542372 140856 542603 140858
rect 542372 140800 542542 140856
rect 542598 140800 542603 140856
rect 542372 140798 542603 140800
rect 542372 140796 542378 140798
rect 542537 140795 542603 140798
rect 57881 140314 57947 140317
rect 57881 140312 60076 140314
rect 57881 140256 57886 140312
rect 57942 140256 60076 140312
rect 57881 140254 60076 140256
rect 57881 140251 57947 140254
rect 57145 139634 57211 139637
rect 540329 139634 540395 139637
rect 541750 139634 541756 139636
rect 57145 139632 60076 139634
rect 57145 139576 57150 139632
rect 57206 139576 60076 139632
rect 57145 139574 60076 139576
rect 540329 139632 541756 139634
rect 540329 139576 540334 139632
rect 540390 139576 541756 139632
rect 540329 139574 541756 139576
rect 57145 139571 57211 139574
rect 540329 139571 540395 139574
rect 541750 139572 541756 139574
rect 541820 139572 541826 139636
rect 50797 139498 50863 139501
rect 50981 139498 51047 139501
rect 50797 139496 51047 139498
rect 50797 139440 50802 139496
rect 50858 139440 50986 139496
rect 51042 139440 51047 139496
rect 50797 139438 51047 139440
rect 50797 139435 50863 139438
rect 50981 139435 51047 139438
rect 540973 139498 541039 139501
rect 541566 139498 541572 139500
rect 540973 139496 541572 139498
rect 540973 139440 540978 139496
rect 541034 139440 541572 139496
rect 540973 139438 541572 139440
rect 540973 139435 541039 139438
rect 541566 139436 541572 139438
rect 541636 139436 541642 139500
rect 580441 139362 580507 139365
rect 583520 139362 584960 139452
rect 580441 139360 584960 139362
rect 580441 139304 580446 139360
rect 580502 139304 584960 139360
rect 580441 139302 584960 139304
rect 580441 139299 580507 139302
rect 583520 139212 584960 139302
rect 50613 138682 50679 138685
rect 58382 138682 58388 138684
rect 50613 138680 58388 138682
rect 50613 138624 50618 138680
rect 50674 138624 58388 138680
rect 50613 138622 58388 138624
rect 50613 138619 50679 138622
rect 58382 138620 58388 138622
rect 58452 138620 58458 138684
rect 543549 138274 543615 138277
rect 539948 138272 543615 138274
rect 539948 138216 543554 138272
rect 543610 138216 543615 138272
rect 539948 138214 543615 138216
rect 543549 138211 543615 138214
rect 58433 138138 58499 138141
rect 541985 138140 542051 138141
rect 58566 138138 58572 138140
rect 58433 138136 58572 138138
rect 58433 138080 58438 138136
rect 58494 138080 58572 138136
rect 58433 138078 58572 138080
rect 58433 138075 58499 138078
rect 58566 138076 58572 138078
rect 58636 138076 58642 138140
rect 541934 138138 541940 138140
rect 541894 138078 541940 138138
rect 542004 138136 542051 138140
rect 542046 138080 542051 138136
rect 541934 138076 541940 138078
rect 542004 138076 542051 138080
rect 541985 138075 542051 138076
rect 57881 137594 57947 137597
rect 57881 137592 60076 137594
rect 57881 137536 57886 137592
rect 57942 137536 60076 137592
rect 57881 137534 60076 137536
rect 57881 137531 57947 137534
rect 545246 137396 545252 137460
rect 545316 137396 545322 137460
rect 543590 137260 543596 137324
rect 543660 137322 543666 137324
rect 543825 137322 543891 137325
rect 543660 137320 543891 137322
rect 543660 137264 543830 137320
rect 543886 137264 543891 137320
rect 543660 137262 543891 137264
rect 543660 137260 543666 137262
rect 543825 137259 543891 137262
rect 545062 137124 545068 137188
rect 545132 137186 545138 137188
rect 545254 137186 545314 137396
rect 545132 137126 545314 137186
rect 545132 137124 545138 137126
rect -960 136778 480 136868
rect 3141 136778 3207 136781
rect -960 136776 3207 136778
rect -960 136720 3146 136776
rect 3202 136720 3207 136776
rect -960 136718 3207 136720
rect -960 136628 480 136718
rect 3141 136715 3207 136718
rect 543549 136234 543615 136237
rect 539948 136232 543615 136234
rect 539948 136176 543554 136232
rect 543610 136176 543615 136232
rect 539948 136174 543615 136176
rect 543549 136171 543615 136174
rect 543641 135554 543707 135557
rect 539948 135552 543707 135554
rect 45134 135220 45140 135284
rect 45204 135282 45210 135284
rect 60046 135282 60106 135524
rect 539948 135496 543646 135552
rect 543702 135496 543707 135552
rect 539948 135494 543707 135496
rect 543641 135491 543707 135494
rect 45204 135222 60106 135282
rect 45204 135220 45210 135222
rect 540789 135146 540855 135149
rect 545021 135148 545087 135149
rect 541014 135146 541020 135148
rect 540789 135144 541020 135146
rect 540789 135088 540794 135144
rect 540850 135088 541020 135144
rect 540789 135086 541020 135088
rect 540789 135083 540855 135086
rect 541014 135084 541020 135086
rect 541084 135084 541090 135148
rect 545021 135146 545068 135148
rect 544976 135144 545068 135146
rect 544976 135088 545026 135144
rect 544976 135086 545068 135088
rect 545021 135084 545068 135086
rect 545132 135084 545138 135148
rect 545021 135083 545087 135084
rect 57881 134874 57947 134877
rect 57881 134872 60076 134874
rect 57881 134816 57886 134872
rect 57942 134816 60076 134872
rect 57881 134814 60076 134816
rect 57881 134811 57947 134814
rect 543406 134404 543412 134468
rect 543476 134466 543482 134468
rect 556981 134466 557047 134469
rect 543476 134464 557047 134466
rect 543476 134408 556986 134464
rect 557042 134408 557047 134464
rect 543476 134406 557047 134408
rect 543476 134404 543482 134406
rect 556981 134403 557047 134406
rect 543549 134194 543615 134197
rect 539948 134192 543615 134194
rect 539948 134136 543554 134192
rect 543610 134136 543615 134192
rect 539948 134134 543615 134136
rect 543549 134131 543615 134134
rect 547638 133860 547644 133924
rect 547708 133922 547714 133924
rect 549897 133922 549963 133925
rect 547708 133920 549963 133922
rect 547708 133864 549902 133920
rect 549958 133864 549963 133920
rect 547708 133862 549963 133864
rect 547708 133860 547714 133862
rect 549897 133859 549963 133862
rect 541433 133514 541499 133517
rect 539948 133512 541499 133514
rect 539948 133456 541438 133512
rect 541494 133456 541499 133512
rect 539948 133454 541499 133456
rect 541433 133451 541499 133454
rect 57881 132834 57947 132837
rect 57881 132832 60076 132834
rect 57881 132776 57886 132832
rect 57942 132776 60076 132832
rect 57881 132774 60076 132776
rect 57881 132771 57947 132774
rect 53373 132562 53439 132565
rect 55438 132562 55444 132564
rect 53373 132560 55444 132562
rect 53373 132504 53378 132560
rect 53434 132504 55444 132560
rect 53373 132502 55444 132504
rect 53373 132499 53439 132502
rect 55438 132500 55444 132502
rect 55508 132500 55514 132564
rect 57053 131474 57119 131477
rect 543549 131474 543615 131477
rect 57053 131472 60076 131474
rect 57053 131416 57058 131472
rect 57114 131416 60076 131472
rect 57053 131414 60076 131416
rect 539948 131472 543615 131474
rect 539948 131416 543554 131472
rect 543610 131416 543615 131472
rect 539948 131414 543615 131416
rect 57053 131411 57119 131414
rect 543549 131411 543615 131414
rect 545021 131066 545087 131069
rect 545246 131066 545252 131068
rect 545021 131064 545252 131066
rect 545021 131008 545026 131064
rect 545082 131008 545252 131064
rect 545021 131006 545252 131008
rect 545021 131003 545087 131006
rect 545246 131004 545252 131006
rect 545316 131004 545322 131068
rect 57237 130794 57303 130797
rect 543549 130794 543615 130797
rect 57237 130792 60076 130794
rect 57237 130736 57242 130792
rect 57298 130736 60076 130792
rect 57237 130734 60076 130736
rect 539948 130792 543615 130794
rect 539948 130736 543554 130792
rect 543610 130736 543615 130792
rect 539948 130734 543615 130736
rect 57237 130731 57303 130734
rect 543549 130731 543615 130734
rect 541566 130188 541572 130252
rect 541636 130250 541642 130252
rect 548006 130250 548012 130252
rect 541636 130190 548012 130250
rect 541636 130188 541642 130190
rect 548006 130188 548012 130190
rect 548076 130188 548082 130252
rect 541750 130052 541756 130116
rect 541820 130114 541826 130116
rect 544101 130114 544167 130117
rect 541820 130112 544167 130114
rect 541820 130056 544106 130112
rect 544162 130056 544167 130112
rect 541820 130054 544167 130056
rect 541820 130052 541826 130054
rect 544101 130051 544167 130054
rect 541382 129916 541388 129980
rect 541452 129978 541458 129980
rect 542813 129978 542879 129981
rect 541452 129976 542879 129978
rect 541452 129920 542818 129976
rect 542874 129920 542879 129976
rect 541452 129918 542879 129920
rect 541452 129916 541458 129918
rect 542813 129915 542879 129918
rect 540881 129842 540947 129845
rect 541750 129842 541756 129844
rect 540881 129840 541756 129842
rect 540881 129784 540886 129840
rect 540942 129784 541756 129840
rect 540881 129782 541756 129784
rect 540881 129779 540947 129782
rect 541750 129780 541756 129782
rect 541820 129780 541826 129844
rect 544326 129434 544332 129436
rect 46238 128828 46244 128892
rect 46308 128890 46314 128892
rect 60046 128890 60106 129404
rect 539948 129374 544332 129434
rect 544326 129372 544332 129374
rect 544396 129372 544402 129436
rect 46308 128830 60106 128890
rect 46308 128828 46314 128830
rect 547505 128482 547571 128485
rect 547822 128482 547828 128484
rect 547505 128480 547828 128482
rect 547505 128424 547510 128480
rect 547566 128424 547828 128480
rect 547505 128422 547828 128424
rect 547505 128419 547571 128422
rect 547822 128420 547828 128422
rect 547892 128420 547898 128484
rect 57237 128074 57303 128077
rect 543549 128074 543615 128077
rect 57237 128072 60076 128074
rect 57237 128016 57242 128072
rect 57298 128016 60076 128072
rect 57237 128014 60076 128016
rect 539948 128072 543615 128074
rect 539948 128016 543554 128072
rect 543610 128016 543615 128072
rect 539948 128014 543615 128016
rect 57237 128011 57303 128014
rect 543549 128011 543615 128014
rect 543089 127666 543155 127669
rect 544510 127666 544516 127668
rect 543089 127664 544516 127666
rect 543089 127608 543094 127664
rect 543150 127608 544516 127664
rect 543089 127606 544516 127608
rect 543089 127603 543155 127606
rect 544510 127604 544516 127606
rect 544580 127604 544586 127668
rect 544878 126924 544884 126988
rect 544948 126986 544954 126988
rect 545614 126986 545620 126988
rect 544948 126926 545620 126986
rect 544948 126924 544954 126926
rect 545614 126924 545620 126926
rect 545684 126924 545690 126988
rect 547454 126924 547460 126988
rect 547524 126986 547530 126988
rect 547781 126986 547847 126989
rect 547524 126984 547847 126986
rect 547524 126928 547786 126984
rect 547842 126928 547847 126984
rect 547524 126926 547847 126928
rect 547524 126924 547530 126926
rect 547781 126923 547847 126926
rect 57237 126714 57303 126717
rect 57237 126712 60076 126714
rect 57237 126656 57242 126712
rect 57298 126656 60076 126712
rect 57237 126654 60076 126656
rect 57237 126651 57303 126654
rect 547638 126244 547644 126308
rect 547708 126306 547714 126308
rect 557073 126306 557139 126309
rect 547708 126304 557139 126306
rect 547708 126248 557078 126304
rect 557134 126248 557139 126304
rect 547708 126246 557139 126248
rect 547708 126244 547714 126246
rect 557073 126243 557139 126246
rect 547505 126170 547571 126173
rect 547638 126170 547644 126172
rect 547505 126168 547644 126170
rect 547505 126112 547510 126168
rect 547566 126112 547644 126168
rect 547505 126110 547644 126112
rect 547505 126107 547571 126110
rect 547638 126108 547644 126110
rect 547708 126108 547714 126172
rect 583520 125884 584960 126124
rect 543825 125626 543891 125629
rect 543958 125626 543964 125628
rect 543825 125624 543964 125626
rect 543825 125568 543830 125624
rect 543886 125568 543964 125624
rect 543825 125566 543964 125568
rect 543825 125563 543891 125566
rect 543958 125564 543964 125566
rect 544028 125564 544034 125628
rect 543406 125428 543412 125492
rect 543476 125490 543482 125492
rect 546585 125490 546651 125493
rect 543476 125488 546651 125490
rect 543476 125432 546590 125488
rect 546646 125432 546651 125488
rect 543476 125430 546651 125432
rect 543476 125428 543482 125430
rect 546585 125427 546651 125430
rect 57237 125354 57303 125357
rect 543549 125354 543615 125357
rect 57237 125352 60076 125354
rect 57237 125296 57242 125352
rect 57298 125296 60076 125352
rect 57237 125294 60076 125296
rect 539948 125352 543615 125354
rect 539948 125296 543554 125352
rect 543610 125296 543615 125352
rect 539948 125294 543615 125296
rect 57237 125291 57303 125294
rect 543549 125291 543615 125294
rect 547270 124674 547276 124676
rect 539948 124614 547276 124674
rect 547270 124612 547276 124614
rect 547340 124612 547346 124676
rect 542854 124068 542860 124132
rect 542924 124130 542930 124132
rect 546217 124130 546283 124133
rect 542924 124128 546283 124130
rect 542924 124072 546222 124128
rect 546278 124072 546283 124128
rect 542924 124070 546283 124072
rect 542924 124068 542930 124070
rect 546217 124067 546283 124070
rect 562174 124068 562180 124132
rect 562244 124130 562250 124132
rect 564709 124130 564775 124133
rect 562244 124128 564775 124130
rect 562244 124072 564714 124128
rect 564770 124072 564775 124128
rect 562244 124070 564775 124072
rect 562244 124068 562250 124070
rect 564709 124067 564775 124070
rect -960 123572 480 123812
rect 57237 123314 57303 123317
rect 57237 123312 60076 123314
rect 57237 123256 57242 123312
rect 57298 123256 60076 123312
rect 57237 123254 60076 123256
rect 57237 123251 57303 123254
rect 539358 122708 539364 122772
rect 539428 122770 539434 122772
rect 540145 122770 540211 122773
rect 539428 122768 540211 122770
rect 539428 122712 540150 122768
rect 540206 122712 540211 122768
rect 539428 122710 540211 122712
rect 539428 122708 539434 122710
rect 540145 122707 540211 122710
rect 543549 121954 543615 121957
rect 539948 121952 543615 121954
rect 539948 121896 543554 121952
rect 543610 121896 543615 121952
rect 539948 121894 543615 121896
rect 543549 121891 543615 121894
rect 57329 120594 57395 120597
rect 543549 120594 543615 120597
rect 57329 120592 60076 120594
rect 57329 120536 57334 120592
rect 57390 120536 60076 120592
rect 57329 120534 60076 120536
rect 539948 120592 543615 120594
rect 539948 120536 543554 120592
rect 543610 120536 543615 120592
rect 539948 120534 543615 120536
rect 57329 120531 57395 120534
rect 543549 120531 543615 120534
rect 57329 119914 57395 119917
rect 57329 119912 60076 119914
rect 57329 119856 57334 119912
rect 57390 119856 60076 119912
rect 57329 119854 60076 119856
rect 57329 119851 57395 119854
rect 56041 119234 56107 119237
rect 56041 119232 60076 119234
rect 56041 119176 56046 119232
rect 56102 119176 60076 119232
rect 56041 119174 60076 119176
rect 56041 119171 56107 119174
rect 548006 118764 548012 118828
rect 548076 118826 548082 118828
rect 549161 118826 549227 118829
rect 548076 118824 549227 118826
rect 548076 118768 549166 118824
rect 549222 118768 549227 118824
rect 548076 118766 549227 118768
rect 548076 118764 548082 118766
rect 549161 118763 549227 118766
rect 544142 117268 544148 117332
rect 544212 117330 544218 117332
rect 544653 117330 544719 117333
rect 544212 117328 544719 117330
rect 544212 117272 544658 117328
rect 544714 117272 544719 117328
rect 544212 117270 544719 117272
rect 544212 117268 544218 117270
rect 544653 117267 544719 117270
rect 57329 117194 57395 117197
rect 57329 117192 60076 117194
rect 57329 117136 57334 117192
rect 57390 117136 60076 117192
rect 57329 117134 60076 117136
rect 57329 117131 57395 117134
rect 543549 116514 543615 116517
rect 539948 116512 543615 116514
rect 539948 116456 543554 116512
rect 543610 116456 543615 116512
rect 539948 116454 543615 116456
rect 543549 116451 543615 116454
rect 57329 115834 57395 115837
rect 543549 115834 543615 115837
rect 57329 115832 60076 115834
rect 57329 115776 57334 115832
rect 57390 115776 60076 115832
rect 57329 115774 60076 115776
rect 539948 115832 543615 115834
rect 539948 115776 543554 115832
rect 543610 115776 543615 115832
rect 539948 115774 543615 115776
rect 57329 115771 57395 115774
rect 543549 115771 543615 115774
rect 58750 115092 58756 115156
rect 58820 115154 58826 115156
rect 58820 115094 60076 115154
rect 58820 115092 58826 115094
rect 544326 115092 544332 115156
rect 544396 115154 544402 115156
rect 552841 115154 552907 115157
rect 544396 115152 552907 115154
rect 544396 115096 552846 115152
rect 552902 115096 552907 115152
rect 544396 115094 552907 115096
rect 544396 115092 544402 115094
rect 552841 115091 552907 115094
rect 58433 114474 58499 114477
rect 58750 114474 58756 114476
rect 58433 114472 58756 114474
rect 58433 114416 58438 114472
rect 58494 114416 58756 114472
rect 58433 114414 58756 114416
rect 58433 114411 58499 114414
rect 58750 114412 58756 114414
rect 58820 114412 58826 114476
rect 543549 114474 543615 114477
rect 539948 114472 543615 114474
rect 57881 114338 57947 114341
rect 60046 114338 60106 114444
rect 539948 114416 543554 114472
rect 543610 114416 543615 114472
rect 539948 114414 543615 114416
rect 543549 114411 543615 114414
rect 57881 114336 60106 114338
rect 57881 114280 57886 114336
rect 57942 114280 60106 114336
rect 57881 114278 60106 114280
rect 57881 114275 57947 114278
rect 539358 114140 539364 114204
rect 539428 114202 539434 114204
rect 540145 114202 540211 114205
rect 539428 114200 540211 114202
rect 539428 114144 540150 114200
rect 540206 114144 540211 114200
rect 539428 114142 540211 114144
rect 539428 114140 539434 114142
rect 540145 114139 540211 114142
rect 543641 113794 543707 113797
rect 539948 113792 543707 113794
rect 539948 113736 543646 113792
rect 543702 113736 543707 113792
rect 539948 113734 543707 113736
rect 543641 113731 543707 113734
rect 57421 113114 57487 113117
rect 542302 113114 542308 113116
rect 57421 113112 60076 113114
rect 57421 113056 57426 113112
rect 57482 113056 60076 113112
rect 57421 113054 60076 113056
rect 539948 113054 542308 113114
rect 57421 113051 57487 113054
rect 542302 113052 542308 113054
rect 542372 113052 542378 113116
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect 48865 112434 48931 112437
rect 59486 112434 59492 112436
rect 48865 112432 59492 112434
rect 48865 112376 48870 112432
rect 48926 112376 59492 112432
rect 48865 112374 59492 112376
rect 48865 112371 48931 112374
rect 59486 112372 59492 112374
rect 59556 112372 59562 112436
rect 556889 112434 556955 112437
rect 566406 112434 566412 112436
rect 556889 112432 566412 112434
rect 556889 112376 556894 112432
rect 556950 112376 566412 112432
rect 556889 112374 566412 112376
rect 556889 112371 556955 112374
rect 566406 112372 566412 112374
rect 566476 112372 566482 112436
rect -960 110516 480 110756
rect 59486 110604 59492 110668
rect 59556 110666 59562 110668
rect 59629 110666 59695 110669
rect 59556 110664 59695 110666
rect 59556 110608 59634 110664
rect 59690 110608 59695 110664
rect 59556 110606 59695 110608
rect 59556 110604 59562 110606
rect 59629 110603 59695 110606
rect 543038 110604 543044 110668
rect 543108 110666 543114 110668
rect 544510 110666 544516 110668
rect 543108 110606 544516 110666
rect 543108 110604 543114 110606
rect 544510 110604 544516 110606
rect 544580 110604 544586 110668
rect 543958 110468 543964 110532
rect 544028 110530 544034 110532
rect 544653 110530 544719 110533
rect 544028 110528 544719 110530
rect 544028 110472 544658 110528
rect 544714 110472 544719 110528
rect 544028 110470 544719 110472
rect 544028 110468 544034 110470
rect 544653 110467 544719 110470
rect 57513 110394 57579 110397
rect 543549 110394 543615 110397
rect 57513 110392 60076 110394
rect 57513 110336 57518 110392
rect 57574 110336 60076 110392
rect 57513 110334 60076 110336
rect 539948 110392 543615 110394
rect 539948 110336 543554 110392
rect 543610 110336 543615 110392
rect 539948 110334 543615 110336
rect 57513 110331 57579 110334
rect 543549 110331 543615 110334
rect 542486 109714 542492 109716
rect 539948 109654 542492 109714
rect 542486 109652 542492 109654
rect 542556 109652 542562 109716
rect 544878 108972 544884 109036
rect 544948 109034 544954 109036
rect 547965 109034 548031 109037
rect 544948 109032 548031 109034
rect 544948 108976 547970 109032
rect 548026 108976 548031 109032
rect 544948 108974 548031 108976
rect 544948 108972 544954 108974
rect 547965 108971 548031 108974
rect 57513 108354 57579 108357
rect 57513 108352 60076 108354
rect 57513 108296 57518 108352
rect 57574 108296 60076 108352
rect 57513 108294 60076 108296
rect 57513 108291 57579 108294
rect 57421 107674 57487 107677
rect 542629 107674 542695 107677
rect 57421 107672 60076 107674
rect 57421 107616 57426 107672
rect 57482 107616 60076 107672
rect 57421 107614 60076 107616
rect 539948 107672 542695 107674
rect 539948 107616 542634 107672
rect 542690 107616 542695 107672
rect 539948 107614 542695 107616
rect 57421 107611 57487 107614
rect 542629 107611 542695 107614
rect 56041 107538 56107 107541
rect 59486 107538 59492 107540
rect 56041 107536 59492 107538
rect 56041 107480 56046 107536
rect 56102 107480 59492 107536
rect 56041 107478 59492 107480
rect 56041 107475 56107 107478
rect 59486 107476 59492 107478
rect 59556 107476 59562 107540
rect 54385 106722 54451 106725
rect 60038 106722 60044 106724
rect 54385 106720 60044 106722
rect 54385 106664 54390 106720
rect 54446 106664 60044 106720
rect 54385 106662 60044 106664
rect 54385 106659 54451 106662
rect 60038 106660 60044 106662
rect 60108 106660 60114 106724
rect 543273 106314 543339 106317
rect 539948 106312 543339 106314
rect 539948 106256 543278 106312
rect 543334 106256 543339 106312
rect 539948 106254 543339 106256
rect 543273 106251 543339 106254
rect 543222 106116 543228 106180
rect 543292 106178 543298 106180
rect 546493 106178 546559 106181
rect 543292 106176 546559 106178
rect 543292 106120 546498 106176
rect 546554 106120 546559 106176
rect 543292 106118 546559 106120
rect 543292 106116 543298 106118
rect 546493 106115 546559 106118
rect 57513 104274 57579 104277
rect 542670 104274 542676 104276
rect 57513 104272 60076 104274
rect 57513 104216 57518 104272
rect 57574 104216 60076 104272
rect 57513 104214 60076 104216
rect 539948 104214 542676 104274
rect 57513 104211 57579 104214
rect 542670 104212 542676 104214
rect 542740 104212 542746 104276
rect 57421 103594 57487 103597
rect 57421 103592 60076 103594
rect 57421 103536 57426 103592
rect 57482 103536 60076 103592
rect 57421 103534 60076 103536
rect 57421 103531 57487 103534
rect 57513 102914 57579 102917
rect 57513 102912 60076 102914
rect 57513 102856 57518 102912
rect 57574 102856 60076 102912
rect 57513 102854 60076 102856
rect 57513 102851 57579 102854
rect 57421 102234 57487 102237
rect 57421 102232 60076 102234
rect 57421 102176 57426 102232
rect 57482 102176 60076 102232
rect 57421 102174 60076 102176
rect 57421 102171 57487 102174
rect 59302 101492 59308 101556
rect 59372 101554 59378 101556
rect 541341 101554 541407 101557
rect 59372 101494 60076 101554
rect 539948 101552 541407 101554
rect 539948 101496 541346 101552
rect 541402 101496 541407 101552
rect 539948 101494 541407 101496
rect 59372 101492 59378 101494
rect 541341 101491 541407 101494
rect 46013 100058 46079 100061
rect 59302 100058 59308 100060
rect 46013 100056 59308 100058
rect 46013 100000 46018 100056
rect 46074 100000 59308 100056
rect 46013 99998 59308 100000
rect 46013 99995 46079 99998
rect 59302 99996 59308 99998
rect 59372 99996 59378 100060
rect 57513 99514 57579 99517
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 57513 99512 60076 99514
rect 57513 99456 57518 99512
rect 57574 99456 60076 99512
rect 57513 99454 60076 99456
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 57513 99451 57579 99454
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect 55949 98154 56015 98157
rect 55949 98152 60076 98154
rect 55949 98096 55954 98152
rect 56010 98096 60076 98152
rect 55949 98094 60076 98096
rect 55949 98091 56015 98094
rect -960 97610 480 97700
rect 2865 97610 2931 97613
rect -960 97608 2931 97610
rect -960 97552 2870 97608
rect 2926 97552 2931 97608
rect -960 97550 2931 97552
rect -960 97460 480 97550
rect 2865 97547 2931 97550
rect 543549 97474 543615 97477
rect 539948 97472 543615 97474
rect 539948 97416 543554 97472
rect 543610 97416 543615 97472
rect 539948 97414 543615 97416
rect 543549 97411 543615 97414
rect 57513 96794 57579 96797
rect 57513 96792 60076 96794
rect 57513 96736 57518 96792
rect 57574 96736 60076 96792
rect 57513 96734 60076 96736
rect 57513 96731 57579 96734
rect 543549 96114 543615 96117
rect 539948 96112 543615 96114
rect 539948 96056 543554 96112
rect 543610 96056 543615 96112
rect 539948 96054 543615 96056
rect 543549 96051 543615 96054
rect 542445 95434 542511 95437
rect 539948 95432 542511 95434
rect 539948 95376 542450 95432
rect 542506 95376 542511 95432
rect 539948 95374 542511 95376
rect 542445 95371 542511 95374
rect 57513 94074 57579 94077
rect 543549 94074 543615 94077
rect 57513 94072 60076 94074
rect 57513 94016 57518 94072
rect 57574 94016 60076 94072
rect 57513 94014 60076 94016
rect 539948 94072 543615 94074
rect 539948 94016 543554 94072
rect 543610 94016 543615 94072
rect 539948 94014 543615 94016
rect 57513 94011 57579 94014
rect 543549 94011 543615 94014
rect 57881 92714 57947 92717
rect 57881 92712 60076 92714
rect 57881 92656 57886 92712
rect 57942 92656 60076 92712
rect 57881 92654 60076 92656
rect 57881 92651 57947 92654
rect 539918 92578 539978 92684
rect 548190 92578 548196 92580
rect 539918 92518 548196 92578
rect 548190 92516 548196 92518
rect 548260 92516 548266 92580
rect 543549 92034 543615 92037
rect 539948 92032 543615 92034
rect 539948 91976 543554 92032
rect 543610 91976 543615 92032
rect 539948 91974 543615 91976
rect 543549 91971 543615 91974
rect 539910 91700 539916 91764
rect 539980 91700 539986 91764
rect 539918 91324 539978 91700
rect 57881 90674 57947 90677
rect 57881 90672 60076 90674
rect 57881 90616 57886 90672
rect 57942 90616 60076 90672
rect 57881 90614 60076 90616
rect 57881 90611 57947 90614
rect 540605 89994 540671 89997
rect 541382 89994 541388 89996
rect 540605 89992 541388 89994
rect 540605 89936 540610 89992
rect 540666 89936 541388 89992
rect 540605 89934 541388 89936
rect 540605 89931 540671 89934
rect 541382 89932 541388 89934
rect 541452 89932 541458 89996
rect 58525 89858 58591 89861
rect 59854 89858 59860 89860
rect 58525 89856 59860 89858
rect 58525 89800 58530 89856
rect 58586 89800 59860 89856
rect 58525 89798 59860 89800
rect 58525 89795 58591 89798
rect 59854 89796 59860 89798
rect 59924 89796 59930 89860
rect 541249 89858 541315 89861
rect 541750 89858 541756 89860
rect 541249 89856 541756 89858
rect 541249 89800 541254 89856
rect 541310 89800 541756 89856
rect 541249 89798 541756 89800
rect 541249 89795 541315 89798
rect 541750 89796 541756 89798
rect 541820 89796 541826 89860
rect 57881 89314 57947 89317
rect 57881 89312 60076 89314
rect 57881 89256 57886 89312
rect 57942 89256 60076 89312
rect 57881 89254 60076 89256
rect 57881 89251 57947 89254
rect 545614 88980 545620 89044
rect 545684 89042 545690 89044
rect 558269 89042 558335 89045
rect 545684 89040 558335 89042
rect 545684 88984 558274 89040
rect 558330 88984 558335 89040
rect 545684 88982 558335 88984
rect 545684 88980 545690 88982
rect 558269 88979 558335 88982
rect 543549 88634 543615 88637
rect 539948 88632 543615 88634
rect 539948 88576 543554 88632
rect 543610 88576 543615 88632
rect 539948 88574 543615 88576
rect 543549 88571 543615 88574
rect 543774 87954 543780 87956
rect 539948 87894 543780 87954
rect 543774 87892 543780 87894
rect 543844 87892 543850 87956
rect 539358 86804 539364 86868
rect 539428 86866 539434 86868
rect 540421 86866 540487 86869
rect 539428 86864 540487 86866
rect 539428 86808 540426 86864
rect 540482 86808 540487 86864
rect 539428 86806 540487 86808
rect 539428 86804 539434 86806
rect 540421 86803 540487 86806
rect 544510 86804 544516 86868
rect 544580 86866 544586 86868
rect 547321 86866 547387 86869
rect 544580 86864 547387 86866
rect 544580 86808 547326 86864
rect 547382 86808 547387 86864
rect 544580 86806 547387 86808
rect 544580 86804 544586 86806
rect 547321 86803 547387 86806
rect 56317 86594 56383 86597
rect 56317 86592 60076 86594
rect 56317 86536 56322 86592
rect 56378 86536 60076 86592
rect 56317 86534 60076 86536
rect 56317 86531 56383 86534
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect 539918 84690 539978 85204
rect 552606 84690 552612 84692
rect 539918 84630 552612 84690
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 552606 84628 552612 84630
rect 552676 84628 552682 84692
rect 542353 84554 542419 84557
rect 539948 84552 542419 84554
rect 539948 84496 542358 84552
rect 542414 84496 542419 84552
rect 539948 84494 542419 84496
rect 542353 84491 542419 84494
rect 543549 83874 543615 83877
rect 539948 83872 543615 83874
rect 539948 83816 543554 83872
rect 543610 83816 543615 83872
rect 539948 83814 543615 83816
rect 543549 83811 543615 83814
rect 544653 82922 544719 82925
rect 547454 82922 547460 82924
rect 544653 82920 547460 82922
rect 544653 82864 544658 82920
rect 544714 82864 547460 82920
rect 544653 82862 547460 82864
rect 544653 82859 544719 82862
rect 547454 82860 547460 82862
rect 547524 82860 547530 82924
rect 57605 82514 57671 82517
rect 543549 82514 543615 82517
rect 57605 82512 60076 82514
rect 57605 82456 57610 82512
rect 57666 82456 60076 82512
rect 57605 82454 60076 82456
rect 539948 82512 543615 82514
rect 539948 82456 543554 82512
rect 543610 82456 543615 82512
rect 539948 82454 543615 82456
rect 57605 82451 57671 82454
rect 543549 82451 543615 82454
rect 57881 81834 57947 81837
rect 57881 81832 60076 81834
rect 57881 81776 57886 81832
rect 57942 81776 60076 81832
rect 57881 81774 60076 81776
rect 57881 81771 57947 81774
rect 57053 81154 57119 81157
rect 57053 81152 60076 81154
rect 57053 81096 57058 81152
rect 57114 81096 60076 81152
rect 57053 81094 60076 81096
rect 57053 81091 57119 81094
rect 543549 78434 543615 78437
rect 539948 78432 543615 78434
rect 539948 78376 543554 78432
rect 543610 78376 543615 78432
rect 539948 78374 543615 78376
rect 543549 78371 543615 78374
rect 543641 77754 543707 77757
rect 539948 77752 543707 77754
rect 539948 77696 543646 77752
rect 543702 77696 543707 77752
rect 539948 77694 543707 77696
rect 543641 77691 543707 77694
rect 56133 77074 56199 77077
rect 56133 77072 60076 77074
rect 56133 77016 56138 77072
rect 56194 77016 60076 77072
rect 56133 77014 60076 77016
rect 56133 77011 56199 77014
rect 543549 76394 543615 76397
rect 539948 76392 543615 76394
rect 539948 76336 543554 76392
rect 543610 76336 543615 76392
rect 539948 76334 543615 76336
rect 543549 76331 543615 76334
rect 540278 75788 540284 75852
rect 540348 75850 540354 75852
rect 541249 75850 541315 75853
rect 540348 75848 541315 75850
rect 540348 75792 541254 75848
rect 541310 75792 541315 75848
rect 540348 75790 541315 75792
rect 540348 75788 540354 75790
rect 541249 75787 541315 75790
rect 57605 75714 57671 75717
rect 543549 75714 543615 75717
rect 57605 75712 60076 75714
rect 57605 75656 57610 75712
rect 57666 75656 60076 75712
rect 57605 75654 60076 75656
rect 539948 75712 543615 75714
rect 539948 75656 543554 75712
rect 543610 75656 543615 75712
rect 539948 75654 543615 75656
rect 57605 75651 57671 75654
rect 543549 75651 543615 75654
rect 57462 74972 57468 75036
rect 57532 75034 57538 75036
rect 542721 75034 542787 75037
rect 57532 74974 60076 75034
rect 539948 75032 542787 75034
rect 539948 74976 542726 75032
rect 542782 74976 542787 75032
rect 539948 74974 542787 74976
rect 57532 74972 57538 74974
rect 542721 74971 542787 74974
rect 545430 72994 545436 72996
rect 539948 72934 545436 72994
rect 545430 72932 545436 72934
rect 545500 72932 545506 72996
rect 580257 72994 580323 72997
rect 583520 72994 584960 73084
rect 580257 72992 584960 72994
rect 580257 72936 580262 72992
rect 580318 72936 584960 72992
rect 580257 72934 584960 72936
rect 580257 72931 580323 72934
rect 583520 72844 584960 72934
rect 547270 72388 547276 72452
rect 547340 72450 547346 72452
rect 547873 72450 547939 72453
rect 547340 72448 547939 72450
rect 547340 72392 547878 72448
rect 547934 72392 547939 72448
rect 547340 72390 547939 72392
rect 547340 72388 547346 72390
rect 547873 72387 547939 72390
rect -960 71484 480 71724
rect 543549 71634 543615 71637
rect 539948 71632 543615 71634
rect 539948 71576 543554 71632
rect 543610 71576 543615 71632
rect 539948 71574 543615 71576
rect 543549 71571 543615 71574
rect 541198 70954 541204 70956
rect 539948 70894 541204 70954
rect 541198 70892 541204 70894
rect 541268 70892 541274 70956
rect 56777 70274 56843 70277
rect 543549 70274 543615 70277
rect 56777 70272 60076 70274
rect 56777 70216 56782 70272
rect 56838 70216 60076 70272
rect 56777 70214 60076 70216
rect 539948 70272 543615 70274
rect 539948 70216 543554 70272
rect 543610 70216 543615 70272
rect 539948 70214 543615 70216
rect 56777 70211 56843 70214
rect 543549 70211 543615 70214
rect 58750 68852 58756 68916
rect 58820 68914 58826 68916
rect 58820 68854 60076 68914
rect 58820 68852 58826 68854
rect 57605 68234 57671 68237
rect 539918 68234 539978 68884
rect 57605 68232 60076 68234
rect 57605 68176 57610 68232
rect 57666 68176 60076 68232
rect 57605 68174 60076 68176
rect 539918 68174 547890 68234
rect 57605 68171 57671 68174
rect 547830 67690 547890 68174
rect 566038 67690 566044 67692
rect 547830 67630 566044 67690
rect 566038 67628 566044 67630
rect 566108 67628 566114 67692
rect 56685 67554 56751 67557
rect 56685 67552 60076 67554
rect 56685 67496 56690 67552
rect 56746 67496 60076 67552
rect 56685 67494 60076 67496
rect 56685 67491 56751 67494
rect 543549 66194 543615 66197
rect 539948 66192 543615 66194
rect 539948 66136 543554 66192
rect 543610 66136 543615 66192
rect 539948 66134 543615 66136
rect 543549 66131 543615 66134
rect 542813 65514 542879 65517
rect 539948 65512 542879 65514
rect 539948 65456 542818 65512
rect 542874 65456 542879 65512
rect 539948 65454 542879 65456
rect 542813 65451 542879 65454
rect 57881 64834 57947 64837
rect 57881 64832 60076 64834
rect 57881 64776 57886 64832
rect 57942 64776 60076 64832
rect 57881 64774 60076 64776
rect 57881 64771 57947 64774
rect 56961 64154 57027 64157
rect 543549 64154 543615 64157
rect 56961 64152 60076 64154
rect 56961 64096 56966 64152
rect 57022 64096 60076 64152
rect 56961 64094 60076 64096
rect 539948 64152 543615 64154
rect 539948 64096 543554 64152
rect 543610 64096 543615 64152
rect 539948 64094 543615 64096
rect 56961 64091 57027 64094
rect 543549 64091 543615 64094
rect 57697 63474 57763 63477
rect 57697 63472 60076 63474
rect 57697 63416 57702 63472
rect 57758 63416 60076 63472
rect 57697 63414 60076 63416
rect 57697 63411 57763 63414
rect 57697 62114 57763 62117
rect 543549 62114 543615 62117
rect 57697 62112 60076 62114
rect 57697 62056 57702 62112
rect 57758 62056 60076 62112
rect 57697 62054 60076 62056
rect 539948 62112 543615 62114
rect 539948 62056 543554 62112
rect 543610 62056 543615 62112
rect 539948 62054 543615 62056
rect 57697 62051 57763 62054
rect 543549 62051 543615 62054
rect 543641 60754 543707 60757
rect 539948 60752 543707 60754
rect 539948 60696 543646 60752
rect 543702 60696 543707 60752
rect 539948 60694 543707 60696
rect 543641 60691 543707 60694
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect 57789 59394 57855 59397
rect 57789 59392 60076 59394
rect 57789 59336 57794 59392
rect 57850 59336 60076 59392
rect 57789 59334 60076 59336
rect 57789 59331 57855 59334
rect 57697 58714 57763 58717
rect 57697 58712 60076 58714
rect -960 58578 480 58668
rect 57697 58656 57702 58712
rect 57758 58656 60076 58712
rect 57697 58654 60076 58656
rect 57697 58651 57763 58654
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 39246 57972 39252 58036
rect 39316 58034 39322 58036
rect 39316 57974 60076 58034
rect 39316 57972 39322 57974
rect 57697 57354 57763 57357
rect 57697 57352 60076 57354
rect 57697 57296 57702 57352
rect 57758 57296 60076 57352
rect 57697 57294 60076 57296
rect 57697 57291 57763 57294
rect 543549 56674 543615 56677
rect 539948 56672 543615 56674
rect 539948 56616 543554 56672
rect 543610 56616 543615 56672
rect 539948 56614 543615 56616
rect 543549 56611 543615 56614
rect 57881 55994 57947 55997
rect 543958 55994 543964 55996
rect 57881 55992 60076 55994
rect 57881 55936 57886 55992
rect 57942 55936 60076 55992
rect 57881 55934 60076 55936
rect 539948 55934 543964 55994
rect 57881 55931 57947 55934
rect 543958 55932 543964 55934
rect 544028 55932 544034 55996
rect 56225 55314 56291 55317
rect 56225 55312 60076 55314
rect 56225 55256 56230 55312
rect 56286 55256 60076 55312
rect 56225 55254 60076 55256
rect 56225 55251 56291 55254
rect 59118 54572 59124 54636
rect 59188 54634 59194 54636
rect 59188 54574 60076 54634
rect 59188 54572 59194 54574
rect 57697 53274 57763 53277
rect 57697 53272 60076 53274
rect 57697 53216 57702 53272
rect 57758 53216 60076 53272
rect 57697 53214 60076 53216
rect 57697 53211 57763 53214
rect 543549 52594 543615 52597
rect 539948 52592 543615 52594
rect 539948 52536 543554 52592
rect 543610 52536 543615 52592
rect 539948 52534 543615 52536
rect 543549 52531 543615 52534
rect 539918 51098 539978 51204
rect 551502 51098 551508 51100
rect 539918 51038 551508 51098
rect 551502 51036 551508 51038
rect 551572 51036 551578 51100
rect 543457 49874 543523 49877
rect 539948 49872 543523 49874
rect 539948 49816 543462 49872
rect 543518 49816 543523 49872
rect 539948 49814 543523 49816
rect 543457 49811 543523 49814
rect 57830 49132 57836 49196
rect 57900 49194 57906 49196
rect 57900 49134 60076 49194
rect 57900 49132 57906 49134
rect 543549 48514 543615 48517
rect 539948 48512 543615 48514
rect 539948 48456 543554 48512
rect 543610 48456 543615 48512
rect 539948 48454 543615 48456
rect 543549 48451 543615 48454
rect 543549 47834 543615 47837
rect 539948 47832 543615 47834
rect 539948 47776 543554 47832
rect 543610 47776 543615 47832
rect 539948 47774 543615 47776
rect 543549 47771 543615 47774
rect 57697 47154 57763 47157
rect 57697 47152 60076 47154
rect 57697 47096 57702 47152
rect 57758 47096 60076 47152
rect 57697 47094 60076 47096
rect 57697 47091 57763 47094
rect 539961 46882 540027 46885
rect 539918 46880 540027 46882
rect 539918 46824 539966 46880
rect 540022 46824 540027 46880
rect 539918 46819 540027 46824
rect 57053 46474 57119 46477
rect 57053 46472 60076 46474
rect 57053 46416 57058 46472
rect 57114 46416 60076 46472
rect 539918 46444 539978 46819
rect 57053 46414 60076 46416
rect 57053 46411 57119 46414
rect 583520 46188 584960 46428
rect 58157 45794 58223 45797
rect 58157 45792 60076 45794
rect 58157 45736 58162 45792
rect 58218 45736 60076 45792
rect 58157 45734 60076 45736
rect 58157 45731 58223 45734
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 58341 45114 58407 45117
rect 543549 45114 543615 45117
rect 58341 45112 60076 45114
rect 58341 45056 58346 45112
rect 58402 45056 60076 45112
rect 58341 45054 60076 45056
rect 539948 45112 543615 45114
rect 539948 45056 543554 45112
rect 543610 45056 543615 45112
rect 539948 45054 543615 45056
rect 58341 45051 58407 45054
rect 543549 45051 543615 45054
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 543641 44434 543707 44437
rect 539948 44432 543707 44434
rect 539948 44376 543646 44432
rect 543702 44376 543707 44432
rect 539948 44374 543707 44376
rect 543641 44371 543707 44374
rect 53046 44298 53052 44300
rect 6870 44238 53052 44298
rect 53046 44236 53052 44238
rect 53116 44236 53122 44300
rect 543549 43754 543615 43757
rect 539948 43752 543615 43754
rect 539948 43696 543554 43752
rect 543610 43696 543615 43752
rect 539948 43694 543615 43696
rect 543549 43691 543615 43694
rect 542353 42394 542419 42397
rect 539948 42392 542419 42394
rect 539948 42336 542358 42392
rect 542414 42336 542419 42392
rect 539948 42334 542419 42336
rect 542353 42331 542419 42334
rect 58249 41714 58315 41717
rect 58249 41712 60076 41714
rect 58249 41656 58254 41712
rect 58310 41656 60076 41712
rect 58249 41654 60076 41656
rect 58249 41651 58315 41654
rect 57697 41034 57763 41037
rect 543549 41034 543615 41037
rect 57697 41032 60076 41034
rect 57697 40976 57702 41032
rect 57758 40976 60076 41032
rect 57697 40974 60076 40976
rect 539948 41032 543615 41034
rect 539948 40976 543554 41032
rect 543610 40976 543615 41032
rect 539948 40974 543615 40976
rect 57697 40971 57763 40974
rect 543549 40971 543615 40974
rect 57145 40354 57211 40357
rect 57145 40352 60076 40354
rect 57145 40296 57150 40352
rect 57206 40296 60076 40352
rect 57145 40294 60076 40296
rect 57145 40291 57211 40294
rect 57697 39674 57763 39677
rect 57697 39672 60076 39674
rect 57697 39616 57702 39672
rect 57758 39616 60076 39672
rect 57697 39614 60076 39616
rect 57697 39611 57763 39614
rect 539542 38524 539548 38588
rect 539612 38524 539618 38588
rect 539550 38284 539610 38524
rect 542353 37634 542419 37637
rect 539948 37632 542419 37634
rect 539948 37576 542358 37632
rect 542414 37576 542419 37632
rect 539948 37574 542419 37576
rect 542353 37571 542419 37574
rect 543549 36274 543615 36277
rect 539948 36272 543615 36274
rect 539948 36216 543554 36272
rect 543610 36216 543615 36272
rect 539948 36214 543615 36216
rect 543549 36211 543615 36214
rect 543549 35594 543615 35597
rect 539948 35592 543615 35594
rect 46606 34988 46612 35052
rect 46676 35050 46682 35052
rect 60046 35050 60106 35564
rect 539948 35536 543554 35592
rect 543610 35536 543615 35592
rect 539948 35534 543615 35536
rect 543549 35531 543615 35534
rect 539726 35260 539732 35324
rect 539796 35260 539802 35324
rect 46676 34990 60106 35050
rect 46676 34988 46682 34990
rect 57278 34852 57284 34916
rect 57348 34914 57354 34916
rect 57348 34854 60076 34914
rect 539734 34884 539794 35260
rect 57348 34852 57354 34854
rect 57697 33554 57763 33557
rect 57697 33552 60076 33554
rect 57697 33496 57702 33552
rect 57758 33496 60076 33552
rect 57697 33494 60076 33496
rect 57697 33491 57763 33494
rect 579797 33146 579863 33149
rect 583520 33146 584960 33236
rect 579797 33144 584960 33146
rect 579797 33088 579802 33144
rect 579858 33088 584960 33144
rect 579797 33086 584960 33088
rect 579797 33083 579863 33086
rect 583520 32996 584960 33086
rect 57697 32874 57763 32877
rect 57697 32872 60076 32874
rect 57697 32816 57702 32872
rect 57758 32816 60076 32872
rect 57697 32814 60076 32816
rect 57697 32811 57763 32814
rect -960 32316 480 32556
rect 57789 32194 57855 32197
rect 57789 32192 60076 32194
rect 57789 32136 57794 32192
rect 57850 32136 60076 32192
rect 57789 32134 60076 32136
rect 57789 32131 57855 32134
rect 539358 31588 539364 31652
rect 539428 31650 539434 31652
rect 540881 31650 540947 31653
rect 539428 31648 540947 31650
rect 539428 31592 540886 31648
rect 540942 31592 540947 31648
rect 539428 31590 540947 31592
rect 539428 31588 539434 31590
rect 540881 31587 540947 31590
rect 57697 31514 57763 31517
rect 57697 31512 60076 31514
rect 57697 31456 57702 31512
rect 57758 31456 60076 31512
rect 57697 31454 60076 31456
rect 57697 31451 57763 31454
rect 44909 31106 44975 31109
rect 60590 31106 60596 31108
rect 44909 31104 60596 31106
rect 44909 31048 44914 31104
rect 44970 31048 60596 31104
rect 44909 31046 60596 31048
rect 44909 31043 44975 31046
rect 60590 31044 60596 31046
rect 60660 31044 60666 31108
rect 539366 30970 539426 31484
rect 539542 31044 539548 31108
rect 539612 31106 539618 31108
rect 539612 31046 547890 31106
rect 539612 31044 539618 31046
rect 547830 30970 547890 31046
rect 582557 30970 582623 30973
rect 539366 30910 543842 30970
rect 547830 30968 582623 30970
rect 547830 30912 582562 30968
rect 582618 30912 582623 30968
rect 547830 30910 582623 30912
rect 57329 30834 57395 30837
rect 543549 30834 543615 30837
rect 57329 30832 60076 30834
rect 57329 30776 57334 30832
rect 57390 30776 60076 30832
rect 57329 30774 60076 30776
rect 539948 30832 543615 30834
rect 539948 30776 543554 30832
rect 543610 30776 543615 30832
rect 539948 30774 543615 30776
rect 543782 30834 543842 30910
rect 582557 30907 582623 30910
rect 552238 30834 552244 30836
rect 543782 30774 552244 30834
rect 57329 30771 57395 30774
rect 543549 30771 543615 30774
rect 552238 30772 552244 30774
rect 552308 30772 552314 30836
rect 59302 30500 59308 30564
rect 59372 30562 59378 30564
rect 59905 30562 59971 30565
rect 59372 30560 59971 30562
rect 59372 30504 59910 30560
rect 59966 30504 59971 30560
rect 59372 30502 59971 30504
rect 59372 30500 59378 30502
rect 59905 30499 59971 30502
rect 539358 30500 539364 30564
rect 539428 30562 539434 30564
rect 541709 30562 541775 30565
rect 539428 30560 541775 30562
rect 539428 30504 541714 30560
rect 541770 30504 541775 30560
rect 539428 30502 541775 30504
rect 539428 30500 539434 30502
rect 541709 30499 541775 30502
rect 59905 29882 59971 29885
rect 66437 29882 66503 29885
rect 59905 29880 66503 29882
rect 59905 29824 59910 29880
rect 59966 29824 66442 29880
rect 66498 29824 66503 29880
rect 59905 29822 66503 29824
rect 59905 29819 59971 29822
rect 66437 29819 66503 29822
rect 539501 29882 539567 29885
rect 561622 29882 561628 29884
rect 539501 29880 561628 29882
rect 539501 29824 539506 29880
rect 539562 29824 561628 29880
rect 539501 29822 561628 29824
rect 539501 29819 539567 29822
rect 561622 29820 561628 29822
rect 561692 29820 561698 29884
rect 54845 29746 54911 29749
rect 82813 29746 82879 29749
rect 54845 29744 82879 29746
rect 54845 29688 54850 29744
rect 54906 29688 82818 29744
rect 82874 29688 82879 29744
rect 54845 29686 82879 29688
rect 54845 29683 54911 29686
rect 82813 29683 82879 29686
rect 49325 29610 49391 29613
rect 61285 29610 61351 29613
rect 49325 29608 61351 29610
rect 49325 29552 49330 29608
rect 49386 29552 61290 29608
rect 61346 29552 61351 29608
rect 49325 29550 61351 29552
rect 49325 29547 49391 29550
rect 61285 29547 61351 29550
rect 521101 29610 521167 29613
rect 552054 29610 552060 29612
rect 521101 29608 552060 29610
rect 521101 29552 521106 29608
rect 521162 29552 552060 29608
rect 521101 29550 552060 29552
rect 521101 29547 521167 29550
rect 552054 29548 552060 29550
rect 552124 29548 552130 29612
rect 41086 29412 41092 29476
rect 41156 29474 41162 29476
rect 284109 29474 284175 29477
rect 41156 29472 284175 29474
rect 41156 29416 284114 29472
rect 284170 29416 284175 29472
rect 41156 29414 284175 29416
rect 41156 29412 41162 29414
rect 284109 29411 284175 29414
rect 519169 29474 519235 29477
rect 564525 29474 564591 29477
rect 519169 29472 564591 29474
rect 519169 29416 519174 29472
rect 519230 29416 564530 29472
rect 564586 29416 564591 29472
rect 519169 29414 564591 29416
rect 519169 29411 519235 29414
rect 564525 29411 564591 29414
rect 48998 29276 49004 29340
rect 49068 29338 49074 29340
rect 300853 29338 300919 29341
rect 49068 29336 300919 29338
rect 49068 29280 300858 29336
rect 300914 29280 300919 29336
rect 49068 29278 300919 29280
rect 49068 29276 49074 29278
rect 300853 29275 300919 29278
rect 314377 29338 314443 29341
rect 561806 29338 561812 29340
rect 314377 29336 561812 29338
rect 314377 29280 314382 29336
rect 314438 29280 561812 29336
rect 314377 29278 561812 29280
rect 314377 29275 314443 29278
rect 561806 29276 561812 29278
rect 561876 29276 561882 29340
rect 49366 29140 49372 29204
rect 49436 29202 49442 29204
rect 59905 29202 59971 29205
rect 49436 29200 59971 29202
rect 49436 29144 59910 29200
rect 59966 29144 59971 29200
rect 49436 29142 59971 29144
rect 49436 29140 49442 29142
rect 59905 29139 59971 29142
rect 182357 29202 182423 29205
rect 550398 29202 550404 29204
rect 182357 29200 550404 29202
rect 182357 29144 182362 29200
rect 182418 29144 550404 29200
rect 182357 29142 550404 29144
rect 182357 29139 182423 29142
rect 550398 29140 550404 29142
rect 550468 29140 550474 29204
rect 23289 29066 23355 29069
rect 416129 29066 416195 29069
rect 23289 29064 416195 29066
rect 23289 29008 23294 29064
rect 23350 29008 416134 29064
rect 416190 29008 416195 29064
rect 23289 29006 416195 29008
rect 23289 29003 23355 29006
rect 416129 29003 416195 29006
rect 481817 29066 481883 29069
rect 565445 29066 565511 29069
rect 481817 29064 565511 29066
rect 481817 29008 481822 29064
rect 481878 29008 565450 29064
rect 565506 29008 565511 29064
rect 481817 29006 565511 29008
rect 481817 29003 481883 29006
rect 565445 29003 565511 29006
rect 30281 28930 30347 28933
rect 117957 28930 118023 28933
rect 539501 28932 539567 28933
rect 539501 28930 539548 28932
rect 30281 28928 118023 28930
rect 30281 28872 30286 28928
rect 30342 28872 117962 28928
rect 118018 28872 118023 28928
rect 30281 28870 118023 28872
rect 539456 28928 539548 28930
rect 539456 28872 539506 28928
rect 539456 28870 539548 28872
rect 30281 28867 30347 28870
rect 117957 28867 118023 28870
rect 539501 28868 539548 28870
rect 539612 28868 539618 28932
rect 539501 28867 539567 28868
rect 38510 28732 38516 28796
rect 38580 28794 38586 28796
rect 479241 28794 479307 28797
rect 38580 28792 479307 28794
rect 38580 28736 479246 28792
rect 479302 28736 479307 28792
rect 38580 28734 479307 28736
rect 38580 28732 38586 28734
rect 479241 28731 479307 28734
rect 487613 28794 487679 28797
rect 563094 28794 563100 28796
rect 487613 28792 563100 28794
rect 487613 28736 487618 28792
rect 487674 28736 563100 28792
rect 487613 28734 563100 28736
rect 487613 28731 487679 28734
rect 563094 28732 563100 28734
rect 563164 28732 563170 28796
rect 173985 28658 174051 28661
rect 561990 28658 561996 28660
rect 173985 28656 561996 28658
rect 173985 28600 173990 28656
rect 174046 28600 561996 28656
rect 173985 28598 561996 28600
rect 173985 28595 174051 28598
rect 561990 28596 561996 28598
rect 562060 28596 562066 28660
rect 58525 28522 58591 28525
rect 188797 28522 188863 28525
rect 58525 28520 188863 28522
rect 58525 28464 58530 28520
rect 58586 28464 188802 28520
rect 188858 28464 188863 28520
rect 58525 28462 188863 28464
rect 58525 28459 58591 28462
rect 188797 28459 188863 28462
rect 234521 28522 234587 28525
rect 527173 28522 527239 28525
rect 234521 28520 527239 28522
rect 234521 28464 234526 28520
rect 234582 28464 527178 28520
rect 527234 28464 527239 28520
rect 234521 28462 527239 28464
rect 234521 28459 234587 28462
rect 527173 28459 527239 28462
rect 528829 28522 528895 28525
rect 560702 28522 560708 28524
rect 528829 28520 560708 28522
rect 528829 28464 528834 28520
rect 528890 28464 560708 28520
rect 528829 28462 560708 28464
rect 528829 28459 528895 28462
rect 560702 28460 560708 28462
rect 560772 28460 560778 28524
rect 48814 28324 48820 28388
rect 48884 28386 48890 28388
rect 166901 28386 166967 28389
rect 48884 28384 166967 28386
rect 48884 28328 166906 28384
rect 166962 28328 166967 28384
rect 48884 28326 166967 28328
rect 48884 28324 48890 28326
rect 166901 28323 166967 28326
rect 333697 28386 333763 28389
rect 562593 28386 562659 28389
rect 333697 28384 562659 28386
rect 333697 28328 333702 28384
rect 333758 28328 562598 28384
rect 562654 28328 562659 28384
rect 333697 28326 562659 28328
rect 333697 28323 333763 28326
rect 562593 28323 562659 28326
rect 54518 28188 54524 28252
rect 54588 28250 54594 28252
rect 67633 28250 67699 28253
rect 54588 28248 67699 28250
rect 54588 28192 67638 28248
rect 67694 28192 67699 28248
rect 54588 28190 67699 28192
rect 54588 28188 54594 28190
rect 67633 28187 67699 28190
rect 69565 28250 69631 28253
rect 186221 28250 186287 28253
rect 69565 28248 186287 28250
rect 69565 28192 69570 28248
rect 69626 28192 186226 28248
rect 186282 28192 186287 28248
rect 69565 28190 186287 28192
rect 69565 28187 69631 28190
rect 186221 28187 186287 28190
rect 359457 28250 359523 28253
rect 559373 28250 559439 28253
rect 359457 28248 559439 28250
rect 359457 28192 359462 28248
rect 359518 28192 559378 28248
rect 559434 28192 559439 28248
rect 359457 28190 559439 28192
rect 359457 28187 359523 28190
rect 559373 28187 559439 28190
rect 99281 28114 99347 28117
rect 583109 28114 583175 28117
rect 99281 28112 583175 28114
rect 99281 28056 99286 28112
rect 99342 28056 583114 28112
rect 583170 28056 583175 28112
rect 99281 28054 583175 28056
rect 99281 28051 99347 28054
rect 583109 28051 583175 28054
rect 44030 27916 44036 27980
rect 44100 27978 44106 27980
rect 175273 27978 175339 27981
rect 44100 27976 175339 27978
rect 44100 27920 175278 27976
rect 175334 27920 175339 27976
rect 44100 27918 175339 27920
rect 44100 27916 44106 27918
rect 175273 27915 175339 27918
rect 536557 27978 536623 27981
rect 552422 27978 552428 27980
rect 536557 27976 552428 27978
rect 536557 27920 536562 27976
rect 536618 27920 552428 27976
rect 536557 27918 552428 27920
rect 536557 27915 536623 27918
rect 552422 27916 552428 27918
rect 552492 27916 552498 27980
rect 50654 27508 50660 27572
rect 50724 27570 50730 27572
rect 65793 27570 65859 27573
rect 50724 27568 65859 27570
rect 50724 27512 65798 27568
rect 65854 27512 65859 27568
rect 50724 27510 65859 27512
rect 50724 27508 50730 27510
rect 65793 27507 65859 27510
rect 71773 27570 71839 27573
rect 72877 27570 72943 27573
rect 71773 27568 72943 27570
rect 71773 27512 71778 27568
rect 71834 27512 72882 27568
rect 72938 27512 72943 27568
rect 71773 27510 72943 27512
rect 71773 27507 71839 27510
rect 72877 27507 72943 27510
rect 525609 27570 525675 27573
rect 575933 27570 575999 27573
rect 525609 27568 575999 27570
rect 525609 27512 525614 27568
rect 525670 27512 575938 27568
rect 575994 27512 575999 27568
rect 525609 27510 575999 27512
rect 525609 27507 525675 27510
rect 575933 27507 575999 27510
rect 65149 27434 65215 27437
rect 549662 27434 549668 27436
rect 65149 27432 549668 27434
rect 65149 27376 65154 27432
rect 65210 27376 549668 27432
rect 65149 27374 549668 27376
rect 65149 27371 65215 27374
rect 549662 27372 549668 27374
rect 549732 27372 549738 27436
rect 53230 27236 53236 27300
rect 53300 27298 53306 27300
rect 85757 27298 85823 27301
rect 53300 27296 85823 27298
rect 53300 27240 85762 27296
rect 85818 27240 85823 27296
rect 53300 27238 85823 27240
rect 53300 27236 53306 27238
rect 85757 27235 85823 27238
rect 532049 27298 532115 27301
rect 565118 27298 565124 27300
rect 532049 27296 565124 27298
rect 532049 27240 532054 27296
rect 532110 27240 565124 27296
rect 532049 27238 565124 27240
rect 532049 27235 532115 27238
rect 565118 27236 565124 27238
rect 565188 27236 565194 27300
rect 40902 27100 40908 27164
rect 40972 27162 40978 27164
rect 385217 27162 385283 27165
rect 40972 27160 385283 27162
rect 40972 27104 385222 27160
rect 385278 27104 385283 27160
rect 40972 27102 385283 27104
rect 40972 27100 40978 27102
rect 385217 27099 385283 27102
rect 421925 27162 421991 27165
rect 565302 27162 565308 27164
rect 421925 27160 565308 27162
rect 421925 27104 421930 27160
rect 421986 27104 565308 27160
rect 421925 27102 565308 27104
rect 421925 27099 421991 27102
rect 565302 27100 565308 27102
rect 565372 27100 565378 27164
rect 41638 26964 41644 27028
rect 41708 27026 41714 27028
rect 373625 27026 373691 27029
rect 41708 27024 373691 27026
rect 41708 26968 373630 27024
rect 373686 26968 373691 27024
rect 41708 26966 373691 26968
rect 41708 26964 41714 26966
rect 373625 26963 373691 26966
rect 452837 27026 452903 27029
rect 548006 27026 548012 27028
rect 452837 27024 548012 27026
rect 452837 26968 452842 27024
rect 452898 26968 548012 27024
rect 452837 26966 548012 26968
rect 452837 26963 452903 26966
rect 548006 26964 548012 26966
rect 548076 26964 548082 27028
rect 43846 26828 43852 26892
rect 43916 26890 43922 26892
rect 369117 26890 369183 26893
rect 43916 26888 369183 26890
rect 43916 26832 369122 26888
rect 369178 26832 369183 26888
rect 43916 26830 369183 26832
rect 43916 26828 43922 26830
rect 369117 26827 369183 26830
rect 41270 26692 41276 26756
rect 41340 26754 41346 26756
rect 71589 26754 71655 26757
rect 41340 26752 71655 26754
rect 41340 26696 71594 26752
rect 71650 26696 71655 26752
rect 41340 26694 71655 26696
rect 41340 26692 41346 26694
rect 71589 26691 71655 26694
rect 71773 26754 71839 26757
rect 542353 26754 542419 26757
rect 71773 26752 542419 26754
rect 71773 26696 71778 26752
rect 71834 26696 542358 26752
rect 542414 26696 542419 26752
rect 71773 26694 542419 26696
rect 71773 26691 71839 26694
rect 542353 26691 542419 26694
rect 31334 26556 31340 26620
rect 31404 26618 31410 26620
rect 524321 26618 524387 26621
rect 31404 26616 524387 26618
rect 31404 26560 524326 26616
rect 524382 26560 524387 26616
rect 31404 26558 524387 26560
rect 31404 26556 31410 26558
rect 524321 26555 524387 26558
rect 480253 26210 480319 26213
rect 556521 26210 556587 26213
rect 480253 26208 556587 26210
rect 480253 26152 480258 26208
rect 480314 26152 556526 26208
rect 556582 26152 556587 26208
rect 480253 26150 556587 26152
rect 480253 26147 480319 26150
rect 556521 26147 556587 26150
rect 47526 26012 47532 26076
rect 47596 26074 47602 26076
rect 367185 26074 367251 26077
rect 47596 26072 367251 26074
rect 47596 26016 367190 26072
rect 367246 26016 367251 26072
rect 47596 26014 367251 26016
rect 47596 26012 47602 26014
rect 367185 26011 367251 26014
rect 378225 26074 378291 26077
rect 577037 26074 577103 26077
rect 378225 26072 577103 26074
rect 378225 26016 378230 26072
rect 378286 26016 577042 26072
rect 577098 26016 577103 26072
rect 378225 26014 577103 26016
rect 378225 26011 378291 26014
rect 577037 26011 577103 26014
rect 54886 25876 54892 25940
rect 54956 25938 54962 25940
rect 70393 25938 70459 25941
rect 54956 25936 70459 25938
rect 54956 25880 70398 25936
rect 70454 25880 70459 25936
rect 54956 25878 70459 25880
rect 54956 25876 54962 25878
rect 70393 25875 70459 25878
rect 354765 25938 354831 25941
rect 579613 25938 579679 25941
rect 354765 25936 579679 25938
rect 354765 25880 354770 25936
rect 354826 25880 579618 25936
rect 579674 25880 579679 25936
rect 354765 25878 579679 25880
rect 354765 25875 354831 25878
rect 579613 25875 579679 25878
rect 53414 25740 53420 25804
rect 53484 25802 53490 25804
rect 74533 25802 74599 25805
rect 53484 25800 74599 25802
rect 53484 25744 74538 25800
rect 74594 25744 74599 25800
rect 53484 25742 74599 25744
rect 53484 25740 53490 25742
rect 74533 25739 74599 25742
rect 385033 25802 385099 25805
rect 575606 25802 575612 25804
rect 385033 25800 575612 25802
rect 385033 25744 385038 25800
rect 385094 25744 575612 25800
rect 385033 25742 575612 25744
rect 385033 25739 385099 25742
rect 575606 25740 575612 25742
rect 575676 25740 575682 25804
rect 52126 25604 52132 25668
rect 52196 25666 52202 25668
rect 85573 25666 85639 25669
rect 52196 25664 85639 25666
rect 52196 25608 85578 25664
rect 85634 25608 85639 25664
rect 52196 25606 85639 25608
rect 52196 25604 52202 25606
rect 85573 25603 85639 25606
rect 231853 25666 231919 25669
rect 566958 25666 566964 25668
rect 231853 25664 566964 25666
rect 231853 25608 231858 25664
rect 231914 25608 566964 25664
rect 231853 25606 566964 25608
rect 231853 25603 231919 25606
rect 566958 25604 566964 25606
rect 567028 25604 567034 25668
rect 54702 25468 54708 25532
rect 54772 25530 54778 25532
rect 88333 25530 88399 25533
rect 54772 25528 88399 25530
rect 54772 25472 88338 25528
rect 88394 25472 88399 25528
rect 54772 25470 88399 25472
rect 54772 25468 54778 25470
rect 88333 25467 88399 25470
rect 184933 25530 184999 25533
rect 553577 25530 553643 25533
rect 184933 25528 553643 25530
rect 184933 25472 184938 25528
rect 184994 25472 553582 25528
rect 553638 25472 553643 25528
rect 184933 25470 553643 25472
rect 184933 25467 184999 25470
rect 553577 25467 553643 25470
rect 32990 25332 32996 25396
rect 33060 25394 33066 25396
rect 484577 25394 484643 25397
rect 33060 25392 484643 25394
rect 33060 25336 484582 25392
rect 484638 25336 484643 25392
rect 33060 25334 484643 25336
rect 33060 25332 33066 25334
rect 484577 25331 484643 25334
rect 52310 24788 52316 24852
rect 52380 24850 52386 24852
rect 91185 24850 91251 24853
rect 52380 24848 91251 24850
rect 52380 24792 91190 24848
rect 91246 24792 91251 24848
rect 52380 24790 91251 24792
rect 52380 24788 52386 24790
rect 91185 24787 91251 24790
rect 44766 24652 44772 24716
rect 44836 24714 44842 24716
rect 255313 24714 255379 24717
rect 44836 24712 255379 24714
rect 44836 24656 255318 24712
rect 255374 24656 255379 24712
rect 44836 24654 255379 24656
rect 44836 24652 44842 24654
rect 255313 24651 255379 24654
rect 274633 24714 274699 24717
rect 565486 24714 565492 24716
rect 274633 24712 565492 24714
rect 274633 24656 274638 24712
rect 274694 24656 565492 24712
rect 274633 24654 565492 24656
rect 274633 24651 274699 24654
rect 565486 24652 565492 24654
rect 565556 24652 565562 24716
rect 304993 24578 305059 24581
rect 563278 24578 563284 24580
rect 304993 24576 563284 24578
rect 304993 24520 304998 24576
rect 305054 24520 563284 24576
rect 304993 24518 563284 24520
rect 304993 24515 305059 24518
rect 563278 24516 563284 24518
rect 563348 24516 563354 24580
rect 50470 24380 50476 24444
rect 50540 24442 50546 24444
rect 77385 24442 77451 24445
rect 50540 24440 77451 24442
rect 50540 24384 77390 24440
rect 77446 24384 77451 24440
rect 50540 24382 77451 24384
rect 50540 24380 50546 24382
rect 77385 24379 77451 24382
rect 224953 24442 225019 24445
rect 567326 24442 567332 24444
rect 224953 24440 567332 24442
rect 224953 24384 224958 24440
rect 225014 24384 567332 24440
rect 224953 24382 567332 24384
rect 224953 24379 225019 24382
rect 567326 24380 567332 24382
rect 567396 24380 567402 24444
rect 207105 24306 207171 24309
rect 567510 24306 567516 24308
rect 207105 24304 567516 24306
rect 207105 24248 207110 24304
rect 207166 24248 567516 24304
rect 207105 24246 567516 24248
rect 207105 24243 207171 24246
rect 567510 24244 567516 24246
rect 567580 24244 567586 24308
rect 164233 24170 164299 24173
rect 568614 24170 568620 24172
rect 164233 24168 568620 24170
rect 164233 24112 164238 24168
rect 164294 24112 568620 24168
rect 164233 24110 568620 24112
rect 164233 24107 164299 24110
rect 568614 24108 568620 24110
rect 568684 24108 568690 24172
rect 44582 23972 44588 24036
rect 44652 24034 44658 24036
rect 303613 24034 303679 24037
rect 44652 24032 303679 24034
rect 44652 23976 303618 24032
rect 303674 23976 303679 24032
rect 44652 23974 303679 23976
rect 44652 23972 44658 23974
rect 303613 23971 303679 23974
rect 347865 24034 347931 24037
rect 565854 24034 565860 24036
rect 347865 24032 565860 24034
rect 347865 23976 347870 24032
rect 347926 23976 565860 24032
rect 347865 23974 565860 23976
rect 347865 23971 347931 23974
rect 565854 23972 565860 23974
rect 565924 23972 565930 24036
rect 578233 24034 578299 24037
rect 578734 24034 578740 24036
rect 578233 24032 578740 24034
rect 578233 23976 578238 24032
rect 578294 23976 578740 24032
rect 578233 23974 578740 23976
rect 578233 23971 578299 23974
rect 578734 23972 578740 23974
rect 578804 23972 578810 24036
rect 36854 23836 36860 23900
rect 36924 23898 36930 23900
rect 321553 23898 321619 23901
rect 36924 23896 321619 23898
rect 36924 23840 321558 23896
rect 321614 23840 321619 23896
rect 36924 23838 321619 23840
rect 36924 23836 36930 23838
rect 321553 23835 321619 23838
rect 165613 23762 165679 23765
rect 578550 23762 578556 23764
rect 165613 23760 578556 23762
rect 165613 23704 165618 23760
rect 165674 23704 578556 23760
rect 165613 23702 578556 23704
rect 165613 23699 165679 23702
rect 578550 23700 578556 23702
rect 578620 23700 578626 23764
rect 22001 23354 22067 23357
rect 468937 23354 469003 23357
rect 22001 23352 469003 23354
rect 22001 23296 22006 23352
rect 22062 23296 468942 23352
rect 468998 23296 469003 23352
rect 22001 23294 469003 23296
rect 22001 23291 22067 23294
rect 468937 23291 469003 23294
rect 518893 23354 518959 23357
rect 547638 23354 547644 23356
rect 518893 23352 547644 23354
rect 518893 23296 518898 23352
rect 518954 23296 547644 23352
rect 518893 23294 547644 23296
rect 518893 23291 518959 23294
rect 547638 23292 547644 23294
rect 547708 23292 547714 23356
rect 48078 23156 48084 23220
rect 48148 23218 48154 23220
rect 107745 23218 107811 23221
rect 48148 23216 107811 23218
rect 48148 23160 107750 23216
rect 107806 23160 107811 23216
rect 48148 23158 107811 23160
rect 48148 23156 48154 23158
rect 107745 23155 107811 23158
rect 107929 23218 107995 23221
rect 542854 23218 542860 23220
rect 107929 23216 542860 23218
rect 107929 23160 107934 23216
rect 107990 23160 542860 23216
rect 107929 23158 542860 23160
rect 107929 23155 107995 23158
rect 542854 23156 542860 23158
rect 542924 23156 542930 23220
rect 35750 23020 35756 23084
rect 35820 23082 35826 23084
rect 408493 23082 408559 23085
rect 35820 23080 408559 23082
rect 35820 23024 408498 23080
rect 408554 23024 408559 23080
rect 35820 23022 408559 23024
rect 35820 23020 35826 23022
rect 408493 23019 408559 23022
rect 444465 23082 444531 23085
rect 544510 23082 544516 23084
rect 444465 23080 544516 23082
rect 444465 23024 444470 23080
rect 444526 23024 544516 23080
rect 444465 23022 544516 23024
rect 444465 23019 444531 23022
rect 544510 23020 544516 23022
rect 544580 23020 544586 23084
rect 37038 22884 37044 22948
rect 37108 22946 37114 22948
rect 318885 22946 318951 22949
rect 37108 22944 318951 22946
rect 37108 22888 318890 22944
rect 318946 22888 318951 22944
rect 37108 22886 318951 22888
rect 37108 22884 37114 22886
rect 318885 22883 318951 22886
rect 358813 22946 358879 22949
rect 560518 22946 560524 22948
rect 358813 22944 560524 22946
rect 358813 22888 358818 22944
rect 358874 22888 560524 22944
rect 358813 22886 560524 22888
rect 358813 22883 358879 22886
rect 560518 22884 560524 22886
rect 560588 22884 560594 22948
rect 391933 22810 391999 22813
rect 545062 22810 545068 22812
rect 391933 22808 545068 22810
rect 391933 22752 391938 22808
rect 391994 22752 545068 22808
rect 391933 22750 545068 22752
rect 391933 22747 391999 22750
rect 545062 22748 545068 22750
rect 545132 22748 545138 22812
rect 49550 22612 49556 22676
rect 49620 22674 49626 22676
rect 124213 22674 124279 22677
rect 49620 22672 124279 22674
rect 49620 22616 124218 22672
rect 124274 22616 124279 22672
rect 49620 22614 124279 22616
rect 49620 22612 49626 22614
rect 124213 22611 124279 22614
rect 178033 22674 178099 22677
rect 553526 22674 553532 22676
rect 178033 22672 553532 22674
rect 178033 22616 178038 22672
rect 178094 22616 553532 22672
rect 178033 22614 553532 22616
rect 178033 22611 178099 22614
rect 553526 22612 553532 22614
rect 553596 22612 553602 22676
rect 491293 22538 491359 22541
rect 553894 22538 553900 22540
rect 491293 22536 553900 22538
rect 491293 22480 491298 22536
rect 491354 22480 553900 22536
rect 491293 22478 553900 22480
rect 491293 22475 491359 22478
rect 553894 22476 553900 22478
rect 553964 22476 553970 22540
rect 59670 21932 59676 21996
rect 59740 21994 59746 21996
rect 74625 21994 74691 21997
rect 59740 21992 74691 21994
rect 59740 21936 74630 21992
rect 74686 21936 74691 21992
rect 59740 21934 74691 21936
rect 59740 21932 59746 21934
rect 74625 21931 74691 21934
rect 528553 21994 528619 21997
rect 538990 21994 538996 21996
rect 528553 21992 538996 21994
rect 528553 21936 528558 21992
rect 528614 21936 538996 21992
rect 528553 21934 538996 21936
rect 528553 21931 528619 21934
rect 538990 21932 538996 21934
rect 539060 21932 539066 21996
rect 46422 21796 46428 21860
rect 46492 21858 46498 21860
rect 318793 21858 318859 21861
rect 46492 21856 318859 21858
rect 46492 21800 318798 21856
rect 318854 21800 318859 21856
rect 46492 21798 318859 21800
rect 46492 21796 46498 21798
rect 318793 21795 318859 21798
rect 463785 21858 463851 21861
rect 540094 21858 540100 21860
rect 463785 21856 540100 21858
rect 463785 21800 463790 21856
rect 463846 21800 540100 21856
rect 463785 21798 540100 21800
rect 463785 21795 463851 21798
rect 540094 21796 540100 21798
rect 540164 21796 540170 21860
rect 58566 21660 58572 21724
rect 58636 21722 58642 21724
rect 207013 21722 207079 21725
rect 58636 21720 207079 21722
rect 58636 21664 207018 21720
rect 207074 21664 207079 21720
rect 58636 21662 207079 21664
rect 58636 21660 58642 21662
rect 207013 21659 207079 21662
rect 476113 21722 476179 21725
rect 544326 21722 544332 21724
rect 476113 21720 544332 21722
rect 476113 21664 476118 21720
rect 476174 21664 544332 21720
rect 476113 21662 544332 21664
rect 476113 21659 476179 21662
rect 544326 21660 544332 21662
rect 544396 21660 544402 21724
rect 55438 21524 55444 21588
rect 55508 21586 55514 21588
rect 125685 21586 125751 21589
rect 55508 21584 125751 21586
rect 55508 21528 125690 21584
rect 125746 21528 125751 21584
rect 55508 21526 125751 21528
rect 55508 21524 55514 21526
rect 125685 21523 125751 21526
rect 183553 21586 183619 21589
rect 547086 21586 547092 21588
rect 183553 21584 547092 21586
rect 183553 21528 183558 21584
rect 183614 21528 547092 21584
rect 183553 21526 547092 21528
rect 183553 21523 183619 21526
rect 547086 21524 547092 21526
rect 547156 21524 547162 21588
rect 146385 21450 146451 21453
rect 567694 21450 567700 21452
rect 146385 21448 567700 21450
rect 146385 21392 146390 21448
rect 146446 21392 567700 21448
rect 146385 21390 567700 21392
rect 146385 21387 146451 21390
rect 567694 21388 567700 21390
rect 567764 21388 567770 21452
rect 128353 21314 128419 21317
rect 553710 21314 553716 21316
rect 128353 21312 553716 21314
rect 128353 21256 128358 21312
rect 128414 21256 553716 21312
rect 128353 21254 553716 21256
rect 128353 21251 128419 21254
rect 553710 21252 553716 21254
rect 553780 21252 553786 21316
rect 50286 21116 50292 21180
rect 50356 21178 50362 21180
rect 459645 21178 459711 21181
rect 50356 21176 459711 21178
rect 50356 21120 459650 21176
rect 459706 21120 459711 21176
rect 50356 21118 459711 21120
rect 50356 21116 50362 21118
rect 459645 21115 459711 21118
rect 484393 21178 484459 21181
rect 563646 21178 563652 21180
rect 484393 21176 563652 21178
rect 484393 21120 484398 21176
rect 484454 21120 563652 21176
rect 484393 21118 563652 21120
rect 484393 21115 484459 21118
rect 563646 21116 563652 21118
rect 563716 21116 563722 21180
rect 560293 20906 560359 20909
rect 561438 20906 561444 20908
rect 560293 20904 561444 20906
rect 560293 20848 560298 20904
rect 560354 20848 561444 20904
rect 560293 20846 561444 20848
rect 560293 20843 560359 20846
rect 561438 20844 561444 20846
rect 561508 20844 561514 20908
rect 569953 20906 570019 20909
rect 570270 20906 570276 20908
rect 569953 20904 570276 20906
rect 569953 20848 569958 20904
rect 570014 20848 570276 20904
rect 569953 20846 570276 20848
rect 569953 20843 570019 20846
rect 570270 20844 570276 20846
rect 570340 20844 570346 20908
rect 571425 20770 571491 20773
rect 571558 20770 571564 20772
rect 571425 20768 571564 20770
rect 571425 20712 571430 20768
rect 571486 20712 571564 20768
rect 571425 20710 571564 20712
rect 571425 20707 571491 20710
rect 571558 20708 571564 20710
rect 571628 20708 571634 20772
rect 32673 20634 32739 20637
rect 538305 20634 538371 20637
rect 32673 20632 538371 20634
rect 32673 20576 32678 20632
rect 32734 20576 538310 20632
rect 538366 20576 538371 20632
rect 32673 20574 538371 20576
rect 32673 20571 32739 20574
rect 538305 20571 538371 20574
rect 20529 20498 20595 20501
rect 525793 20498 525859 20501
rect 20529 20496 525859 20498
rect 20529 20440 20534 20496
rect 20590 20440 525798 20496
rect 525854 20440 525859 20496
rect 20529 20438 525859 20440
rect 20529 20435 20595 20438
rect 525793 20435 525859 20438
rect 436093 20362 436159 20365
rect 573357 20362 573423 20365
rect 436093 20360 573423 20362
rect 436093 20304 436098 20360
rect 436154 20304 573362 20360
rect 573418 20304 573423 20360
rect 436093 20302 573423 20304
rect 436093 20299 436159 20302
rect 573357 20299 573423 20302
rect 324313 20226 324379 20229
rect 543038 20226 543044 20228
rect 324313 20224 543044 20226
rect 324313 20168 324318 20224
rect 324374 20168 543044 20224
rect 324313 20166 543044 20168
rect 324313 20163 324379 20166
rect 543038 20164 543044 20166
rect 543108 20164 543114 20228
rect 60038 20028 60044 20092
rect 60108 20090 60114 20092
rect 139393 20090 139459 20093
rect 60108 20088 139459 20090
rect 60108 20032 139398 20088
rect 139454 20032 139459 20088
rect 60108 20030 139459 20032
rect 60108 20028 60114 20030
rect 139393 20027 139459 20030
rect 310513 20090 310579 20093
rect 561070 20090 561076 20092
rect 310513 20088 561076 20090
rect 310513 20032 310518 20088
rect 310574 20032 561076 20088
rect 310513 20030 561076 20032
rect 310513 20027 310579 20030
rect 561070 20028 561076 20030
rect 561140 20028 561146 20092
rect 99373 19954 99439 19957
rect 559230 19954 559236 19956
rect 99373 19952 559236 19954
rect 99373 19896 99378 19952
rect 99434 19896 559236 19952
rect 99373 19894 559236 19896
rect 99373 19891 99439 19894
rect 559230 19892 559236 19894
rect 559300 19892 559306 19956
rect 17861 19818 17927 19821
rect 445845 19818 445911 19821
rect 556286 19818 556292 19820
rect 17861 19816 431970 19818
rect 17861 19760 17866 19816
rect 17922 19760 431970 19816
rect 17861 19758 431970 19760
rect 17861 19755 17927 19758
rect 431910 19682 431970 19758
rect 445845 19816 556292 19818
rect 445845 19760 445850 19816
rect 445906 19760 556292 19816
rect 445845 19758 556292 19760
rect 445845 19755 445911 19758
rect 556286 19756 556292 19758
rect 556356 19756 556362 19820
rect 578877 19818 578943 19821
rect 583520 19818 584960 19908
rect 578877 19816 584960 19818
rect 578877 19760 578882 19816
rect 578938 19760 584960 19816
rect 578877 19758 584960 19760
rect 578877 19755 578943 19758
rect 446029 19682 446095 19685
rect 431910 19680 446095 19682
rect 431910 19624 446034 19680
rect 446090 19624 446095 19680
rect 583520 19668 584960 19758
rect 431910 19622 446095 19624
rect 446029 19619 446095 19622
rect -960 19410 480 19500
rect 28206 19410 28212 19412
rect -960 19350 28212 19410
rect -960 19260 480 19350
rect 28206 19348 28212 19350
rect 28276 19348 28282 19412
rect 50797 19274 50863 19277
rect 367093 19274 367159 19277
rect 50797 19272 367159 19274
rect 50797 19216 50802 19272
rect 50858 19216 367098 19272
rect 367154 19216 367159 19272
rect 50797 19214 367159 19216
rect 50797 19211 50863 19214
rect 367093 19211 367159 19214
rect 57605 19138 57671 19141
rect 168373 19138 168439 19141
rect 57605 19136 168439 19138
rect 57605 19080 57610 19136
rect 57666 19080 168378 19136
rect 168434 19080 168439 19136
rect 57605 19078 168439 19080
rect 57605 19075 57671 19078
rect 168373 19075 168439 19078
rect 289813 19138 289879 19141
rect 572662 19138 572668 19140
rect 289813 19136 572668 19138
rect 289813 19080 289818 19136
rect 289874 19080 572668 19136
rect 289813 19078 572668 19080
rect 289813 19075 289879 19078
rect 572662 19076 572668 19078
rect 572732 19076 572738 19140
rect 19241 19002 19307 19005
rect 95417 19002 95483 19005
rect 19241 19000 95483 19002
rect 19241 18944 19246 19000
rect 19302 18944 95422 19000
rect 95478 18944 95483 19000
rect 19241 18942 95483 18944
rect 19241 18939 19307 18942
rect 95417 18939 95483 18942
rect 260833 19002 260899 19005
rect 554814 19002 554820 19004
rect 260833 19000 554820 19002
rect 260833 18944 260838 19000
rect 260894 18944 554820 19000
rect 260833 18942 554820 18944
rect 260833 18939 260899 18942
rect 554814 18940 554820 18942
rect 554884 18940 554890 19004
rect 278773 18866 278839 18869
rect 574134 18866 574140 18868
rect 278773 18864 574140 18866
rect 278773 18808 278778 18864
rect 278834 18808 574140 18864
rect 278773 18806 574140 18808
rect 278773 18803 278839 18806
rect 574134 18804 574140 18806
rect 574204 18804 574210 18868
rect 113173 18730 113239 18733
rect 549478 18730 549484 18732
rect 113173 18728 549484 18730
rect 113173 18672 113178 18728
rect 113234 18672 549484 18728
rect 113173 18670 549484 18672
rect 113173 18667 113239 18670
rect 549478 18668 549484 18670
rect 549548 18668 549554 18732
rect 106273 18594 106339 18597
rect 576894 18594 576900 18596
rect 106273 18592 576900 18594
rect 106273 18536 106278 18592
rect 106334 18536 576900 18592
rect 106273 18534 576900 18536
rect 106273 18531 106339 18534
rect 576894 18532 576900 18534
rect 576964 18532 576970 18596
rect 58934 18396 58940 18460
rect 59004 18458 59010 18460
rect 329833 18458 329899 18461
rect 59004 18456 329899 18458
rect 59004 18400 329838 18456
rect 329894 18400 329899 18456
rect 59004 18398 329899 18400
rect 59004 18396 59010 18398
rect 329833 18395 329899 18398
rect 335353 18458 335419 18461
rect 557574 18458 557580 18460
rect 335353 18456 557580 18458
rect 335353 18400 335358 18456
rect 335414 18400 557580 18456
rect 335353 18398 557580 18400
rect 335353 18395 335419 18398
rect 557574 18396 557580 18398
rect 557644 18396 557650 18460
rect 84193 17914 84259 17917
rect 572253 17914 572319 17917
rect 84193 17912 572319 17914
rect 84193 17856 84198 17912
rect 84254 17856 572258 17912
rect 572314 17856 572319 17912
rect 84193 17854 572319 17856
rect 84193 17851 84259 17854
rect 572253 17851 572319 17854
rect 106365 17778 106431 17781
rect 579838 17778 579844 17780
rect 106365 17776 579844 17778
rect 106365 17720 106370 17776
rect 106426 17720 579844 17776
rect 106365 17718 579844 17720
rect 106365 17715 106431 17718
rect 579838 17716 579844 17718
rect 579908 17716 579914 17780
rect 178125 17642 178191 17645
rect 580942 17642 580948 17644
rect 178125 17640 580948 17642
rect 178125 17584 178130 17640
rect 178186 17584 580948 17640
rect 178125 17582 580948 17584
rect 178125 17579 178191 17582
rect 580942 17580 580948 17582
rect 581012 17580 581018 17644
rect 35249 17506 35315 17509
rect 153193 17506 153259 17509
rect 35249 17504 153259 17506
rect 35249 17448 35254 17504
rect 35310 17448 153198 17504
rect 153254 17448 153259 17504
rect 35249 17446 153259 17448
rect 35249 17443 35315 17446
rect 153193 17443 153259 17446
rect 212625 17506 212691 17509
rect 545614 17506 545620 17508
rect 212625 17504 545620 17506
rect 212625 17448 212630 17504
rect 212686 17448 545620 17504
rect 212625 17446 545620 17448
rect 212625 17443 212691 17446
rect 545614 17444 545620 17446
rect 545684 17444 545690 17508
rect 58617 17370 58683 17373
rect 222193 17370 222259 17373
rect 58617 17368 222259 17370
rect 58617 17312 58622 17368
rect 58678 17312 222198 17368
rect 222254 17312 222259 17368
rect 58617 17310 222259 17312
rect 58617 17307 58683 17310
rect 222193 17307 222259 17310
rect 282913 17370 282979 17373
rect 570086 17370 570092 17372
rect 282913 17368 570092 17370
rect 282913 17312 282918 17368
rect 282974 17312 570092 17368
rect 282913 17310 570092 17312
rect 282913 17307 282979 17310
rect 570086 17308 570092 17310
rect 570156 17308 570162 17372
rect 136633 17234 136699 17237
rect 556470 17234 556476 17236
rect 136633 17232 556476 17234
rect 136633 17176 136638 17232
rect 136694 17176 556476 17232
rect 136633 17174 556476 17176
rect 136633 17171 136699 17174
rect 556470 17172 556476 17174
rect 556540 17172 556546 17236
rect 24761 17098 24827 17101
rect 180793 17098 180859 17101
rect 24761 17096 180859 17098
rect 24761 17040 24766 17096
rect 24822 17040 180798 17096
rect 180854 17040 180859 17096
rect 24761 17038 180859 17040
rect 24761 17035 24827 17038
rect 180793 17035 180859 17038
rect 242985 16554 243051 16557
rect 541382 16554 541388 16556
rect 242985 16552 541388 16554
rect 242985 16496 242990 16552
rect 243046 16496 541388 16552
rect 242985 16494 541388 16496
rect 242985 16491 243051 16494
rect 541382 16492 541388 16494
rect 541452 16492 541458 16556
rect 431953 16418 432019 16421
rect 543222 16418 543228 16420
rect 431953 16416 543228 16418
rect 431953 16360 431958 16416
rect 432014 16360 543228 16416
rect 431953 16358 543228 16360
rect 431953 16355 432019 16358
rect 543222 16356 543228 16358
rect 543292 16356 543298 16420
rect 378409 16146 378475 16149
rect 545246 16146 545252 16148
rect 378409 16144 545252 16146
rect 378409 16088 378414 16144
rect 378470 16088 545252 16144
rect 378409 16086 545252 16088
rect 378409 16083 378475 16086
rect 545246 16084 545252 16086
rect 545316 16084 545322 16148
rect 144729 16010 144795 16013
rect 558126 16010 558132 16012
rect 144729 16008 558132 16010
rect 144729 15952 144734 16008
rect 144790 15952 558132 16008
rect 144729 15950 558132 15952
rect 144729 15947 144795 15950
rect 558126 15948 558132 15950
rect 558196 15948 558202 16012
rect 92473 15874 92539 15877
rect 548374 15874 548380 15876
rect 92473 15872 548380 15874
rect 92473 15816 92478 15872
rect 92534 15816 548380 15872
rect 92473 15814 548380 15816
rect 92473 15811 92539 15814
rect 548374 15812 548380 15814
rect 548444 15812 548450 15876
rect 251173 15058 251239 15061
rect 547270 15058 547276 15060
rect 251173 15056 547276 15058
rect 251173 15000 251178 15056
rect 251234 15000 547276 15056
rect 251173 14998 547276 15000
rect 251173 14995 251239 14998
rect 547270 14996 547276 14998
rect 547340 14996 547346 15060
rect 203425 14922 203491 14925
rect 540278 14922 540284 14924
rect 203425 14920 540284 14922
rect 203425 14864 203430 14920
rect 203486 14864 540284 14920
rect 203425 14862 540284 14864
rect 203425 14859 203491 14862
rect 540278 14860 540284 14862
rect 540348 14860 540354 14924
rect 226333 14786 226399 14789
rect 569902 14786 569908 14788
rect 226333 14784 569908 14786
rect 226333 14728 226338 14784
rect 226394 14728 569908 14784
rect 226333 14726 569908 14728
rect 226333 14723 226399 14726
rect 569902 14724 569908 14726
rect 569972 14724 569978 14788
rect 214465 14650 214531 14653
rect 579654 14650 579660 14652
rect 214465 14648 579660 14650
rect 214465 14592 214470 14648
rect 214526 14592 579660 14648
rect 214465 14590 579660 14592
rect 214465 14587 214531 14590
rect 579654 14588 579660 14590
rect 579724 14588 579730 14652
rect 46657 14514 46723 14517
rect 557942 14514 557948 14516
rect 46657 14512 557948 14514
rect 46657 14456 46662 14512
rect 46718 14456 557948 14512
rect 46657 14454 557948 14456
rect 46657 14451 46723 14454
rect 557942 14452 557948 14454
rect 558012 14452 558018 14516
rect 231945 13698 232011 13701
rect 549897 13698 549963 13701
rect 231945 13696 549963 13698
rect 231945 13640 231950 13696
rect 232006 13640 549902 13696
rect 549958 13640 549963 13696
rect 231945 13638 549963 13640
rect 231945 13635 232011 13638
rect 549897 13635 549963 13638
rect 303889 13154 303955 13157
rect 557625 13154 557691 13157
rect 303889 13152 557691 13154
rect 303889 13096 303894 13152
rect 303950 13096 557630 13152
rect 557686 13096 557691 13152
rect 303889 13094 557691 13096
rect 303889 13091 303955 13094
rect 557625 13091 557691 13094
rect 208577 13018 208643 13021
rect 555049 13018 555115 13021
rect 208577 13016 555115 13018
rect 208577 12960 208582 13016
rect 208638 12960 555054 13016
rect 555110 12960 555115 13016
rect 208577 12958 555115 12960
rect 208577 12955 208643 12958
rect 555049 12955 555115 12958
rect 328729 12066 328795 12069
rect 557758 12066 557764 12068
rect 328729 12064 557764 12066
rect 328729 12008 328734 12064
rect 328790 12008 557764 12064
rect 328729 12006 557764 12008
rect 328729 12003 328795 12006
rect 557758 12004 557764 12006
rect 557828 12004 557834 12068
rect 242893 11930 242959 11933
rect 553342 11930 553348 11932
rect 242893 11928 553348 11930
rect 242893 11872 242898 11928
rect 242954 11872 553348 11928
rect 242893 11870 553348 11872
rect 242893 11867 242959 11870
rect 553342 11868 553348 11870
rect 553412 11868 553418 11932
rect 222745 11794 222811 11797
rect 541014 11794 541020 11796
rect 222745 11792 541020 11794
rect 222745 11736 222750 11792
rect 222806 11736 541020 11792
rect 222745 11734 541020 11736
rect 222745 11731 222811 11734
rect 541014 11732 541020 11734
rect 541084 11732 541090 11796
rect 218053 11658 218119 11661
rect 556102 11658 556108 11660
rect 218053 11656 556108 11658
rect 218053 11600 218058 11656
rect 218114 11600 556108 11656
rect 218053 11598 556108 11600
rect 218053 11595 218119 11598
rect 556102 11596 556108 11598
rect 556172 11596 556178 11660
rect 276013 10978 276079 10981
rect 538806 10978 538812 10980
rect 276013 10976 538812 10978
rect 276013 10920 276018 10976
rect 276074 10920 538812 10976
rect 276013 10918 538812 10920
rect 276013 10915 276079 10918
rect 538806 10916 538812 10918
rect 538876 10916 538882 10980
rect 205081 10298 205147 10301
rect 556654 10298 556660 10300
rect 205081 10296 556660 10298
rect 205081 10240 205086 10296
rect 205142 10240 556660 10296
rect 205081 10238 556660 10240
rect 205081 10235 205147 10238
rect 556654 10236 556660 10238
rect 556724 10236 556730 10300
rect 1669 7578 1735 7581
rect 554998 7578 555004 7580
rect 1669 7576 555004 7578
rect 1669 7520 1674 7576
rect 1730 7520 555004 7576
rect 1669 7518 555004 7520
rect 1669 7515 1735 7518
rect 554998 7516 555004 7518
rect 555068 7516 555074 7580
rect 474549 6626 474615 6629
rect 541566 6626 541572 6628
rect 474549 6624 541572 6626
rect -960 6490 480 6580
rect 474549 6568 474554 6624
rect 474610 6568 541572 6624
rect 474549 6566 541572 6568
rect 474549 6563 474615 6566
rect 541566 6564 541572 6566
rect 541636 6564 541642 6628
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 481725 6490 481791 6493
rect 563462 6490 563468 6492
rect 481725 6488 563468 6490
rect 481725 6432 481730 6488
rect 481786 6432 563468 6488
rect 481725 6430 563468 6432
rect 481725 6427 481791 6430
rect 563462 6428 563468 6430
rect 563532 6428 563538 6492
rect 583520 6476 584960 6716
rect 240501 6354 240567 6357
rect 550582 6354 550588 6356
rect 240501 6352 550588 6354
rect 240501 6296 240506 6352
rect 240562 6296 550588 6352
rect 240501 6294 550588 6296
rect 240501 6291 240567 6294
rect 550582 6292 550588 6294
rect 550652 6292 550658 6356
rect 19425 6218 19491 6221
rect 559046 6218 559052 6220
rect 19425 6216 559052 6218
rect 19425 6160 19430 6216
rect 19486 6160 559052 6216
rect 19425 6158 559052 6160
rect 19425 6155 19491 6158
rect 559046 6156 559052 6158
rect 559116 6156 559122 6220
rect 155401 4994 155467 4997
rect 558862 4994 558868 4996
rect 155401 4992 558868 4994
rect 155401 4936 155406 4992
rect 155462 4936 558868 4992
rect 155401 4934 558868 4936
rect 155401 4931 155467 4934
rect 558862 4932 558868 4934
rect 558932 4932 558938 4996
rect 64321 4858 64387 4861
rect 550214 4858 550220 4860
rect 64321 4856 550220 4858
rect 64321 4800 64326 4856
rect 64382 4800 550220 4856
rect 64321 4798 550220 4800
rect 64321 4795 64387 4798
rect 550214 4796 550220 4798
rect 550284 4796 550290 4860
rect 53598 3980 53604 4044
rect 53668 4042 53674 4044
rect 197905 4042 197971 4045
rect 53668 4040 197971 4042
rect 53668 3984 197910 4040
rect 197966 3984 197971 4040
rect 53668 3982 197971 3984
rect 53668 3980 53674 3982
rect 197905 3979 197971 3982
rect 549069 4042 549135 4045
rect 571333 4042 571399 4045
rect 549069 4040 571399 4042
rect 549069 3984 549074 4040
rect 549130 3984 571338 4040
rect 571394 3984 571399 4040
rect 549069 3982 571399 3984
rect 549069 3979 549135 3982
rect 571333 3979 571399 3982
rect 55622 3844 55628 3908
rect 55692 3906 55698 3908
rect 200297 3906 200363 3909
rect 55692 3904 200363 3906
rect 55692 3848 200302 3904
rect 200358 3848 200363 3904
rect 55692 3846 200363 3848
rect 55692 3844 55698 3846
rect 200297 3843 200363 3846
rect 531313 3906 531379 3909
rect 566222 3906 566228 3908
rect 531313 3904 566228 3906
rect 531313 3848 531318 3904
rect 531374 3848 566228 3904
rect 531313 3846 566228 3848
rect 531313 3843 531379 3846
rect 566222 3844 566228 3846
rect 566292 3844 566298 3908
rect 169569 3770 169635 3773
rect 574318 3770 574324 3772
rect 169569 3768 574324 3770
rect 169569 3712 169574 3768
rect 169630 3712 574324 3768
rect 169569 3710 574324 3712
rect 169569 3707 169635 3710
rect 574318 3708 574324 3710
rect 574388 3708 574394 3772
rect 157793 3634 157859 3637
rect 575422 3634 575428 3636
rect 157793 3632 575428 3634
rect 157793 3576 157798 3632
rect 157854 3576 575428 3632
rect 157793 3574 575428 3576
rect 157793 3571 157859 3574
rect 575422 3572 575428 3574
rect 575492 3572 575498 3636
rect 24209 3498 24275 3501
rect 25446 3498 25452 3500
rect 24209 3496 25452 3498
rect 24209 3440 24214 3496
rect 24270 3440 25452 3496
rect 24209 3438 25452 3440
rect 24209 3435 24275 3438
rect 25446 3436 25452 3438
rect 25516 3436 25522 3500
rect 43069 3498 43135 3501
rect 43662 3498 43668 3500
rect 43069 3496 43668 3498
rect 43069 3440 43074 3496
rect 43130 3440 43668 3496
rect 43069 3438 43668 3440
rect 43069 3435 43135 3438
rect 43662 3436 43668 3438
rect 43732 3436 43738 3500
rect 50153 3498 50219 3501
rect 50838 3498 50844 3500
rect 50153 3496 50844 3498
rect 50153 3440 50158 3496
rect 50214 3440 50844 3496
rect 50153 3438 50844 3440
rect 50153 3435 50219 3438
rect 50838 3436 50844 3438
rect 50908 3436 50914 3500
rect 60825 3498 60891 3501
rect 61142 3498 61148 3500
rect 60825 3496 61148 3498
rect 60825 3440 60830 3496
rect 60886 3440 61148 3496
rect 60825 3438 61148 3440
rect 60825 3435 60891 3438
rect 61142 3436 61148 3438
rect 61212 3436 61218 3500
rect 150617 3498 150683 3501
rect 570229 3498 570295 3501
rect 150617 3496 570295 3498
rect 150617 3440 150622 3496
rect 150678 3440 570234 3496
rect 570290 3440 570295 3496
rect 150617 3438 570295 3440
rect 150617 3435 150683 3438
rect 570229 3435 570295 3438
rect 55070 3300 55076 3364
rect 55140 3362 55146 3364
rect 103329 3362 103395 3365
rect 55140 3360 103395 3362
rect 55140 3304 103334 3360
rect 103390 3304 103395 3360
rect 55140 3302 103395 3304
rect 55140 3300 55146 3302
rect 103329 3299 103395 3302
rect 126973 3362 127039 3365
rect 571374 3362 571380 3364
rect 126973 3360 571380 3362
rect 126973 3304 126978 3360
rect 127034 3304 571380 3360
rect 126973 3302 571380 3304
rect 126973 3299 127039 3302
rect 571374 3300 571380 3302
rect 571444 3300 571450 3364
rect 39798 3164 39804 3228
rect 39868 3226 39874 3228
rect 182541 3226 182607 3229
rect 39868 3224 182607 3226
rect 39868 3168 182546 3224
rect 182602 3168 182607 3224
rect 39868 3166 182607 3168
rect 39868 3164 39874 3166
rect 182541 3163 182607 3166
<< via3 >>
rect 566044 700300 566108 700364
rect 359412 687244 359476 687308
rect 28212 685884 28276 685948
rect 552060 685884 552124 685948
rect 382780 685204 382844 685268
rect 575428 685204 575492 685268
rect 355180 685068 355244 685132
rect 579660 685068 579724 685132
rect 551692 684932 551756 684996
rect 569908 684796 569972 684860
rect 361436 684660 361500 684724
rect 25452 684524 25516 684588
rect 551508 684524 551572 684588
rect 409828 683844 409892 683908
rect 393084 683708 393148 683772
rect 402100 683572 402164 683636
rect 375052 683436 375116 683500
rect 400812 682620 400876 682684
rect 371740 682484 371804 682548
rect 400996 682348 401060 682412
rect 566964 682348 567028 682412
rect 383516 682212 383580 682276
rect 560524 682212 560588 682276
rect 356652 682076 356716 682140
rect 389772 681940 389836 682004
rect 574140 681940 574204 682004
rect 406516 681804 406580 681868
rect 570092 681124 570156 681188
rect 363460 680988 363524 681052
rect 368980 680852 369044 680916
rect 370636 680716 370700 680780
rect 410012 680580 410076 680644
rect 578556 680444 578620 680508
rect 403572 680308 403636 680372
rect 388300 679900 388364 679964
rect 409644 679764 409708 679828
rect 552428 679628 552492 679692
rect 565124 679492 565188 679556
rect 409828 678268 409892 678332
rect 164924 678132 164988 678196
rect 153700 677724 153764 677788
rect 346900 677724 346964 677788
rect 152412 677588 152476 677652
rect 324452 677588 324516 677652
rect 336780 677588 336844 677652
rect 409828 677588 409892 677652
rect 325740 677104 325804 677108
rect 325740 677048 325790 677104
rect 325790 677048 325804 677104
rect 325740 677044 325804 677048
rect 552060 673916 552124 673980
rect 551508 673372 551572 673436
rect 552244 673372 552308 673436
rect 580948 669836 581012 669900
rect 557580 668476 557644 668540
rect 563100 667796 563164 667860
rect 570276 666436 570340 666500
rect 565308 663716 565372 663780
rect 391060 660996 391124 661060
rect 405596 658956 405660 659020
rect 377260 657596 377324 657660
rect 561628 650796 561692 650860
rect 558868 649436 558932 649500
rect 408356 646716 408420 646780
rect 578740 646036 578804 646100
rect 552060 641276 552124 641340
rect 406332 637876 406396 637940
rect 364932 635836 364996 635900
rect 557764 633796 557828 633860
rect 391796 628356 391860 628420
rect 553348 628356 553412 628420
rect 406148 627676 406212 627740
rect 576900 626996 576964 627060
rect 572668 625228 572732 625292
rect 401364 624276 401428 624340
rect 395844 619516 395908 619580
rect 575612 612716 575676 612780
rect 559052 612036 559116 612100
rect 388484 611356 388548 611420
rect 556292 607956 556356 608020
rect 387564 604420 387628 604484
rect 563284 602516 563348 602580
rect 571380 601836 571444 601900
rect 31524 599388 31588 599452
rect 560708 599796 560772 599860
rect 556108 599116 556172 599180
rect 378732 598436 378796 598500
rect 371924 593676 371988 593740
rect 397316 590956 397380 591020
rect 50108 590608 50172 590612
rect 50108 590552 50122 590608
rect 50122 590552 50172 590608
rect 50108 590548 50172 590552
rect 55812 590608 55876 590612
rect 55812 590552 55862 590608
rect 55862 590552 55876 590608
rect 55812 590548 55876 590552
rect 60412 590608 60476 590612
rect 60412 590552 60426 590608
rect 60426 590552 60476 590608
rect 60412 590548 60476 590552
rect 69796 590548 69860 590612
rect 74764 590608 74828 590612
rect 74764 590552 74814 590608
rect 74814 590552 74828 590608
rect 74764 590548 74828 590552
rect 77524 590548 77588 590612
rect 99972 590608 100036 590612
rect 99972 590552 99986 590608
rect 99986 590552 100036 590608
rect 99972 590548 100036 590552
rect 107516 590608 107580 590612
rect 107516 590552 107566 590608
rect 107566 590552 107580 590608
rect 107516 590548 107580 590552
rect 127388 590608 127452 590612
rect 127388 590552 127402 590608
rect 127402 590552 127452 590608
rect 127388 590548 127452 590552
rect 129780 590608 129844 590612
rect 129780 590552 129794 590608
rect 129794 590552 129844 590608
rect 129780 590548 129844 590552
rect 221964 590548 222028 590612
rect 223068 590608 223132 590612
rect 223068 590552 223082 590608
rect 223082 590552 223132 590608
rect 223068 590548 223132 590552
rect 238340 590608 238404 590612
rect 238340 590552 238390 590608
rect 238390 590552 238404 590608
rect 238340 590548 238404 590552
rect 241836 590548 241900 590612
rect 246620 590608 246684 590612
rect 246620 590552 246670 590608
rect 246670 590552 246684 590608
rect 246620 590548 246684 590552
rect 252324 590608 252388 590612
rect 252324 590552 252374 590608
rect 252374 590552 252388 590608
rect 252324 590548 252388 590552
rect 274220 590548 274284 590612
rect 289492 590608 289556 590612
rect 289492 590552 289542 590608
rect 289542 590552 289556 590608
rect 289492 590548 289556 590552
rect 292068 590608 292132 590612
rect 292068 590552 292118 590608
rect 292118 590552 292132 590608
rect 292068 590548 292132 590552
rect 311940 590548 312004 590612
rect 48452 590412 48516 590476
rect 77892 590412 77956 590476
rect 79916 590412 79980 590476
rect 93164 590412 93228 590476
rect 97580 590412 97644 590476
rect 351132 590412 351196 590476
rect 43484 590276 43548 590340
rect 43852 590140 43916 590204
rect 85252 589732 85316 589796
rect 122604 589792 122668 589796
rect 122604 589736 122618 589792
rect 122618 589736 122668 589792
rect 122604 589732 122668 589736
rect 240548 589792 240612 589796
rect 240548 589736 240598 589792
rect 240598 589736 240612 589792
rect 240548 589732 240612 589736
rect 255820 589732 255884 589796
rect 304580 589732 304644 589796
rect 350580 589732 350644 589796
rect 68508 589596 68572 589660
rect 137324 589656 137388 589660
rect 137324 589600 137338 589656
rect 137338 589600 137388 589656
rect 137324 589596 137388 589600
rect 279372 589596 279436 589660
rect 329236 589596 329300 589660
rect 52132 589460 52196 589524
rect 54524 589460 54588 589524
rect 59492 589460 59556 589524
rect 62620 589460 62684 589524
rect 72188 589460 72252 589524
rect 75684 589460 75748 589524
rect 79180 589460 79244 589524
rect 80468 589460 80532 589524
rect 82308 589460 82372 589524
rect 84884 589460 84948 589524
rect 87276 589460 87340 589524
rect 88380 589460 88444 589524
rect 90036 589460 90100 589524
rect 104940 589520 105004 589524
rect 104940 589464 104954 589520
rect 104954 589464 105004 589520
rect 104940 589460 105004 589464
rect 229140 589460 229204 589524
rect 231348 589460 231412 589524
rect 234292 589460 234356 589524
rect 237236 589460 237300 589524
rect 239628 589460 239692 589524
rect 242204 589460 242268 589524
rect 244412 589460 244476 589524
rect 248828 589460 248892 589524
rect 251220 589520 251284 589524
rect 251220 589464 251234 589520
rect 251234 589464 251284 589520
rect 251220 589460 251284 589464
rect 254716 589460 254780 589524
rect 256924 589460 256988 589524
rect 260420 589460 260484 589524
rect 262076 589460 262140 589524
rect 264100 589460 264164 589524
rect 266860 589460 266924 589524
rect 294460 589460 294524 589524
rect 297036 589460 297100 589524
rect 299428 589520 299492 589524
rect 299428 589464 299478 589520
rect 299478 589464 299492 589520
rect 299428 589460 299492 589464
rect 301820 589460 301884 589524
rect 306972 589460 307036 589524
rect 309364 589460 309428 589524
rect 329420 589460 329484 589524
rect 51212 589384 51276 589388
rect 51212 589328 51226 589384
rect 51226 589328 51276 589384
rect 51212 589324 51276 589328
rect 53604 589324 53668 589388
rect 57100 589324 57164 589388
rect 58204 589324 58268 589388
rect 61516 589324 61580 589388
rect 62252 589324 62316 589388
rect 64092 589324 64156 589388
rect 64828 589384 64892 589388
rect 64828 589328 64842 589384
rect 64842 589328 64892 589384
rect 64828 589324 64892 589328
rect 65380 589384 65444 589388
rect 65380 589328 65430 589384
rect 65430 589328 65444 589384
rect 65380 589324 65444 589328
rect 66300 589384 66364 589388
rect 66300 589328 66314 589384
rect 66314 589328 66364 589384
rect 66300 589324 66364 589328
rect 67404 589324 67468 589388
rect 67772 589384 67836 589388
rect 67772 589328 67786 589384
rect 67786 589328 67836 589384
rect 67772 589324 67836 589328
rect 70164 589324 70228 589388
rect 71084 589384 71148 589388
rect 71084 589328 71134 589384
rect 71134 589328 71148 589384
rect 71084 589324 71148 589328
rect 72372 589324 72436 589388
rect 73476 589324 73540 589388
rect 75132 589324 75196 589388
rect 76788 589324 76852 589388
rect 81572 589324 81636 589388
rect 82676 589384 82740 589388
rect 82676 589328 82690 589384
rect 82690 589328 82740 589384
rect 82676 589324 82740 589328
rect 83780 589324 83844 589388
rect 86172 589324 86236 589388
rect 87644 589324 87708 589388
rect 89852 589324 89916 589388
rect 90956 589384 91020 589388
rect 90956 589328 90970 589384
rect 90970 589328 91020 589384
rect 90956 589324 91020 589328
rect 92060 589324 92124 589388
rect 92428 589324 92492 589388
rect 95004 589324 95068 589388
rect 102364 589324 102428 589388
rect 109908 589324 109972 589388
rect 112484 589324 112548 589388
rect 114876 589324 114940 589388
rect 117452 589324 117516 589388
rect 120028 589384 120092 589388
rect 120028 589328 120042 589384
rect 120042 589328 120092 589384
rect 120028 589324 120092 589328
rect 124996 589324 125060 589388
rect 132540 589384 132604 589388
rect 132540 589328 132554 589384
rect 132554 589328 132604 589384
rect 132540 589324 132604 589328
rect 134932 589324 134996 589388
rect 139900 589324 139964 589388
rect 157196 589384 157260 589388
rect 157196 589328 157246 589384
rect 157246 589328 157260 589384
rect 157196 589324 157260 589328
rect 157380 589324 157444 589388
rect 224172 589324 224236 589388
rect 225644 589324 225708 589388
rect 226564 589384 226628 589388
rect 226564 589328 226614 589384
rect 226614 589328 226628 589384
rect 226564 589324 226628 589328
rect 227852 589324 227916 589388
rect 230244 589324 230308 589388
rect 232452 589324 232516 589388
rect 233556 589324 233620 589388
rect 234660 589384 234724 589388
rect 234660 589328 234674 589384
rect 234674 589328 234724 589384
rect 234660 589324 234724 589328
rect 236132 589384 236196 589388
rect 236132 589328 236146 589384
rect 236146 589328 236196 589384
rect 236132 589324 236196 589328
rect 236684 589324 236748 589388
rect 239444 589324 239508 589388
rect 242940 589384 243004 589388
rect 242940 589328 242954 589384
rect 242954 589328 243004 589384
rect 242940 589324 243004 589328
rect 244044 589324 244108 589388
rect 245516 589384 245580 589388
rect 245516 589328 245566 589384
rect 245566 589328 245580 589384
rect 245516 589324 245580 589328
rect 246988 589384 247052 589388
rect 246988 589328 247038 589384
rect 247038 589328 247052 589384
rect 246988 589324 247052 589328
rect 247724 589324 247788 589388
rect 249564 589324 249628 589388
rect 249932 589324 249996 589388
rect 251956 589324 252020 589388
rect 253612 589324 253676 589388
rect 254164 589384 254228 589388
rect 254164 589328 254178 589384
rect 254178 589328 254228 589384
rect 254164 589324 254228 589328
rect 257292 589324 257356 589388
rect 258212 589324 258276 589388
rect 259316 589384 259380 589388
rect 259316 589328 259330 589384
rect 259330 589328 259380 589384
rect 259316 589324 259380 589328
rect 259684 589324 259748 589388
rect 261708 589324 261772 589388
rect 262996 589324 263060 589388
rect 264468 589324 264532 589388
rect 265204 589324 265268 589388
rect 269620 589324 269684 589388
rect 272012 589324 272076 589388
rect 276980 589324 277044 589388
rect 281948 589324 282012 589388
rect 284524 589324 284588 589388
rect 286916 589324 286980 589388
rect 347084 589324 347148 589388
rect 348004 588508 348068 588572
rect 567332 586196 567396 586260
rect 46796 585652 46860 585716
rect 381676 584836 381740 584900
rect 349476 584428 349540 584492
rect 399708 584292 399772 584356
rect 354444 582932 354508 582996
rect 571564 582116 571628 582180
rect 385540 581436 385604 581500
rect 373396 580756 373460 580820
rect 567516 580756 567580 580820
rect 359596 578716 359660 578780
rect 561812 576676 561876 576740
rect 45140 575996 45204 576060
rect 47164 574772 47228 574836
rect 46612 574636 46676 574700
rect 46980 572188 47044 572252
rect 346348 572052 346412 572116
rect 46428 571916 46492 571980
rect 550772 569876 550836 569940
rect 352052 568788 352116 568852
rect 376892 568652 376956 568716
rect 347084 568244 347148 568308
rect 347084 567972 347148 568036
rect 45324 567836 45388 567900
rect 378916 567292 378980 567356
rect 381492 567156 381556 567220
rect 369164 566748 369228 566812
rect 390140 566612 390204 566676
rect 347820 566476 347884 566540
rect 568620 566476 568684 566540
rect 349108 566340 349172 566404
rect 360700 566204 360764 566268
rect 351868 566068 351932 566132
rect 373212 565932 373276 565996
rect 365116 565796 365180 565860
rect 346900 565116 346964 565180
rect 347636 565116 347700 565180
rect 395292 564844 395356 564908
rect 396580 564436 396644 564500
rect 350948 563620 351012 563684
rect 41276 563212 41340 563276
rect 399524 563212 399588 563276
rect 48452 562668 48516 562732
rect 27476 562532 27540 562596
rect 346348 562532 346412 562596
rect 347452 562532 347516 562596
rect 41644 562396 41708 562460
rect 374500 561988 374564 562052
rect 367140 561716 367204 561780
rect 348372 561580 348436 561644
rect 349292 561036 349356 561100
rect 399340 560900 399404 560964
rect 46244 560492 46308 560556
rect 389956 560356 390020 560420
rect 347636 558860 347700 558924
rect 349660 558860 349724 558924
rect 385724 557636 385788 557700
rect 347636 557228 347700 557292
rect 48268 556140 48332 556204
rect 561996 552876 562060 552940
rect 565860 552060 565924 552124
rect 37596 546484 37660 546548
rect 560892 546756 560956 546820
rect 574324 544716 574388 544780
rect 349292 540908 349356 540972
rect 405412 537916 405476 537980
rect 35756 534108 35820 534172
rect 556476 534516 556540 534580
rect 557948 531796 558012 531860
rect 44036 530708 44100 530772
rect 407620 529076 407684 529140
rect 35572 527308 35636 527372
rect 39804 527172 39868 527236
rect 358124 527036 358188 527100
rect 47900 524588 47964 524652
rect 350580 522956 350644 523020
rect 391244 521596 391308 521660
rect 552428 520916 552492 520980
rect 353524 518876 353588 518940
rect 36676 514932 36740 514996
rect 348372 511940 348436 512004
rect 387012 510716 387076 510780
rect 350580 507860 350644 507924
rect 41092 506908 41156 506972
rect 356836 506636 356900 506700
rect 554820 505956 554884 506020
rect 392532 502420 392596 502484
rect 38516 499700 38580 499764
rect 40724 498748 40788 498812
rect 558132 497116 558196 497180
rect 350764 494532 350828 494596
rect 556660 494396 556724 494460
rect 553532 491676 553596 491740
rect 348372 487188 348436 487252
rect 44772 486508 44836 486572
rect 41828 485148 41892 485212
rect 349108 482972 349172 483036
rect 37044 480388 37108 480452
rect 559236 479436 559300 479500
rect 43852 476172 43916 476236
rect 565492 472636 565556 472700
rect 35388 470868 35452 470932
rect 350948 469236 351012 469300
rect 42012 466516 42076 466580
rect 36492 465156 36556 465220
rect 350948 463932 351012 463996
rect 43852 456860 43916 456924
rect 46244 455772 46308 455836
rect 39620 450468 39684 450532
rect 43668 449108 43732 449172
rect 349292 441900 349356 441964
rect 551508 441356 551572 441420
rect 579844 435916 579908 435980
rect 349108 434828 349172 434892
rect 44956 429252 45020 429316
rect 43484 424492 43548 424556
rect 35204 418372 35268 418436
rect 46428 412932 46492 412996
rect 367692 407356 367756 407420
rect 353708 407084 353772 407148
rect 555004 404636 555068 404700
rect 39436 402052 39500 402116
rect 32996 400828 33060 400892
rect 40908 396612 40972 396676
rect 36860 390628 36924 390692
rect 349660 385732 349724 385796
rect 349476 383692 349540 383756
rect 43484 382332 43548 382396
rect 351132 379476 351196 379540
rect 47716 378184 47780 378248
rect 407804 378116 407868 378180
rect 32812 374036 32876 374100
rect 403756 369276 403820 369340
rect 409460 357716 409524 357780
rect 550220 336636 550284 336700
rect 395476 331196 395540 331260
rect 348188 330652 348252 330716
rect 44772 321600 44836 321604
rect 44772 321544 44786 321600
rect 44786 321544 44836 321600
rect 44772 321540 44836 321544
rect 553716 315556 553780 315620
rect 409276 306036 409340 306100
rect 41644 304948 41708 305012
rect 41644 303588 41708 303652
rect 349476 295488 349540 295492
rect 349476 295432 349490 295488
rect 349490 295432 349540 295488
rect 349476 295428 349540 295432
rect 404860 293116 404924 293180
rect 566228 293116 566292 293180
rect 44772 292572 44836 292636
rect 47532 288424 47596 288488
rect 348004 286724 348068 286788
rect 567700 286316 567764 286380
rect 46244 284276 46308 284340
rect 46428 282916 46492 282980
rect 354444 278700 354508 278764
rect 409644 277476 409708 277540
rect 403940 272716 404004 272780
rect 355364 264964 355428 265028
rect 362908 262924 362972 262988
rect 31340 262244 31404 262308
rect 550404 262516 550468 262580
rect 27476 253948 27540 254012
rect 566044 249596 566108 249660
rect 46612 247284 46676 247348
rect 46060 247012 46124 247076
rect 46612 244352 46676 244356
rect 46612 244296 46626 244352
rect 46626 244296 46676 244352
rect 46612 244292 46676 244296
rect 46796 244292 46860 244356
rect 409828 242796 409892 242860
rect 410012 242388 410076 242452
rect 410012 242252 410076 242316
rect 44404 241436 44468 241500
rect 45140 240892 45204 240956
rect 409460 240348 409524 240412
rect 386460 239804 386524 239868
rect 548380 239668 548444 239732
rect 547092 239532 547156 239596
rect 551508 238580 551572 238644
rect 399708 238444 399772 238508
rect 549484 238308 549548 238372
rect 545068 238172 545132 238236
rect 552244 237220 552308 237284
rect 551692 237084 551756 237148
rect 409644 236948 409708 237012
rect 538812 236540 538876 236604
rect 393084 235452 393148 235516
rect 402100 235316 402164 235380
rect 561076 235180 561140 235244
rect 401364 234092 401428 234156
rect 538996 234092 539060 234156
rect 545252 232868 545316 232932
rect 387564 232732 387628 232796
rect 562180 232596 562244 232660
rect 357020 232460 357084 232524
rect 539180 230284 539244 230348
rect 47900 229740 47964 229804
rect 391796 229740 391860 229804
rect 47164 229332 47228 229396
rect 44772 224844 44836 224908
rect 44588 224164 44652 224228
rect 47164 220764 47228 220828
rect 46980 220492 47044 220556
rect 348556 214508 348620 214572
rect 44588 212604 44652 212668
rect 44772 211788 44836 211852
rect 44588 210428 44652 210492
rect 45324 210292 45388 210356
rect 48084 209612 48148 209676
rect 47164 209476 47228 209540
rect 406148 206212 406212 206276
rect 542676 204852 542740 204916
rect 37596 201376 37660 201380
rect 37596 201320 37646 201376
rect 37646 201320 37660 201376
rect 37596 201316 37660 201320
rect 347636 201316 347700 201380
rect 352052 201316 352116 201380
rect 47900 201180 47964 201244
rect 48268 200908 48332 200972
rect 347636 200908 347700 200972
rect 48268 200500 48332 200564
rect 347820 200288 347884 200292
rect 347820 200232 347834 200288
rect 347834 200232 347884 200288
rect 347820 200228 347884 200232
rect 48268 200092 48332 200156
rect 347636 199684 347700 199748
rect 356652 199548 356716 199612
rect 359412 199412 359476 199476
rect 346900 199276 346964 199340
rect 347636 199140 347700 199204
rect 560708 198596 560772 198660
rect 403572 198188 403636 198252
rect 364932 198052 364996 198116
rect 368980 197916 369044 197980
rect 561444 197372 561508 197436
rect 560892 197236 560956 197300
rect 400996 197100 401060 197164
rect 31524 196964 31588 197028
rect 348372 196828 348436 196892
rect 59124 196556 59188 196620
rect 407804 196556 407868 196620
rect 347636 195876 347700 195940
rect 363460 195604 363524 195668
rect 48084 195468 48148 195532
rect 387012 194516 387076 194580
rect 57652 193972 57716 194036
rect 53052 193836 53116 193900
rect 49188 192884 49252 192948
rect 53420 192748 53484 192812
rect 373396 192748 373460 192812
rect 44404 192612 44468 192676
rect 54892 190980 54956 191044
rect 350948 189892 351012 189956
rect 54524 189756 54588 189820
rect 395476 189756 395540 189820
rect 350580 188804 350644 188868
rect 41828 188668 41892 188732
rect 381676 188532 381740 188596
rect 54708 188396 54772 188460
rect 371924 188396 371988 188460
rect 378732 188260 378796 188324
rect 55076 187308 55140 187372
rect 367692 187308 367756 187372
rect 385724 187172 385788 187236
rect 43668 187036 43732 187100
rect 61332 185812 61396 185876
rect 36676 185676 36740 185740
rect 46244 185540 46308 185604
rect 539548 185540 539612 185604
rect 61516 184860 61580 184924
rect 349476 184724 349540 184788
rect 58572 184588 58636 184652
rect 407620 184588 407684 184652
rect 392532 184452 392596 184516
rect 43484 184316 43548 184380
rect 50844 184180 50908 184244
rect 350764 184044 350828 184108
rect 383516 183636 383580 183700
rect 349292 183228 349356 183292
rect 49556 183092 49620 183156
rect 382780 183092 382844 183156
rect 404860 182956 404924 183020
rect 35572 182820 35636 182884
rect 371740 182004 371804 182068
rect 348556 181868 348620 181932
rect 57836 181732 57900 181796
rect 365116 181732 365180 181796
rect 52316 181596 52380 181660
rect 47716 181460 47780 181524
rect 385540 181324 385604 181388
rect 59860 180508 59924 180572
rect 50660 180372 50724 180436
rect 358124 180372 358188 180436
rect 39804 180236 39868 180300
rect 539732 180100 539796 180164
rect 46244 179964 46308 180028
rect 552060 179964 552124 180028
rect 353524 179148 353588 179212
rect 49372 179012 49436 179076
rect 386460 179012 386524 179076
rect 388484 178876 388548 178940
rect 403756 178740 403820 178804
rect 39252 178604 39316 178668
rect 60412 177652 60476 177716
rect 52132 177516 52196 177580
rect 391060 177516 391124 177580
rect 44956 177380 45020 177444
rect 45140 177244 45204 177308
rect 353708 176564 353772 176628
rect 48084 176428 48148 176492
rect 367140 176428 367204 176492
rect 53236 176292 53300 176356
rect 39804 176156 39868 176220
rect 391244 176020 391308 176084
rect 541204 175884 541268 175948
rect 400812 175748 400876 175812
rect 53604 174796 53668 174860
rect 43668 174660 43732 174724
rect 55628 174524 55692 174588
rect 39436 173164 39500 173228
rect 403940 171668 404004 171732
rect 50476 170308 50540 170372
rect 389772 170308 389836 170372
rect 356836 168948 356900 169012
rect 58756 167860 58820 167924
rect 349108 167860 349172 167924
rect 40724 167724 40788 167788
rect 542676 167724 542740 167788
rect 42012 167588 42076 167652
rect 405412 166364 405476 166428
rect 547644 166364 547708 166428
rect 405596 166228 405660 166292
rect 560708 166228 560772 166292
rect 543964 165140 544028 165204
rect 397316 165004 397380 165068
rect 35204 164868 35268 164932
rect 390140 163508 390204 163572
rect 552060 163508 552124 163572
rect 369164 163372 369228 163436
rect 551508 163372 551572 163436
rect 409644 162420 409708 162484
rect 39620 162012 39684 162076
rect 399524 160924 399588 160988
rect 552612 160924 552676 160988
rect 378916 160788 378980 160852
rect 373212 160652 373276 160716
rect 552244 160652 552308 160716
rect 410012 159700 410076 159764
rect 563468 159700 563532 159764
rect 540100 159564 540164 159628
rect 57468 159428 57532 159492
rect 362908 159428 362972 159492
rect 395292 159428 395356 159492
rect 395844 158612 395908 158676
rect 541020 158476 541084 158540
rect 545436 158340 545500 158404
rect 60044 158204 60108 158268
rect 553900 158204 553964 158268
rect 46060 158068 46124 158132
rect 539916 158068 539980 158132
rect 32812 157932 32876 157996
rect 547276 157932 547340 157996
rect 375052 156980 375116 157044
rect 548012 156980 548076 157044
rect 542860 156844 542924 156908
rect 36492 156572 36556 156636
rect 406332 156572 406396 156636
rect 355364 155892 355428 155956
rect 544332 155892 544396 155956
rect 50292 155756 50356 155820
rect 376892 155756 376956 155820
rect 543044 155756 543108 155820
rect 35388 155620 35452 155684
rect 59308 155484 59372 155548
rect 46612 155348 46676 155412
rect 543780 155348 543844 155412
rect 566044 155212 566108 155276
rect 410196 155076 410260 155140
rect 406516 153988 406580 154052
rect 381492 153852 381556 153916
rect 541388 153852 541452 153916
rect 57284 153716 57348 153780
rect 359596 153716 359660 153780
rect 360700 153716 360764 153780
rect 552428 153716 552492 153780
rect 347084 153036 347148 153100
rect 370636 153096 370700 153100
rect 370636 153040 370650 153096
rect 370650 153040 370700 153096
rect 370636 153036 370700 153040
rect 396580 153036 396644 153100
rect 355180 152900 355244 152964
rect 357020 152764 357084 152828
rect 389956 152764 390020 152828
rect 388300 152628 388364 152692
rect 399340 152628 399404 152692
rect 346900 152492 346964 152556
rect 374500 152492 374564 152556
rect 563652 152492 563716 152556
rect 377260 152356 377324 152420
rect 408540 152356 408604 152420
rect 409828 152356 409892 152420
rect 351868 152220 351932 152284
rect 361436 152220 361500 152284
rect 541572 151676 541636 151740
rect 60964 151540 61028 151604
rect 566412 151404 566476 151468
rect 548196 151268 548260 151332
rect 544148 151132 544212 151196
rect 46612 150452 46676 150516
rect 545620 150044 545684 150108
rect 549668 149092 549732 149156
rect 542124 148956 542188 149020
rect 539364 148820 539428 148884
rect 539364 147868 539428 147932
rect 541388 147868 541452 147932
rect 60596 147460 60660 147524
rect 541940 147596 542004 147660
rect 539364 147324 539428 147388
rect 59676 147188 59740 147252
rect 60596 147188 60660 147252
rect 539364 147188 539428 147252
rect 541020 146916 541084 146980
rect 58940 146780 59004 146844
rect 60044 146780 60108 146844
rect 60596 146508 60660 146572
rect 542860 144740 542924 144804
rect 543596 144740 543660 144804
rect 57652 142972 57716 143036
rect 59492 141340 59556 141404
rect 542124 141204 542188 141268
rect 541388 141068 541452 141132
rect 543044 141068 543108 141132
rect 60412 140932 60476 140996
rect 542308 140796 542372 140860
rect 541756 139572 541820 139636
rect 541572 139436 541636 139500
rect 58388 138620 58452 138684
rect 58572 138076 58636 138140
rect 541940 138136 542004 138140
rect 541940 138080 541990 138136
rect 541990 138080 542004 138136
rect 541940 138076 542004 138080
rect 545252 137396 545316 137460
rect 543596 137260 543660 137324
rect 545068 137124 545132 137188
rect 45140 135220 45204 135284
rect 541020 135084 541084 135148
rect 545068 135144 545132 135148
rect 545068 135088 545082 135144
rect 545082 135088 545132 135144
rect 545068 135084 545132 135088
rect 543412 134404 543476 134468
rect 547644 133860 547708 133924
rect 55444 132500 55508 132564
rect 545252 131004 545316 131068
rect 541572 130188 541636 130252
rect 548012 130188 548076 130252
rect 541756 130052 541820 130116
rect 541388 129916 541452 129980
rect 541756 129780 541820 129844
rect 46244 128828 46308 128892
rect 544332 129372 544396 129436
rect 547828 128420 547892 128484
rect 544516 127604 544580 127668
rect 544884 126924 544948 126988
rect 545620 126924 545684 126988
rect 547460 126924 547524 126988
rect 547644 126244 547708 126308
rect 547644 126108 547708 126172
rect 543964 125564 544028 125628
rect 543412 125428 543476 125492
rect 547276 124612 547340 124676
rect 542860 124068 542924 124132
rect 562180 124068 562244 124132
rect 539364 122708 539428 122772
rect 548012 118764 548076 118828
rect 544148 117268 544212 117332
rect 58756 115092 58820 115156
rect 544332 115092 544396 115156
rect 58756 114412 58820 114476
rect 539364 114140 539428 114204
rect 542308 113052 542372 113116
rect 59492 112372 59556 112436
rect 566412 112372 566476 112436
rect 59492 110604 59556 110668
rect 543044 110604 543108 110668
rect 544516 110604 544580 110668
rect 543964 110468 544028 110532
rect 542492 109652 542556 109716
rect 544884 108972 544948 109036
rect 59492 107476 59556 107540
rect 60044 106660 60108 106724
rect 543228 106116 543292 106180
rect 542676 104212 542740 104276
rect 59308 101492 59372 101556
rect 59308 99996 59372 100060
rect 548196 92516 548260 92580
rect 539916 91700 539980 91764
rect 541388 89932 541452 89996
rect 59860 89796 59924 89860
rect 541756 89796 541820 89860
rect 545620 88980 545684 89044
rect 543780 87892 543844 87956
rect 539364 86804 539428 86868
rect 544516 86804 544580 86868
rect 552612 84628 552676 84692
rect 547460 82860 547524 82924
rect 540284 75788 540348 75852
rect 57468 74972 57532 75036
rect 545436 72932 545500 72996
rect 547276 72388 547340 72452
rect 541204 70892 541268 70956
rect 58756 68852 58820 68916
rect 566044 67628 566108 67692
rect 39252 57972 39316 58036
rect 543964 55932 544028 55996
rect 59124 54572 59188 54636
rect 551508 51036 551572 51100
rect 57836 49132 57900 49196
rect 53052 44236 53116 44300
rect 539548 38524 539612 38588
rect 46612 34988 46676 35052
rect 539732 35260 539796 35324
rect 57284 34852 57348 34916
rect 539364 31588 539428 31652
rect 60596 31044 60660 31108
rect 539548 31044 539612 31108
rect 552244 30772 552308 30836
rect 59308 30500 59372 30564
rect 539364 30500 539428 30564
rect 561628 29820 561692 29884
rect 552060 29548 552124 29612
rect 41092 29412 41156 29476
rect 49004 29276 49068 29340
rect 561812 29276 561876 29340
rect 49372 29140 49436 29204
rect 550404 29140 550468 29204
rect 539548 28928 539612 28932
rect 539548 28872 539562 28928
rect 539562 28872 539612 28928
rect 539548 28868 539612 28872
rect 38516 28732 38580 28796
rect 563100 28732 563164 28796
rect 561996 28596 562060 28660
rect 560708 28460 560772 28524
rect 48820 28324 48884 28388
rect 54524 28188 54588 28252
rect 44036 27916 44100 27980
rect 552428 27916 552492 27980
rect 50660 27508 50724 27572
rect 549668 27372 549732 27436
rect 53236 27236 53300 27300
rect 565124 27236 565188 27300
rect 40908 27100 40972 27164
rect 565308 27100 565372 27164
rect 41644 26964 41708 27028
rect 548012 26964 548076 27028
rect 43852 26828 43916 26892
rect 41276 26692 41340 26756
rect 31340 26556 31404 26620
rect 47532 26012 47596 26076
rect 54892 25876 54956 25940
rect 53420 25740 53484 25804
rect 575612 25740 575676 25804
rect 52132 25604 52196 25668
rect 566964 25604 567028 25668
rect 54708 25468 54772 25532
rect 32996 25332 33060 25396
rect 52316 24788 52380 24852
rect 44772 24652 44836 24716
rect 565492 24652 565556 24716
rect 563284 24516 563348 24580
rect 50476 24380 50540 24444
rect 567332 24380 567396 24444
rect 567516 24244 567580 24308
rect 568620 24108 568684 24172
rect 44588 23972 44652 24036
rect 565860 23972 565924 24036
rect 578740 23972 578804 24036
rect 36860 23836 36924 23900
rect 578556 23700 578620 23764
rect 547644 23292 547708 23356
rect 48084 23156 48148 23220
rect 542860 23156 542924 23220
rect 35756 23020 35820 23084
rect 544516 23020 544580 23084
rect 37044 22884 37108 22948
rect 560524 22884 560588 22948
rect 545068 22748 545132 22812
rect 49556 22612 49620 22676
rect 553532 22612 553596 22676
rect 553900 22476 553964 22540
rect 59676 21932 59740 21996
rect 538996 21932 539060 21996
rect 46428 21796 46492 21860
rect 540100 21796 540164 21860
rect 58572 21660 58636 21724
rect 544332 21660 544396 21724
rect 55444 21524 55508 21588
rect 547092 21524 547156 21588
rect 567700 21388 567764 21452
rect 553716 21252 553780 21316
rect 50292 21116 50356 21180
rect 563652 21116 563716 21180
rect 561444 20844 561508 20908
rect 570276 20844 570340 20908
rect 571564 20708 571628 20772
rect 543044 20164 543108 20228
rect 60044 20028 60108 20092
rect 561076 20028 561140 20092
rect 559236 19892 559300 19956
rect 556292 19756 556356 19820
rect 28212 19348 28276 19412
rect 572668 19076 572732 19140
rect 554820 18940 554884 19004
rect 574140 18804 574204 18868
rect 549484 18668 549548 18732
rect 576900 18532 576964 18596
rect 58940 18396 59004 18460
rect 557580 18396 557644 18460
rect 579844 17716 579908 17780
rect 580948 17580 581012 17644
rect 545620 17444 545684 17508
rect 570092 17308 570156 17372
rect 556476 17172 556540 17236
rect 541388 16492 541452 16556
rect 543228 16356 543292 16420
rect 545252 16084 545316 16148
rect 558132 15948 558196 16012
rect 548380 15812 548444 15876
rect 547276 14996 547340 15060
rect 540284 14860 540348 14924
rect 569908 14724 569972 14788
rect 579660 14588 579724 14652
rect 557948 14452 558012 14516
rect 557764 12004 557828 12068
rect 553348 11868 553412 11932
rect 541020 11732 541084 11796
rect 556108 11596 556172 11660
rect 538812 10916 538876 10980
rect 556660 10236 556724 10300
rect 555004 7516 555068 7580
rect 541572 6564 541636 6628
rect 563468 6428 563532 6492
rect 550588 6292 550652 6356
rect 559052 6156 559116 6220
rect 558868 4932 558932 4996
rect 550220 4796 550284 4860
rect 53604 3980 53668 4044
rect 55628 3844 55692 3908
rect 566228 3844 566292 3908
rect 574324 3708 574388 3772
rect 575428 3572 575492 3636
rect 25452 3436 25516 3500
rect 43668 3436 43732 3500
rect 50844 3436 50908 3500
rect 61148 3436 61212 3500
rect 55076 3300 55140 3364
rect 571380 3300 571444 3364
rect 39804 3164 39868 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28211 685948 28277 685949
rect 28211 685884 28212 685948
rect 28276 685884 28277 685948
rect 28211 685883 28277 685884
rect 25451 684588 25517 684589
rect 25451 684524 25452 684588
rect 25516 684524 25517 684588
rect 25451 684523 25517 684524
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 25454 3501 25514 684523
rect 27475 562596 27541 562597
rect 27475 562532 27476 562596
rect 27540 562532 27541 562596
rect 27475 562531 27541 562532
rect 27478 254013 27538 562531
rect 27475 254012 27541 254013
rect 27475 253948 27476 254012
rect 27540 253948 27541 254012
rect 27475 253947 27541 253948
rect 28214 19413 28274 685883
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 677308 33914 682398
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 677308 38414 686898
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 677308 42914 691398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 677308 47414 695898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 677308 51914 700398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 677308 65414 677898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 677308 69914 682398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 677308 74414 686898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 677308 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 677308 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 677308 87914 700398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 677308 101414 677898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 677308 105914 682398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 677308 110414 686898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 677308 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 677308 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 677308 123914 700398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 677308 137414 677898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 677308 141914 682398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 677308 146414 686898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 677308 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 153699 677788 153765 677789
rect 153699 677724 153700 677788
rect 153764 677724 153765 677788
rect 153699 677723 153765 677724
rect 152411 677652 152477 677653
rect 152411 677588 152412 677652
rect 152476 677588 152477 677652
rect 152411 677587 152477 677588
rect 152414 675610 152474 677587
rect 153702 675610 153762 677723
rect 154794 677308 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 677308 159914 700398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 164923 678196 164989 678197
rect 164923 678132 164924 678196
rect 164988 678132 164989 678196
rect 164923 678131 164989 678132
rect 172794 678134 173414 678218
rect 164926 675610 164986 678131
rect 152414 675550 152524 675610
rect 152464 675240 152524 675550
rect 153688 675550 153762 675610
rect 164840 675550 164986 675610
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 153688 675240 153748 675550
rect 164840 675240 164900 675550
rect 34272 655954 34620 655986
rect 34272 655718 34328 655954
rect 34564 655718 34620 655954
rect 34272 655634 34620 655718
rect 34272 655398 34328 655634
rect 34564 655398 34620 655634
rect 34272 655366 34620 655398
rect 170000 655954 170348 655986
rect 170000 655718 170056 655954
rect 170292 655718 170348 655954
rect 170000 655634 170348 655718
rect 170000 655398 170056 655634
rect 170292 655398 170348 655634
rect 170000 655366 170348 655398
rect 34952 651454 35300 651486
rect 34952 651218 35008 651454
rect 35244 651218 35300 651454
rect 34952 651134 35300 651218
rect 34952 650898 35008 651134
rect 35244 650898 35300 651134
rect 34952 650866 35300 650898
rect 169320 651454 169668 651486
rect 169320 651218 169376 651454
rect 169612 651218 169668 651454
rect 169320 651134 169668 651218
rect 169320 650898 169376 651134
rect 169612 650898 169668 651134
rect 169320 650866 169668 650898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 34272 619954 34620 619986
rect 34272 619718 34328 619954
rect 34564 619718 34620 619954
rect 34272 619634 34620 619718
rect 34272 619398 34328 619634
rect 34564 619398 34620 619634
rect 34272 619366 34620 619398
rect 170000 619954 170348 619986
rect 170000 619718 170056 619954
rect 170292 619718 170348 619954
rect 170000 619634 170348 619718
rect 170000 619398 170056 619634
rect 170292 619398 170348 619634
rect 170000 619366 170348 619398
rect 34952 615454 35300 615486
rect 34952 615218 35008 615454
rect 35244 615218 35300 615454
rect 34952 615134 35300 615218
rect 34952 614898 35008 615134
rect 35244 614898 35300 615134
rect 34952 614866 35300 614898
rect 169320 615454 169668 615486
rect 169320 615218 169376 615454
rect 169612 615218 169668 615454
rect 169320 615134 169668 615218
rect 169320 614898 169376 615134
rect 169612 614898 169668 615134
rect 169320 614866 169668 614898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 31523 599452 31589 599453
rect 31523 599388 31524 599452
rect 31588 599388 31589 599452
rect 31523 599387 31589 599388
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 31339 262308 31405 262309
rect 31339 262244 31340 262308
rect 31404 262244 31405 262308
rect 31339 262243 31405 262244
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28211 19412 28277 19413
rect 28211 19348 28212 19412
rect 28276 19348 28277 19412
rect 28211 19347 28277 19348
rect 25451 3500 25517 3501
rect 25451 3436 25452 3500
rect 25516 3436 25517 3500
rect 25451 3435 25517 3436
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 -6106 29414 29898
rect 31342 26621 31402 262243
rect 31526 197029 31586 599387
rect 50056 591290 50116 592106
rect 51144 591290 51204 592106
rect 52232 591290 52292 592106
rect 50056 591230 50170 591290
rect 51144 591230 51274 591290
rect 50110 590613 50170 591230
rect 50107 590612 50173 590613
rect 50107 590548 50108 590612
rect 50172 590548 50173 590612
rect 50107 590547 50173 590548
rect 48451 590476 48517 590477
rect 48451 590412 48452 590476
rect 48516 590412 48517 590476
rect 48451 590411 48517 590412
rect 43483 590340 43549 590341
rect 43483 590276 43484 590340
rect 43548 590276 43549 590340
rect 43483 590275 43549 590276
rect 33294 574954 33914 590000
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 37794 579454 38414 590000
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37595 546548 37661 546549
rect 37595 546484 37596 546548
rect 37660 546484 37661 546548
rect 37595 546483 37661 546484
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 35755 534172 35821 534173
rect 35755 534108 35756 534172
rect 35820 534108 35821 534172
rect 35755 534107 35821 534108
rect 35571 527372 35637 527373
rect 35571 527308 35572 527372
rect 35636 527308 35637 527372
rect 35571 527307 35637 527308
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 35387 470932 35453 470933
rect 35387 470868 35388 470932
rect 35452 470868 35453 470932
rect 35387 470867 35453 470868
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 32995 400892 33061 400893
rect 32995 400828 32996 400892
rect 33060 400828 33061 400892
rect 32995 400827 33061 400828
rect 32811 374100 32877 374101
rect 32811 374036 32812 374100
rect 32876 374036 32877 374100
rect 32811 374035 32877 374036
rect 31523 197028 31589 197029
rect 31523 196964 31524 197028
rect 31588 196964 31589 197028
rect 31523 196963 31589 196964
rect 32814 157997 32874 374035
rect 32811 157996 32877 157997
rect 32811 157932 32812 157996
rect 32876 157932 32877 157996
rect 32811 157931 32877 157932
rect 31339 26620 31405 26621
rect 31339 26556 31340 26620
rect 31404 26556 31405 26620
rect 31339 26555 31405 26556
rect 32998 25397 33058 400827
rect 33294 394954 33914 430398
rect 35203 418436 35269 418437
rect 35203 418372 35204 418436
rect 35268 418372 35269 418436
rect 35203 418371 35269 418372
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 35206 164933 35266 418371
rect 35203 164932 35269 164933
rect 35203 164868 35204 164932
rect 35268 164868 35269 164932
rect 35203 164867 35269 164868
rect 35390 155685 35450 470867
rect 35574 182885 35634 527307
rect 35571 182884 35637 182885
rect 35571 182820 35572 182884
rect 35636 182820 35637 182884
rect 35571 182819 35637 182820
rect 35387 155684 35453 155685
rect 35387 155620 35388 155684
rect 35452 155620 35453 155684
rect 35387 155619 35453 155620
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 32995 25396 33061 25397
rect 32995 25332 32996 25396
rect 33060 25332 33061 25396
rect 32995 25331 33061 25332
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 -7066 33914 34398
rect 35758 23085 35818 534107
rect 36675 514996 36741 514997
rect 36675 514932 36676 514996
rect 36740 514932 36741 514996
rect 36675 514931 36741 514932
rect 36491 465220 36557 465221
rect 36491 465156 36492 465220
rect 36556 465156 36557 465220
rect 36491 465155 36557 465156
rect 36494 156637 36554 465155
rect 36678 185741 36738 514931
rect 37043 480452 37109 480453
rect 37043 480388 37044 480452
rect 37108 480388 37109 480452
rect 37043 480387 37109 480388
rect 36859 390692 36925 390693
rect 36859 390628 36860 390692
rect 36924 390628 36925 390692
rect 36859 390627 36925 390628
rect 36675 185740 36741 185741
rect 36675 185676 36676 185740
rect 36740 185676 36741 185740
rect 36675 185675 36741 185676
rect 36491 156636 36557 156637
rect 36491 156572 36492 156636
rect 36556 156572 36557 156636
rect 36491 156571 36557 156572
rect 36862 23901 36922 390627
rect 36859 23900 36925 23901
rect 36859 23836 36860 23900
rect 36924 23836 36925 23900
rect 36859 23835 36925 23836
rect 35755 23084 35821 23085
rect 35755 23020 35756 23084
rect 35820 23020 35821 23084
rect 35755 23019 35821 23020
rect 37046 22949 37106 480387
rect 37598 201381 37658 546483
rect 37794 543454 38414 578898
rect 42294 583954 42914 590000
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 41275 563276 41341 563277
rect 41275 563212 41276 563276
rect 41340 563212 41341 563276
rect 41275 563211 41341 563212
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 39803 527236 39869 527237
rect 39803 527172 39804 527236
rect 39868 527172 39869 527236
rect 39803 527171 39869 527172
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 38515 499764 38581 499765
rect 38515 499700 38516 499764
rect 38580 499700 38581 499764
rect 38515 499699 38581 499700
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37595 201380 37661 201381
rect 37595 201316 37596 201380
rect 37660 201316 37661 201380
rect 37595 201315 37661 201316
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37043 22948 37109 22949
rect 37043 22884 37044 22948
rect 37108 22884 37109 22948
rect 37043 22883 37109 22884
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 3454 38414 38898
rect 38518 28797 38578 499699
rect 39619 450532 39685 450533
rect 39619 450468 39620 450532
rect 39684 450468 39685 450532
rect 39619 450467 39685 450468
rect 39435 402116 39501 402117
rect 39435 402052 39436 402116
rect 39500 402052 39501 402116
rect 39435 402051 39501 402052
rect 39251 178668 39317 178669
rect 39251 178604 39252 178668
rect 39316 178604 39317 178668
rect 39251 178603 39317 178604
rect 39254 58037 39314 178603
rect 39438 173229 39498 402051
rect 39435 173228 39501 173229
rect 39435 173164 39436 173228
rect 39500 173164 39501 173228
rect 39435 173163 39501 173164
rect 39622 162077 39682 450467
rect 39806 180301 39866 527171
rect 41091 506972 41157 506973
rect 41091 506908 41092 506972
rect 41156 506908 41157 506972
rect 41091 506907 41157 506908
rect 40723 498812 40789 498813
rect 40723 498748 40724 498812
rect 40788 498748 40789 498812
rect 40723 498747 40789 498748
rect 39803 180300 39869 180301
rect 39803 180236 39804 180300
rect 39868 180236 39869 180300
rect 39803 180235 39869 180236
rect 39803 176220 39869 176221
rect 39803 176156 39804 176220
rect 39868 176156 39869 176220
rect 39803 176155 39869 176156
rect 39619 162076 39685 162077
rect 39619 162012 39620 162076
rect 39684 162012 39685 162076
rect 39619 162011 39685 162012
rect 39251 58036 39317 58037
rect 39251 57972 39252 58036
rect 39316 57972 39317 58036
rect 39251 57971 39317 57972
rect 38515 28796 38581 28797
rect 38515 28732 38516 28796
rect 38580 28732 38581 28796
rect 38515 28731 38581 28732
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 39806 3229 39866 176155
rect 40726 167789 40786 498747
rect 40907 396676 40973 396677
rect 40907 396612 40908 396676
rect 40972 396612 40973 396676
rect 40907 396611 40973 396612
rect 40723 167788 40789 167789
rect 40723 167724 40724 167788
rect 40788 167724 40789 167788
rect 40723 167723 40789 167724
rect 40910 27165 40970 396611
rect 41094 29477 41154 506907
rect 41091 29476 41157 29477
rect 41091 29412 41092 29476
rect 41156 29412 41157 29476
rect 41091 29411 41157 29412
rect 40907 27164 40973 27165
rect 40907 27100 40908 27164
rect 40972 27100 40973 27164
rect 40907 27099 40973 27100
rect 41278 26757 41338 563211
rect 41643 562460 41709 562461
rect 41643 562396 41644 562460
rect 41708 562396 41709 562460
rect 41643 562395 41709 562396
rect 41646 305013 41706 562395
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 41827 485212 41893 485213
rect 41827 485148 41828 485212
rect 41892 485148 41893 485212
rect 41827 485147 41893 485148
rect 41643 305012 41709 305013
rect 41643 304948 41644 305012
rect 41708 304948 41709 305012
rect 41643 304947 41709 304948
rect 41643 303652 41709 303653
rect 41643 303588 41644 303652
rect 41708 303588 41709 303652
rect 41643 303587 41709 303588
rect 41646 27029 41706 303587
rect 41830 188733 41890 485147
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42011 466580 42077 466581
rect 42011 466516 42012 466580
rect 42076 466516 42077 466580
rect 42011 466515 42077 466516
rect 41827 188732 41893 188733
rect 41827 188668 41828 188732
rect 41892 188668 41893 188732
rect 41827 188667 41893 188668
rect 42014 167653 42074 466515
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 43486 424557 43546 590275
rect 43851 590204 43917 590205
rect 43851 590140 43852 590204
rect 43916 590140 43917 590204
rect 43851 590139 43917 590140
rect 43854 476237 43914 590139
rect 46795 585716 46861 585717
rect 46795 585652 46796 585716
rect 46860 585652 46861 585716
rect 46795 585651 46861 585652
rect 45139 576060 45205 576061
rect 45139 575996 45140 576060
rect 45204 575996 45205 576060
rect 45139 575995 45205 575996
rect 44035 530772 44101 530773
rect 44035 530708 44036 530772
rect 44100 530708 44101 530772
rect 44035 530707 44101 530708
rect 43851 476236 43917 476237
rect 43851 476172 43852 476236
rect 43916 476172 43917 476236
rect 43851 476171 43917 476172
rect 43851 456924 43917 456925
rect 43851 456860 43852 456924
rect 43916 456860 43917 456924
rect 43851 456859 43917 456860
rect 43667 449172 43733 449173
rect 43667 449108 43668 449172
rect 43732 449108 43733 449172
rect 43667 449107 43733 449108
rect 43483 424556 43549 424557
rect 43483 424492 43484 424556
rect 43548 424492 43549 424556
rect 43483 424491 43549 424492
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 43483 382396 43549 382397
rect 43483 382332 43484 382396
rect 43548 382332 43549 382396
rect 43483 382331 43549 382332
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42011 167652 42077 167653
rect 42011 167588 42012 167652
rect 42076 167588 42077 167652
rect 42011 167587 42077 167588
rect 42294 151954 42914 187398
rect 43486 184381 43546 382331
rect 43670 187101 43730 449107
rect 43667 187100 43733 187101
rect 43667 187036 43668 187100
rect 43732 187036 43733 187100
rect 43667 187035 43733 187036
rect 43483 184380 43549 184381
rect 43483 184316 43484 184380
rect 43548 184316 43549 184380
rect 43483 184315 43549 184316
rect 43667 174724 43733 174725
rect 43667 174660 43668 174724
rect 43732 174660 43733 174724
rect 43667 174659 43733 174660
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 41643 27028 41709 27029
rect 41643 26964 41644 27028
rect 41708 26964 41709 27028
rect 41643 26963 41709 26964
rect 41275 26756 41341 26757
rect 41275 26692 41276 26756
rect 41340 26692 41341 26756
rect 41275 26691 41341 26692
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 37794 3134 38414 3218
rect 39803 3228 39869 3229
rect 39803 3164 39804 3228
rect 39868 3164 39869 3228
rect 39803 3163 39869 3164
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 -1306 42914 7398
rect 43670 3501 43730 174659
rect 43854 26893 43914 456859
rect 44038 27981 44098 530707
rect 44771 486572 44837 486573
rect 44771 486508 44772 486572
rect 44836 486508 44837 486572
rect 44771 486507 44837 486508
rect 44774 321605 44834 486507
rect 44955 429316 45021 429317
rect 44955 429252 44956 429316
rect 45020 429252 45021 429316
rect 44955 429251 45021 429252
rect 44771 321604 44837 321605
rect 44771 321540 44772 321604
rect 44836 321540 44837 321604
rect 44771 321539 44837 321540
rect 44771 292636 44837 292637
rect 44771 292572 44772 292636
rect 44836 292572 44837 292636
rect 44771 292571 44837 292572
rect 44403 241500 44469 241501
rect 44403 241436 44404 241500
rect 44468 241436 44469 241500
rect 44403 241435 44469 241436
rect 44406 192677 44466 241435
rect 44774 224909 44834 292571
rect 44771 224908 44837 224909
rect 44771 224844 44772 224908
rect 44836 224844 44837 224908
rect 44771 224843 44837 224844
rect 44587 224228 44653 224229
rect 44587 224164 44588 224228
rect 44652 224164 44653 224228
rect 44587 224163 44653 224164
rect 44590 212669 44650 224163
rect 44587 212668 44653 212669
rect 44587 212604 44588 212668
rect 44652 212604 44653 212668
rect 44587 212603 44653 212604
rect 44771 211852 44837 211853
rect 44771 211788 44772 211852
rect 44836 211788 44837 211852
rect 44771 211787 44837 211788
rect 44587 210492 44653 210493
rect 44587 210428 44588 210492
rect 44652 210428 44653 210492
rect 44587 210427 44653 210428
rect 44403 192676 44469 192677
rect 44403 192612 44404 192676
rect 44468 192612 44469 192676
rect 44403 192611 44469 192612
rect 44035 27980 44101 27981
rect 44035 27916 44036 27980
rect 44100 27916 44101 27980
rect 44035 27915 44101 27916
rect 43851 26892 43917 26893
rect 43851 26828 43852 26892
rect 43916 26828 43917 26892
rect 43851 26827 43917 26828
rect 44590 24037 44650 210427
rect 44774 24717 44834 211787
rect 44958 177445 45018 429251
rect 45142 240957 45202 575995
rect 46611 574700 46677 574701
rect 46611 574636 46612 574700
rect 46676 574636 46677 574700
rect 46611 574635 46677 574636
rect 46427 571980 46493 571981
rect 46427 571916 46428 571980
rect 46492 571916 46493 571980
rect 46427 571915 46493 571916
rect 45323 567900 45389 567901
rect 45323 567836 45324 567900
rect 45388 567836 45389 567900
rect 45323 567835 45389 567836
rect 45139 240956 45205 240957
rect 45139 240892 45140 240956
rect 45204 240892 45205 240956
rect 45139 240891 45205 240892
rect 45326 210357 45386 567835
rect 46243 560556 46309 560557
rect 46243 560492 46244 560556
rect 46308 560492 46309 560556
rect 46243 560491 46309 560492
rect 46246 455837 46306 560491
rect 46243 455836 46309 455837
rect 46243 455772 46244 455836
rect 46308 455772 46309 455836
rect 46243 455771 46309 455772
rect 46430 412997 46490 571915
rect 46427 412996 46493 412997
rect 46427 412932 46428 412996
rect 46492 412932 46493 412996
rect 46427 412931 46493 412932
rect 46243 284340 46309 284341
rect 46243 284276 46244 284340
rect 46308 284276 46309 284340
rect 46243 284275 46309 284276
rect 46059 247076 46125 247077
rect 46059 247012 46060 247076
rect 46124 247012 46125 247076
rect 46059 247011 46125 247012
rect 45323 210356 45389 210357
rect 45323 210292 45324 210356
rect 45388 210292 45389 210356
rect 45323 210291 45389 210292
rect 44955 177444 45021 177445
rect 44955 177380 44956 177444
rect 45020 177380 45021 177444
rect 44955 177379 45021 177380
rect 45139 177308 45205 177309
rect 45139 177244 45140 177308
rect 45204 177244 45205 177308
rect 45139 177243 45205 177244
rect 45142 135285 45202 177243
rect 46062 158133 46122 247011
rect 46246 185605 46306 284275
rect 46427 282980 46493 282981
rect 46427 282916 46428 282980
rect 46492 282916 46493 282980
rect 46427 282915 46493 282916
rect 46243 185604 46309 185605
rect 46243 185540 46244 185604
rect 46308 185540 46309 185604
rect 46243 185539 46309 185540
rect 46243 180028 46309 180029
rect 46243 179964 46244 180028
rect 46308 179964 46309 180028
rect 46243 179963 46309 179964
rect 46059 158132 46125 158133
rect 46059 158068 46060 158132
rect 46124 158068 46125 158132
rect 46059 158067 46125 158068
rect 45139 135284 45205 135285
rect 45139 135220 45140 135284
rect 45204 135220 45205 135284
rect 45139 135219 45205 135220
rect 46246 128893 46306 179963
rect 46243 128892 46309 128893
rect 46243 128828 46244 128892
rect 46308 128828 46309 128892
rect 46243 128827 46309 128828
rect 44771 24716 44837 24717
rect 44771 24652 44772 24716
rect 44836 24652 44837 24716
rect 44771 24651 44837 24652
rect 44587 24036 44653 24037
rect 44587 23972 44588 24036
rect 44652 23972 44653 24036
rect 44587 23971 44653 23972
rect 46430 21861 46490 282915
rect 46614 247349 46674 574635
rect 46611 247348 46677 247349
rect 46611 247284 46612 247348
rect 46676 247284 46677 247348
rect 46611 247283 46677 247284
rect 46798 244357 46858 585651
rect 48454 576870 48514 590411
rect 51214 589389 51274 591230
rect 52134 591230 52292 591290
rect 53592 591290 53652 592106
rect 54544 591290 54604 592106
rect 53592 591230 53666 591290
rect 52134 589525 52194 591230
rect 52131 589524 52197 589525
rect 52131 589460 52132 589524
rect 52196 589460 52197 589524
rect 52131 589459 52197 589460
rect 53606 589389 53666 591230
rect 54526 591230 54604 591290
rect 55768 591290 55828 592106
rect 57128 591290 57188 592106
rect 58216 591290 58276 592106
rect 55768 591230 55874 591290
rect 54526 589525 54586 591230
rect 55814 590613 55874 591230
rect 57102 591230 57188 591290
rect 58206 591230 58276 591290
rect 59440 591290 59500 592106
rect 60528 591290 60588 592106
rect 61616 592050 61676 592106
rect 62296 592050 62356 592106
rect 62704 592050 62764 592106
rect 59440 591230 59554 591290
rect 55811 590612 55877 590613
rect 55811 590548 55812 590612
rect 55876 590548 55877 590612
rect 55811 590547 55877 590548
rect 54523 589524 54589 589525
rect 54523 589460 54524 589524
rect 54588 589460 54589 589524
rect 54523 589459 54589 589460
rect 57102 589389 57162 591230
rect 58206 589389 58266 591230
rect 59494 589525 59554 591230
rect 60414 591230 60588 591290
rect 61518 591990 61676 592050
rect 62254 591990 62356 592050
rect 62622 591990 62764 592050
rect 64064 592050 64124 592106
rect 64744 592050 64804 592106
rect 65288 592050 65348 592106
rect 66376 592050 66436 592106
rect 67464 592050 67524 592106
rect 64064 591990 64154 592050
rect 64744 591990 64890 592050
rect 65288 591990 65442 592050
rect 60414 590613 60474 591230
rect 60411 590612 60477 590613
rect 60411 590548 60412 590612
rect 60476 590548 60477 590612
rect 60411 590547 60477 590548
rect 59491 589524 59557 589525
rect 59491 589460 59492 589524
rect 59556 589460 59557 589524
rect 59491 589459 59557 589460
rect 61518 589389 61578 591990
rect 62254 589389 62314 591990
rect 62622 589525 62682 591990
rect 62619 589524 62685 589525
rect 62619 589460 62620 589524
rect 62684 589460 62685 589524
rect 62619 589459 62685 589460
rect 64094 589389 64154 591990
rect 64830 589389 64890 591990
rect 65382 589389 65442 591990
rect 66302 591990 66436 592050
rect 67406 591990 67524 592050
rect 67600 592050 67660 592106
rect 68552 592050 68612 592106
rect 69912 592050 69972 592106
rect 67600 591990 67834 592050
rect 66302 589389 66362 591990
rect 67406 589389 67466 591990
rect 67774 589389 67834 591990
rect 68510 591990 68612 592050
rect 69798 591990 69972 592050
rect 70048 592050 70108 592106
rect 71000 592050 71060 592106
rect 72088 592050 72148 592106
rect 72496 592050 72556 592106
rect 70048 591990 70226 592050
rect 71000 591990 71146 592050
rect 72088 591990 72250 592050
rect 68510 589661 68570 591990
rect 69798 590613 69858 591990
rect 69795 590612 69861 590613
rect 69795 590548 69796 590612
rect 69860 590548 69861 590612
rect 69795 590547 69861 590548
rect 68507 589660 68573 589661
rect 68507 589596 68508 589660
rect 68572 589596 68573 589660
rect 68507 589595 68573 589596
rect 70166 589389 70226 591990
rect 71086 589389 71146 591990
rect 72190 589525 72250 591990
rect 72374 591990 72556 592050
rect 73448 592050 73508 592106
rect 74672 592050 74732 592106
rect 75080 592050 75140 592106
rect 75760 592050 75820 592106
rect 76848 592050 76908 592106
rect 77528 592050 77588 592106
rect 77936 592050 77996 592106
rect 79296 592050 79356 592106
rect 79976 592050 80036 592106
rect 73448 591990 73538 592050
rect 74672 591990 74826 592050
rect 75080 591990 75194 592050
rect 72187 589524 72253 589525
rect 72187 589460 72188 589524
rect 72252 589460 72253 589524
rect 72187 589459 72253 589460
rect 72374 589389 72434 591990
rect 73478 589389 73538 591990
rect 74766 590613 74826 591990
rect 74763 590612 74829 590613
rect 74763 590548 74764 590612
rect 74828 590548 74829 590612
rect 74763 590547 74829 590548
rect 75134 589389 75194 591990
rect 75686 591990 75820 592050
rect 76790 591990 76908 592050
rect 77526 591990 77588 592050
rect 77894 591990 77996 592050
rect 79182 591990 79356 592050
rect 79918 591990 80036 592050
rect 80384 592050 80444 592106
rect 81608 592050 81668 592106
rect 80384 591990 80530 592050
rect 75686 589525 75746 591990
rect 75683 589524 75749 589525
rect 75683 589460 75684 589524
rect 75748 589460 75749 589524
rect 75683 589459 75749 589460
rect 76790 589389 76850 591990
rect 77526 590613 77586 591990
rect 77523 590612 77589 590613
rect 77523 590548 77524 590612
rect 77588 590548 77589 590612
rect 77523 590547 77589 590548
rect 77894 590477 77954 591990
rect 77891 590476 77957 590477
rect 77891 590412 77892 590476
rect 77956 590412 77957 590476
rect 77891 590411 77957 590412
rect 79182 589525 79242 591990
rect 79918 590477 79978 591990
rect 79915 590476 79981 590477
rect 79915 590412 79916 590476
rect 79980 590412 79981 590476
rect 79915 590411 79981 590412
rect 80470 589525 80530 591990
rect 81574 591990 81668 592050
rect 82288 592050 82348 592106
rect 82696 592050 82756 592106
rect 83784 592050 83844 592106
rect 85008 592050 85068 592106
rect 82288 591990 82370 592050
rect 79179 589524 79245 589525
rect 79179 589460 79180 589524
rect 79244 589460 79245 589524
rect 79179 589459 79245 589460
rect 80467 589524 80533 589525
rect 80467 589460 80468 589524
rect 80532 589460 80533 589524
rect 80467 589459 80533 589460
rect 81574 589389 81634 591990
rect 82310 589525 82370 591990
rect 82678 591990 82756 592050
rect 83782 591990 83844 592050
rect 84886 591990 85068 592050
rect 85144 592050 85204 592106
rect 86232 592050 86292 592106
rect 87320 592050 87380 592106
rect 85144 591990 85314 592050
rect 82307 589524 82373 589525
rect 82307 589460 82308 589524
rect 82372 589460 82373 589524
rect 82307 589459 82373 589460
rect 82678 589389 82738 591990
rect 83782 589389 83842 591990
rect 84886 589525 84946 591990
rect 85254 589797 85314 591990
rect 86174 591990 86292 592050
rect 87278 591990 87380 592050
rect 87592 592050 87652 592106
rect 88408 592050 88468 592106
rect 87592 591990 87706 592050
rect 85251 589796 85317 589797
rect 85251 589732 85252 589796
rect 85316 589732 85317 589796
rect 85251 589731 85317 589732
rect 84883 589524 84949 589525
rect 84883 589460 84884 589524
rect 84948 589460 84949 589524
rect 84883 589459 84949 589460
rect 86174 589389 86234 591990
rect 87278 589525 87338 591990
rect 87275 589524 87341 589525
rect 87275 589460 87276 589524
rect 87340 589460 87341 589524
rect 87275 589459 87341 589460
rect 87646 589389 87706 591990
rect 88382 591990 88468 592050
rect 89768 592050 89828 592106
rect 90040 592050 90100 592106
rect 90992 592050 91052 592106
rect 92080 592050 92140 592106
rect 92488 592050 92548 592106
rect 93168 592050 93228 592106
rect 89768 591990 89914 592050
rect 88382 589525 88442 591990
rect 88379 589524 88445 589525
rect 88379 589460 88380 589524
rect 88444 589460 88445 589524
rect 88379 589459 88445 589460
rect 89854 589389 89914 591990
rect 90038 591990 90100 592050
rect 90958 591990 91052 592050
rect 92062 591990 92140 592050
rect 92430 591990 92548 592050
rect 93166 591990 93228 592050
rect 94936 592050 94996 592106
rect 97520 592050 97580 592106
rect 94936 591990 95066 592050
rect 97520 591990 97642 592050
rect 90038 589525 90098 591990
rect 90035 589524 90101 589525
rect 90035 589460 90036 589524
rect 90100 589460 90101 589524
rect 90035 589459 90101 589460
rect 90958 589389 91018 591990
rect 92062 589389 92122 591990
rect 92430 589389 92490 591990
rect 93166 590477 93226 591990
rect 93163 590476 93229 590477
rect 93163 590412 93164 590476
rect 93228 590412 93229 590476
rect 93163 590411 93229 590412
rect 95006 589389 95066 591990
rect 97582 590477 97642 591990
rect 99968 591290 100028 592106
rect 102280 591290 102340 592106
rect 105000 591290 105060 592106
rect 99968 591230 100034 591290
rect 102280 591230 102426 591290
rect 99974 590613 100034 591230
rect 99971 590612 100037 590613
rect 99971 590548 99972 590612
rect 100036 590548 100037 590612
rect 99971 590547 100037 590548
rect 97579 590476 97645 590477
rect 97579 590412 97580 590476
rect 97644 590412 97645 590476
rect 97579 590411 97645 590412
rect 102366 589389 102426 591230
rect 104942 591230 105060 591290
rect 107448 591290 107508 592106
rect 109896 591290 109956 592106
rect 112480 591290 112540 592106
rect 114928 591290 114988 592106
rect 117512 591290 117572 592106
rect 107448 591230 107578 591290
rect 109896 591230 109970 591290
rect 112480 591230 112546 591290
rect 104942 589525 105002 591230
rect 107518 590613 107578 591230
rect 107515 590612 107581 590613
rect 107515 590548 107516 590612
rect 107580 590548 107581 590612
rect 107515 590547 107581 590548
rect 104939 589524 105005 589525
rect 104939 589460 104940 589524
rect 105004 589460 105005 589524
rect 104939 589459 105005 589460
rect 109910 589389 109970 591230
rect 112486 589389 112546 591230
rect 114878 591230 114988 591290
rect 117454 591230 117572 591290
rect 119960 591290 120020 592106
rect 122544 591290 122604 592106
rect 124992 591290 125052 592106
rect 127440 591290 127500 592106
rect 129888 591290 129948 592106
rect 119960 591230 120090 591290
rect 122544 591230 122666 591290
rect 124992 591230 125058 591290
rect 114878 589389 114938 591230
rect 117454 589389 117514 591230
rect 120030 589389 120090 591230
rect 122606 589797 122666 591230
rect 122603 589796 122669 589797
rect 122603 589732 122604 589796
rect 122668 589732 122669 589796
rect 122603 589731 122669 589732
rect 124998 589389 125058 591230
rect 127390 591230 127500 591290
rect 129782 591230 129948 591290
rect 132472 591290 132532 592106
rect 134920 591290 134980 592106
rect 137368 591290 137428 592106
rect 139952 591290 140012 592106
rect 157224 591290 157284 592106
rect 132472 591230 132602 591290
rect 134920 591230 134994 591290
rect 127390 590613 127450 591230
rect 129782 590613 129842 591230
rect 127387 590612 127453 590613
rect 127387 590548 127388 590612
rect 127452 590548 127453 590612
rect 127387 590547 127453 590548
rect 129779 590612 129845 590613
rect 129779 590548 129780 590612
rect 129844 590548 129845 590612
rect 129779 590547 129845 590548
rect 132542 589389 132602 591230
rect 134934 589389 134994 591230
rect 137326 591230 137428 591290
rect 139902 591230 140012 591290
rect 157198 591230 157284 591290
rect 157360 591290 157420 592106
rect 157360 591230 157442 591290
rect 137326 589661 137386 591230
rect 137323 589660 137389 589661
rect 137323 589596 137324 589660
rect 137388 589596 137389 589660
rect 137323 589595 137389 589596
rect 139902 589389 139962 591230
rect 157198 589389 157258 591230
rect 157382 589389 157442 591230
rect 51211 589388 51277 589389
rect 51211 589324 51212 589388
rect 51276 589324 51277 589388
rect 51211 589323 51277 589324
rect 53603 589388 53669 589389
rect 53603 589324 53604 589388
rect 53668 589324 53669 589388
rect 53603 589323 53669 589324
rect 57099 589388 57165 589389
rect 57099 589324 57100 589388
rect 57164 589324 57165 589388
rect 57099 589323 57165 589324
rect 58203 589388 58269 589389
rect 58203 589324 58204 589388
rect 58268 589324 58269 589388
rect 58203 589323 58269 589324
rect 61515 589388 61581 589389
rect 61515 589324 61516 589388
rect 61580 589324 61581 589388
rect 61515 589323 61581 589324
rect 62251 589388 62317 589389
rect 62251 589324 62252 589388
rect 62316 589324 62317 589388
rect 62251 589323 62317 589324
rect 64091 589388 64157 589389
rect 64091 589324 64092 589388
rect 64156 589324 64157 589388
rect 64091 589323 64157 589324
rect 64827 589388 64893 589389
rect 64827 589324 64828 589388
rect 64892 589324 64893 589388
rect 64827 589323 64893 589324
rect 65379 589388 65445 589389
rect 65379 589324 65380 589388
rect 65444 589324 65445 589388
rect 65379 589323 65445 589324
rect 66299 589388 66365 589389
rect 66299 589324 66300 589388
rect 66364 589324 66365 589388
rect 66299 589323 66365 589324
rect 67403 589388 67469 589389
rect 67403 589324 67404 589388
rect 67468 589324 67469 589388
rect 67403 589323 67469 589324
rect 67771 589388 67837 589389
rect 67771 589324 67772 589388
rect 67836 589324 67837 589388
rect 67771 589323 67837 589324
rect 70163 589388 70229 589389
rect 70163 589324 70164 589388
rect 70228 589324 70229 589388
rect 70163 589323 70229 589324
rect 71083 589388 71149 589389
rect 71083 589324 71084 589388
rect 71148 589324 71149 589388
rect 71083 589323 71149 589324
rect 72371 589388 72437 589389
rect 72371 589324 72372 589388
rect 72436 589324 72437 589388
rect 72371 589323 72437 589324
rect 73475 589388 73541 589389
rect 73475 589324 73476 589388
rect 73540 589324 73541 589388
rect 73475 589323 73541 589324
rect 75131 589388 75197 589389
rect 75131 589324 75132 589388
rect 75196 589324 75197 589388
rect 75131 589323 75197 589324
rect 76787 589388 76853 589389
rect 76787 589324 76788 589388
rect 76852 589324 76853 589388
rect 76787 589323 76853 589324
rect 81571 589388 81637 589389
rect 81571 589324 81572 589388
rect 81636 589324 81637 589388
rect 81571 589323 81637 589324
rect 82675 589388 82741 589389
rect 82675 589324 82676 589388
rect 82740 589324 82741 589388
rect 82675 589323 82741 589324
rect 83779 589388 83845 589389
rect 83779 589324 83780 589388
rect 83844 589324 83845 589388
rect 83779 589323 83845 589324
rect 86171 589388 86237 589389
rect 86171 589324 86172 589388
rect 86236 589324 86237 589388
rect 86171 589323 86237 589324
rect 87643 589388 87709 589389
rect 87643 589324 87644 589388
rect 87708 589324 87709 589388
rect 87643 589323 87709 589324
rect 89851 589388 89917 589389
rect 89851 589324 89852 589388
rect 89916 589324 89917 589388
rect 89851 589323 89917 589324
rect 90955 589388 91021 589389
rect 90955 589324 90956 589388
rect 91020 589324 91021 589388
rect 90955 589323 91021 589324
rect 92059 589388 92125 589389
rect 92059 589324 92060 589388
rect 92124 589324 92125 589388
rect 92059 589323 92125 589324
rect 92427 589388 92493 589389
rect 92427 589324 92428 589388
rect 92492 589324 92493 589388
rect 92427 589323 92493 589324
rect 95003 589388 95069 589389
rect 95003 589324 95004 589388
rect 95068 589324 95069 589388
rect 95003 589323 95069 589324
rect 102363 589388 102429 589389
rect 102363 589324 102364 589388
rect 102428 589324 102429 589388
rect 102363 589323 102429 589324
rect 109907 589388 109973 589389
rect 109907 589324 109908 589388
rect 109972 589324 109973 589388
rect 109907 589323 109973 589324
rect 112483 589388 112549 589389
rect 112483 589324 112484 589388
rect 112548 589324 112549 589388
rect 112483 589323 112549 589324
rect 114875 589388 114941 589389
rect 114875 589324 114876 589388
rect 114940 589324 114941 589388
rect 114875 589323 114941 589324
rect 117451 589388 117517 589389
rect 117451 589324 117452 589388
rect 117516 589324 117517 589388
rect 117451 589323 117517 589324
rect 120027 589388 120093 589389
rect 120027 589324 120028 589388
rect 120092 589324 120093 589388
rect 120027 589323 120093 589324
rect 124995 589388 125061 589389
rect 124995 589324 124996 589388
rect 125060 589324 125061 589388
rect 124995 589323 125061 589324
rect 132539 589388 132605 589389
rect 132539 589324 132540 589388
rect 132604 589324 132605 589388
rect 132539 589323 132605 589324
rect 134931 589388 134997 589389
rect 134931 589324 134932 589388
rect 134996 589324 134997 589388
rect 134931 589323 134997 589324
rect 139899 589388 139965 589389
rect 139899 589324 139900 589388
rect 139964 589324 139965 589388
rect 139899 589323 139965 589324
rect 157195 589388 157261 589389
rect 157195 589324 157196 589388
rect 157260 589324 157261 589388
rect 157195 589323 157261 589324
rect 157379 589388 157445 589389
rect 157379 589324 157380 589388
rect 157444 589324 157445 589388
rect 157379 589323 157445 589324
rect 48454 576810 48698 576870
rect 47163 574836 47229 574837
rect 47163 574772 47164 574836
rect 47228 574772 47229 574836
rect 47163 574771 47229 574772
rect 46979 572252 47045 572253
rect 46979 572188 46980 572252
rect 47044 572188 47045 572252
rect 46979 572187 47045 572188
rect 46611 244356 46677 244357
rect 46611 244292 46612 244356
rect 46676 244292 46677 244356
rect 46611 244291 46677 244292
rect 46795 244356 46861 244357
rect 46795 244292 46796 244356
rect 46860 244292 46861 244356
rect 46795 244291 46861 244292
rect 46614 155413 46674 244291
rect 46982 220557 47042 572187
rect 47166 229397 47226 574771
rect 48638 563070 48698 576810
rect 48270 563010 48698 563070
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 48270 556205 48330 563010
rect 48451 562732 48517 562733
rect 48451 562668 48452 562732
rect 48516 562668 48517 562732
rect 48451 562667 48517 562668
rect 48267 556204 48333 556205
rect 48267 556140 48268 556204
rect 48332 556140 48333 556204
rect 48267 556139 48333 556140
rect 48454 555930 48514 562667
rect 172794 562000 173414 569898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 562000 177914 574398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 562000 182414 578898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 562000 186914 583398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 562000 191414 587898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 562000 195914 592398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 677308 209414 677898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 677308 213914 682398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 677308 218414 686898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 677308 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 677308 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 677308 231914 700398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 677308 245414 677898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 677308 249914 682398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 677308 254414 686898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 677308 258914 691398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 677308 263414 695898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 677308 267914 700398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 677308 281414 677898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 677308 285914 682398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 677308 290414 686898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 677308 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 677308 299414 695898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 677308 303914 700398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 677308 317414 677898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 677308 321914 682398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 324451 677652 324517 677653
rect 324451 677588 324452 677652
rect 324516 677588 324517 677652
rect 324451 677587 324517 677588
rect 324454 675610 324514 677587
rect 325794 677308 326414 686898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 677308 330914 691398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 677308 335414 695898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 336779 677652 336845 677653
rect 336779 677588 336780 677652
rect 336844 677588 336845 677652
rect 336779 677587 336845 677588
rect 325739 677108 325805 677109
rect 325739 677044 325740 677108
rect 325804 677044 325805 677108
rect 325739 677043 325805 677044
rect 325742 675610 325802 677043
rect 324454 675550 324524 675610
rect 324464 675240 324524 675550
rect 325688 675550 325802 675610
rect 336782 675610 336842 677587
rect 339294 677308 339914 700398
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 346899 677788 346965 677789
rect 346899 677724 346900 677788
rect 346964 677724 346965 677788
rect 346899 677723 346965 677724
rect 336782 675550 336900 675610
rect 325688 675240 325748 675550
rect 336840 675240 336900 675550
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 206272 655954 206620 655986
rect 206272 655718 206328 655954
rect 206564 655718 206620 655954
rect 206272 655634 206620 655718
rect 206272 655398 206328 655634
rect 206564 655398 206620 655634
rect 206272 655366 206620 655398
rect 342000 655954 342348 655986
rect 342000 655718 342056 655954
rect 342292 655718 342348 655954
rect 342000 655634 342348 655718
rect 342000 655398 342056 655634
rect 342292 655398 342348 655634
rect 342000 655366 342348 655398
rect 206952 651454 207300 651486
rect 206952 651218 207008 651454
rect 207244 651218 207300 651454
rect 206952 651134 207300 651218
rect 206952 650898 207008 651134
rect 207244 650898 207300 651134
rect 206952 650866 207300 650898
rect 341320 651454 341668 651486
rect 341320 651218 341376 651454
rect 341612 651218 341668 651454
rect 341320 651134 341668 651218
rect 341320 650898 341376 651134
rect 341612 650898 341668 651134
rect 341320 650866 341668 650898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 206272 619954 206620 619986
rect 206272 619718 206328 619954
rect 206564 619718 206620 619954
rect 206272 619634 206620 619718
rect 206272 619398 206328 619634
rect 206564 619398 206620 619634
rect 206272 619366 206620 619398
rect 342000 619954 342348 619986
rect 342000 619718 342056 619954
rect 342292 619718 342348 619954
rect 342000 619634 342348 619718
rect 342000 619398 342056 619634
rect 342292 619398 342348 619634
rect 342000 619366 342348 619398
rect 206952 615454 207300 615486
rect 206952 615218 207008 615454
rect 207244 615218 207300 615454
rect 206952 615134 207300 615218
rect 206952 614898 207008 615134
rect 207244 614898 207300 615134
rect 206952 614866 207300 614898
rect 341320 615454 341668 615486
rect 341320 615218 341376 615454
rect 341612 615218 341668 615454
rect 341320 615134 341668 615218
rect 341320 614898 341376 615134
rect 341612 614898 341668 615134
rect 341320 614866 341668 614898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 562000 200414 596898
rect 222056 591290 222116 592106
rect 223144 591290 223204 592106
rect 224232 591290 224292 592106
rect 225592 592050 225652 592106
rect 226544 592050 226604 592106
rect 227768 592050 227828 592106
rect 229128 592050 229188 592106
rect 230216 592050 230276 592106
rect 231440 592050 231500 592106
rect 232528 592050 232588 592106
rect 233616 592050 233676 592106
rect 234296 592050 234356 592106
rect 234704 592050 234764 592106
rect 225592 591990 225706 592050
rect 226544 591990 226626 592050
rect 227768 591990 227914 592050
rect 229128 591990 229202 592050
rect 230216 591990 230306 592050
rect 221966 591230 222116 591290
rect 223070 591230 223204 591290
rect 224174 591230 224292 591290
rect 221966 590613 222026 591230
rect 223070 590613 223130 591230
rect 221963 590612 222029 590613
rect 221963 590548 221964 590612
rect 222028 590548 222029 590612
rect 221963 590547 222029 590548
rect 223067 590612 223133 590613
rect 223067 590548 223068 590612
rect 223132 590548 223133 590612
rect 223067 590547 223133 590548
rect 224174 589389 224234 591230
rect 225646 589389 225706 591990
rect 226566 589389 226626 591990
rect 227854 589389 227914 591990
rect 229142 589525 229202 591990
rect 229139 589524 229205 589525
rect 229139 589460 229140 589524
rect 229204 589460 229205 589524
rect 229139 589459 229205 589460
rect 230246 589389 230306 591990
rect 231350 591990 231500 592050
rect 232454 591990 232588 592050
rect 233558 591990 233676 592050
rect 234294 591990 234356 592050
rect 234662 591990 234764 592050
rect 236064 592050 236124 592106
rect 236744 592050 236804 592106
rect 237288 592050 237348 592106
rect 238376 592050 238436 592106
rect 239464 592050 239524 592106
rect 236064 591990 236194 592050
rect 231350 589525 231410 591990
rect 231347 589524 231413 589525
rect 231347 589460 231348 589524
rect 231412 589460 231413 589524
rect 231347 589459 231413 589460
rect 232454 589389 232514 591990
rect 233558 589389 233618 591990
rect 234294 589525 234354 591990
rect 234291 589524 234357 589525
rect 234291 589460 234292 589524
rect 234356 589460 234357 589524
rect 234291 589459 234357 589460
rect 234662 589389 234722 591990
rect 236134 589389 236194 591990
rect 236686 591990 236804 592050
rect 237238 591990 237348 592050
rect 238342 591990 238436 592050
rect 239446 591990 239524 592050
rect 239600 592050 239660 592106
rect 240552 592050 240612 592106
rect 241912 592050 241972 592106
rect 239600 591990 239690 592050
rect 236686 589389 236746 591990
rect 237238 589525 237298 591990
rect 238342 590613 238402 591990
rect 238339 590612 238405 590613
rect 238339 590548 238340 590612
rect 238404 590548 238405 590612
rect 238339 590547 238405 590548
rect 237235 589524 237301 589525
rect 237235 589460 237236 589524
rect 237300 589460 237301 589524
rect 237235 589459 237301 589460
rect 239446 589389 239506 591990
rect 239630 589525 239690 591990
rect 240550 591990 240612 592050
rect 241838 591990 241972 592050
rect 242048 592050 242108 592106
rect 243000 592050 243060 592106
rect 244088 592050 244148 592106
rect 244496 592050 244556 592106
rect 242048 591990 242266 592050
rect 240550 589797 240610 591990
rect 241838 590613 241898 591990
rect 241835 590612 241901 590613
rect 241835 590548 241836 590612
rect 241900 590548 241901 590612
rect 241835 590547 241901 590548
rect 240547 589796 240613 589797
rect 240547 589732 240548 589796
rect 240612 589732 240613 589796
rect 240547 589731 240613 589732
rect 242206 589525 242266 591990
rect 242942 591990 243060 592050
rect 244046 591990 244148 592050
rect 244414 591990 244556 592050
rect 245448 592050 245508 592106
rect 246672 592050 246732 592106
rect 247080 592050 247140 592106
rect 247760 592050 247820 592106
rect 248848 592050 248908 592106
rect 245448 591990 245578 592050
rect 239627 589524 239693 589525
rect 239627 589460 239628 589524
rect 239692 589460 239693 589524
rect 239627 589459 239693 589460
rect 242203 589524 242269 589525
rect 242203 589460 242204 589524
rect 242268 589460 242269 589524
rect 242203 589459 242269 589460
rect 242942 589389 243002 591990
rect 244046 589389 244106 591990
rect 244414 589525 244474 591990
rect 244411 589524 244477 589525
rect 244411 589460 244412 589524
rect 244476 589460 244477 589524
rect 244411 589459 244477 589460
rect 245518 589389 245578 591990
rect 246622 591990 246732 592050
rect 246990 591990 247140 592050
rect 247726 591990 247820 592050
rect 248830 591990 248908 592050
rect 249528 592050 249588 592106
rect 249936 592050 249996 592106
rect 251296 592050 251356 592106
rect 251976 592050 252036 592106
rect 252384 592050 252444 592106
rect 249528 591990 249626 592050
rect 246622 590613 246682 591990
rect 246619 590612 246685 590613
rect 246619 590548 246620 590612
rect 246684 590548 246685 590612
rect 246619 590547 246685 590548
rect 246990 589389 247050 591990
rect 247726 589389 247786 591990
rect 248830 589525 248890 591990
rect 248827 589524 248893 589525
rect 248827 589460 248828 589524
rect 248892 589460 248893 589524
rect 248827 589459 248893 589460
rect 249566 589389 249626 591990
rect 249934 591990 249996 592050
rect 251222 591990 251356 592050
rect 251958 591990 252036 592050
rect 252326 591990 252444 592050
rect 253608 592050 253668 592106
rect 254288 592050 254348 592106
rect 253608 591990 253674 592050
rect 249934 589389 249994 591990
rect 251222 589525 251282 591990
rect 251219 589524 251285 589525
rect 251219 589460 251220 589524
rect 251284 589460 251285 589524
rect 251219 589459 251285 589460
rect 251958 589389 252018 591990
rect 252326 590613 252386 591990
rect 252323 590612 252389 590613
rect 252323 590548 252324 590612
rect 252388 590548 252389 590612
rect 252323 590547 252389 590548
rect 253614 589389 253674 591990
rect 254166 591990 254348 592050
rect 254696 592050 254756 592106
rect 255784 592050 255844 592106
rect 257008 592050 257068 592106
rect 254696 591990 254778 592050
rect 255784 591990 255882 592050
rect 254166 589389 254226 591990
rect 254718 589525 254778 591990
rect 255822 589797 255882 591990
rect 256926 591990 257068 592050
rect 257144 592050 257204 592106
rect 258232 592050 258292 592106
rect 259320 592050 259380 592106
rect 257144 591990 257354 592050
rect 255819 589796 255885 589797
rect 255819 589732 255820 589796
rect 255884 589732 255885 589796
rect 255819 589731 255885 589732
rect 256926 589525 256986 591990
rect 254715 589524 254781 589525
rect 254715 589460 254716 589524
rect 254780 589460 254781 589524
rect 254715 589459 254781 589460
rect 256923 589524 256989 589525
rect 256923 589460 256924 589524
rect 256988 589460 256989 589524
rect 256923 589459 256989 589460
rect 257294 589389 257354 591990
rect 258214 591990 258292 592050
rect 259318 591990 259380 592050
rect 259592 592050 259652 592106
rect 260408 592050 260468 592106
rect 261768 592050 261828 592106
rect 259592 591990 259746 592050
rect 260408 591990 260482 592050
rect 258214 589389 258274 591990
rect 259318 589389 259378 591990
rect 259686 589389 259746 591990
rect 260422 589525 260482 591990
rect 261710 591990 261828 592050
rect 262040 592050 262100 592106
rect 262992 592050 263052 592106
rect 264080 592050 264140 592106
rect 264488 592050 264548 592106
rect 262040 591990 262138 592050
rect 262992 591990 263058 592050
rect 264080 591990 264162 592050
rect 260419 589524 260485 589525
rect 260419 589460 260420 589524
rect 260484 589460 260485 589524
rect 260419 589459 260485 589460
rect 261710 589389 261770 591990
rect 262078 589525 262138 591990
rect 262075 589524 262141 589525
rect 262075 589460 262076 589524
rect 262140 589460 262141 589524
rect 262075 589459 262141 589460
rect 262998 589389 263058 591990
rect 264102 589525 264162 591990
rect 264470 591990 264548 592050
rect 265168 592050 265228 592106
rect 266936 592050 266996 592106
rect 265168 591990 265266 592050
rect 264099 589524 264165 589525
rect 264099 589460 264100 589524
rect 264164 589460 264165 589524
rect 264099 589459 264165 589460
rect 264470 589389 264530 591990
rect 265206 589389 265266 591990
rect 266862 591990 266996 592050
rect 269520 592050 269580 592106
rect 271968 592050 272028 592106
rect 269520 591990 269682 592050
rect 271968 591990 272074 592050
rect 266862 589525 266922 591990
rect 266859 589524 266925 589525
rect 266859 589460 266860 589524
rect 266924 589460 266925 589524
rect 266859 589459 266925 589460
rect 269622 589389 269682 591990
rect 272014 589389 272074 591990
rect 274280 591290 274340 592106
rect 277000 591290 277060 592106
rect 279448 591290 279508 592106
rect 274222 591230 274340 591290
rect 276982 591230 277060 591290
rect 279374 591230 279508 591290
rect 281896 591290 281956 592106
rect 284480 591290 284540 592106
rect 286928 591290 286988 592106
rect 289512 591290 289572 592106
rect 281896 591230 282010 591290
rect 284480 591230 284586 591290
rect 274222 590613 274282 591230
rect 274219 590612 274285 590613
rect 274219 590548 274220 590612
rect 274284 590548 274285 590612
rect 274219 590547 274285 590548
rect 276982 589389 277042 591230
rect 279374 589661 279434 591230
rect 279371 589660 279437 589661
rect 279371 589596 279372 589660
rect 279436 589596 279437 589660
rect 279371 589595 279437 589596
rect 281950 589389 282010 591230
rect 284526 589389 284586 591230
rect 286918 591230 286988 591290
rect 289494 591230 289572 591290
rect 291960 591290 292020 592106
rect 294544 592050 294604 592106
rect 294462 591990 294604 592050
rect 296992 592050 297052 592106
rect 299440 592050 299500 592106
rect 301888 592050 301948 592106
rect 296992 591990 297098 592050
rect 291960 591230 292130 591290
rect 286918 589389 286978 591230
rect 289494 590613 289554 591230
rect 292070 590613 292130 591230
rect 289491 590612 289557 590613
rect 289491 590548 289492 590612
rect 289556 590548 289557 590612
rect 289491 590547 289557 590548
rect 292067 590612 292133 590613
rect 292067 590548 292068 590612
rect 292132 590548 292133 590612
rect 292067 590547 292133 590548
rect 294462 589525 294522 591990
rect 297038 589525 297098 591990
rect 299430 591990 299500 592050
rect 301822 591990 301948 592050
rect 299430 589525 299490 591990
rect 301822 589525 301882 591990
rect 304472 591290 304532 592106
rect 306920 591290 306980 592106
rect 309368 591290 309428 592106
rect 311952 591290 312012 592106
rect 304472 591230 304642 591290
rect 306920 591230 307034 591290
rect 304582 589797 304642 591230
rect 304579 589796 304645 589797
rect 304579 589732 304580 589796
rect 304644 589732 304645 589796
rect 304579 589731 304645 589732
rect 306974 589525 307034 591230
rect 309366 591230 309428 591290
rect 311942 591230 312012 591290
rect 329224 591290 329284 592106
rect 329360 591290 329420 592106
rect 329224 591230 329298 591290
rect 329360 591230 329482 591290
rect 309366 589525 309426 591230
rect 311942 590613 312002 591230
rect 311939 590612 312005 590613
rect 311939 590548 311940 590612
rect 312004 590548 312005 590612
rect 311939 590547 312005 590548
rect 329238 589661 329298 591230
rect 329235 589660 329301 589661
rect 329235 589596 329236 589660
rect 329300 589596 329301 589660
rect 329235 589595 329301 589596
rect 329422 589525 329482 591230
rect 294459 589524 294525 589525
rect 294459 589460 294460 589524
rect 294524 589460 294525 589524
rect 294459 589459 294525 589460
rect 297035 589524 297101 589525
rect 297035 589460 297036 589524
rect 297100 589460 297101 589524
rect 297035 589459 297101 589460
rect 299427 589524 299493 589525
rect 299427 589460 299428 589524
rect 299492 589460 299493 589524
rect 299427 589459 299493 589460
rect 301819 589524 301885 589525
rect 301819 589460 301820 589524
rect 301884 589460 301885 589524
rect 301819 589459 301885 589460
rect 306971 589524 307037 589525
rect 306971 589460 306972 589524
rect 307036 589460 307037 589524
rect 306971 589459 307037 589460
rect 309363 589524 309429 589525
rect 309363 589460 309364 589524
rect 309428 589460 309429 589524
rect 309363 589459 309429 589460
rect 329419 589524 329485 589525
rect 329419 589460 329420 589524
rect 329484 589460 329485 589524
rect 329419 589459 329485 589460
rect 224171 589388 224237 589389
rect 224171 589324 224172 589388
rect 224236 589324 224237 589388
rect 224171 589323 224237 589324
rect 225643 589388 225709 589389
rect 225643 589324 225644 589388
rect 225708 589324 225709 589388
rect 225643 589323 225709 589324
rect 226563 589388 226629 589389
rect 226563 589324 226564 589388
rect 226628 589324 226629 589388
rect 226563 589323 226629 589324
rect 227851 589388 227917 589389
rect 227851 589324 227852 589388
rect 227916 589324 227917 589388
rect 227851 589323 227917 589324
rect 230243 589388 230309 589389
rect 230243 589324 230244 589388
rect 230308 589324 230309 589388
rect 230243 589323 230309 589324
rect 232451 589388 232517 589389
rect 232451 589324 232452 589388
rect 232516 589324 232517 589388
rect 232451 589323 232517 589324
rect 233555 589388 233621 589389
rect 233555 589324 233556 589388
rect 233620 589324 233621 589388
rect 233555 589323 233621 589324
rect 234659 589388 234725 589389
rect 234659 589324 234660 589388
rect 234724 589324 234725 589388
rect 234659 589323 234725 589324
rect 236131 589388 236197 589389
rect 236131 589324 236132 589388
rect 236196 589324 236197 589388
rect 236131 589323 236197 589324
rect 236683 589388 236749 589389
rect 236683 589324 236684 589388
rect 236748 589324 236749 589388
rect 236683 589323 236749 589324
rect 239443 589388 239509 589389
rect 239443 589324 239444 589388
rect 239508 589324 239509 589388
rect 239443 589323 239509 589324
rect 242939 589388 243005 589389
rect 242939 589324 242940 589388
rect 243004 589324 243005 589388
rect 242939 589323 243005 589324
rect 244043 589388 244109 589389
rect 244043 589324 244044 589388
rect 244108 589324 244109 589388
rect 244043 589323 244109 589324
rect 245515 589388 245581 589389
rect 245515 589324 245516 589388
rect 245580 589324 245581 589388
rect 245515 589323 245581 589324
rect 246987 589388 247053 589389
rect 246987 589324 246988 589388
rect 247052 589324 247053 589388
rect 246987 589323 247053 589324
rect 247723 589388 247789 589389
rect 247723 589324 247724 589388
rect 247788 589324 247789 589388
rect 247723 589323 247789 589324
rect 249563 589388 249629 589389
rect 249563 589324 249564 589388
rect 249628 589324 249629 589388
rect 249563 589323 249629 589324
rect 249931 589388 249997 589389
rect 249931 589324 249932 589388
rect 249996 589324 249997 589388
rect 249931 589323 249997 589324
rect 251955 589388 252021 589389
rect 251955 589324 251956 589388
rect 252020 589324 252021 589388
rect 251955 589323 252021 589324
rect 253611 589388 253677 589389
rect 253611 589324 253612 589388
rect 253676 589324 253677 589388
rect 253611 589323 253677 589324
rect 254163 589388 254229 589389
rect 254163 589324 254164 589388
rect 254228 589324 254229 589388
rect 254163 589323 254229 589324
rect 257291 589388 257357 589389
rect 257291 589324 257292 589388
rect 257356 589324 257357 589388
rect 257291 589323 257357 589324
rect 258211 589388 258277 589389
rect 258211 589324 258212 589388
rect 258276 589324 258277 589388
rect 258211 589323 258277 589324
rect 259315 589388 259381 589389
rect 259315 589324 259316 589388
rect 259380 589324 259381 589388
rect 259315 589323 259381 589324
rect 259683 589388 259749 589389
rect 259683 589324 259684 589388
rect 259748 589324 259749 589388
rect 259683 589323 259749 589324
rect 261707 589388 261773 589389
rect 261707 589324 261708 589388
rect 261772 589324 261773 589388
rect 261707 589323 261773 589324
rect 262995 589388 263061 589389
rect 262995 589324 262996 589388
rect 263060 589324 263061 589388
rect 262995 589323 263061 589324
rect 264467 589388 264533 589389
rect 264467 589324 264468 589388
rect 264532 589324 264533 589388
rect 264467 589323 264533 589324
rect 265203 589388 265269 589389
rect 265203 589324 265204 589388
rect 265268 589324 265269 589388
rect 265203 589323 265269 589324
rect 269619 589388 269685 589389
rect 269619 589324 269620 589388
rect 269684 589324 269685 589388
rect 269619 589323 269685 589324
rect 272011 589388 272077 589389
rect 272011 589324 272012 589388
rect 272076 589324 272077 589388
rect 272011 589323 272077 589324
rect 276979 589388 277045 589389
rect 276979 589324 276980 589388
rect 277044 589324 277045 589388
rect 276979 589323 277045 589324
rect 281947 589388 282013 589389
rect 281947 589324 281948 589388
rect 282012 589324 282013 589388
rect 281947 589323 282013 589324
rect 284523 589388 284589 589389
rect 284523 589324 284524 589388
rect 284588 589324 284589 589388
rect 284523 589323 284589 589324
rect 286915 589388 286981 589389
rect 286915 589324 286916 589388
rect 286980 589324 286981 589388
rect 286915 589323 286981 589324
rect 346347 572116 346413 572117
rect 346347 572052 346348 572116
rect 346412 572052 346413 572116
rect 346347 572051 346413 572052
rect 346350 562597 346410 572051
rect 346902 565181 346962 677723
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 347083 589388 347149 589389
rect 347083 589324 347084 589388
rect 347148 589324 347149 589388
rect 347083 589323 347149 589324
rect 347086 568309 347146 589323
rect 348003 588572 348069 588573
rect 348003 588508 348004 588572
rect 348068 588508 348069 588572
rect 348003 588507 348069 588508
rect 347083 568308 347149 568309
rect 347083 568244 347084 568308
rect 347148 568244 347149 568308
rect 347083 568243 347149 568244
rect 347083 568036 347149 568037
rect 347083 567972 347084 568036
rect 347148 567972 347149 568036
rect 347083 567971 347149 567972
rect 346899 565180 346965 565181
rect 346899 565116 346900 565180
rect 346964 565116 346965 565180
rect 346899 565115 346965 565116
rect 346347 562596 346413 562597
rect 346347 562532 346348 562596
rect 346412 562532 346413 562596
rect 346347 562531 346413 562532
rect 347086 556610 347146 567971
rect 347819 566540 347885 566541
rect 347819 566476 347820 566540
rect 347884 566476 347885 566540
rect 347819 566475 347885 566476
rect 347635 565180 347701 565181
rect 347635 565116 347636 565180
rect 347700 565116 347701 565180
rect 347635 565115 347701 565116
rect 347451 562596 347517 562597
rect 347451 562532 347452 562596
rect 347516 562532 347517 562596
rect 347451 562531 347517 562532
rect 347454 557550 347514 562531
rect 347638 558925 347698 565115
rect 347635 558924 347701 558925
rect 347635 558860 347636 558924
rect 347700 558860 347701 558924
rect 347635 558859 347701 558860
rect 347822 557550 347882 566475
rect 348006 561370 348066 588507
rect 348294 565954 348914 601398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 355179 685132 355245 685133
rect 355179 685068 355180 685132
rect 355244 685068 355245 685132
rect 355179 685067 355245 685068
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 351131 590476 351197 590477
rect 351131 590412 351132 590476
rect 351196 590412 351197 590476
rect 351131 590411 351197 590412
rect 350579 589796 350645 589797
rect 350579 589732 350580 589796
rect 350644 589732 350645 589796
rect 350579 589731 350645 589732
rect 349475 584492 349541 584493
rect 349475 584428 349476 584492
rect 349540 584428 349541 584492
rect 349475 584427 349541 584428
rect 349107 566404 349173 566405
rect 349107 566340 349108 566404
rect 349172 566340 349173 566404
rect 349107 566339 349173 566340
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 562000 348914 565398
rect 348371 561644 348437 561645
rect 348371 561580 348372 561644
rect 348436 561580 348437 561644
rect 348371 561579 348437 561580
rect 348006 561310 348250 561370
rect 347454 557490 347698 557550
rect 347822 557490 348066 557550
rect 347638 557293 347698 557490
rect 347635 557292 347701 557293
rect 347635 557228 347636 557292
rect 347700 557228 347701 557292
rect 347635 557227 347701 557228
rect 347086 556550 347882 556610
rect 48086 555870 48514 555930
rect 48086 528570 48146 555870
rect 67568 547954 67888 547986
rect 67568 547718 67610 547954
rect 67846 547718 67888 547954
rect 67568 547634 67888 547718
rect 67568 547398 67610 547634
rect 67846 547398 67888 547634
rect 67568 547366 67888 547398
rect 98288 547954 98608 547986
rect 98288 547718 98330 547954
rect 98566 547718 98608 547954
rect 98288 547634 98608 547718
rect 98288 547398 98330 547634
rect 98566 547398 98608 547634
rect 98288 547366 98608 547398
rect 129008 547954 129328 547986
rect 129008 547718 129050 547954
rect 129286 547718 129328 547954
rect 129008 547634 129328 547718
rect 129008 547398 129050 547634
rect 129286 547398 129328 547634
rect 129008 547366 129328 547398
rect 159728 547954 160048 547986
rect 159728 547718 159770 547954
rect 160006 547718 160048 547954
rect 159728 547634 160048 547718
rect 159728 547398 159770 547634
rect 160006 547398 160048 547634
rect 159728 547366 160048 547398
rect 190448 547954 190768 547986
rect 190448 547718 190490 547954
rect 190726 547718 190768 547954
rect 190448 547634 190768 547718
rect 190448 547398 190490 547634
rect 190726 547398 190768 547634
rect 190448 547366 190768 547398
rect 221168 547954 221488 547986
rect 221168 547718 221210 547954
rect 221446 547718 221488 547954
rect 221168 547634 221488 547718
rect 221168 547398 221210 547634
rect 221446 547398 221488 547634
rect 221168 547366 221488 547398
rect 251888 547954 252208 547986
rect 251888 547718 251930 547954
rect 252166 547718 252208 547954
rect 251888 547634 252208 547718
rect 251888 547398 251930 547634
rect 252166 547398 252208 547634
rect 251888 547366 252208 547398
rect 282608 547954 282928 547986
rect 282608 547718 282650 547954
rect 282886 547718 282928 547954
rect 282608 547634 282928 547718
rect 282608 547398 282650 547634
rect 282886 547398 282928 547634
rect 282608 547366 282928 547398
rect 313328 547954 313648 547986
rect 313328 547718 313370 547954
rect 313606 547718 313648 547954
rect 313328 547634 313648 547718
rect 313328 547398 313370 547634
rect 313606 547398 313648 547634
rect 313328 547366 313648 547398
rect 344048 547954 344368 547986
rect 344048 547718 344090 547954
rect 344326 547718 344368 547954
rect 344048 547634 344368 547718
rect 344048 547398 344090 547634
rect 344326 547398 344368 547634
rect 344048 547366 344368 547398
rect 52208 543454 52528 543486
rect 52208 543218 52250 543454
rect 52486 543218 52528 543454
rect 52208 543134 52528 543218
rect 52208 542898 52250 543134
rect 52486 542898 52528 543134
rect 52208 542866 52528 542898
rect 82928 543454 83248 543486
rect 82928 543218 82970 543454
rect 83206 543218 83248 543454
rect 82928 543134 83248 543218
rect 82928 542898 82970 543134
rect 83206 542898 83248 543134
rect 82928 542866 83248 542898
rect 113648 543454 113968 543486
rect 113648 543218 113690 543454
rect 113926 543218 113968 543454
rect 113648 543134 113968 543218
rect 113648 542898 113690 543134
rect 113926 542898 113968 543134
rect 113648 542866 113968 542898
rect 144368 543454 144688 543486
rect 144368 543218 144410 543454
rect 144646 543218 144688 543454
rect 144368 543134 144688 543218
rect 144368 542898 144410 543134
rect 144646 542898 144688 543134
rect 144368 542866 144688 542898
rect 175088 543454 175408 543486
rect 175088 543218 175130 543454
rect 175366 543218 175408 543454
rect 175088 543134 175408 543218
rect 175088 542898 175130 543134
rect 175366 542898 175408 543134
rect 175088 542866 175408 542898
rect 205808 543454 206128 543486
rect 205808 543218 205850 543454
rect 206086 543218 206128 543454
rect 205808 543134 206128 543218
rect 205808 542898 205850 543134
rect 206086 542898 206128 543134
rect 205808 542866 206128 542898
rect 236528 543454 236848 543486
rect 236528 543218 236570 543454
rect 236806 543218 236848 543454
rect 236528 543134 236848 543218
rect 236528 542898 236570 543134
rect 236806 542898 236848 543134
rect 236528 542866 236848 542898
rect 267248 543454 267568 543486
rect 267248 543218 267290 543454
rect 267526 543218 267568 543454
rect 267248 543134 267568 543218
rect 267248 542898 267290 543134
rect 267526 542898 267568 543134
rect 267248 542866 267568 542898
rect 297968 543454 298288 543486
rect 297968 543218 298010 543454
rect 298246 543218 298288 543454
rect 297968 543134 298288 543218
rect 297968 542898 298010 543134
rect 298246 542898 298288 543134
rect 297968 542866 298288 542898
rect 328688 543454 329008 543486
rect 328688 543218 328730 543454
rect 328966 543218 329008 543454
rect 328688 543134 329008 543218
rect 328688 542898 328730 543134
rect 328966 542898 329008 543134
rect 328688 542866 329008 542898
rect 47902 528510 48146 528570
rect 47902 524653 47962 528510
rect 47899 524652 47965 524653
rect 47899 524588 47900 524652
rect 47964 524588 47965 524652
rect 47899 524587 47965 524588
rect 67568 511954 67888 511986
rect 67568 511718 67610 511954
rect 67846 511718 67888 511954
rect 67568 511634 67888 511718
rect 67568 511398 67610 511634
rect 67846 511398 67888 511634
rect 67568 511366 67888 511398
rect 98288 511954 98608 511986
rect 98288 511718 98330 511954
rect 98566 511718 98608 511954
rect 98288 511634 98608 511718
rect 98288 511398 98330 511634
rect 98566 511398 98608 511634
rect 98288 511366 98608 511398
rect 129008 511954 129328 511986
rect 129008 511718 129050 511954
rect 129286 511718 129328 511954
rect 129008 511634 129328 511718
rect 129008 511398 129050 511634
rect 129286 511398 129328 511634
rect 129008 511366 129328 511398
rect 159728 511954 160048 511986
rect 159728 511718 159770 511954
rect 160006 511718 160048 511954
rect 159728 511634 160048 511718
rect 159728 511398 159770 511634
rect 160006 511398 160048 511634
rect 159728 511366 160048 511398
rect 190448 511954 190768 511986
rect 190448 511718 190490 511954
rect 190726 511718 190768 511954
rect 190448 511634 190768 511718
rect 190448 511398 190490 511634
rect 190726 511398 190768 511634
rect 190448 511366 190768 511398
rect 221168 511954 221488 511986
rect 221168 511718 221210 511954
rect 221446 511718 221488 511954
rect 221168 511634 221488 511718
rect 221168 511398 221210 511634
rect 221446 511398 221488 511634
rect 221168 511366 221488 511398
rect 251888 511954 252208 511986
rect 251888 511718 251930 511954
rect 252166 511718 252208 511954
rect 251888 511634 252208 511718
rect 251888 511398 251930 511634
rect 252166 511398 252208 511634
rect 251888 511366 252208 511398
rect 282608 511954 282928 511986
rect 282608 511718 282650 511954
rect 282886 511718 282928 511954
rect 282608 511634 282928 511718
rect 282608 511398 282650 511634
rect 282886 511398 282928 511634
rect 282608 511366 282928 511398
rect 313328 511954 313648 511986
rect 313328 511718 313370 511954
rect 313606 511718 313648 511954
rect 313328 511634 313648 511718
rect 313328 511398 313370 511634
rect 313606 511398 313648 511634
rect 313328 511366 313648 511398
rect 344048 511954 344368 511986
rect 344048 511718 344090 511954
rect 344326 511718 344368 511954
rect 344048 511634 344368 511718
rect 344048 511398 344090 511634
rect 344326 511398 344368 511634
rect 344048 511366 344368 511398
rect 52208 507454 52528 507486
rect 52208 507218 52250 507454
rect 52486 507218 52528 507454
rect 52208 507134 52528 507218
rect 52208 506898 52250 507134
rect 52486 506898 52528 507134
rect 52208 506866 52528 506898
rect 82928 507454 83248 507486
rect 82928 507218 82970 507454
rect 83206 507218 83248 507454
rect 82928 507134 83248 507218
rect 82928 506898 82970 507134
rect 83206 506898 83248 507134
rect 82928 506866 83248 506898
rect 113648 507454 113968 507486
rect 113648 507218 113690 507454
rect 113926 507218 113968 507454
rect 113648 507134 113968 507218
rect 113648 506898 113690 507134
rect 113926 506898 113968 507134
rect 113648 506866 113968 506898
rect 144368 507454 144688 507486
rect 144368 507218 144410 507454
rect 144646 507218 144688 507454
rect 144368 507134 144688 507218
rect 144368 506898 144410 507134
rect 144646 506898 144688 507134
rect 144368 506866 144688 506898
rect 175088 507454 175408 507486
rect 175088 507218 175130 507454
rect 175366 507218 175408 507454
rect 175088 507134 175408 507218
rect 175088 506898 175130 507134
rect 175366 506898 175408 507134
rect 175088 506866 175408 506898
rect 205808 507454 206128 507486
rect 205808 507218 205850 507454
rect 206086 507218 206128 507454
rect 205808 507134 206128 507218
rect 205808 506898 205850 507134
rect 206086 506898 206128 507134
rect 205808 506866 206128 506898
rect 236528 507454 236848 507486
rect 236528 507218 236570 507454
rect 236806 507218 236848 507454
rect 236528 507134 236848 507218
rect 236528 506898 236570 507134
rect 236806 506898 236848 507134
rect 236528 506866 236848 506898
rect 267248 507454 267568 507486
rect 267248 507218 267290 507454
rect 267526 507218 267568 507454
rect 267248 507134 267568 507218
rect 267248 506898 267290 507134
rect 267526 506898 267568 507134
rect 267248 506866 267568 506898
rect 297968 507454 298288 507486
rect 297968 507218 298010 507454
rect 298246 507218 298288 507454
rect 297968 507134 298288 507218
rect 297968 506898 298010 507134
rect 298246 506898 298288 507134
rect 297968 506866 298288 506898
rect 328688 507454 329008 507486
rect 328688 507218 328730 507454
rect 328966 507218 329008 507454
rect 328688 507134 329008 507218
rect 328688 506898 328730 507134
rect 328966 506898 329008 507134
rect 328688 506866 329008 506898
rect 67568 475954 67888 475986
rect 67568 475718 67610 475954
rect 67846 475718 67888 475954
rect 67568 475634 67888 475718
rect 67568 475398 67610 475634
rect 67846 475398 67888 475634
rect 67568 475366 67888 475398
rect 98288 475954 98608 475986
rect 98288 475718 98330 475954
rect 98566 475718 98608 475954
rect 98288 475634 98608 475718
rect 98288 475398 98330 475634
rect 98566 475398 98608 475634
rect 98288 475366 98608 475398
rect 129008 475954 129328 475986
rect 129008 475718 129050 475954
rect 129286 475718 129328 475954
rect 129008 475634 129328 475718
rect 129008 475398 129050 475634
rect 129286 475398 129328 475634
rect 129008 475366 129328 475398
rect 159728 475954 160048 475986
rect 159728 475718 159770 475954
rect 160006 475718 160048 475954
rect 159728 475634 160048 475718
rect 159728 475398 159770 475634
rect 160006 475398 160048 475634
rect 159728 475366 160048 475398
rect 190448 475954 190768 475986
rect 190448 475718 190490 475954
rect 190726 475718 190768 475954
rect 190448 475634 190768 475718
rect 190448 475398 190490 475634
rect 190726 475398 190768 475634
rect 190448 475366 190768 475398
rect 221168 475954 221488 475986
rect 221168 475718 221210 475954
rect 221446 475718 221488 475954
rect 221168 475634 221488 475718
rect 221168 475398 221210 475634
rect 221446 475398 221488 475634
rect 221168 475366 221488 475398
rect 251888 475954 252208 475986
rect 251888 475718 251930 475954
rect 252166 475718 252208 475954
rect 251888 475634 252208 475718
rect 251888 475398 251930 475634
rect 252166 475398 252208 475634
rect 251888 475366 252208 475398
rect 282608 475954 282928 475986
rect 282608 475718 282650 475954
rect 282886 475718 282928 475954
rect 282608 475634 282928 475718
rect 282608 475398 282650 475634
rect 282886 475398 282928 475634
rect 282608 475366 282928 475398
rect 313328 475954 313648 475986
rect 313328 475718 313370 475954
rect 313606 475718 313648 475954
rect 313328 475634 313648 475718
rect 313328 475398 313370 475634
rect 313606 475398 313648 475634
rect 313328 475366 313648 475398
rect 344048 475954 344368 475986
rect 344048 475718 344090 475954
rect 344326 475718 344368 475954
rect 344048 475634 344368 475718
rect 344048 475398 344090 475634
rect 344326 475398 344368 475634
rect 344048 475366 344368 475398
rect 52208 471454 52528 471486
rect 52208 471218 52250 471454
rect 52486 471218 52528 471454
rect 52208 471134 52528 471218
rect 52208 470898 52250 471134
rect 52486 470898 52528 471134
rect 52208 470866 52528 470898
rect 82928 471454 83248 471486
rect 82928 471218 82970 471454
rect 83206 471218 83248 471454
rect 82928 471134 83248 471218
rect 82928 470898 82970 471134
rect 83206 470898 83248 471134
rect 82928 470866 83248 470898
rect 113648 471454 113968 471486
rect 113648 471218 113690 471454
rect 113926 471218 113968 471454
rect 113648 471134 113968 471218
rect 113648 470898 113690 471134
rect 113926 470898 113968 471134
rect 113648 470866 113968 470898
rect 144368 471454 144688 471486
rect 144368 471218 144410 471454
rect 144646 471218 144688 471454
rect 144368 471134 144688 471218
rect 144368 470898 144410 471134
rect 144646 470898 144688 471134
rect 144368 470866 144688 470898
rect 175088 471454 175408 471486
rect 175088 471218 175130 471454
rect 175366 471218 175408 471454
rect 175088 471134 175408 471218
rect 175088 470898 175130 471134
rect 175366 470898 175408 471134
rect 175088 470866 175408 470898
rect 205808 471454 206128 471486
rect 205808 471218 205850 471454
rect 206086 471218 206128 471454
rect 205808 471134 206128 471218
rect 205808 470898 205850 471134
rect 206086 470898 206128 471134
rect 205808 470866 206128 470898
rect 236528 471454 236848 471486
rect 236528 471218 236570 471454
rect 236806 471218 236848 471454
rect 236528 471134 236848 471218
rect 236528 470898 236570 471134
rect 236806 470898 236848 471134
rect 236528 470866 236848 470898
rect 267248 471454 267568 471486
rect 267248 471218 267290 471454
rect 267526 471218 267568 471454
rect 267248 471134 267568 471218
rect 267248 470898 267290 471134
rect 267526 470898 267568 471134
rect 267248 470866 267568 470898
rect 297968 471454 298288 471486
rect 297968 471218 298010 471454
rect 298246 471218 298288 471454
rect 297968 471134 298288 471218
rect 297968 470898 298010 471134
rect 298246 470898 298288 471134
rect 297968 470866 298288 470898
rect 328688 471454 329008 471486
rect 328688 471218 328730 471454
rect 328966 471218 329008 471454
rect 328688 471134 329008 471218
rect 328688 470898 328730 471134
rect 328966 470898 329008 471134
rect 328688 470866 329008 470898
rect 67568 439954 67888 439986
rect 67568 439718 67610 439954
rect 67846 439718 67888 439954
rect 67568 439634 67888 439718
rect 67568 439398 67610 439634
rect 67846 439398 67888 439634
rect 67568 439366 67888 439398
rect 98288 439954 98608 439986
rect 98288 439718 98330 439954
rect 98566 439718 98608 439954
rect 98288 439634 98608 439718
rect 98288 439398 98330 439634
rect 98566 439398 98608 439634
rect 98288 439366 98608 439398
rect 129008 439954 129328 439986
rect 129008 439718 129050 439954
rect 129286 439718 129328 439954
rect 129008 439634 129328 439718
rect 129008 439398 129050 439634
rect 129286 439398 129328 439634
rect 129008 439366 129328 439398
rect 159728 439954 160048 439986
rect 159728 439718 159770 439954
rect 160006 439718 160048 439954
rect 159728 439634 160048 439718
rect 159728 439398 159770 439634
rect 160006 439398 160048 439634
rect 159728 439366 160048 439398
rect 190448 439954 190768 439986
rect 190448 439718 190490 439954
rect 190726 439718 190768 439954
rect 190448 439634 190768 439718
rect 190448 439398 190490 439634
rect 190726 439398 190768 439634
rect 190448 439366 190768 439398
rect 221168 439954 221488 439986
rect 221168 439718 221210 439954
rect 221446 439718 221488 439954
rect 221168 439634 221488 439718
rect 221168 439398 221210 439634
rect 221446 439398 221488 439634
rect 221168 439366 221488 439398
rect 251888 439954 252208 439986
rect 251888 439718 251930 439954
rect 252166 439718 252208 439954
rect 251888 439634 252208 439718
rect 251888 439398 251930 439634
rect 252166 439398 252208 439634
rect 251888 439366 252208 439398
rect 282608 439954 282928 439986
rect 282608 439718 282650 439954
rect 282886 439718 282928 439954
rect 282608 439634 282928 439718
rect 282608 439398 282650 439634
rect 282886 439398 282928 439634
rect 282608 439366 282928 439398
rect 313328 439954 313648 439986
rect 313328 439718 313370 439954
rect 313606 439718 313648 439954
rect 313328 439634 313648 439718
rect 313328 439398 313370 439634
rect 313606 439398 313648 439634
rect 313328 439366 313648 439398
rect 344048 439954 344368 439986
rect 344048 439718 344090 439954
rect 344326 439718 344368 439954
rect 344048 439634 344368 439718
rect 344048 439398 344090 439634
rect 344326 439398 344368 439634
rect 344048 439366 344368 439398
rect 52208 435454 52528 435486
rect 52208 435218 52250 435454
rect 52486 435218 52528 435454
rect 52208 435134 52528 435218
rect 52208 434898 52250 435134
rect 52486 434898 52528 435134
rect 52208 434866 52528 434898
rect 82928 435454 83248 435486
rect 82928 435218 82970 435454
rect 83206 435218 83248 435454
rect 82928 435134 83248 435218
rect 82928 434898 82970 435134
rect 83206 434898 83248 435134
rect 82928 434866 83248 434898
rect 113648 435454 113968 435486
rect 113648 435218 113690 435454
rect 113926 435218 113968 435454
rect 113648 435134 113968 435218
rect 113648 434898 113690 435134
rect 113926 434898 113968 435134
rect 113648 434866 113968 434898
rect 144368 435454 144688 435486
rect 144368 435218 144410 435454
rect 144646 435218 144688 435454
rect 144368 435134 144688 435218
rect 144368 434898 144410 435134
rect 144646 434898 144688 435134
rect 144368 434866 144688 434898
rect 175088 435454 175408 435486
rect 175088 435218 175130 435454
rect 175366 435218 175408 435454
rect 175088 435134 175408 435218
rect 175088 434898 175130 435134
rect 175366 434898 175408 435134
rect 175088 434866 175408 434898
rect 205808 435454 206128 435486
rect 205808 435218 205850 435454
rect 206086 435218 206128 435454
rect 205808 435134 206128 435218
rect 205808 434898 205850 435134
rect 206086 434898 206128 435134
rect 205808 434866 206128 434898
rect 236528 435454 236848 435486
rect 236528 435218 236570 435454
rect 236806 435218 236848 435454
rect 236528 435134 236848 435218
rect 236528 434898 236570 435134
rect 236806 434898 236848 435134
rect 236528 434866 236848 434898
rect 267248 435454 267568 435486
rect 267248 435218 267290 435454
rect 267526 435218 267568 435454
rect 267248 435134 267568 435218
rect 267248 434898 267290 435134
rect 267526 434898 267568 435134
rect 267248 434866 267568 434898
rect 297968 435454 298288 435486
rect 297968 435218 298010 435454
rect 298246 435218 298288 435454
rect 297968 435134 298288 435218
rect 297968 434898 298010 435134
rect 298246 434898 298288 435134
rect 297968 434866 298288 434898
rect 328688 435454 329008 435486
rect 328688 435218 328730 435454
rect 328966 435218 329008 435454
rect 328688 435134 329008 435218
rect 328688 434898 328730 435134
rect 328966 434898 329008 435134
rect 328688 434866 329008 434898
rect 67568 403954 67888 403986
rect 67568 403718 67610 403954
rect 67846 403718 67888 403954
rect 67568 403634 67888 403718
rect 67568 403398 67610 403634
rect 67846 403398 67888 403634
rect 67568 403366 67888 403398
rect 98288 403954 98608 403986
rect 98288 403718 98330 403954
rect 98566 403718 98608 403954
rect 98288 403634 98608 403718
rect 98288 403398 98330 403634
rect 98566 403398 98608 403634
rect 98288 403366 98608 403398
rect 129008 403954 129328 403986
rect 129008 403718 129050 403954
rect 129286 403718 129328 403954
rect 129008 403634 129328 403718
rect 129008 403398 129050 403634
rect 129286 403398 129328 403634
rect 129008 403366 129328 403398
rect 159728 403954 160048 403986
rect 159728 403718 159770 403954
rect 160006 403718 160048 403954
rect 159728 403634 160048 403718
rect 159728 403398 159770 403634
rect 160006 403398 160048 403634
rect 159728 403366 160048 403398
rect 190448 403954 190768 403986
rect 190448 403718 190490 403954
rect 190726 403718 190768 403954
rect 190448 403634 190768 403718
rect 190448 403398 190490 403634
rect 190726 403398 190768 403634
rect 190448 403366 190768 403398
rect 221168 403954 221488 403986
rect 221168 403718 221210 403954
rect 221446 403718 221488 403954
rect 221168 403634 221488 403718
rect 221168 403398 221210 403634
rect 221446 403398 221488 403634
rect 221168 403366 221488 403398
rect 251888 403954 252208 403986
rect 251888 403718 251930 403954
rect 252166 403718 252208 403954
rect 251888 403634 252208 403718
rect 251888 403398 251930 403634
rect 252166 403398 252208 403634
rect 251888 403366 252208 403398
rect 282608 403954 282928 403986
rect 282608 403718 282650 403954
rect 282886 403718 282928 403954
rect 282608 403634 282928 403718
rect 282608 403398 282650 403634
rect 282886 403398 282928 403634
rect 282608 403366 282928 403398
rect 313328 403954 313648 403986
rect 313328 403718 313370 403954
rect 313606 403718 313648 403954
rect 313328 403634 313648 403718
rect 313328 403398 313370 403634
rect 313606 403398 313648 403634
rect 313328 403366 313648 403398
rect 344048 403954 344368 403986
rect 344048 403718 344090 403954
rect 344326 403718 344368 403954
rect 344048 403634 344368 403718
rect 344048 403398 344090 403634
rect 344326 403398 344368 403634
rect 344048 403366 344368 403398
rect 52208 399454 52528 399486
rect 52208 399218 52250 399454
rect 52486 399218 52528 399454
rect 52208 399134 52528 399218
rect 52208 398898 52250 399134
rect 52486 398898 52528 399134
rect 52208 398866 52528 398898
rect 82928 399454 83248 399486
rect 82928 399218 82970 399454
rect 83206 399218 83248 399454
rect 82928 399134 83248 399218
rect 82928 398898 82970 399134
rect 83206 398898 83248 399134
rect 82928 398866 83248 398898
rect 113648 399454 113968 399486
rect 113648 399218 113690 399454
rect 113926 399218 113968 399454
rect 113648 399134 113968 399218
rect 113648 398898 113690 399134
rect 113926 398898 113968 399134
rect 113648 398866 113968 398898
rect 144368 399454 144688 399486
rect 144368 399218 144410 399454
rect 144646 399218 144688 399454
rect 144368 399134 144688 399218
rect 144368 398898 144410 399134
rect 144646 398898 144688 399134
rect 144368 398866 144688 398898
rect 175088 399454 175408 399486
rect 175088 399218 175130 399454
rect 175366 399218 175408 399454
rect 175088 399134 175408 399218
rect 175088 398898 175130 399134
rect 175366 398898 175408 399134
rect 175088 398866 175408 398898
rect 205808 399454 206128 399486
rect 205808 399218 205850 399454
rect 206086 399218 206128 399454
rect 205808 399134 206128 399218
rect 205808 398898 205850 399134
rect 206086 398898 206128 399134
rect 205808 398866 206128 398898
rect 236528 399454 236848 399486
rect 236528 399218 236570 399454
rect 236806 399218 236848 399454
rect 236528 399134 236848 399218
rect 236528 398898 236570 399134
rect 236806 398898 236848 399134
rect 236528 398866 236848 398898
rect 267248 399454 267568 399486
rect 267248 399218 267290 399454
rect 267526 399218 267568 399454
rect 267248 399134 267568 399218
rect 267248 398898 267290 399134
rect 267526 398898 267568 399134
rect 267248 398866 267568 398898
rect 297968 399454 298288 399486
rect 297968 399218 298010 399454
rect 298246 399218 298288 399454
rect 297968 399134 298288 399218
rect 297968 398898 298010 399134
rect 298246 398898 298288 399134
rect 297968 398866 298288 398898
rect 328688 399454 329008 399486
rect 328688 399218 328730 399454
rect 328966 399218 329008 399454
rect 328688 399134 329008 399218
rect 328688 398898 328730 399134
rect 328966 398898 329008 399134
rect 328688 398866 329008 398898
rect 47715 378248 47781 378249
rect 47715 378184 47716 378248
rect 47780 378184 47781 378248
rect 47715 378183 47781 378184
rect 47531 288488 47597 288489
rect 47531 288424 47532 288488
rect 47596 288424 47597 288488
rect 47531 288423 47597 288424
rect 47163 229396 47229 229397
rect 47163 229332 47164 229396
rect 47228 229332 47229 229396
rect 47163 229331 47229 229332
rect 47163 220828 47229 220829
rect 47163 220764 47164 220828
rect 47228 220764 47229 220828
rect 47163 220763 47229 220764
rect 46979 220556 47045 220557
rect 46979 220492 46980 220556
rect 47044 220492 47045 220556
rect 46979 220491 47045 220492
rect 47166 209541 47226 220763
rect 47163 209540 47229 209541
rect 47163 209476 47164 209540
rect 47228 209476 47229 209540
rect 47163 209475 47229 209476
rect 46794 192454 47414 198000
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46611 155412 46677 155413
rect 46611 155348 46612 155412
rect 46676 155348 46677 155412
rect 46611 155347 46677 155348
rect 46611 150516 46677 150517
rect 46611 150452 46612 150516
rect 46676 150452 46677 150516
rect 46611 150451 46677 150452
rect 46614 35053 46674 150451
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46611 35052 46677 35053
rect 46611 34988 46612 35052
rect 46676 34988 46677 35052
rect 46611 34987 46677 34988
rect 46427 21860 46493 21861
rect 46427 21796 46428 21860
rect 46492 21796 46493 21860
rect 46427 21795 46493 21796
rect 46794 12454 47414 47898
rect 47534 26077 47594 288423
rect 47718 181525 47778 378183
rect 67568 367954 67888 367986
rect 67568 367718 67610 367954
rect 67846 367718 67888 367954
rect 67568 367634 67888 367718
rect 67568 367398 67610 367634
rect 67846 367398 67888 367634
rect 67568 367366 67888 367398
rect 98288 367954 98608 367986
rect 98288 367718 98330 367954
rect 98566 367718 98608 367954
rect 98288 367634 98608 367718
rect 98288 367398 98330 367634
rect 98566 367398 98608 367634
rect 98288 367366 98608 367398
rect 129008 367954 129328 367986
rect 129008 367718 129050 367954
rect 129286 367718 129328 367954
rect 129008 367634 129328 367718
rect 129008 367398 129050 367634
rect 129286 367398 129328 367634
rect 129008 367366 129328 367398
rect 159728 367954 160048 367986
rect 159728 367718 159770 367954
rect 160006 367718 160048 367954
rect 159728 367634 160048 367718
rect 159728 367398 159770 367634
rect 160006 367398 160048 367634
rect 159728 367366 160048 367398
rect 190448 367954 190768 367986
rect 190448 367718 190490 367954
rect 190726 367718 190768 367954
rect 190448 367634 190768 367718
rect 190448 367398 190490 367634
rect 190726 367398 190768 367634
rect 190448 367366 190768 367398
rect 221168 367954 221488 367986
rect 221168 367718 221210 367954
rect 221446 367718 221488 367954
rect 221168 367634 221488 367718
rect 221168 367398 221210 367634
rect 221446 367398 221488 367634
rect 221168 367366 221488 367398
rect 251888 367954 252208 367986
rect 251888 367718 251930 367954
rect 252166 367718 252208 367954
rect 251888 367634 252208 367718
rect 251888 367398 251930 367634
rect 252166 367398 252208 367634
rect 251888 367366 252208 367398
rect 282608 367954 282928 367986
rect 282608 367718 282650 367954
rect 282886 367718 282928 367954
rect 282608 367634 282928 367718
rect 282608 367398 282650 367634
rect 282886 367398 282928 367634
rect 282608 367366 282928 367398
rect 313328 367954 313648 367986
rect 313328 367718 313370 367954
rect 313606 367718 313648 367954
rect 313328 367634 313648 367718
rect 313328 367398 313370 367634
rect 313606 367398 313648 367634
rect 313328 367366 313648 367398
rect 344048 367954 344368 367986
rect 344048 367718 344090 367954
rect 344326 367718 344368 367954
rect 344048 367634 344368 367718
rect 344048 367398 344090 367634
rect 344326 367398 344368 367634
rect 344048 367366 344368 367398
rect 52208 363454 52528 363486
rect 52208 363218 52250 363454
rect 52486 363218 52528 363454
rect 52208 363134 52528 363218
rect 52208 362898 52250 363134
rect 52486 362898 52528 363134
rect 52208 362866 52528 362898
rect 82928 363454 83248 363486
rect 82928 363218 82970 363454
rect 83206 363218 83248 363454
rect 82928 363134 83248 363218
rect 82928 362898 82970 363134
rect 83206 362898 83248 363134
rect 82928 362866 83248 362898
rect 113648 363454 113968 363486
rect 113648 363218 113690 363454
rect 113926 363218 113968 363454
rect 113648 363134 113968 363218
rect 113648 362898 113690 363134
rect 113926 362898 113968 363134
rect 113648 362866 113968 362898
rect 144368 363454 144688 363486
rect 144368 363218 144410 363454
rect 144646 363218 144688 363454
rect 144368 363134 144688 363218
rect 144368 362898 144410 363134
rect 144646 362898 144688 363134
rect 144368 362866 144688 362898
rect 175088 363454 175408 363486
rect 175088 363218 175130 363454
rect 175366 363218 175408 363454
rect 175088 363134 175408 363218
rect 175088 362898 175130 363134
rect 175366 362898 175408 363134
rect 175088 362866 175408 362898
rect 205808 363454 206128 363486
rect 205808 363218 205850 363454
rect 206086 363218 206128 363454
rect 205808 363134 206128 363218
rect 205808 362898 205850 363134
rect 206086 362898 206128 363134
rect 205808 362866 206128 362898
rect 236528 363454 236848 363486
rect 236528 363218 236570 363454
rect 236806 363218 236848 363454
rect 236528 363134 236848 363218
rect 236528 362898 236570 363134
rect 236806 362898 236848 363134
rect 236528 362866 236848 362898
rect 267248 363454 267568 363486
rect 267248 363218 267290 363454
rect 267526 363218 267568 363454
rect 267248 363134 267568 363218
rect 267248 362898 267290 363134
rect 267526 362898 267568 363134
rect 267248 362866 267568 362898
rect 297968 363454 298288 363486
rect 297968 363218 298010 363454
rect 298246 363218 298288 363454
rect 297968 363134 298288 363218
rect 297968 362898 298010 363134
rect 298246 362898 298288 363134
rect 297968 362866 298288 362898
rect 328688 363454 329008 363486
rect 328688 363218 328730 363454
rect 328966 363218 329008 363454
rect 328688 363134 329008 363218
rect 328688 362898 328730 363134
rect 328966 362898 329008 363134
rect 328688 362866 329008 362898
rect 67568 331954 67888 331986
rect 67568 331718 67610 331954
rect 67846 331718 67888 331954
rect 67568 331634 67888 331718
rect 67568 331398 67610 331634
rect 67846 331398 67888 331634
rect 67568 331366 67888 331398
rect 98288 331954 98608 331986
rect 98288 331718 98330 331954
rect 98566 331718 98608 331954
rect 98288 331634 98608 331718
rect 98288 331398 98330 331634
rect 98566 331398 98608 331634
rect 98288 331366 98608 331398
rect 129008 331954 129328 331986
rect 129008 331718 129050 331954
rect 129286 331718 129328 331954
rect 129008 331634 129328 331718
rect 129008 331398 129050 331634
rect 129286 331398 129328 331634
rect 129008 331366 129328 331398
rect 159728 331954 160048 331986
rect 159728 331718 159770 331954
rect 160006 331718 160048 331954
rect 159728 331634 160048 331718
rect 159728 331398 159770 331634
rect 160006 331398 160048 331634
rect 159728 331366 160048 331398
rect 190448 331954 190768 331986
rect 190448 331718 190490 331954
rect 190726 331718 190768 331954
rect 190448 331634 190768 331718
rect 190448 331398 190490 331634
rect 190726 331398 190768 331634
rect 190448 331366 190768 331398
rect 221168 331954 221488 331986
rect 221168 331718 221210 331954
rect 221446 331718 221488 331954
rect 221168 331634 221488 331718
rect 221168 331398 221210 331634
rect 221446 331398 221488 331634
rect 221168 331366 221488 331398
rect 251888 331954 252208 331986
rect 251888 331718 251930 331954
rect 252166 331718 252208 331954
rect 251888 331634 252208 331718
rect 251888 331398 251930 331634
rect 252166 331398 252208 331634
rect 251888 331366 252208 331398
rect 282608 331954 282928 331986
rect 282608 331718 282650 331954
rect 282886 331718 282928 331954
rect 282608 331634 282928 331718
rect 282608 331398 282650 331634
rect 282886 331398 282928 331634
rect 282608 331366 282928 331398
rect 313328 331954 313648 331986
rect 313328 331718 313370 331954
rect 313606 331718 313648 331954
rect 313328 331634 313648 331718
rect 313328 331398 313370 331634
rect 313606 331398 313648 331634
rect 313328 331366 313648 331398
rect 344048 331954 344368 331986
rect 344048 331718 344090 331954
rect 344326 331718 344368 331954
rect 344048 331634 344368 331718
rect 344048 331398 344090 331634
rect 344326 331398 344368 331634
rect 344048 331366 344368 331398
rect 52208 327454 52528 327486
rect 52208 327218 52250 327454
rect 52486 327218 52528 327454
rect 52208 327134 52528 327218
rect 52208 326898 52250 327134
rect 52486 326898 52528 327134
rect 52208 326866 52528 326898
rect 82928 327454 83248 327486
rect 82928 327218 82970 327454
rect 83206 327218 83248 327454
rect 82928 327134 83248 327218
rect 82928 326898 82970 327134
rect 83206 326898 83248 327134
rect 82928 326866 83248 326898
rect 113648 327454 113968 327486
rect 113648 327218 113690 327454
rect 113926 327218 113968 327454
rect 113648 327134 113968 327218
rect 113648 326898 113690 327134
rect 113926 326898 113968 327134
rect 113648 326866 113968 326898
rect 144368 327454 144688 327486
rect 144368 327218 144410 327454
rect 144646 327218 144688 327454
rect 144368 327134 144688 327218
rect 144368 326898 144410 327134
rect 144646 326898 144688 327134
rect 144368 326866 144688 326898
rect 175088 327454 175408 327486
rect 175088 327218 175130 327454
rect 175366 327218 175408 327454
rect 175088 327134 175408 327218
rect 175088 326898 175130 327134
rect 175366 326898 175408 327134
rect 175088 326866 175408 326898
rect 205808 327454 206128 327486
rect 205808 327218 205850 327454
rect 206086 327218 206128 327454
rect 205808 327134 206128 327218
rect 205808 326898 205850 327134
rect 206086 326898 206128 327134
rect 205808 326866 206128 326898
rect 236528 327454 236848 327486
rect 236528 327218 236570 327454
rect 236806 327218 236848 327454
rect 236528 327134 236848 327218
rect 236528 326898 236570 327134
rect 236806 326898 236848 327134
rect 236528 326866 236848 326898
rect 267248 327454 267568 327486
rect 267248 327218 267290 327454
rect 267526 327218 267568 327454
rect 267248 327134 267568 327218
rect 267248 326898 267290 327134
rect 267526 326898 267568 327134
rect 267248 326866 267568 326898
rect 297968 327454 298288 327486
rect 297968 327218 298010 327454
rect 298246 327218 298288 327454
rect 297968 327134 298288 327218
rect 297968 326898 298010 327134
rect 298246 326898 298288 327134
rect 297968 326866 298288 326898
rect 328688 327454 329008 327486
rect 328688 327218 328730 327454
rect 328966 327218 329008 327454
rect 328688 327134 329008 327218
rect 328688 326898 328730 327134
rect 328966 326898 329008 327134
rect 328688 326866 329008 326898
rect 67568 295954 67888 295986
rect 67568 295718 67610 295954
rect 67846 295718 67888 295954
rect 67568 295634 67888 295718
rect 67568 295398 67610 295634
rect 67846 295398 67888 295634
rect 67568 295366 67888 295398
rect 98288 295954 98608 295986
rect 98288 295718 98330 295954
rect 98566 295718 98608 295954
rect 98288 295634 98608 295718
rect 98288 295398 98330 295634
rect 98566 295398 98608 295634
rect 98288 295366 98608 295398
rect 129008 295954 129328 295986
rect 129008 295718 129050 295954
rect 129286 295718 129328 295954
rect 129008 295634 129328 295718
rect 129008 295398 129050 295634
rect 129286 295398 129328 295634
rect 129008 295366 129328 295398
rect 159728 295954 160048 295986
rect 159728 295718 159770 295954
rect 160006 295718 160048 295954
rect 159728 295634 160048 295718
rect 159728 295398 159770 295634
rect 160006 295398 160048 295634
rect 159728 295366 160048 295398
rect 190448 295954 190768 295986
rect 190448 295718 190490 295954
rect 190726 295718 190768 295954
rect 190448 295634 190768 295718
rect 190448 295398 190490 295634
rect 190726 295398 190768 295634
rect 190448 295366 190768 295398
rect 221168 295954 221488 295986
rect 221168 295718 221210 295954
rect 221446 295718 221488 295954
rect 221168 295634 221488 295718
rect 221168 295398 221210 295634
rect 221446 295398 221488 295634
rect 221168 295366 221488 295398
rect 251888 295954 252208 295986
rect 251888 295718 251930 295954
rect 252166 295718 252208 295954
rect 251888 295634 252208 295718
rect 251888 295398 251930 295634
rect 252166 295398 252208 295634
rect 251888 295366 252208 295398
rect 282608 295954 282928 295986
rect 282608 295718 282650 295954
rect 282886 295718 282928 295954
rect 282608 295634 282928 295718
rect 282608 295398 282650 295634
rect 282886 295398 282928 295634
rect 282608 295366 282928 295398
rect 313328 295954 313648 295986
rect 313328 295718 313370 295954
rect 313606 295718 313648 295954
rect 313328 295634 313648 295718
rect 313328 295398 313370 295634
rect 313606 295398 313648 295634
rect 313328 295366 313648 295398
rect 344048 295954 344368 295986
rect 344048 295718 344090 295954
rect 344326 295718 344368 295954
rect 344048 295634 344368 295718
rect 344048 295398 344090 295634
rect 344326 295398 344368 295634
rect 344048 295366 344368 295398
rect 52208 291454 52528 291486
rect 52208 291218 52250 291454
rect 52486 291218 52528 291454
rect 52208 291134 52528 291218
rect 52208 290898 52250 291134
rect 52486 290898 52528 291134
rect 52208 290866 52528 290898
rect 82928 291454 83248 291486
rect 82928 291218 82970 291454
rect 83206 291218 83248 291454
rect 82928 291134 83248 291218
rect 82928 290898 82970 291134
rect 83206 290898 83248 291134
rect 82928 290866 83248 290898
rect 113648 291454 113968 291486
rect 113648 291218 113690 291454
rect 113926 291218 113968 291454
rect 113648 291134 113968 291218
rect 113648 290898 113690 291134
rect 113926 290898 113968 291134
rect 113648 290866 113968 290898
rect 144368 291454 144688 291486
rect 144368 291218 144410 291454
rect 144646 291218 144688 291454
rect 144368 291134 144688 291218
rect 144368 290898 144410 291134
rect 144646 290898 144688 291134
rect 144368 290866 144688 290898
rect 175088 291454 175408 291486
rect 175088 291218 175130 291454
rect 175366 291218 175408 291454
rect 175088 291134 175408 291218
rect 175088 290898 175130 291134
rect 175366 290898 175408 291134
rect 175088 290866 175408 290898
rect 205808 291454 206128 291486
rect 205808 291218 205850 291454
rect 206086 291218 206128 291454
rect 205808 291134 206128 291218
rect 205808 290898 205850 291134
rect 206086 290898 206128 291134
rect 205808 290866 206128 290898
rect 236528 291454 236848 291486
rect 236528 291218 236570 291454
rect 236806 291218 236848 291454
rect 236528 291134 236848 291218
rect 236528 290898 236570 291134
rect 236806 290898 236848 291134
rect 236528 290866 236848 290898
rect 267248 291454 267568 291486
rect 267248 291218 267290 291454
rect 267526 291218 267568 291454
rect 267248 291134 267568 291218
rect 267248 290898 267290 291134
rect 267526 290898 267568 291134
rect 267248 290866 267568 290898
rect 297968 291454 298288 291486
rect 297968 291218 298010 291454
rect 298246 291218 298288 291454
rect 297968 291134 298288 291218
rect 297968 290898 298010 291134
rect 298246 290898 298288 291134
rect 297968 290866 298288 290898
rect 328688 291454 329008 291486
rect 328688 291218 328730 291454
rect 328966 291218 329008 291454
rect 328688 291134 329008 291218
rect 328688 290898 328730 291134
rect 328966 290898 329008 291134
rect 328688 290866 329008 290898
rect 67568 259954 67888 259986
rect 67568 259718 67610 259954
rect 67846 259718 67888 259954
rect 67568 259634 67888 259718
rect 67568 259398 67610 259634
rect 67846 259398 67888 259634
rect 67568 259366 67888 259398
rect 98288 259954 98608 259986
rect 98288 259718 98330 259954
rect 98566 259718 98608 259954
rect 98288 259634 98608 259718
rect 98288 259398 98330 259634
rect 98566 259398 98608 259634
rect 98288 259366 98608 259398
rect 129008 259954 129328 259986
rect 129008 259718 129050 259954
rect 129286 259718 129328 259954
rect 129008 259634 129328 259718
rect 129008 259398 129050 259634
rect 129286 259398 129328 259634
rect 129008 259366 129328 259398
rect 159728 259954 160048 259986
rect 159728 259718 159770 259954
rect 160006 259718 160048 259954
rect 159728 259634 160048 259718
rect 159728 259398 159770 259634
rect 160006 259398 160048 259634
rect 159728 259366 160048 259398
rect 190448 259954 190768 259986
rect 190448 259718 190490 259954
rect 190726 259718 190768 259954
rect 190448 259634 190768 259718
rect 190448 259398 190490 259634
rect 190726 259398 190768 259634
rect 190448 259366 190768 259398
rect 221168 259954 221488 259986
rect 221168 259718 221210 259954
rect 221446 259718 221488 259954
rect 221168 259634 221488 259718
rect 221168 259398 221210 259634
rect 221446 259398 221488 259634
rect 221168 259366 221488 259398
rect 251888 259954 252208 259986
rect 251888 259718 251930 259954
rect 252166 259718 252208 259954
rect 251888 259634 252208 259718
rect 251888 259398 251930 259634
rect 252166 259398 252208 259634
rect 251888 259366 252208 259398
rect 282608 259954 282928 259986
rect 282608 259718 282650 259954
rect 282886 259718 282928 259954
rect 282608 259634 282928 259718
rect 282608 259398 282650 259634
rect 282886 259398 282928 259634
rect 282608 259366 282928 259398
rect 313328 259954 313648 259986
rect 313328 259718 313370 259954
rect 313606 259718 313648 259954
rect 313328 259634 313648 259718
rect 313328 259398 313370 259634
rect 313606 259398 313648 259634
rect 313328 259366 313648 259398
rect 344048 259954 344368 259986
rect 344048 259718 344090 259954
rect 344326 259718 344368 259954
rect 344048 259634 344368 259718
rect 344048 259398 344090 259634
rect 344326 259398 344368 259634
rect 344048 259366 344368 259398
rect 52208 255454 52528 255486
rect 52208 255218 52250 255454
rect 52486 255218 52528 255454
rect 52208 255134 52528 255218
rect 52208 254898 52250 255134
rect 52486 254898 52528 255134
rect 52208 254866 52528 254898
rect 82928 255454 83248 255486
rect 82928 255218 82970 255454
rect 83206 255218 83248 255454
rect 82928 255134 83248 255218
rect 82928 254898 82970 255134
rect 83206 254898 83248 255134
rect 82928 254866 83248 254898
rect 113648 255454 113968 255486
rect 113648 255218 113690 255454
rect 113926 255218 113968 255454
rect 113648 255134 113968 255218
rect 113648 254898 113690 255134
rect 113926 254898 113968 255134
rect 113648 254866 113968 254898
rect 144368 255454 144688 255486
rect 144368 255218 144410 255454
rect 144646 255218 144688 255454
rect 144368 255134 144688 255218
rect 144368 254898 144410 255134
rect 144646 254898 144688 255134
rect 144368 254866 144688 254898
rect 175088 255454 175408 255486
rect 175088 255218 175130 255454
rect 175366 255218 175408 255454
rect 175088 255134 175408 255218
rect 175088 254898 175130 255134
rect 175366 254898 175408 255134
rect 175088 254866 175408 254898
rect 205808 255454 206128 255486
rect 205808 255218 205850 255454
rect 206086 255218 206128 255454
rect 205808 255134 206128 255218
rect 205808 254898 205850 255134
rect 206086 254898 206128 255134
rect 205808 254866 206128 254898
rect 236528 255454 236848 255486
rect 236528 255218 236570 255454
rect 236806 255218 236848 255454
rect 236528 255134 236848 255218
rect 236528 254898 236570 255134
rect 236806 254898 236848 255134
rect 236528 254866 236848 254898
rect 267248 255454 267568 255486
rect 267248 255218 267290 255454
rect 267526 255218 267568 255454
rect 267248 255134 267568 255218
rect 267248 254898 267290 255134
rect 267526 254898 267568 255134
rect 267248 254866 267568 254898
rect 297968 255454 298288 255486
rect 297968 255218 298010 255454
rect 298246 255218 298288 255454
rect 297968 255134 298288 255218
rect 297968 254898 298010 255134
rect 298246 254898 298288 255134
rect 297968 254866 298288 254898
rect 328688 255454 329008 255486
rect 328688 255218 328730 255454
rect 328966 255218 329008 255454
rect 328688 255134 329008 255218
rect 328688 254898 328730 255134
rect 328966 254898 329008 255134
rect 328688 254866 329008 254898
rect 47899 229804 47965 229805
rect 47899 229740 47900 229804
rect 47964 229740 47965 229804
rect 47899 229739 47965 229740
rect 47902 201245 47962 229739
rect 67568 223954 67888 223986
rect 67568 223718 67610 223954
rect 67846 223718 67888 223954
rect 67568 223634 67888 223718
rect 67568 223398 67610 223634
rect 67846 223398 67888 223634
rect 67568 223366 67888 223398
rect 98288 223954 98608 223986
rect 98288 223718 98330 223954
rect 98566 223718 98608 223954
rect 98288 223634 98608 223718
rect 98288 223398 98330 223634
rect 98566 223398 98608 223634
rect 98288 223366 98608 223398
rect 129008 223954 129328 223986
rect 129008 223718 129050 223954
rect 129286 223718 129328 223954
rect 129008 223634 129328 223718
rect 129008 223398 129050 223634
rect 129286 223398 129328 223634
rect 129008 223366 129328 223398
rect 159728 223954 160048 223986
rect 159728 223718 159770 223954
rect 160006 223718 160048 223954
rect 159728 223634 160048 223718
rect 159728 223398 159770 223634
rect 160006 223398 160048 223634
rect 159728 223366 160048 223398
rect 190448 223954 190768 223986
rect 190448 223718 190490 223954
rect 190726 223718 190768 223954
rect 190448 223634 190768 223718
rect 190448 223398 190490 223634
rect 190726 223398 190768 223634
rect 190448 223366 190768 223398
rect 221168 223954 221488 223986
rect 221168 223718 221210 223954
rect 221446 223718 221488 223954
rect 221168 223634 221488 223718
rect 221168 223398 221210 223634
rect 221446 223398 221488 223634
rect 221168 223366 221488 223398
rect 251888 223954 252208 223986
rect 251888 223718 251930 223954
rect 252166 223718 252208 223954
rect 251888 223634 252208 223718
rect 251888 223398 251930 223634
rect 252166 223398 252208 223634
rect 251888 223366 252208 223398
rect 282608 223954 282928 223986
rect 282608 223718 282650 223954
rect 282886 223718 282928 223954
rect 282608 223634 282928 223718
rect 282608 223398 282650 223634
rect 282886 223398 282928 223634
rect 282608 223366 282928 223398
rect 313328 223954 313648 223986
rect 313328 223718 313370 223954
rect 313606 223718 313648 223954
rect 313328 223634 313648 223718
rect 313328 223398 313370 223634
rect 313606 223398 313648 223634
rect 313328 223366 313648 223398
rect 344048 223954 344368 223986
rect 344048 223718 344090 223954
rect 344326 223718 344368 223954
rect 344048 223634 344368 223718
rect 344048 223398 344090 223634
rect 344326 223398 344368 223634
rect 344048 223366 344368 223398
rect 52208 219454 52528 219486
rect 52208 219218 52250 219454
rect 52486 219218 52528 219454
rect 52208 219134 52528 219218
rect 52208 218898 52250 219134
rect 52486 218898 52528 219134
rect 52208 218866 52528 218898
rect 82928 219454 83248 219486
rect 82928 219218 82970 219454
rect 83206 219218 83248 219454
rect 82928 219134 83248 219218
rect 82928 218898 82970 219134
rect 83206 218898 83248 219134
rect 82928 218866 83248 218898
rect 113648 219454 113968 219486
rect 113648 219218 113690 219454
rect 113926 219218 113968 219454
rect 113648 219134 113968 219218
rect 113648 218898 113690 219134
rect 113926 218898 113968 219134
rect 113648 218866 113968 218898
rect 144368 219454 144688 219486
rect 144368 219218 144410 219454
rect 144646 219218 144688 219454
rect 144368 219134 144688 219218
rect 144368 218898 144410 219134
rect 144646 218898 144688 219134
rect 144368 218866 144688 218898
rect 175088 219454 175408 219486
rect 175088 219218 175130 219454
rect 175366 219218 175408 219454
rect 175088 219134 175408 219218
rect 175088 218898 175130 219134
rect 175366 218898 175408 219134
rect 175088 218866 175408 218898
rect 205808 219454 206128 219486
rect 205808 219218 205850 219454
rect 206086 219218 206128 219454
rect 205808 219134 206128 219218
rect 205808 218898 205850 219134
rect 206086 218898 206128 219134
rect 205808 218866 206128 218898
rect 236528 219454 236848 219486
rect 236528 219218 236570 219454
rect 236806 219218 236848 219454
rect 236528 219134 236848 219218
rect 236528 218898 236570 219134
rect 236806 218898 236848 219134
rect 236528 218866 236848 218898
rect 267248 219454 267568 219486
rect 267248 219218 267290 219454
rect 267526 219218 267568 219454
rect 267248 219134 267568 219218
rect 267248 218898 267290 219134
rect 267526 218898 267568 219134
rect 267248 218866 267568 218898
rect 297968 219454 298288 219486
rect 297968 219218 298010 219454
rect 298246 219218 298288 219454
rect 297968 219134 298288 219218
rect 297968 218898 298010 219134
rect 298246 218898 298288 219134
rect 297968 218866 298288 218898
rect 328688 219454 329008 219486
rect 328688 219218 328730 219454
rect 328966 219218 329008 219454
rect 328688 219134 329008 219218
rect 328688 218898 328730 219134
rect 328966 218898 329008 219134
rect 328688 218866 329008 218898
rect 48083 209676 48149 209677
rect 48083 209612 48084 209676
rect 48148 209612 48149 209676
rect 48083 209611 48149 209612
rect 47899 201244 47965 201245
rect 47899 201180 47900 201244
rect 47964 201180 47965 201244
rect 47899 201179 47965 201180
rect 48086 195533 48146 209611
rect 347454 201590 347698 201650
rect 48267 200972 48333 200973
rect 48267 200908 48268 200972
rect 48332 200970 48333 200972
rect 48332 200910 49250 200970
rect 48332 200908 48333 200910
rect 48267 200907 48333 200908
rect 48267 200564 48333 200565
rect 48267 200500 48268 200564
rect 48332 200500 48333 200564
rect 48267 200499 48333 200500
rect 48270 200290 48330 200499
rect 48270 200230 49066 200290
rect 48267 200156 48333 200157
rect 48267 200092 48268 200156
rect 48332 200130 48333 200156
rect 48332 200092 48882 200130
rect 48267 200091 48882 200092
rect 48270 200070 48882 200091
rect 48083 195532 48149 195533
rect 48083 195468 48084 195532
rect 48148 195468 48149 195532
rect 48083 195467 48149 195468
rect 47715 181524 47781 181525
rect 47715 181460 47716 181524
rect 47780 181460 47781 181524
rect 47715 181459 47781 181460
rect 48083 176492 48149 176493
rect 48083 176428 48084 176492
rect 48148 176428 48149 176492
rect 48083 176427 48149 176428
rect 47531 26076 47597 26077
rect 47531 26012 47532 26076
rect 47596 26012 47597 26076
rect 47531 26011 47597 26012
rect 48086 23221 48146 176427
rect 48822 28389 48882 200070
rect 49006 29341 49066 200230
rect 49190 192949 49250 200910
rect 346899 199340 346965 199341
rect 346899 199276 346900 199340
rect 346964 199276 346965 199340
rect 346899 199275 346965 199276
rect 51294 196954 51914 198000
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 49187 192948 49253 192949
rect 49187 192884 49188 192948
rect 49252 192884 49253 192948
rect 49187 192883 49253 192884
rect 50843 184244 50909 184245
rect 50843 184180 50844 184244
rect 50908 184180 50909 184244
rect 50843 184179 50909 184180
rect 49555 183156 49621 183157
rect 49555 183092 49556 183156
rect 49620 183092 49621 183156
rect 49555 183091 49621 183092
rect 49371 179076 49437 179077
rect 49371 179012 49372 179076
rect 49436 179012 49437 179076
rect 49371 179011 49437 179012
rect 49003 29340 49069 29341
rect 49003 29276 49004 29340
rect 49068 29276 49069 29340
rect 49003 29275 49069 29276
rect 49374 29205 49434 179011
rect 49371 29204 49437 29205
rect 49371 29140 49372 29204
rect 49436 29140 49437 29204
rect 49371 29139 49437 29140
rect 48819 28388 48885 28389
rect 48819 28324 48820 28388
rect 48884 28324 48885 28388
rect 48819 28323 48885 28324
rect 48083 23220 48149 23221
rect 48083 23156 48084 23220
rect 48148 23156 48149 23220
rect 48083 23155 48149 23156
rect 49558 22677 49618 183091
rect 50659 180436 50725 180437
rect 50659 180372 50660 180436
rect 50724 180372 50725 180436
rect 50659 180371 50725 180372
rect 50475 170372 50541 170373
rect 50475 170308 50476 170372
rect 50540 170308 50541 170372
rect 50475 170307 50541 170308
rect 50291 155820 50357 155821
rect 50291 155756 50292 155820
rect 50356 155756 50357 155820
rect 50291 155755 50357 155756
rect 49555 22676 49621 22677
rect 49555 22612 49556 22676
rect 49620 22612 49621 22676
rect 49555 22611 49621 22612
rect 50294 21181 50354 155755
rect 50478 24445 50538 170307
rect 50662 27573 50722 180371
rect 50659 27572 50725 27573
rect 50659 27508 50660 27572
rect 50724 27508 50725 27572
rect 50659 27507 50725 27508
rect 50475 24444 50541 24445
rect 50475 24380 50476 24444
rect 50540 24380 50541 24444
rect 50475 24379 50541 24380
rect 50291 21180 50357 21181
rect 50291 21116 50292 21180
rect 50356 21116 50357 21180
rect 50291 21115 50357 21116
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 43667 3500 43733 3501
rect 43667 3436 43668 3500
rect 43732 3436 43733 3500
rect 43667 3435 43733 3436
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 -2266 47414 11898
rect 50846 3501 50906 184179
rect 51294 160954 51914 196398
rect 53051 193900 53117 193901
rect 53051 193836 53052 193900
rect 53116 193836 53117 193900
rect 53051 193835 53117 193836
rect 52315 181660 52381 181661
rect 52315 181596 52316 181660
rect 52380 181596 52381 181660
rect 52315 181595 52381 181596
rect 52131 177580 52197 177581
rect 52131 177516 52132 177580
rect 52196 177516 52197 177580
rect 52131 177515 52197 177516
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 52134 25669 52194 177515
rect 52131 25668 52197 25669
rect 52131 25604 52132 25668
rect 52196 25604 52197 25668
rect 52131 25603 52197 25604
rect 52318 24853 52378 181595
rect 53054 44301 53114 193835
rect 53419 192812 53485 192813
rect 53419 192748 53420 192812
rect 53484 192748 53485 192812
rect 53419 192747 53485 192748
rect 53235 176356 53301 176357
rect 53235 176292 53236 176356
rect 53300 176292 53301 176356
rect 53235 176291 53301 176292
rect 53051 44300 53117 44301
rect 53051 44236 53052 44300
rect 53116 44236 53117 44300
rect 53051 44235 53117 44236
rect 53238 27301 53298 176291
rect 53235 27300 53301 27301
rect 53235 27236 53236 27300
rect 53300 27236 53301 27300
rect 53235 27235 53301 27236
rect 53422 25805 53482 192747
rect 54891 191044 54957 191045
rect 54891 190980 54892 191044
rect 54956 190980 54957 191044
rect 54891 190979 54957 190980
rect 54523 189820 54589 189821
rect 54523 189756 54524 189820
rect 54588 189756 54589 189820
rect 54523 189755 54589 189756
rect 53603 174860 53669 174861
rect 53603 174796 53604 174860
rect 53668 174796 53669 174860
rect 53603 174795 53669 174796
rect 53419 25804 53485 25805
rect 53419 25740 53420 25804
rect 53484 25740 53485 25804
rect 53419 25739 53485 25740
rect 52315 24852 52381 24853
rect 52315 24788 52316 24852
rect 52380 24788 52381 24852
rect 52315 24787 52381 24788
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 50843 3500 50909 3501
rect 50843 3436 50844 3500
rect 50908 3436 50909 3500
rect 50843 3435 50909 3436
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 -3226 51914 16398
rect 53606 4045 53666 174795
rect 54526 28253 54586 189755
rect 54707 188460 54773 188461
rect 54707 188396 54708 188460
rect 54772 188396 54773 188460
rect 54707 188395 54773 188396
rect 54523 28252 54589 28253
rect 54523 28188 54524 28252
rect 54588 28188 54589 28252
rect 54523 28187 54589 28188
rect 54710 25533 54770 188395
rect 54894 25941 54954 190979
rect 55075 187372 55141 187373
rect 55075 187308 55076 187372
rect 55140 187308 55141 187372
rect 55075 187307 55141 187308
rect 54891 25940 54957 25941
rect 54891 25876 54892 25940
rect 54956 25876 54957 25940
rect 54891 25875 54957 25876
rect 54707 25532 54773 25533
rect 54707 25468 54708 25532
rect 54772 25468 54773 25532
rect 54707 25467 54773 25468
rect 53603 4044 53669 4045
rect 53603 3980 53604 4044
rect 53668 3980 53669 4044
rect 53603 3979 53669 3980
rect 55078 3365 55138 187307
rect 55627 174588 55693 174589
rect 55627 174524 55628 174588
rect 55692 174524 55693 174588
rect 55627 174523 55693 174524
rect 55443 132564 55509 132565
rect 55443 132500 55444 132564
rect 55508 132500 55509 132564
rect 55443 132499 55509 132500
rect 55446 21589 55506 132499
rect 55443 21588 55509 21589
rect 55443 21524 55444 21588
rect 55508 21524 55509 21588
rect 55443 21523 55509 21524
rect 55630 3909 55690 174523
rect 55794 165454 56414 198000
rect 59123 196620 59189 196621
rect 59123 196556 59124 196620
rect 59188 196556 59189 196620
rect 59123 196555 59189 196556
rect 57651 194036 57717 194037
rect 57651 193972 57652 194036
rect 57716 193972 57717 194036
rect 57651 193971 57717 193972
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57467 159492 57533 159493
rect 57467 159428 57468 159492
rect 57532 159428 57533 159492
rect 57467 159427 57533 159428
rect 57283 153780 57349 153781
rect 57283 153716 57284 153780
rect 57348 153716 57349 153780
rect 57283 153715 57349 153716
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 57286 34917 57346 153715
rect 57470 75037 57530 159427
rect 57654 143037 57714 193971
rect 58571 184652 58637 184653
rect 58571 184588 58572 184652
rect 58636 184588 58637 184652
rect 58571 184587 58637 184588
rect 57835 181796 57901 181797
rect 57835 181732 57836 181796
rect 57900 181732 57901 181796
rect 57835 181731 57901 181732
rect 57651 143036 57717 143037
rect 57651 142972 57652 143036
rect 57716 142972 57717 143036
rect 57651 142971 57717 142972
rect 57467 75036 57533 75037
rect 57467 74972 57468 75036
rect 57532 74972 57533 75036
rect 57467 74971 57533 74972
rect 57838 49197 57898 181731
rect 58387 138684 58453 138685
rect 58387 138620 58388 138684
rect 58452 138620 58453 138684
rect 58387 138619 58453 138620
rect 58390 132510 58450 138619
rect 58574 138141 58634 184587
rect 58755 167924 58821 167925
rect 58755 167860 58756 167924
rect 58820 167860 58821 167924
rect 58755 167859 58821 167860
rect 58571 138140 58637 138141
rect 58571 138076 58572 138140
rect 58636 138076 58637 138140
rect 58571 138075 58637 138076
rect 58390 132450 58634 132510
rect 57835 49196 57901 49197
rect 57835 49132 57836 49196
rect 57900 49132 57901 49196
rect 57835 49131 57901 49132
rect 57283 34916 57349 34917
rect 57283 34852 57284 34916
rect 57348 34852 57349 34916
rect 57283 34851 57349 34852
rect 58574 21725 58634 132450
rect 58758 115157 58818 167859
rect 58939 146844 59005 146845
rect 58939 146780 58940 146844
rect 59004 146780 59005 146844
rect 58939 146779 59005 146780
rect 58755 115156 58821 115157
rect 58755 115092 58756 115156
rect 58820 115092 58821 115156
rect 58755 115091 58821 115092
rect 58755 114476 58821 114477
rect 58755 114412 58756 114476
rect 58820 114412 58821 114476
rect 58755 114411 58821 114412
rect 58758 68917 58818 114411
rect 58755 68916 58821 68917
rect 58755 68852 58756 68916
rect 58820 68852 58821 68916
rect 58755 68851 58821 68852
rect 58571 21724 58637 21725
rect 58571 21660 58572 21724
rect 58636 21660 58637 21724
rect 58571 21659 58637 21660
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55627 3908 55693 3909
rect 55627 3844 55628 3908
rect 55692 3844 55693 3908
rect 55627 3843 55693 3844
rect 55075 3364 55141 3365
rect 55075 3300 55076 3364
rect 55140 3300 55141 3364
rect 55075 3299 55141 3300
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 -4186 56414 20898
rect 58942 18461 59002 146779
rect 59126 54637 59186 196555
rect 82794 192454 83414 198000
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 61331 185876 61397 185877
rect 61331 185812 61332 185876
rect 61396 185812 61397 185876
rect 61331 185811 61397 185812
rect 59859 180572 59925 180573
rect 59859 180508 59860 180572
rect 59924 180508 59925 180572
rect 59859 180507 59925 180508
rect 59307 155548 59373 155549
rect 59307 155484 59308 155548
rect 59372 155484 59373 155548
rect 59307 155483 59373 155484
rect 59310 101557 59370 155483
rect 59675 147252 59741 147253
rect 59675 147188 59676 147252
rect 59740 147188 59741 147252
rect 59675 147187 59741 147188
rect 59491 141404 59557 141405
rect 59491 141340 59492 141404
rect 59556 141340 59557 141404
rect 59491 141339 59557 141340
rect 59494 112437 59554 141339
rect 59491 112436 59557 112437
rect 59491 112372 59492 112436
rect 59556 112372 59557 112436
rect 59491 112371 59557 112372
rect 59491 110668 59557 110669
rect 59491 110604 59492 110668
rect 59556 110604 59557 110668
rect 59491 110603 59557 110604
rect 59494 107541 59554 110603
rect 59491 107540 59557 107541
rect 59491 107476 59492 107540
rect 59556 107476 59557 107540
rect 59491 107475 59557 107476
rect 59307 101556 59373 101557
rect 59307 101492 59308 101556
rect 59372 101492 59373 101556
rect 59307 101491 59373 101492
rect 59307 100060 59373 100061
rect 59307 99996 59308 100060
rect 59372 99996 59373 100060
rect 59307 99995 59373 99996
rect 59123 54636 59189 54637
rect 59123 54572 59124 54636
rect 59188 54572 59189 54636
rect 59123 54571 59189 54572
rect 59310 30565 59370 99995
rect 59307 30564 59373 30565
rect 59307 30500 59308 30564
rect 59372 30500 59373 30564
rect 59307 30499 59373 30500
rect 59678 21997 59738 147187
rect 59862 89861 59922 180507
rect 60411 177716 60477 177717
rect 60411 177652 60412 177716
rect 60476 177652 60477 177716
rect 60411 177651 60477 177652
rect 60043 158268 60109 158269
rect 60043 158204 60044 158268
rect 60108 158204 60109 158268
rect 60043 158203 60109 158204
rect 60046 146845 60106 158203
rect 60043 146844 60109 146845
rect 60043 146780 60044 146844
rect 60108 146780 60109 146844
rect 60043 146779 60109 146780
rect 60414 140997 60474 177651
rect 61334 151830 61394 185811
rect 61515 184924 61581 184925
rect 61515 184860 61516 184924
rect 61580 184860 61581 184924
rect 61515 184859 61581 184860
rect 61150 151770 61394 151830
rect 60963 151604 61029 151605
rect 60963 151540 60964 151604
rect 61028 151540 61029 151604
rect 60963 151539 61029 151540
rect 60966 147930 61026 151539
rect 60598 147870 61026 147930
rect 60598 147525 60658 147870
rect 60595 147524 60661 147525
rect 60595 147460 60596 147524
rect 60660 147460 60661 147524
rect 60595 147459 60661 147460
rect 60595 147252 60661 147253
rect 60595 147188 60596 147252
rect 60660 147250 60661 147252
rect 61150 147250 61210 151770
rect 60660 147190 61210 147250
rect 60660 147188 60661 147190
rect 60595 147187 60661 147188
rect 60595 146572 60661 146573
rect 60595 146508 60596 146572
rect 60660 146570 60661 146572
rect 61518 146570 61578 184859
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 152000 83414 155898
rect 87294 196954 87914 198000
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 152000 87914 160398
rect 118794 192454 119414 198000
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 152000 119414 155898
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 152000 123914 160398
rect 154794 192454 155414 198000
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 152000 155414 155898
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 152000 159914 160398
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 152000 191414 155898
rect 195294 196954 195914 198000
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 152000 195914 160398
rect 226794 192454 227414 198000
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 152000 227414 155898
rect 231294 196954 231914 198000
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 152000 231914 160398
rect 262794 192454 263414 198000
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 152000 263414 155898
rect 267294 196954 267914 198000
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 152000 267914 160398
rect 298794 192454 299414 198000
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 152000 299414 155898
rect 303294 196954 303914 198000
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 152000 303914 160398
rect 334794 192454 335414 198000
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 152000 335414 155898
rect 339294 196954 339914 198000
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 152000 339914 160398
rect 346902 152557 346962 199275
rect 347454 180810 347514 201590
rect 347638 201381 347698 201590
rect 347635 201380 347701 201381
rect 347635 201316 347636 201380
rect 347700 201316 347701 201380
rect 347635 201315 347701 201316
rect 347635 200972 347701 200973
rect 347635 200908 347636 200972
rect 347700 200908 347701 200972
rect 347635 200907 347701 200908
rect 347638 199749 347698 200907
rect 347822 200293 347882 556550
rect 348006 286789 348066 557490
rect 348190 330717 348250 561310
rect 348374 512005 348434 561579
rect 348371 512004 348437 512005
rect 348371 511940 348372 512004
rect 348436 511940 348437 512004
rect 348371 511939 348437 511940
rect 348371 487252 348437 487253
rect 348371 487188 348372 487252
rect 348436 487188 348437 487252
rect 348371 487187 348437 487188
rect 348187 330716 348253 330717
rect 348187 330652 348188 330716
rect 348252 330652 348253 330716
rect 348187 330651 348253 330652
rect 348003 286788 348069 286789
rect 348003 286724 348004 286788
rect 348068 286724 348069 286788
rect 348003 286723 348069 286724
rect 347819 200292 347885 200293
rect 347819 200228 347820 200292
rect 347884 200228 347885 200292
rect 347819 200227 347885 200228
rect 347635 199748 347701 199749
rect 347635 199684 347636 199748
rect 347700 199684 347701 199748
rect 347635 199683 347701 199684
rect 347635 199204 347701 199205
rect 347635 199140 347636 199204
rect 347700 199140 347701 199204
rect 347635 199139 347701 199140
rect 347638 195941 347698 199139
rect 348374 196893 348434 487187
rect 349110 483037 349170 566339
rect 349291 561100 349357 561101
rect 349291 561036 349292 561100
rect 349356 561036 349357 561100
rect 349291 561035 349357 561036
rect 349294 540973 349354 561035
rect 349291 540972 349357 540973
rect 349291 540908 349292 540972
rect 349356 540908 349357 540972
rect 349291 540907 349357 540908
rect 349107 483036 349173 483037
rect 349107 482972 349108 483036
rect 349172 482972 349173 483036
rect 349107 482971 349173 482972
rect 349291 441964 349357 441965
rect 349291 441900 349292 441964
rect 349356 441900 349357 441964
rect 349291 441899 349357 441900
rect 349107 434892 349173 434893
rect 349107 434828 349108 434892
rect 349172 434828 349173 434892
rect 349107 434827 349173 434828
rect 348555 214572 348621 214573
rect 348555 214508 348556 214572
rect 348620 214508 348621 214572
rect 348555 214507 348621 214508
rect 348371 196892 348437 196893
rect 348371 196828 348372 196892
rect 348436 196828 348437 196892
rect 348371 196827 348437 196828
rect 347635 195940 347701 195941
rect 347635 195876 347636 195940
rect 347700 195876 347701 195940
rect 347635 195875 347701 195876
rect 348558 181933 348618 214507
rect 348555 181932 348621 181933
rect 348555 181868 348556 181932
rect 348620 181868 348621 181932
rect 348555 181867 348621 181868
rect 347086 180750 347514 180810
rect 347086 153101 347146 180750
rect 349110 167925 349170 434827
rect 349294 183293 349354 441899
rect 349478 383757 349538 584427
rect 349659 558924 349725 558925
rect 349659 558860 349660 558924
rect 349724 558860 349725 558924
rect 349659 558859 349725 558860
rect 349662 385797 349722 558859
rect 350582 523021 350642 589731
rect 350947 563684 351013 563685
rect 350947 563620 350948 563684
rect 351012 563620 351013 563684
rect 350947 563619 351013 563620
rect 350579 523020 350645 523021
rect 350579 522956 350580 523020
rect 350644 522956 350645 523020
rect 350579 522955 350645 522956
rect 350579 507924 350645 507925
rect 350579 507860 350580 507924
rect 350644 507860 350645 507924
rect 350579 507859 350645 507860
rect 349659 385796 349725 385797
rect 349659 385732 349660 385796
rect 349724 385732 349725 385796
rect 349659 385731 349725 385732
rect 349475 383756 349541 383757
rect 349475 383692 349476 383756
rect 349540 383692 349541 383756
rect 349475 383691 349541 383692
rect 349475 295492 349541 295493
rect 349475 295428 349476 295492
rect 349540 295428 349541 295492
rect 349475 295427 349541 295428
rect 349478 184789 349538 295427
rect 350582 188869 350642 507859
rect 350763 494596 350829 494597
rect 350763 494532 350764 494596
rect 350828 494532 350829 494596
rect 350763 494531 350829 494532
rect 350579 188868 350645 188869
rect 350579 188804 350580 188868
rect 350644 188804 350645 188868
rect 350579 188803 350645 188804
rect 349475 184788 349541 184789
rect 349475 184724 349476 184788
rect 349540 184724 349541 184788
rect 349475 184723 349541 184724
rect 350766 184109 350826 494531
rect 350950 469301 351010 563619
rect 350947 469300 351013 469301
rect 350947 469236 350948 469300
rect 351012 469236 351013 469300
rect 350947 469235 351013 469236
rect 350947 463996 351013 463997
rect 350947 463932 350948 463996
rect 351012 463932 351013 463996
rect 350947 463931 351013 463932
rect 350950 189957 351010 463931
rect 351134 379541 351194 590411
rect 352794 570454 353414 605898
rect 354443 582996 354509 582997
rect 354443 582932 354444 582996
rect 354508 582932 354509 582996
rect 354443 582931 354509 582932
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352051 568852 352117 568853
rect 352051 568788 352052 568852
rect 352116 568788 352117 568852
rect 352051 568787 352117 568788
rect 351867 566132 351933 566133
rect 351867 566068 351868 566132
rect 351932 566068 351933 566132
rect 351867 566067 351933 566068
rect 351131 379540 351197 379541
rect 351131 379476 351132 379540
rect 351196 379476 351197 379540
rect 351131 379475 351197 379476
rect 350947 189956 351013 189957
rect 350947 189892 350948 189956
rect 351012 189892 351013 189956
rect 350947 189891 351013 189892
rect 350763 184108 350829 184109
rect 350763 184044 350764 184108
rect 350828 184044 350829 184108
rect 350763 184043 350829 184044
rect 349291 183292 349357 183293
rect 349291 183228 349292 183292
rect 349356 183228 349357 183292
rect 349291 183227 349357 183228
rect 349107 167924 349173 167925
rect 349107 167860 349108 167924
rect 349172 167860 349173 167924
rect 349107 167859 349173 167860
rect 347083 153100 347149 153101
rect 347083 153036 347084 153100
rect 347148 153036 347149 153100
rect 347083 153035 347149 153036
rect 346899 152556 346965 152557
rect 346899 152492 346900 152556
rect 346964 152492 346965 152556
rect 346899 152491 346965 152492
rect 351870 152285 351930 566067
rect 352054 201381 352114 568787
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 353523 518940 353589 518941
rect 353523 518876 353524 518940
rect 353588 518876 353589 518940
rect 353523 518875 353589 518876
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352051 201380 352117 201381
rect 352051 201316 352052 201380
rect 352116 201316 352117 201380
rect 352051 201315 352117 201316
rect 352794 174454 353414 209898
rect 353526 179213 353586 518875
rect 353707 407148 353773 407149
rect 353707 407084 353708 407148
rect 353772 407084 353773 407148
rect 353707 407083 353773 407084
rect 353523 179212 353589 179213
rect 353523 179148 353524 179212
rect 353588 179148 353589 179212
rect 353523 179147 353589 179148
rect 353710 176629 353770 407083
rect 354446 278765 354506 582931
rect 354443 278764 354509 278765
rect 354443 278700 354444 278764
rect 354508 278700 354509 278764
rect 354443 278699 354509 278700
rect 353707 176628 353773 176629
rect 353707 176564 353708 176628
rect 353772 176564 353773 176628
rect 353707 176563 353773 176564
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 351867 152284 351933 152285
rect 351867 152220 351868 152284
rect 351932 152220 351933 152284
rect 351867 152219 351933 152220
rect 352794 152000 353414 173898
rect 355182 152965 355242 685067
rect 357294 682954 357914 711002
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 359411 687308 359477 687309
rect 359411 687244 359412 687308
rect 359476 687244 359477 687308
rect 359411 687243 359477 687244
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 356651 682140 356717 682141
rect 356651 682076 356652 682140
rect 356716 682076 356717 682140
rect 356651 682075 356717 682076
rect 355363 265028 355429 265029
rect 355363 264964 355364 265028
rect 355428 264964 355429 265028
rect 355363 264963 355429 264964
rect 355366 155957 355426 264963
rect 356654 199613 356714 682075
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 356835 506700 356901 506701
rect 356835 506636 356836 506700
rect 356900 506636 356901 506700
rect 356835 506635 356901 506636
rect 356651 199612 356717 199613
rect 356651 199548 356652 199612
rect 356716 199548 356717 199612
rect 356651 199547 356717 199548
rect 356838 169013 356898 506635
rect 357294 502954 357914 538398
rect 358123 527100 358189 527101
rect 358123 527036 358124 527100
rect 358188 527036 358189 527100
rect 358123 527035 358189 527036
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357019 232524 357085 232525
rect 357019 232460 357020 232524
rect 357084 232460 357085 232524
rect 357019 232459 357085 232460
rect 356835 169012 356901 169013
rect 356835 168948 356836 169012
rect 356900 168948 356901 169012
rect 356835 168947 356901 168948
rect 355363 155956 355429 155957
rect 355363 155892 355364 155956
rect 355428 155892 355429 155956
rect 355363 155891 355429 155892
rect 355179 152964 355245 152965
rect 355179 152900 355180 152964
rect 355244 152900 355245 152964
rect 355179 152899 355245 152900
rect 357022 152829 357082 232459
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 358126 180437 358186 527035
rect 359414 199477 359474 687243
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361435 684724 361501 684725
rect 361435 684660 361436 684724
rect 361500 684660 361501 684724
rect 361435 684659 361501 684660
rect 359595 578780 359661 578781
rect 359595 578716 359596 578780
rect 359660 578716 359661 578780
rect 359595 578715 359661 578716
rect 359411 199476 359477 199477
rect 359411 199412 359412 199476
rect 359476 199412 359477 199476
rect 359411 199411 359477 199412
rect 358123 180436 358189 180437
rect 358123 180372 358124 180436
rect 358188 180372 358189 180436
rect 358123 180371 358189 180372
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357019 152828 357085 152829
rect 357019 152764 357020 152828
rect 357084 152764 357085 152828
rect 357019 152763 357085 152764
rect 357294 152000 357914 178398
rect 359598 153781 359658 578715
rect 360699 566268 360765 566269
rect 360699 566204 360700 566268
rect 360764 566204 360765 566268
rect 360699 566203 360765 566204
rect 360702 153781 360762 566203
rect 359595 153780 359661 153781
rect 359595 153716 359596 153780
rect 359660 153716 359661 153780
rect 359595 153715 359661 153716
rect 360699 153780 360765 153781
rect 360699 153716 360700 153780
rect 360764 153716 360765 153780
rect 360699 153715 360765 153716
rect 361438 152285 361498 684659
rect 361794 651454 362414 686898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 363459 681052 363525 681053
rect 363459 680988 363460 681052
rect 363524 680988 363525 681052
rect 363459 680987 363525 680988
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 362907 262988 362973 262989
rect 362907 262924 362908 262988
rect 362972 262924 362973 262988
rect 362907 262923 362973 262924
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361435 152284 361501 152285
rect 361435 152220 361436 152284
rect 361500 152220 361501 152284
rect 361435 152219 361501 152220
rect 361794 152000 362414 182898
rect 362910 159493 362970 262923
rect 363462 195669 363522 680987
rect 366294 655954 366914 691398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 368979 680916 369045 680917
rect 368979 680852 368980 680916
rect 369044 680852 369045 680916
rect 368979 680851 369045 680852
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 364931 635900 364997 635901
rect 364931 635836 364932 635900
rect 364996 635836 364997 635900
rect 364931 635835 364997 635836
rect 364934 198117 364994 635835
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 365115 565860 365181 565861
rect 365115 565796 365116 565860
rect 365180 565796 365181 565860
rect 365115 565795 365181 565796
rect 364931 198116 364997 198117
rect 364931 198052 364932 198116
rect 364996 198052 364997 198116
rect 364931 198051 364997 198052
rect 363459 195668 363525 195669
rect 363459 195604 363460 195668
rect 363524 195604 363525 195668
rect 363459 195603 363525 195604
rect 365118 181797 365178 565795
rect 366294 547954 366914 583398
rect 367139 561780 367205 561781
rect 367139 561716 367140 561780
rect 367204 561716 367205 561780
rect 367139 561715 367205 561716
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 365115 181796 365181 181797
rect 365115 181732 365116 181796
rect 365180 181732 365181 181796
rect 365115 181731 365181 181732
rect 362907 159492 362973 159493
rect 362907 159428 362908 159492
rect 362972 159428 362973 159492
rect 362907 159427 362973 159428
rect 366294 152000 366914 187398
rect 367142 176493 367202 561715
rect 367691 407420 367757 407421
rect 367691 407356 367692 407420
rect 367756 407356 367757 407420
rect 367691 407355 367757 407356
rect 367694 187373 367754 407355
rect 368982 197981 369042 680851
rect 370635 680780 370701 680781
rect 370635 680716 370636 680780
rect 370700 680716 370701 680780
rect 370635 680715 370701 680716
rect 369163 566812 369229 566813
rect 369163 566748 369164 566812
rect 369228 566748 369229 566812
rect 369163 566747 369229 566748
rect 368979 197980 369045 197981
rect 368979 197916 368980 197980
rect 369044 197916 369045 197980
rect 368979 197915 369045 197916
rect 367691 187372 367757 187373
rect 367691 187308 367692 187372
rect 367756 187308 367757 187372
rect 367691 187307 367757 187308
rect 367139 176492 367205 176493
rect 367139 176428 367140 176492
rect 367204 176428 367205 176492
rect 367139 176427 367205 176428
rect 369166 163437 369226 566747
rect 369163 163436 369229 163437
rect 369163 163372 369164 163436
rect 369228 163372 369229 163436
rect 369163 163371 369229 163372
rect 370638 153101 370698 680715
rect 370794 660454 371414 695898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375051 683500 375117 683501
rect 375051 683436 375052 683500
rect 375116 683436 375117 683500
rect 375051 683435 375117 683436
rect 371739 682548 371805 682549
rect 371739 682484 371740 682548
rect 371804 682484 371805 682548
rect 371739 682483 371805 682484
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 371742 182069 371802 682483
rect 371923 593740 371989 593741
rect 371923 593676 371924 593740
rect 371988 593676 371989 593740
rect 371923 593675 371989 593676
rect 371926 188461 371986 593675
rect 373395 580820 373461 580821
rect 373395 580756 373396 580820
rect 373460 580756 373461 580820
rect 373395 580755 373461 580756
rect 373211 565996 373277 565997
rect 373211 565932 373212 565996
rect 373276 565932 373277 565996
rect 373211 565931 373277 565932
rect 371923 188460 371989 188461
rect 371923 188396 371924 188460
rect 371988 188396 371989 188460
rect 371923 188395 371989 188396
rect 371739 182068 371805 182069
rect 371739 182004 371740 182068
rect 371804 182004 371805 182068
rect 371739 182003 371805 182004
rect 373214 160717 373274 565931
rect 373398 192813 373458 580755
rect 374499 562052 374565 562053
rect 374499 561988 374500 562052
rect 374564 561988 374565 562052
rect 374499 561987 374565 561988
rect 373395 192812 373461 192813
rect 373395 192748 373396 192812
rect 373460 192748 373461 192812
rect 373395 192747 373461 192748
rect 373211 160716 373277 160717
rect 373211 160652 373212 160716
rect 373276 160652 373277 160716
rect 373211 160651 373277 160652
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370635 153100 370701 153101
rect 370635 153036 370636 153100
rect 370700 153036 370701 153100
rect 370635 153035 370701 153036
rect 370794 152000 371414 155898
rect 374502 152557 374562 561987
rect 375054 157045 375114 683435
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 382779 685268 382845 685269
rect 382779 685204 382780 685268
rect 382844 685204 382845 685268
rect 382779 685203 382845 685204
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 377259 657660 377325 657661
rect 377259 657596 377260 657660
rect 377324 657596 377325 657660
rect 377259 657595 377325 657596
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 376891 568716 376957 568717
rect 376891 568652 376892 568716
rect 376956 568652 376957 568716
rect 376891 568651 376957 568652
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375051 157044 375117 157045
rect 375051 156980 375052 157044
rect 375116 156980 375117 157044
rect 375051 156979 375117 156980
rect 374499 152556 374565 152557
rect 374499 152492 374500 152556
rect 374564 152492 374565 152556
rect 374499 152491 374565 152492
rect 375294 152000 375914 160398
rect 376894 155821 376954 568651
rect 376891 155820 376957 155821
rect 376891 155756 376892 155820
rect 376956 155756 376957 155820
rect 376891 155755 376957 155756
rect 377262 152421 377322 657595
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 378731 598500 378797 598501
rect 378731 598436 378732 598500
rect 378796 598436 378797 598500
rect 378731 598435 378797 598436
rect 378734 188325 378794 598435
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 378915 567356 378981 567357
rect 378915 567292 378916 567356
rect 378980 567292 378981 567356
rect 378915 567291 378981 567292
rect 378731 188324 378797 188325
rect 378731 188260 378732 188324
rect 378796 188260 378797 188324
rect 378731 188259 378797 188260
rect 378918 160853 378978 567291
rect 379794 561454 380414 596898
rect 381675 584900 381741 584901
rect 381675 584836 381676 584900
rect 381740 584836 381741 584900
rect 381675 584835 381741 584836
rect 381491 567220 381557 567221
rect 381491 567156 381492 567220
rect 381556 567156 381557 567220
rect 381491 567155 381557 567156
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 378915 160852 378981 160853
rect 378915 160788 378916 160852
rect 378980 160788 378981 160852
rect 378915 160787 378981 160788
rect 377259 152420 377325 152421
rect 377259 152356 377260 152420
rect 377324 152356 377325 152420
rect 377259 152355 377325 152356
rect 379794 152000 380414 164898
rect 381494 153917 381554 567155
rect 381678 188597 381738 584835
rect 381675 188596 381741 188597
rect 381675 188532 381676 188596
rect 381740 188532 381741 188596
rect 381675 188531 381741 188532
rect 382782 183157 382842 685203
rect 383515 682276 383581 682277
rect 383515 682212 383516 682276
rect 383580 682212 383581 682276
rect 383515 682211 383581 682212
rect 383518 183701 383578 682211
rect 384294 673954 384914 709082
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388299 679964 388365 679965
rect 388299 679900 388300 679964
rect 388364 679900 388365 679964
rect 388299 679899 388365 679900
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 387563 604484 387629 604485
rect 387563 604420 387564 604484
rect 387628 604420 387629 604484
rect 387563 604419 387629 604420
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 385539 581500 385605 581501
rect 385539 581436 385540 581500
rect 385604 581436 385605 581500
rect 385539 581435 385605 581436
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 383515 183700 383581 183701
rect 383515 183636 383516 183700
rect 383580 183636 383581 183700
rect 383515 183635 383581 183636
rect 382779 183156 382845 183157
rect 382779 183092 382780 183156
rect 382844 183092 382845 183156
rect 382779 183091 382845 183092
rect 384294 169954 384914 205398
rect 385542 181389 385602 581435
rect 385723 557700 385789 557701
rect 385723 557636 385724 557700
rect 385788 557636 385789 557700
rect 385723 557635 385789 557636
rect 385726 187237 385786 557635
rect 387011 510780 387077 510781
rect 387011 510716 387012 510780
rect 387076 510716 387077 510780
rect 387011 510715 387077 510716
rect 386459 239868 386525 239869
rect 386459 239804 386460 239868
rect 386524 239804 386525 239868
rect 386459 239803 386525 239804
rect 385723 187236 385789 187237
rect 385723 187172 385724 187236
rect 385788 187172 385789 187236
rect 385723 187171 385789 187172
rect 385539 181388 385605 181389
rect 385539 181324 385540 181388
rect 385604 181324 385605 181388
rect 385539 181323 385605 181324
rect 386462 179077 386522 239803
rect 387014 194581 387074 510715
rect 387566 232797 387626 604419
rect 387563 232796 387629 232797
rect 387563 232732 387564 232796
rect 387628 232732 387629 232796
rect 387563 232731 387629 232732
rect 387011 194580 387077 194581
rect 387011 194516 387012 194580
rect 387076 194516 387077 194580
rect 387011 194515 387077 194516
rect 386459 179076 386525 179077
rect 386459 179012 386460 179076
rect 386524 179012 386525 179076
rect 386459 179011 386525 179012
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 381491 153916 381557 153917
rect 381491 153852 381492 153916
rect 381556 153852 381557 153916
rect 381491 153851 381557 153852
rect 384294 152000 384914 169398
rect 388302 152693 388362 679899
rect 388794 678454 389414 710042
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393083 683772 393149 683773
rect 393083 683708 393084 683772
rect 393148 683708 393149 683772
rect 393083 683707 393149 683708
rect 389771 682004 389837 682005
rect 389771 681940 389772 682004
rect 389836 681940 389837 682004
rect 389771 681939 389837 681940
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388483 611420 388549 611421
rect 388483 611356 388484 611420
rect 388548 611356 388549 611420
rect 388483 611355 388549 611356
rect 388486 178941 388546 611355
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388483 178940 388549 178941
rect 388483 178876 388484 178940
rect 388548 178876 388549 178940
rect 388483 178875 388549 178876
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388299 152692 388365 152693
rect 388299 152628 388300 152692
rect 388364 152628 388365 152692
rect 388299 152627 388365 152628
rect 388794 152000 389414 173898
rect 389774 170373 389834 681939
rect 391059 661060 391125 661061
rect 391059 660996 391060 661060
rect 391124 660996 391125 661060
rect 391059 660995 391125 660996
rect 390139 566676 390205 566677
rect 390139 566612 390140 566676
rect 390204 566612 390205 566676
rect 390139 566611 390205 566612
rect 389955 560420 390021 560421
rect 389955 560356 389956 560420
rect 390020 560356 390021 560420
rect 389955 560355 390021 560356
rect 389771 170372 389837 170373
rect 389771 170308 389772 170372
rect 389836 170308 389837 170372
rect 389771 170307 389837 170308
rect 389958 152829 390018 560355
rect 390142 163573 390202 566611
rect 391062 177581 391122 660995
rect 391795 628420 391861 628421
rect 391795 628356 391796 628420
rect 391860 628356 391861 628420
rect 391795 628355 391861 628356
rect 391243 521660 391309 521661
rect 391243 521596 391244 521660
rect 391308 521596 391309 521660
rect 391243 521595 391309 521596
rect 391059 177580 391125 177581
rect 391059 177516 391060 177580
rect 391124 177516 391125 177580
rect 391059 177515 391125 177516
rect 391246 176085 391306 521595
rect 391798 229805 391858 628355
rect 392531 502484 392597 502485
rect 392531 502420 392532 502484
rect 392596 502420 392597 502484
rect 392531 502419 392597 502420
rect 391795 229804 391861 229805
rect 391795 229740 391796 229804
rect 391860 229740 391861 229804
rect 391795 229739 391861 229740
rect 392534 184517 392594 502419
rect 393086 235517 393146 683707
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402099 683636 402165 683637
rect 402099 683572 402100 683636
rect 402164 683572 402165 683636
rect 402099 683571 402165 683572
rect 400811 682684 400877 682685
rect 400811 682620 400812 682684
rect 400876 682620 400877 682684
rect 400811 682619 400877 682620
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 395843 619580 395909 619581
rect 395843 619516 395844 619580
rect 395908 619516 395909 619580
rect 395843 619515 395909 619516
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 395291 564908 395357 564909
rect 395291 564844 395292 564908
rect 395356 564844 395357 564908
rect 395291 564843 395357 564844
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393083 235516 393149 235517
rect 393083 235452 393084 235516
rect 393148 235452 393149 235516
rect 393083 235451 393149 235452
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 392531 184516 392597 184517
rect 392531 184452 392532 184516
rect 392596 184452 392597 184516
rect 392531 184451 392597 184452
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 391243 176084 391309 176085
rect 391243 176020 391244 176084
rect 391308 176020 391309 176084
rect 391243 176019 391309 176020
rect 390139 163572 390205 163573
rect 390139 163508 390140 163572
rect 390204 163508 390205 163572
rect 390139 163507 390205 163508
rect 389955 152828 390021 152829
rect 389955 152764 389956 152828
rect 390020 152764 390021 152828
rect 389955 152763 390021 152764
rect 393294 152000 393914 178398
rect 395294 159493 395354 564843
rect 395475 331260 395541 331261
rect 395475 331196 395476 331260
rect 395540 331196 395541 331260
rect 395475 331195 395541 331196
rect 395478 189821 395538 331195
rect 395475 189820 395541 189821
rect 395475 189756 395476 189820
rect 395540 189756 395541 189820
rect 395475 189755 395541 189756
rect 395291 159492 395357 159493
rect 395291 159428 395292 159492
rect 395356 159428 395357 159492
rect 395291 159427 395357 159428
rect 395846 158677 395906 619515
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397315 591020 397381 591021
rect 397315 590956 397316 591020
rect 397380 590956 397381 591020
rect 397315 590955 397381 590956
rect 396579 564500 396645 564501
rect 396579 564436 396580 564500
rect 396644 564436 396645 564500
rect 396579 564435 396645 564436
rect 395843 158676 395909 158677
rect 395843 158612 395844 158676
rect 395908 158612 395909 158676
rect 395843 158611 395909 158612
rect 396582 153101 396642 564435
rect 397318 165069 397378 590955
rect 397794 579454 398414 614898
rect 399707 584356 399773 584357
rect 399707 584292 399708 584356
rect 399772 584292 399773 584356
rect 399707 584291 399773 584292
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 399523 563276 399589 563277
rect 399523 563212 399524 563276
rect 399588 563212 399589 563276
rect 399523 563211 399589 563212
rect 399339 560964 399405 560965
rect 399339 560900 399340 560964
rect 399404 560900 399405 560964
rect 399339 560899 399405 560900
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397315 165068 397381 165069
rect 397315 165004 397316 165068
rect 397380 165004 397381 165068
rect 397315 165003 397381 165004
rect 396579 153100 396645 153101
rect 396579 153036 396580 153100
rect 396644 153036 396645 153100
rect 396579 153035 396645 153036
rect 397794 152000 398414 182898
rect 399342 152693 399402 560899
rect 399526 160989 399586 563211
rect 399710 238509 399770 584291
rect 399707 238508 399773 238509
rect 399707 238444 399708 238508
rect 399772 238444 399773 238508
rect 399707 238443 399773 238444
rect 400814 175813 400874 682619
rect 400995 682412 401061 682413
rect 400995 682348 400996 682412
rect 401060 682348 401061 682412
rect 400995 682347 401061 682348
rect 400998 197165 401058 682347
rect 401363 624340 401429 624341
rect 401363 624276 401364 624340
rect 401428 624276 401429 624340
rect 401363 624275 401429 624276
rect 401366 234157 401426 624275
rect 402102 235381 402162 683571
rect 402294 655954 402914 691398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406515 681868 406581 681869
rect 406515 681804 406516 681868
rect 406580 681804 406581 681868
rect 406515 681803 406581 681804
rect 403571 680372 403637 680373
rect 403571 680308 403572 680372
rect 403636 680308 403637 680372
rect 403571 680307 403637 680308
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402099 235380 402165 235381
rect 402099 235316 402100 235380
rect 402164 235316 402165 235380
rect 402099 235315 402165 235316
rect 401363 234156 401429 234157
rect 401363 234092 401364 234156
rect 401428 234092 401429 234156
rect 401363 234091 401429 234092
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 400995 197164 401061 197165
rect 400995 197100 400996 197164
rect 401060 197100 401061 197164
rect 400995 197099 401061 197100
rect 402294 187954 402914 223398
rect 403574 198253 403634 680307
rect 405595 659020 405661 659021
rect 405595 658956 405596 659020
rect 405660 658956 405661 659020
rect 405595 658955 405661 658956
rect 405411 537980 405477 537981
rect 405411 537916 405412 537980
rect 405476 537916 405477 537980
rect 405411 537915 405477 537916
rect 403755 369340 403821 369341
rect 403755 369276 403756 369340
rect 403820 369276 403821 369340
rect 403755 369275 403821 369276
rect 403571 198252 403637 198253
rect 403571 198188 403572 198252
rect 403636 198188 403637 198252
rect 403571 198187 403637 198188
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 400811 175812 400877 175813
rect 400811 175748 400812 175812
rect 400876 175748 400877 175812
rect 400811 175747 400877 175748
rect 399523 160988 399589 160989
rect 399523 160924 399524 160988
rect 399588 160924 399589 160988
rect 399523 160923 399589 160924
rect 399339 152692 399405 152693
rect 399339 152628 399340 152692
rect 399404 152628 399405 152692
rect 399339 152627 399405 152628
rect 402294 152000 402914 187398
rect 403758 178805 403818 369275
rect 404859 293180 404925 293181
rect 404859 293116 404860 293180
rect 404924 293116 404925 293180
rect 404859 293115 404925 293116
rect 403939 272780 404005 272781
rect 403939 272716 403940 272780
rect 404004 272716 404005 272780
rect 403939 272715 404005 272716
rect 403755 178804 403821 178805
rect 403755 178740 403756 178804
rect 403820 178740 403821 178804
rect 403755 178739 403821 178740
rect 403942 171733 404002 272715
rect 404862 183021 404922 293115
rect 404859 183020 404925 183021
rect 404859 182956 404860 183020
rect 404924 182956 404925 183020
rect 404859 182955 404925 182956
rect 403939 171732 404005 171733
rect 403939 171668 403940 171732
rect 404004 171668 404005 171732
rect 403939 171667 404005 171668
rect 405414 166429 405474 537915
rect 405411 166428 405477 166429
rect 405411 166364 405412 166428
rect 405476 166364 405477 166428
rect 405411 166363 405477 166364
rect 405598 166293 405658 658955
rect 406331 637940 406397 637941
rect 406331 637876 406332 637940
rect 406396 637876 406397 637940
rect 406331 637875 406397 637876
rect 406147 627740 406213 627741
rect 406147 627676 406148 627740
rect 406212 627676 406213 627740
rect 406147 627675 406213 627676
rect 406150 206277 406210 627675
rect 406147 206276 406213 206277
rect 406147 206212 406148 206276
rect 406212 206212 406213 206276
rect 406147 206211 406213 206212
rect 405595 166292 405661 166293
rect 405595 166228 405596 166292
rect 405660 166228 405661 166292
rect 405595 166227 405661 166228
rect 406334 156637 406394 637875
rect 406331 156636 406397 156637
rect 406331 156572 406332 156636
rect 406396 156572 406397 156636
rect 406331 156571 406397 156572
rect 406518 154053 406578 681803
rect 406794 660454 407414 695898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 409827 683908 409893 683909
rect 409827 683844 409828 683908
rect 409892 683844 409893 683908
rect 409827 683843 409893 683844
rect 409643 679828 409709 679829
rect 409643 679764 409644 679828
rect 409708 679764 409709 679828
rect 409643 679763 409709 679764
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 408355 646780 408421 646781
rect 408355 646716 408356 646780
rect 408420 646716 408421 646780
rect 408355 646715 408421 646716
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 407619 529140 407685 529141
rect 407619 529076 407620 529140
rect 407684 529076 407685 529140
rect 407619 529075 407685 529076
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 407622 184653 407682 529075
rect 408358 428090 408418 646715
rect 408358 428030 408602 428090
rect 407803 378180 407869 378181
rect 407803 378116 407804 378180
rect 407868 378116 407869 378180
rect 407803 378115 407869 378116
rect 407806 196621 407866 378115
rect 407803 196620 407869 196621
rect 407803 196556 407804 196620
rect 407868 196556 407869 196620
rect 407803 196555 407869 196556
rect 407619 184652 407685 184653
rect 407619 184588 407620 184652
rect 407684 184588 407685 184652
rect 407619 184587 407685 184588
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406515 154052 406581 154053
rect 406515 153988 406516 154052
rect 406580 153988 406581 154052
rect 406515 153987 406581 153988
rect 406794 152000 407414 155898
rect 408542 152421 408602 428030
rect 409459 357780 409525 357781
rect 409459 357716 409460 357780
rect 409524 357716 409525 357780
rect 409459 357715 409525 357716
rect 409275 306100 409341 306101
rect 409275 306036 409276 306100
rect 409340 306036 409341 306100
rect 409275 306035 409341 306036
rect 409278 238770 409338 306035
rect 409462 240413 409522 357715
rect 409646 277541 409706 679763
rect 409830 678333 409890 683843
rect 411294 682000 411914 700398
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 682000 429914 682398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 682000 434414 686898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 682000 438914 691398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 682000 443414 695898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 682000 447914 700398
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 682000 465914 682398
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 682000 470414 686898
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 682000 474914 691398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 682000 479414 695898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 682000 483914 700398
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 682000 501914 682398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 682000 506414 686898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 682000 510914 691398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 682000 515414 695898
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 682000 519914 700398
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 682000 537914 682398
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 682000 542414 686898
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 682000 546914 691398
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 682000 551414 695898
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 552059 685948 552125 685949
rect 552059 685884 552060 685948
rect 552124 685884 552125 685948
rect 552059 685883 552125 685884
rect 551691 684996 551757 684997
rect 551691 684932 551692 684996
rect 551756 684932 551757 684996
rect 551691 684931 551757 684932
rect 551507 684588 551573 684589
rect 551507 684524 551508 684588
rect 551572 684524 551573 684588
rect 551507 684523 551573 684524
rect 410011 680644 410077 680645
rect 410011 680580 410012 680644
rect 410076 680580 410077 680644
rect 410011 680579 410077 680580
rect 409827 678332 409893 678333
rect 409827 678268 409828 678332
rect 409892 678268 409893 678332
rect 409827 678267 409893 678268
rect 409827 677652 409893 677653
rect 409827 677588 409828 677652
rect 409892 677650 409893 677652
rect 410014 677650 410074 680579
rect 409892 677590 410074 677650
rect 409892 677588 409893 677590
rect 409827 677587 409893 677588
rect 551510 673437 551570 684523
rect 551507 673436 551573 673437
rect 551507 673372 551508 673436
rect 551572 673372 551573 673436
rect 551507 673371 551573 673372
rect 429568 655954 429888 655986
rect 429568 655718 429610 655954
rect 429846 655718 429888 655954
rect 429568 655634 429888 655718
rect 429568 655398 429610 655634
rect 429846 655398 429888 655634
rect 429568 655366 429888 655398
rect 460288 655954 460608 655986
rect 460288 655718 460330 655954
rect 460566 655718 460608 655954
rect 460288 655634 460608 655718
rect 460288 655398 460330 655634
rect 460566 655398 460608 655634
rect 460288 655366 460608 655398
rect 491008 655954 491328 655986
rect 491008 655718 491050 655954
rect 491286 655718 491328 655954
rect 491008 655634 491328 655718
rect 491008 655398 491050 655634
rect 491286 655398 491328 655634
rect 491008 655366 491328 655398
rect 521728 655954 522048 655986
rect 521728 655718 521770 655954
rect 522006 655718 522048 655954
rect 521728 655634 522048 655718
rect 521728 655398 521770 655634
rect 522006 655398 522048 655634
rect 521728 655366 522048 655398
rect 414208 651454 414528 651486
rect 414208 651218 414250 651454
rect 414486 651218 414528 651454
rect 414208 651134 414528 651218
rect 414208 650898 414250 651134
rect 414486 650898 414528 651134
rect 414208 650866 414528 650898
rect 444928 651454 445248 651486
rect 444928 651218 444970 651454
rect 445206 651218 445248 651454
rect 444928 651134 445248 651218
rect 444928 650898 444970 651134
rect 445206 650898 445248 651134
rect 444928 650866 445248 650898
rect 475648 651454 475968 651486
rect 475648 651218 475690 651454
rect 475926 651218 475968 651454
rect 475648 651134 475968 651218
rect 475648 650898 475690 651134
rect 475926 650898 475968 651134
rect 475648 650866 475968 650898
rect 506368 651454 506688 651486
rect 506368 651218 506410 651454
rect 506646 651218 506688 651454
rect 506368 651134 506688 651218
rect 506368 650898 506410 651134
rect 506646 650898 506688 651134
rect 506368 650866 506688 650898
rect 537088 651454 537408 651486
rect 537088 651218 537130 651454
rect 537366 651218 537408 651454
rect 537088 651134 537408 651218
rect 537088 650898 537130 651134
rect 537366 650898 537408 651134
rect 537088 650866 537408 650898
rect 429568 619954 429888 619986
rect 429568 619718 429610 619954
rect 429846 619718 429888 619954
rect 429568 619634 429888 619718
rect 429568 619398 429610 619634
rect 429846 619398 429888 619634
rect 429568 619366 429888 619398
rect 460288 619954 460608 619986
rect 460288 619718 460330 619954
rect 460566 619718 460608 619954
rect 460288 619634 460608 619718
rect 460288 619398 460330 619634
rect 460566 619398 460608 619634
rect 460288 619366 460608 619398
rect 491008 619954 491328 619986
rect 491008 619718 491050 619954
rect 491286 619718 491328 619954
rect 491008 619634 491328 619718
rect 491008 619398 491050 619634
rect 491286 619398 491328 619634
rect 491008 619366 491328 619398
rect 521728 619954 522048 619986
rect 521728 619718 521770 619954
rect 522006 619718 522048 619954
rect 521728 619634 522048 619718
rect 521728 619398 521770 619634
rect 522006 619398 522048 619634
rect 521728 619366 522048 619398
rect 414208 615454 414528 615486
rect 414208 615218 414250 615454
rect 414486 615218 414528 615454
rect 414208 615134 414528 615218
rect 414208 614898 414250 615134
rect 414486 614898 414528 615134
rect 414208 614866 414528 614898
rect 444928 615454 445248 615486
rect 444928 615218 444970 615454
rect 445206 615218 445248 615454
rect 444928 615134 445248 615218
rect 444928 614898 444970 615134
rect 445206 614898 445248 615134
rect 444928 614866 445248 614898
rect 475648 615454 475968 615486
rect 475648 615218 475690 615454
rect 475926 615218 475968 615454
rect 475648 615134 475968 615218
rect 475648 614898 475690 615134
rect 475926 614898 475968 615134
rect 475648 614866 475968 614898
rect 506368 615454 506688 615486
rect 506368 615218 506410 615454
rect 506646 615218 506688 615454
rect 506368 615134 506688 615218
rect 506368 614898 506410 615134
rect 506646 614898 506688 615134
rect 506368 614866 506688 614898
rect 537088 615454 537408 615486
rect 537088 615218 537130 615454
rect 537366 615218 537408 615454
rect 537088 615134 537408 615218
rect 537088 614898 537130 615134
rect 537366 614898 537408 615134
rect 537088 614866 537408 614898
rect 429568 583954 429888 583986
rect 429568 583718 429610 583954
rect 429846 583718 429888 583954
rect 429568 583634 429888 583718
rect 429568 583398 429610 583634
rect 429846 583398 429888 583634
rect 429568 583366 429888 583398
rect 460288 583954 460608 583986
rect 460288 583718 460330 583954
rect 460566 583718 460608 583954
rect 460288 583634 460608 583718
rect 460288 583398 460330 583634
rect 460566 583398 460608 583634
rect 460288 583366 460608 583398
rect 491008 583954 491328 583986
rect 491008 583718 491050 583954
rect 491286 583718 491328 583954
rect 491008 583634 491328 583718
rect 491008 583398 491050 583634
rect 491286 583398 491328 583634
rect 491008 583366 491328 583398
rect 521728 583954 522048 583986
rect 521728 583718 521770 583954
rect 522006 583718 522048 583954
rect 521728 583634 522048 583718
rect 521728 583398 521770 583634
rect 522006 583398 522048 583634
rect 521728 583366 522048 583398
rect 414208 579454 414528 579486
rect 414208 579218 414250 579454
rect 414486 579218 414528 579454
rect 414208 579134 414528 579218
rect 414208 578898 414250 579134
rect 414486 578898 414528 579134
rect 414208 578866 414528 578898
rect 444928 579454 445248 579486
rect 444928 579218 444970 579454
rect 445206 579218 445248 579454
rect 444928 579134 445248 579218
rect 444928 578898 444970 579134
rect 445206 578898 445248 579134
rect 444928 578866 445248 578898
rect 475648 579454 475968 579486
rect 475648 579218 475690 579454
rect 475926 579218 475968 579454
rect 475648 579134 475968 579218
rect 475648 578898 475690 579134
rect 475926 578898 475968 579134
rect 475648 578866 475968 578898
rect 506368 579454 506688 579486
rect 506368 579218 506410 579454
rect 506646 579218 506688 579454
rect 506368 579134 506688 579218
rect 506368 578898 506410 579134
rect 506646 578898 506688 579134
rect 506368 578866 506688 578898
rect 537088 579454 537408 579486
rect 537088 579218 537130 579454
rect 537366 579218 537408 579454
rect 537088 579134 537408 579218
rect 537088 578898 537130 579134
rect 537366 578898 537408 579134
rect 537088 578866 537408 578898
rect 550771 569940 550837 569941
rect 550771 569876 550772 569940
rect 550836 569876 550837 569940
rect 550771 569875 550837 569876
rect 429568 547954 429888 547986
rect 429568 547718 429610 547954
rect 429846 547718 429888 547954
rect 429568 547634 429888 547718
rect 429568 547398 429610 547634
rect 429846 547398 429888 547634
rect 429568 547366 429888 547398
rect 460288 547954 460608 547986
rect 460288 547718 460330 547954
rect 460566 547718 460608 547954
rect 460288 547634 460608 547718
rect 460288 547398 460330 547634
rect 460566 547398 460608 547634
rect 460288 547366 460608 547398
rect 491008 547954 491328 547986
rect 491008 547718 491050 547954
rect 491286 547718 491328 547954
rect 491008 547634 491328 547718
rect 491008 547398 491050 547634
rect 491286 547398 491328 547634
rect 491008 547366 491328 547398
rect 521728 547954 522048 547986
rect 521728 547718 521770 547954
rect 522006 547718 522048 547954
rect 521728 547634 522048 547718
rect 521728 547398 521770 547634
rect 522006 547398 522048 547634
rect 521728 547366 522048 547398
rect 414208 543454 414528 543486
rect 414208 543218 414250 543454
rect 414486 543218 414528 543454
rect 414208 543134 414528 543218
rect 414208 542898 414250 543134
rect 414486 542898 414528 543134
rect 414208 542866 414528 542898
rect 444928 543454 445248 543486
rect 444928 543218 444970 543454
rect 445206 543218 445248 543454
rect 444928 543134 445248 543218
rect 444928 542898 444970 543134
rect 445206 542898 445248 543134
rect 444928 542866 445248 542898
rect 475648 543454 475968 543486
rect 475648 543218 475690 543454
rect 475926 543218 475968 543454
rect 475648 543134 475968 543218
rect 475648 542898 475690 543134
rect 475926 542898 475968 543134
rect 475648 542866 475968 542898
rect 506368 543454 506688 543486
rect 506368 543218 506410 543454
rect 506646 543218 506688 543454
rect 506368 543134 506688 543218
rect 506368 542898 506410 543134
rect 506646 542898 506688 543134
rect 506368 542866 506688 542898
rect 537088 543454 537408 543486
rect 537088 543218 537130 543454
rect 537366 543218 537408 543454
rect 537088 543134 537408 543218
rect 537088 542898 537130 543134
rect 537366 542898 537408 543134
rect 537088 542866 537408 542898
rect 429568 511954 429888 511986
rect 429568 511718 429610 511954
rect 429846 511718 429888 511954
rect 429568 511634 429888 511718
rect 429568 511398 429610 511634
rect 429846 511398 429888 511634
rect 429568 511366 429888 511398
rect 460288 511954 460608 511986
rect 460288 511718 460330 511954
rect 460566 511718 460608 511954
rect 460288 511634 460608 511718
rect 460288 511398 460330 511634
rect 460566 511398 460608 511634
rect 460288 511366 460608 511398
rect 491008 511954 491328 511986
rect 491008 511718 491050 511954
rect 491286 511718 491328 511954
rect 491008 511634 491328 511718
rect 491008 511398 491050 511634
rect 491286 511398 491328 511634
rect 491008 511366 491328 511398
rect 521728 511954 522048 511986
rect 521728 511718 521770 511954
rect 522006 511718 522048 511954
rect 521728 511634 522048 511718
rect 521728 511398 521770 511634
rect 522006 511398 522048 511634
rect 521728 511366 522048 511398
rect 414208 507454 414528 507486
rect 414208 507218 414250 507454
rect 414486 507218 414528 507454
rect 414208 507134 414528 507218
rect 414208 506898 414250 507134
rect 414486 506898 414528 507134
rect 414208 506866 414528 506898
rect 444928 507454 445248 507486
rect 444928 507218 444970 507454
rect 445206 507218 445248 507454
rect 444928 507134 445248 507218
rect 444928 506898 444970 507134
rect 445206 506898 445248 507134
rect 444928 506866 445248 506898
rect 475648 507454 475968 507486
rect 475648 507218 475690 507454
rect 475926 507218 475968 507454
rect 475648 507134 475968 507218
rect 475648 506898 475690 507134
rect 475926 506898 475968 507134
rect 475648 506866 475968 506898
rect 506368 507454 506688 507486
rect 506368 507218 506410 507454
rect 506646 507218 506688 507454
rect 506368 507134 506688 507218
rect 506368 506898 506410 507134
rect 506646 506898 506688 507134
rect 506368 506866 506688 506898
rect 537088 507454 537408 507486
rect 537088 507218 537130 507454
rect 537366 507218 537408 507454
rect 537088 507134 537408 507218
rect 537088 506898 537130 507134
rect 537366 506898 537408 507134
rect 537088 506866 537408 506898
rect 429568 475954 429888 475986
rect 429568 475718 429610 475954
rect 429846 475718 429888 475954
rect 429568 475634 429888 475718
rect 429568 475398 429610 475634
rect 429846 475398 429888 475634
rect 429568 475366 429888 475398
rect 460288 475954 460608 475986
rect 460288 475718 460330 475954
rect 460566 475718 460608 475954
rect 460288 475634 460608 475718
rect 460288 475398 460330 475634
rect 460566 475398 460608 475634
rect 460288 475366 460608 475398
rect 491008 475954 491328 475986
rect 491008 475718 491050 475954
rect 491286 475718 491328 475954
rect 491008 475634 491328 475718
rect 491008 475398 491050 475634
rect 491286 475398 491328 475634
rect 491008 475366 491328 475398
rect 521728 475954 522048 475986
rect 521728 475718 521770 475954
rect 522006 475718 522048 475954
rect 521728 475634 522048 475718
rect 521728 475398 521770 475634
rect 522006 475398 522048 475634
rect 521728 475366 522048 475398
rect 414208 471454 414528 471486
rect 414208 471218 414250 471454
rect 414486 471218 414528 471454
rect 414208 471134 414528 471218
rect 414208 470898 414250 471134
rect 414486 470898 414528 471134
rect 414208 470866 414528 470898
rect 444928 471454 445248 471486
rect 444928 471218 444970 471454
rect 445206 471218 445248 471454
rect 444928 471134 445248 471218
rect 444928 470898 444970 471134
rect 445206 470898 445248 471134
rect 444928 470866 445248 470898
rect 475648 471454 475968 471486
rect 475648 471218 475690 471454
rect 475926 471218 475968 471454
rect 475648 471134 475968 471218
rect 475648 470898 475690 471134
rect 475926 470898 475968 471134
rect 475648 470866 475968 470898
rect 506368 471454 506688 471486
rect 506368 471218 506410 471454
rect 506646 471218 506688 471454
rect 506368 471134 506688 471218
rect 506368 470898 506410 471134
rect 506646 470898 506688 471134
rect 506368 470866 506688 470898
rect 537088 471454 537408 471486
rect 537088 471218 537130 471454
rect 537366 471218 537408 471454
rect 537088 471134 537408 471218
rect 537088 470898 537130 471134
rect 537366 470898 537408 471134
rect 537088 470866 537408 470898
rect 429568 439954 429888 439986
rect 429568 439718 429610 439954
rect 429846 439718 429888 439954
rect 429568 439634 429888 439718
rect 429568 439398 429610 439634
rect 429846 439398 429888 439634
rect 429568 439366 429888 439398
rect 460288 439954 460608 439986
rect 460288 439718 460330 439954
rect 460566 439718 460608 439954
rect 460288 439634 460608 439718
rect 460288 439398 460330 439634
rect 460566 439398 460608 439634
rect 460288 439366 460608 439398
rect 491008 439954 491328 439986
rect 491008 439718 491050 439954
rect 491286 439718 491328 439954
rect 491008 439634 491328 439718
rect 491008 439398 491050 439634
rect 491286 439398 491328 439634
rect 491008 439366 491328 439398
rect 521728 439954 522048 439986
rect 521728 439718 521770 439954
rect 522006 439718 522048 439954
rect 521728 439634 522048 439718
rect 521728 439398 521770 439634
rect 522006 439398 522048 439634
rect 521728 439366 522048 439398
rect 414208 435454 414528 435486
rect 414208 435218 414250 435454
rect 414486 435218 414528 435454
rect 414208 435134 414528 435218
rect 414208 434898 414250 435134
rect 414486 434898 414528 435134
rect 414208 434866 414528 434898
rect 444928 435454 445248 435486
rect 444928 435218 444970 435454
rect 445206 435218 445248 435454
rect 444928 435134 445248 435218
rect 444928 434898 444970 435134
rect 445206 434898 445248 435134
rect 444928 434866 445248 434898
rect 475648 435454 475968 435486
rect 475648 435218 475690 435454
rect 475926 435218 475968 435454
rect 475648 435134 475968 435218
rect 475648 434898 475690 435134
rect 475926 434898 475968 435134
rect 475648 434866 475968 434898
rect 506368 435454 506688 435486
rect 506368 435218 506410 435454
rect 506646 435218 506688 435454
rect 506368 435134 506688 435218
rect 506368 434898 506410 435134
rect 506646 434898 506688 435134
rect 506368 434866 506688 434898
rect 537088 435454 537408 435486
rect 537088 435218 537130 435454
rect 537366 435218 537408 435454
rect 537088 435134 537408 435218
rect 537088 434898 537130 435134
rect 537366 434898 537408 435134
rect 537088 434866 537408 434898
rect 429568 403954 429888 403986
rect 429568 403718 429610 403954
rect 429846 403718 429888 403954
rect 429568 403634 429888 403718
rect 429568 403398 429610 403634
rect 429846 403398 429888 403634
rect 429568 403366 429888 403398
rect 460288 403954 460608 403986
rect 460288 403718 460330 403954
rect 460566 403718 460608 403954
rect 460288 403634 460608 403718
rect 460288 403398 460330 403634
rect 460566 403398 460608 403634
rect 460288 403366 460608 403398
rect 491008 403954 491328 403986
rect 491008 403718 491050 403954
rect 491286 403718 491328 403954
rect 491008 403634 491328 403718
rect 491008 403398 491050 403634
rect 491286 403398 491328 403634
rect 491008 403366 491328 403398
rect 521728 403954 522048 403986
rect 521728 403718 521770 403954
rect 522006 403718 522048 403954
rect 521728 403634 522048 403718
rect 521728 403398 521770 403634
rect 522006 403398 522048 403634
rect 521728 403366 522048 403398
rect 414208 399454 414528 399486
rect 414208 399218 414250 399454
rect 414486 399218 414528 399454
rect 414208 399134 414528 399218
rect 414208 398898 414250 399134
rect 414486 398898 414528 399134
rect 414208 398866 414528 398898
rect 444928 399454 445248 399486
rect 444928 399218 444970 399454
rect 445206 399218 445248 399454
rect 444928 399134 445248 399218
rect 444928 398898 444970 399134
rect 445206 398898 445248 399134
rect 444928 398866 445248 398898
rect 475648 399454 475968 399486
rect 475648 399218 475690 399454
rect 475926 399218 475968 399454
rect 475648 399134 475968 399218
rect 475648 398898 475690 399134
rect 475926 398898 475968 399134
rect 475648 398866 475968 398898
rect 506368 399454 506688 399486
rect 506368 399218 506410 399454
rect 506646 399218 506688 399454
rect 506368 399134 506688 399218
rect 506368 398898 506410 399134
rect 506646 398898 506688 399134
rect 506368 398866 506688 398898
rect 537088 399454 537408 399486
rect 537088 399218 537130 399454
rect 537366 399218 537408 399454
rect 537088 399134 537408 399218
rect 537088 398898 537130 399134
rect 537366 398898 537408 399134
rect 537088 398866 537408 398898
rect 429568 367954 429888 367986
rect 429568 367718 429610 367954
rect 429846 367718 429888 367954
rect 429568 367634 429888 367718
rect 429568 367398 429610 367634
rect 429846 367398 429888 367634
rect 429568 367366 429888 367398
rect 460288 367954 460608 367986
rect 460288 367718 460330 367954
rect 460566 367718 460608 367954
rect 460288 367634 460608 367718
rect 460288 367398 460330 367634
rect 460566 367398 460608 367634
rect 460288 367366 460608 367398
rect 491008 367954 491328 367986
rect 491008 367718 491050 367954
rect 491286 367718 491328 367954
rect 491008 367634 491328 367718
rect 491008 367398 491050 367634
rect 491286 367398 491328 367634
rect 491008 367366 491328 367398
rect 521728 367954 522048 367986
rect 521728 367718 521770 367954
rect 522006 367718 522048 367954
rect 521728 367634 522048 367718
rect 521728 367398 521770 367634
rect 522006 367398 522048 367634
rect 521728 367366 522048 367398
rect 414208 363454 414528 363486
rect 414208 363218 414250 363454
rect 414486 363218 414528 363454
rect 414208 363134 414528 363218
rect 414208 362898 414250 363134
rect 414486 362898 414528 363134
rect 414208 362866 414528 362898
rect 444928 363454 445248 363486
rect 444928 363218 444970 363454
rect 445206 363218 445248 363454
rect 444928 363134 445248 363218
rect 444928 362898 444970 363134
rect 445206 362898 445248 363134
rect 444928 362866 445248 362898
rect 475648 363454 475968 363486
rect 475648 363218 475690 363454
rect 475926 363218 475968 363454
rect 475648 363134 475968 363218
rect 475648 362898 475690 363134
rect 475926 362898 475968 363134
rect 475648 362866 475968 362898
rect 506368 363454 506688 363486
rect 506368 363218 506410 363454
rect 506646 363218 506688 363454
rect 506368 363134 506688 363218
rect 506368 362898 506410 363134
rect 506646 362898 506688 363134
rect 506368 362866 506688 362898
rect 537088 363454 537408 363486
rect 537088 363218 537130 363454
rect 537366 363218 537408 363454
rect 537088 363134 537408 363218
rect 537088 362898 537130 363134
rect 537366 362898 537408 363134
rect 537088 362866 537408 362898
rect 550219 336700 550285 336701
rect 550219 336636 550220 336700
rect 550284 336636 550285 336700
rect 550219 336635 550285 336636
rect 429568 331954 429888 331986
rect 429568 331718 429610 331954
rect 429846 331718 429888 331954
rect 429568 331634 429888 331718
rect 429568 331398 429610 331634
rect 429846 331398 429888 331634
rect 429568 331366 429888 331398
rect 460288 331954 460608 331986
rect 460288 331718 460330 331954
rect 460566 331718 460608 331954
rect 460288 331634 460608 331718
rect 460288 331398 460330 331634
rect 460566 331398 460608 331634
rect 460288 331366 460608 331398
rect 491008 331954 491328 331986
rect 491008 331718 491050 331954
rect 491286 331718 491328 331954
rect 491008 331634 491328 331718
rect 491008 331398 491050 331634
rect 491286 331398 491328 331634
rect 491008 331366 491328 331398
rect 521728 331954 522048 331986
rect 521728 331718 521770 331954
rect 522006 331718 522048 331954
rect 521728 331634 522048 331718
rect 521728 331398 521770 331634
rect 522006 331398 522048 331634
rect 521728 331366 522048 331398
rect 414208 327454 414528 327486
rect 414208 327218 414250 327454
rect 414486 327218 414528 327454
rect 414208 327134 414528 327218
rect 414208 326898 414250 327134
rect 414486 326898 414528 327134
rect 414208 326866 414528 326898
rect 444928 327454 445248 327486
rect 444928 327218 444970 327454
rect 445206 327218 445248 327454
rect 444928 327134 445248 327218
rect 444928 326898 444970 327134
rect 445206 326898 445248 327134
rect 444928 326866 445248 326898
rect 475648 327454 475968 327486
rect 475648 327218 475690 327454
rect 475926 327218 475968 327454
rect 475648 327134 475968 327218
rect 475648 326898 475690 327134
rect 475926 326898 475968 327134
rect 475648 326866 475968 326898
rect 506368 327454 506688 327486
rect 506368 327218 506410 327454
rect 506646 327218 506688 327454
rect 506368 327134 506688 327218
rect 506368 326898 506410 327134
rect 506646 326898 506688 327134
rect 506368 326866 506688 326898
rect 537088 327454 537408 327486
rect 537088 327218 537130 327454
rect 537366 327218 537408 327454
rect 537088 327134 537408 327218
rect 537088 326898 537130 327134
rect 537366 326898 537408 327134
rect 537088 326866 537408 326898
rect 429568 295954 429888 295986
rect 429568 295718 429610 295954
rect 429846 295718 429888 295954
rect 429568 295634 429888 295718
rect 429568 295398 429610 295634
rect 429846 295398 429888 295634
rect 429568 295366 429888 295398
rect 460288 295954 460608 295986
rect 460288 295718 460330 295954
rect 460566 295718 460608 295954
rect 460288 295634 460608 295718
rect 460288 295398 460330 295634
rect 460566 295398 460608 295634
rect 460288 295366 460608 295398
rect 491008 295954 491328 295986
rect 491008 295718 491050 295954
rect 491286 295718 491328 295954
rect 491008 295634 491328 295718
rect 491008 295398 491050 295634
rect 491286 295398 491328 295634
rect 491008 295366 491328 295398
rect 521728 295954 522048 295986
rect 521728 295718 521770 295954
rect 522006 295718 522048 295954
rect 521728 295634 522048 295718
rect 521728 295398 521770 295634
rect 522006 295398 522048 295634
rect 521728 295366 522048 295398
rect 414208 291454 414528 291486
rect 414208 291218 414250 291454
rect 414486 291218 414528 291454
rect 414208 291134 414528 291218
rect 414208 290898 414250 291134
rect 414486 290898 414528 291134
rect 414208 290866 414528 290898
rect 444928 291454 445248 291486
rect 444928 291218 444970 291454
rect 445206 291218 445248 291454
rect 444928 291134 445248 291218
rect 444928 290898 444970 291134
rect 445206 290898 445248 291134
rect 444928 290866 445248 290898
rect 475648 291454 475968 291486
rect 475648 291218 475690 291454
rect 475926 291218 475968 291454
rect 475648 291134 475968 291218
rect 475648 290898 475690 291134
rect 475926 290898 475968 291134
rect 475648 290866 475968 290898
rect 506368 291454 506688 291486
rect 506368 291218 506410 291454
rect 506646 291218 506688 291454
rect 506368 291134 506688 291218
rect 506368 290898 506410 291134
rect 506646 290898 506688 291134
rect 506368 290866 506688 290898
rect 537088 291454 537408 291486
rect 537088 291218 537130 291454
rect 537366 291218 537408 291454
rect 537088 291134 537408 291218
rect 537088 290898 537130 291134
rect 537366 290898 537408 291134
rect 537088 290866 537408 290898
rect 409643 277540 409709 277541
rect 409643 277476 409644 277540
rect 409708 277476 409709 277540
rect 409643 277475 409709 277476
rect 429568 259954 429888 259986
rect 429568 259718 429610 259954
rect 429846 259718 429888 259954
rect 429568 259634 429888 259718
rect 429568 259398 429610 259634
rect 429846 259398 429888 259634
rect 429568 259366 429888 259398
rect 460288 259954 460608 259986
rect 460288 259718 460330 259954
rect 460566 259718 460608 259954
rect 460288 259634 460608 259718
rect 460288 259398 460330 259634
rect 460566 259398 460608 259634
rect 460288 259366 460608 259398
rect 491008 259954 491328 259986
rect 491008 259718 491050 259954
rect 491286 259718 491328 259954
rect 491008 259634 491328 259718
rect 491008 259398 491050 259634
rect 491286 259398 491328 259634
rect 491008 259366 491328 259398
rect 521728 259954 522048 259986
rect 521728 259718 521770 259954
rect 522006 259718 522048 259954
rect 521728 259634 522048 259718
rect 521728 259398 521770 259634
rect 522006 259398 522048 259634
rect 521728 259366 522048 259398
rect 414208 255454 414528 255486
rect 414208 255218 414250 255454
rect 414486 255218 414528 255454
rect 414208 255134 414528 255218
rect 414208 254898 414250 255134
rect 414486 254898 414528 255134
rect 414208 254866 414528 254898
rect 444928 255454 445248 255486
rect 444928 255218 444970 255454
rect 445206 255218 445248 255454
rect 444928 255134 445248 255218
rect 444928 254898 444970 255134
rect 445206 254898 445248 255134
rect 444928 254866 445248 254898
rect 475648 255454 475968 255486
rect 475648 255218 475690 255454
rect 475926 255218 475968 255454
rect 475648 255134 475968 255218
rect 475648 254898 475690 255134
rect 475926 254898 475968 255134
rect 475648 254866 475968 254898
rect 506368 255454 506688 255486
rect 506368 255218 506410 255454
rect 506646 255218 506688 255454
rect 506368 255134 506688 255218
rect 506368 254898 506410 255134
rect 506646 254898 506688 255134
rect 506368 254866 506688 254898
rect 537088 255454 537408 255486
rect 537088 255218 537130 255454
rect 537366 255218 537408 255454
rect 537088 255134 537408 255218
rect 537088 254898 537130 255134
rect 537366 254898 537408 255134
rect 537088 254866 537408 254898
rect 409827 242860 409893 242861
rect 409827 242796 409828 242860
rect 409892 242796 409893 242860
rect 409827 242795 409893 242796
rect 409459 240412 409525 240413
rect 409459 240348 409460 240412
rect 409524 240348 409525 240412
rect 409459 240347 409525 240348
rect 409278 238710 409706 238770
rect 409646 237013 409706 238710
rect 409643 237012 409709 237013
rect 409643 236948 409644 237012
rect 409708 236948 409709 237012
rect 409643 236947 409709 236948
rect 409646 162485 409706 236947
rect 409643 162484 409709 162485
rect 409643 162420 409644 162484
rect 409708 162420 409709 162484
rect 409643 162419 409709 162420
rect 409830 152421 409890 242795
rect 410011 242452 410077 242453
rect 410011 242388 410012 242452
rect 410076 242450 410077 242452
rect 410076 242390 410258 242450
rect 410076 242388 410077 242390
rect 410011 242387 410077 242388
rect 410011 242316 410077 242317
rect 410011 242252 410012 242316
rect 410076 242252 410077 242316
rect 410011 242251 410077 242252
rect 410014 159765 410074 242251
rect 410011 159764 410077 159765
rect 410011 159700 410012 159764
rect 410076 159700 410077 159764
rect 410011 159699 410077 159700
rect 410198 155141 410258 242390
rect 548379 239732 548445 239733
rect 548379 239668 548380 239732
rect 548444 239668 548445 239732
rect 548379 239667 548445 239668
rect 547091 239596 547157 239597
rect 547091 239532 547092 239596
rect 547156 239532 547157 239596
rect 547091 239531 547157 239532
rect 545067 238236 545133 238237
rect 545067 238172 545068 238236
rect 545132 238172 545133 238236
rect 545067 238171 545133 238172
rect 411294 232954 411914 238000
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 410195 155140 410261 155141
rect 410195 155076 410196 155140
rect 410260 155076 410261 155140
rect 410195 155075 410261 155076
rect 408539 152420 408605 152421
rect 408539 152356 408540 152420
rect 408604 152356 408605 152420
rect 408539 152355 408605 152356
rect 409827 152420 409893 152421
rect 409827 152356 409828 152420
rect 409892 152356 409893 152420
rect 409827 152355 409893 152356
rect 411294 152000 411914 160398
rect 415794 237454 416414 238000
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 152000 416414 164898
rect 420294 205954 420914 238000
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 152000 420914 169398
rect 424794 210454 425414 238000
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 152000 425414 173898
rect 429294 214954 429914 238000
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 152000 429914 178398
rect 433794 219454 434414 238000
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 152000 434414 182898
rect 438294 223954 438914 238000
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 152000 438914 187398
rect 442794 228454 443414 238000
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 152000 443414 155898
rect 447294 232954 447914 238000
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 152000 447914 160398
rect 451794 237454 452414 238000
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 152000 452414 164898
rect 456294 205954 456914 238000
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 152000 456914 169398
rect 460794 210454 461414 238000
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 152000 461414 173898
rect 465294 214954 465914 238000
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 152000 465914 178398
rect 469794 219454 470414 238000
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 152000 470414 182898
rect 474294 223954 474914 238000
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 152000 474914 187398
rect 478794 228454 479414 238000
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 152000 479414 155898
rect 483294 232954 483914 238000
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 152000 483914 160398
rect 487794 237454 488414 238000
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 152000 488414 164898
rect 492294 205954 492914 238000
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 152000 492914 169398
rect 496794 210454 497414 238000
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 152000 497414 173898
rect 501294 214954 501914 238000
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 152000 501914 178398
rect 505794 219454 506414 238000
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 152000 506414 182898
rect 510294 223954 510914 238000
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 152000 510914 187398
rect 514794 228454 515414 238000
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 152000 515414 155898
rect 519294 232954 519914 238000
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 152000 519914 160398
rect 523794 237454 524414 238000
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 152000 524414 164898
rect 528294 205954 528914 238000
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 152000 528914 169398
rect 532794 210454 533414 238000
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 152000 533414 173898
rect 537294 214954 537914 238000
rect 538811 236604 538877 236605
rect 538811 236540 538812 236604
rect 538876 236540 538877 236604
rect 538811 236539 538877 236540
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 152000 537914 178398
rect 538814 147690 538874 236539
rect 538995 234156 539061 234157
rect 538995 234092 538996 234156
rect 539060 234092 539061 234156
rect 538995 234091 539061 234092
rect 538998 147930 539058 234091
rect 539179 230348 539245 230349
rect 539179 230284 539180 230348
rect 539244 230284 539245 230348
rect 539179 230283 539245 230284
rect 539182 157350 539242 230283
rect 541794 219454 542414 238000
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 539547 185604 539613 185605
rect 539547 185540 539548 185604
rect 539612 185540 539613 185604
rect 539547 185539 539613 185540
rect 539182 157290 539426 157350
rect 539366 148885 539426 157290
rect 539363 148884 539429 148885
rect 539363 148820 539364 148884
rect 539428 148820 539429 148884
rect 539363 148819 539429 148820
rect 539363 147932 539429 147933
rect 539363 147930 539364 147932
rect 538998 147870 539364 147930
rect 539363 147868 539364 147870
rect 539428 147868 539429 147932
rect 539363 147867 539429 147868
rect 538814 147630 539426 147690
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 248528 147454 248848 147486
rect 248528 147218 248570 147454
rect 248806 147218 248848 147454
rect 248528 147134 248848 147218
rect 248528 146898 248570 147134
rect 248806 146898 248848 147134
rect 248528 146866 248848 146898
rect 279248 147454 279568 147486
rect 279248 147218 279290 147454
rect 279526 147218 279568 147454
rect 279248 147134 279568 147218
rect 279248 146898 279290 147134
rect 279526 146898 279568 147134
rect 279248 146866 279568 146898
rect 309968 147454 310288 147486
rect 309968 147218 310010 147454
rect 310246 147218 310288 147454
rect 309968 147134 310288 147218
rect 309968 146898 310010 147134
rect 310246 146898 310288 147134
rect 309968 146866 310288 146898
rect 340688 147454 341008 147486
rect 340688 147218 340730 147454
rect 340966 147218 341008 147454
rect 340688 147134 341008 147218
rect 340688 146898 340730 147134
rect 340966 146898 341008 147134
rect 340688 146866 341008 146898
rect 371408 147454 371728 147486
rect 371408 147218 371450 147454
rect 371686 147218 371728 147454
rect 371408 147134 371728 147218
rect 371408 146898 371450 147134
rect 371686 146898 371728 147134
rect 371408 146866 371728 146898
rect 402128 147454 402448 147486
rect 402128 147218 402170 147454
rect 402406 147218 402448 147454
rect 402128 147134 402448 147218
rect 402128 146898 402170 147134
rect 402406 146898 402448 147134
rect 402128 146866 402448 146898
rect 432848 147454 433168 147486
rect 432848 147218 432890 147454
rect 433126 147218 433168 147454
rect 432848 147134 433168 147218
rect 432848 146898 432890 147134
rect 433126 146898 433168 147134
rect 432848 146866 433168 146898
rect 463568 147454 463888 147486
rect 463568 147218 463610 147454
rect 463846 147218 463888 147454
rect 463568 147134 463888 147218
rect 463568 146898 463610 147134
rect 463846 146898 463888 147134
rect 463568 146866 463888 146898
rect 494288 147454 494608 147486
rect 494288 147218 494330 147454
rect 494566 147218 494608 147454
rect 494288 147134 494608 147218
rect 494288 146898 494330 147134
rect 494566 146898 494608 147134
rect 494288 146866 494608 146898
rect 525008 147454 525328 147486
rect 525008 147218 525050 147454
rect 525286 147218 525328 147454
rect 539366 147389 539426 147630
rect 539363 147388 539429 147389
rect 539363 147324 539364 147388
rect 539428 147324 539429 147388
rect 539363 147323 539429 147324
rect 525008 147134 525328 147218
rect 539363 147252 539429 147253
rect 539363 147188 539364 147252
rect 539428 147188 539429 147252
rect 539363 147187 539429 147188
rect 525008 146898 525050 147134
rect 525286 146898 525328 147134
rect 525008 146866 525328 146898
rect 60660 146510 61578 146570
rect 60660 146508 60661 146510
rect 60595 146507 60661 146508
rect 539366 142170 539426 147187
rect 539182 142110 539426 142170
rect 60411 140996 60477 140997
rect 60411 140932 60412 140996
rect 60476 140932 60477 140996
rect 60411 140931 60477 140932
rect 539182 132510 539242 142110
rect 539182 132450 539426 132510
rect 539366 122773 539426 132450
rect 539363 122772 539429 122773
rect 539363 122708 539364 122772
rect 539428 122708 539429 122772
rect 539363 122707 539429 122708
rect 79568 115954 79888 115986
rect 79568 115718 79610 115954
rect 79846 115718 79888 115954
rect 79568 115634 79888 115718
rect 79568 115398 79610 115634
rect 79846 115398 79888 115634
rect 79568 115366 79888 115398
rect 110288 115954 110608 115986
rect 110288 115718 110330 115954
rect 110566 115718 110608 115954
rect 110288 115634 110608 115718
rect 110288 115398 110330 115634
rect 110566 115398 110608 115634
rect 110288 115366 110608 115398
rect 141008 115954 141328 115986
rect 141008 115718 141050 115954
rect 141286 115718 141328 115954
rect 141008 115634 141328 115718
rect 141008 115398 141050 115634
rect 141286 115398 141328 115634
rect 141008 115366 141328 115398
rect 171728 115954 172048 115986
rect 171728 115718 171770 115954
rect 172006 115718 172048 115954
rect 171728 115634 172048 115718
rect 171728 115398 171770 115634
rect 172006 115398 172048 115634
rect 171728 115366 172048 115398
rect 202448 115954 202768 115986
rect 202448 115718 202490 115954
rect 202726 115718 202768 115954
rect 202448 115634 202768 115718
rect 202448 115398 202490 115634
rect 202726 115398 202768 115634
rect 202448 115366 202768 115398
rect 233168 115954 233488 115986
rect 233168 115718 233210 115954
rect 233446 115718 233488 115954
rect 233168 115634 233488 115718
rect 233168 115398 233210 115634
rect 233446 115398 233488 115634
rect 233168 115366 233488 115398
rect 263888 115954 264208 115986
rect 263888 115718 263930 115954
rect 264166 115718 264208 115954
rect 263888 115634 264208 115718
rect 263888 115398 263930 115634
rect 264166 115398 264208 115634
rect 263888 115366 264208 115398
rect 294608 115954 294928 115986
rect 294608 115718 294650 115954
rect 294886 115718 294928 115954
rect 294608 115634 294928 115718
rect 294608 115398 294650 115634
rect 294886 115398 294928 115634
rect 294608 115366 294928 115398
rect 325328 115954 325648 115986
rect 325328 115718 325370 115954
rect 325606 115718 325648 115954
rect 325328 115634 325648 115718
rect 325328 115398 325370 115634
rect 325606 115398 325648 115634
rect 325328 115366 325648 115398
rect 356048 115954 356368 115986
rect 356048 115718 356090 115954
rect 356326 115718 356368 115954
rect 356048 115634 356368 115718
rect 356048 115398 356090 115634
rect 356326 115398 356368 115634
rect 356048 115366 356368 115398
rect 386768 115954 387088 115986
rect 386768 115718 386810 115954
rect 387046 115718 387088 115954
rect 386768 115634 387088 115718
rect 386768 115398 386810 115634
rect 387046 115398 387088 115634
rect 386768 115366 387088 115398
rect 417488 115954 417808 115986
rect 417488 115718 417530 115954
rect 417766 115718 417808 115954
rect 417488 115634 417808 115718
rect 417488 115398 417530 115634
rect 417766 115398 417808 115634
rect 417488 115366 417808 115398
rect 448208 115954 448528 115986
rect 448208 115718 448250 115954
rect 448486 115718 448528 115954
rect 448208 115634 448528 115718
rect 448208 115398 448250 115634
rect 448486 115398 448528 115634
rect 448208 115366 448528 115398
rect 478928 115954 479248 115986
rect 478928 115718 478970 115954
rect 479206 115718 479248 115954
rect 478928 115634 479248 115718
rect 478928 115398 478970 115634
rect 479206 115398 479248 115634
rect 478928 115366 479248 115398
rect 509648 115954 509968 115986
rect 509648 115718 509690 115954
rect 509926 115718 509968 115954
rect 509648 115634 509968 115718
rect 509648 115398 509690 115634
rect 509926 115398 509968 115634
rect 509648 115366 509968 115398
rect 539363 114204 539429 114205
rect 539363 114140 539364 114204
rect 539428 114140 539429 114204
rect 539363 114139 539429 114140
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 248528 111454 248848 111486
rect 248528 111218 248570 111454
rect 248806 111218 248848 111454
rect 248528 111134 248848 111218
rect 248528 110898 248570 111134
rect 248806 110898 248848 111134
rect 248528 110866 248848 110898
rect 279248 111454 279568 111486
rect 279248 111218 279290 111454
rect 279526 111218 279568 111454
rect 279248 111134 279568 111218
rect 279248 110898 279290 111134
rect 279526 110898 279568 111134
rect 279248 110866 279568 110898
rect 309968 111454 310288 111486
rect 309968 111218 310010 111454
rect 310246 111218 310288 111454
rect 309968 111134 310288 111218
rect 309968 110898 310010 111134
rect 310246 110898 310288 111134
rect 309968 110866 310288 110898
rect 340688 111454 341008 111486
rect 340688 111218 340730 111454
rect 340966 111218 341008 111454
rect 340688 111134 341008 111218
rect 340688 110898 340730 111134
rect 340966 110898 341008 111134
rect 340688 110866 341008 110898
rect 371408 111454 371728 111486
rect 371408 111218 371450 111454
rect 371686 111218 371728 111454
rect 371408 111134 371728 111218
rect 371408 110898 371450 111134
rect 371686 110898 371728 111134
rect 371408 110866 371728 110898
rect 402128 111454 402448 111486
rect 402128 111218 402170 111454
rect 402406 111218 402448 111454
rect 402128 111134 402448 111218
rect 402128 110898 402170 111134
rect 402406 110898 402448 111134
rect 402128 110866 402448 110898
rect 432848 111454 433168 111486
rect 432848 111218 432890 111454
rect 433126 111218 433168 111454
rect 432848 111134 433168 111218
rect 432848 110898 432890 111134
rect 433126 110898 433168 111134
rect 432848 110866 433168 110898
rect 463568 111454 463888 111486
rect 463568 111218 463610 111454
rect 463846 111218 463888 111454
rect 463568 111134 463888 111218
rect 463568 110898 463610 111134
rect 463846 110898 463888 111134
rect 463568 110866 463888 110898
rect 494288 111454 494608 111486
rect 494288 111218 494330 111454
rect 494566 111218 494608 111454
rect 494288 111134 494608 111218
rect 494288 110898 494330 111134
rect 494566 110898 494608 111134
rect 494288 110866 494608 110898
rect 525008 111454 525328 111486
rect 525008 111218 525050 111454
rect 525286 111218 525328 111454
rect 525008 111134 525328 111218
rect 525008 110898 525050 111134
rect 525286 110898 525328 111134
rect 525008 110866 525328 110898
rect 60043 106724 60109 106725
rect 60043 106660 60044 106724
rect 60108 106660 60109 106724
rect 60043 106659 60109 106660
rect 59859 89860 59925 89861
rect 59859 89796 59860 89860
rect 59924 89796 59925 89860
rect 59859 89795 59925 89796
rect 59675 21996 59741 21997
rect 59675 21932 59676 21996
rect 59740 21932 59741 21996
rect 59675 21931 59741 21932
rect 60046 20093 60106 106659
rect 539366 86869 539426 114139
rect 539363 86868 539429 86869
rect 539363 86804 539364 86868
rect 539428 86804 539429 86868
rect 539363 86803 539429 86804
rect 79568 79954 79888 79986
rect 79568 79718 79610 79954
rect 79846 79718 79888 79954
rect 79568 79634 79888 79718
rect 79568 79398 79610 79634
rect 79846 79398 79888 79634
rect 79568 79366 79888 79398
rect 110288 79954 110608 79986
rect 110288 79718 110330 79954
rect 110566 79718 110608 79954
rect 110288 79634 110608 79718
rect 110288 79398 110330 79634
rect 110566 79398 110608 79634
rect 110288 79366 110608 79398
rect 141008 79954 141328 79986
rect 141008 79718 141050 79954
rect 141286 79718 141328 79954
rect 141008 79634 141328 79718
rect 141008 79398 141050 79634
rect 141286 79398 141328 79634
rect 141008 79366 141328 79398
rect 171728 79954 172048 79986
rect 171728 79718 171770 79954
rect 172006 79718 172048 79954
rect 171728 79634 172048 79718
rect 171728 79398 171770 79634
rect 172006 79398 172048 79634
rect 171728 79366 172048 79398
rect 202448 79954 202768 79986
rect 202448 79718 202490 79954
rect 202726 79718 202768 79954
rect 202448 79634 202768 79718
rect 202448 79398 202490 79634
rect 202726 79398 202768 79634
rect 202448 79366 202768 79398
rect 233168 79954 233488 79986
rect 233168 79718 233210 79954
rect 233446 79718 233488 79954
rect 233168 79634 233488 79718
rect 233168 79398 233210 79634
rect 233446 79398 233488 79634
rect 233168 79366 233488 79398
rect 263888 79954 264208 79986
rect 263888 79718 263930 79954
rect 264166 79718 264208 79954
rect 263888 79634 264208 79718
rect 263888 79398 263930 79634
rect 264166 79398 264208 79634
rect 263888 79366 264208 79398
rect 294608 79954 294928 79986
rect 294608 79718 294650 79954
rect 294886 79718 294928 79954
rect 294608 79634 294928 79718
rect 294608 79398 294650 79634
rect 294886 79398 294928 79634
rect 294608 79366 294928 79398
rect 325328 79954 325648 79986
rect 325328 79718 325370 79954
rect 325606 79718 325648 79954
rect 325328 79634 325648 79718
rect 325328 79398 325370 79634
rect 325606 79398 325648 79634
rect 325328 79366 325648 79398
rect 356048 79954 356368 79986
rect 356048 79718 356090 79954
rect 356326 79718 356368 79954
rect 356048 79634 356368 79718
rect 356048 79398 356090 79634
rect 356326 79398 356368 79634
rect 356048 79366 356368 79398
rect 386768 79954 387088 79986
rect 386768 79718 386810 79954
rect 387046 79718 387088 79954
rect 386768 79634 387088 79718
rect 386768 79398 386810 79634
rect 387046 79398 387088 79634
rect 386768 79366 387088 79398
rect 417488 79954 417808 79986
rect 417488 79718 417530 79954
rect 417766 79718 417808 79954
rect 417488 79634 417808 79718
rect 417488 79398 417530 79634
rect 417766 79398 417808 79634
rect 417488 79366 417808 79398
rect 448208 79954 448528 79986
rect 448208 79718 448250 79954
rect 448486 79718 448528 79954
rect 448208 79634 448528 79718
rect 448208 79398 448250 79634
rect 448486 79398 448528 79634
rect 448208 79366 448528 79398
rect 478928 79954 479248 79986
rect 478928 79718 478970 79954
rect 479206 79718 479248 79954
rect 478928 79634 479248 79718
rect 478928 79398 478970 79634
rect 479206 79398 479248 79634
rect 478928 79366 479248 79398
rect 509648 79954 509968 79986
rect 509648 79718 509690 79954
rect 509926 79718 509968 79954
rect 509648 79634 509968 79718
rect 509648 79398 509690 79634
rect 509926 79398 509968 79634
rect 509648 79366 509968 79398
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 248528 75454 248848 75486
rect 248528 75218 248570 75454
rect 248806 75218 248848 75454
rect 248528 75134 248848 75218
rect 248528 74898 248570 75134
rect 248806 74898 248848 75134
rect 248528 74866 248848 74898
rect 279248 75454 279568 75486
rect 279248 75218 279290 75454
rect 279526 75218 279568 75454
rect 279248 75134 279568 75218
rect 279248 74898 279290 75134
rect 279526 74898 279568 75134
rect 279248 74866 279568 74898
rect 309968 75454 310288 75486
rect 309968 75218 310010 75454
rect 310246 75218 310288 75454
rect 309968 75134 310288 75218
rect 309968 74898 310010 75134
rect 310246 74898 310288 75134
rect 309968 74866 310288 74898
rect 340688 75454 341008 75486
rect 340688 75218 340730 75454
rect 340966 75218 341008 75454
rect 340688 75134 341008 75218
rect 340688 74898 340730 75134
rect 340966 74898 341008 75134
rect 340688 74866 341008 74898
rect 371408 75454 371728 75486
rect 371408 75218 371450 75454
rect 371686 75218 371728 75454
rect 371408 75134 371728 75218
rect 371408 74898 371450 75134
rect 371686 74898 371728 75134
rect 371408 74866 371728 74898
rect 402128 75454 402448 75486
rect 402128 75218 402170 75454
rect 402406 75218 402448 75454
rect 402128 75134 402448 75218
rect 402128 74898 402170 75134
rect 402406 74898 402448 75134
rect 402128 74866 402448 74898
rect 432848 75454 433168 75486
rect 432848 75218 432890 75454
rect 433126 75218 433168 75454
rect 432848 75134 433168 75218
rect 432848 74898 432890 75134
rect 433126 74898 433168 75134
rect 432848 74866 433168 74898
rect 463568 75454 463888 75486
rect 463568 75218 463610 75454
rect 463846 75218 463888 75454
rect 463568 75134 463888 75218
rect 463568 74898 463610 75134
rect 463846 74898 463888 75134
rect 463568 74866 463888 74898
rect 494288 75454 494608 75486
rect 494288 75218 494330 75454
rect 494566 75218 494608 75454
rect 494288 75134 494608 75218
rect 494288 74898 494330 75134
rect 494566 74898 494608 75134
rect 494288 74866 494608 74898
rect 525008 75454 525328 75486
rect 525008 75218 525050 75454
rect 525286 75218 525328 75454
rect 525008 75134 525328 75218
rect 525008 74898 525050 75134
rect 525286 74898 525328 75134
rect 525008 74866 525328 74898
rect 79568 43954 79888 43986
rect 79568 43718 79610 43954
rect 79846 43718 79888 43954
rect 79568 43634 79888 43718
rect 79568 43398 79610 43634
rect 79846 43398 79888 43634
rect 79568 43366 79888 43398
rect 110288 43954 110608 43986
rect 110288 43718 110330 43954
rect 110566 43718 110608 43954
rect 110288 43634 110608 43718
rect 110288 43398 110330 43634
rect 110566 43398 110608 43634
rect 110288 43366 110608 43398
rect 141008 43954 141328 43986
rect 141008 43718 141050 43954
rect 141286 43718 141328 43954
rect 141008 43634 141328 43718
rect 141008 43398 141050 43634
rect 141286 43398 141328 43634
rect 141008 43366 141328 43398
rect 171728 43954 172048 43986
rect 171728 43718 171770 43954
rect 172006 43718 172048 43954
rect 171728 43634 172048 43718
rect 171728 43398 171770 43634
rect 172006 43398 172048 43634
rect 171728 43366 172048 43398
rect 202448 43954 202768 43986
rect 202448 43718 202490 43954
rect 202726 43718 202768 43954
rect 202448 43634 202768 43718
rect 202448 43398 202490 43634
rect 202726 43398 202768 43634
rect 202448 43366 202768 43398
rect 233168 43954 233488 43986
rect 233168 43718 233210 43954
rect 233446 43718 233488 43954
rect 233168 43634 233488 43718
rect 233168 43398 233210 43634
rect 233446 43398 233488 43634
rect 233168 43366 233488 43398
rect 263888 43954 264208 43986
rect 263888 43718 263930 43954
rect 264166 43718 264208 43954
rect 263888 43634 264208 43718
rect 263888 43398 263930 43634
rect 264166 43398 264208 43634
rect 263888 43366 264208 43398
rect 294608 43954 294928 43986
rect 294608 43718 294650 43954
rect 294886 43718 294928 43954
rect 294608 43634 294928 43718
rect 294608 43398 294650 43634
rect 294886 43398 294928 43634
rect 294608 43366 294928 43398
rect 325328 43954 325648 43986
rect 325328 43718 325370 43954
rect 325606 43718 325648 43954
rect 325328 43634 325648 43718
rect 325328 43398 325370 43634
rect 325606 43398 325648 43634
rect 325328 43366 325648 43398
rect 356048 43954 356368 43986
rect 356048 43718 356090 43954
rect 356326 43718 356368 43954
rect 356048 43634 356368 43718
rect 356048 43398 356090 43634
rect 356326 43398 356368 43634
rect 356048 43366 356368 43398
rect 386768 43954 387088 43986
rect 386768 43718 386810 43954
rect 387046 43718 387088 43954
rect 386768 43634 387088 43718
rect 386768 43398 386810 43634
rect 387046 43398 387088 43634
rect 386768 43366 387088 43398
rect 417488 43954 417808 43986
rect 417488 43718 417530 43954
rect 417766 43718 417808 43954
rect 417488 43634 417808 43718
rect 417488 43398 417530 43634
rect 417766 43398 417808 43634
rect 417488 43366 417808 43398
rect 448208 43954 448528 43986
rect 448208 43718 448250 43954
rect 448486 43718 448528 43954
rect 448208 43634 448528 43718
rect 448208 43398 448250 43634
rect 448486 43398 448528 43634
rect 448208 43366 448528 43398
rect 478928 43954 479248 43986
rect 478928 43718 478970 43954
rect 479206 43718 479248 43954
rect 478928 43634 479248 43718
rect 478928 43398 478970 43634
rect 479206 43398 479248 43634
rect 478928 43366 479248 43398
rect 509648 43954 509968 43986
rect 509648 43718 509690 43954
rect 509926 43718 509968 43954
rect 509648 43634 509968 43718
rect 509648 43398 509690 43634
rect 509926 43398 509968 43634
rect 509648 43366 509968 43398
rect 64208 39454 64528 39486
rect 64208 39218 64250 39454
rect 64486 39218 64528 39454
rect 64208 39134 64528 39218
rect 64208 38898 64250 39134
rect 64486 38898 64528 39134
rect 64208 38866 64528 38898
rect 94928 39454 95248 39486
rect 94928 39218 94970 39454
rect 95206 39218 95248 39454
rect 94928 39134 95248 39218
rect 94928 38898 94970 39134
rect 95206 38898 95248 39134
rect 94928 38866 95248 38898
rect 125648 39454 125968 39486
rect 125648 39218 125690 39454
rect 125926 39218 125968 39454
rect 125648 39134 125968 39218
rect 125648 38898 125690 39134
rect 125926 38898 125968 39134
rect 125648 38866 125968 38898
rect 156368 39454 156688 39486
rect 156368 39218 156410 39454
rect 156646 39218 156688 39454
rect 156368 39134 156688 39218
rect 156368 38898 156410 39134
rect 156646 38898 156688 39134
rect 156368 38866 156688 38898
rect 187088 39454 187408 39486
rect 187088 39218 187130 39454
rect 187366 39218 187408 39454
rect 187088 39134 187408 39218
rect 187088 38898 187130 39134
rect 187366 38898 187408 39134
rect 187088 38866 187408 38898
rect 217808 39454 218128 39486
rect 217808 39218 217850 39454
rect 218086 39218 218128 39454
rect 217808 39134 218128 39218
rect 217808 38898 217850 39134
rect 218086 38898 218128 39134
rect 217808 38866 218128 38898
rect 248528 39454 248848 39486
rect 248528 39218 248570 39454
rect 248806 39218 248848 39454
rect 248528 39134 248848 39218
rect 248528 38898 248570 39134
rect 248806 38898 248848 39134
rect 248528 38866 248848 38898
rect 279248 39454 279568 39486
rect 279248 39218 279290 39454
rect 279526 39218 279568 39454
rect 279248 39134 279568 39218
rect 279248 38898 279290 39134
rect 279526 38898 279568 39134
rect 279248 38866 279568 38898
rect 309968 39454 310288 39486
rect 309968 39218 310010 39454
rect 310246 39218 310288 39454
rect 309968 39134 310288 39218
rect 309968 38898 310010 39134
rect 310246 38898 310288 39134
rect 309968 38866 310288 38898
rect 340688 39454 341008 39486
rect 340688 39218 340730 39454
rect 340966 39218 341008 39454
rect 340688 39134 341008 39218
rect 340688 38898 340730 39134
rect 340966 38898 341008 39134
rect 340688 38866 341008 38898
rect 371408 39454 371728 39486
rect 371408 39218 371450 39454
rect 371686 39218 371728 39454
rect 371408 39134 371728 39218
rect 371408 38898 371450 39134
rect 371686 38898 371728 39134
rect 371408 38866 371728 38898
rect 402128 39454 402448 39486
rect 402128 39218 402170 39454
rect 402406 39218 402448 39454
rect 402128 39134 402448 39218
rect 402128 38898 402170 39134
rect 402406 38898 402448 39134
rect 402128 38866 402448 38898
rect 432848 39454 433168 39486
rect 432848 39218 432890 39454
rect 433126 39218 433168 39454
rect 432848 39134 433168 39218
rect 432848 38898 432890 39134
rect 433126 38898 433168 39134
rect 432848 38866 433168 38898
rect 463568 39454 463888 39486
rect 463568 39218 463610 39454
rect 463846 39218 463888 39454
rect 463568 39134 463888 39218
rect 463568 38898 463610 39134
rect 463846 38898 463888 39134
rect 463568 38866 463888 38898
rect 494288 39454 494608 39486
rect 494288 39218 494330 39454
rect 494566 39218 494608 39454
rect 494288 39134 494608 39218
rect 494288 38898 494330 39134
rect 494566 38898 494608 39134
rect 494288 38866 494608 38898
rect 525008 39454 525328 39486
rect 525008 39218 525050 39454
rect 525286 39218 525328 39454
rect 525008 39134 525328 39218
rect 525008 38898 525050 39134
rect 525286 38898 525328 39134
rect 525008 38866 525328 38898
rect 539550 38589 539610 185539
rect 541794 183454 542414 218898
rect 542675 204916 542741 204917
rect 542675 204852 542676 204916
rect 542740 204852 542741 204916
rect 542675 204851 542741 204852
rect 542678 200130 542738 204851
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 539731 180164 539797 180165
rect 539731 180100 539732 180164
rect 539796 180100 539797 180164
rect 539731 180099 539797 180100
rect 539547 38588 539613 38589
rect 539547 38524 539548 38588
rect 539612 38524 539613 38588
rect 539547 38523 539613 38524
rect 539734 35325 539794 180099
rect 541203 175948 541269 175949
rect 541203 175884 541204 175948
rect 541268 175884 541269 175948
rect 541203 175883 541269 175884
rect 540099 159628 540165 159629
rect 540099 159564 540100 159628
rect 540164 159564 540165 159628
rect 540099 159563 540165 159564
rect 539915 158132 539981 158133
rect 539915 158068 539916 158132
rect 539980 158068 539981 158132
rect 539915 158067 539981 158068
rect 539918 91765 539978 158067
rect 539915 91764 539981 91765
rect 539915 91700 539916 91764
rect 539980 91700 539981 91764
rect 539915 91699 539981 91700
rect 539731 35324 539797 35325
rect 539731 35260 539732 35324
rect 539796 35260 539797 35324
rect 539731 35259 539797 35260
rect 539363 31652 539429 31653
rect 539363 31650 539364 31652
rect 538814 31590 539364 31650
rect 60595 31108 60661 31109
rect 60595 31044 60596 31108
rect 60660 31044 60661 31108
rect 60595 31043 60661 31044
rect 60598 30970 60658 31043
rect 60598 30910 60842 30970
rect 60782 29610 60842 30910
rect 60782 29550 61210 29610
rect 60294 25954 60914 28000
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60043 20092 60109 20093
rect 60043 20028 60044 20092
rect 60108 20028 60109 20092
rect 60043 20027 60109 20028
rect 58939 18460 59005 18461
rect 58939 18396 58940 18460
rect 59004 18396 59005 18460
rect 58939 18395 59005 18396
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 -5146 60914 25398
rect 61150 3501 61210 29550
rect 61147 3500 61213 3501
rect 61147 3436 61148 3500
rect 61212 3436 61213 3500
rect 61147 3435 61213 3436
rect 73794 3454 74414 28000
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 7954 78914 28000
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 12454 83414 28000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 16954 87914 28000
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 21454 92414 28000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 25954 96914 28000
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 109794 3454 110414 28000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 7954 114914 28000
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 28000
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 16954 123914 28000
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 21454 128414 28000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 25954 132914 28000
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 145794 3454 146414 28000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 28000
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 28000
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 28000
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 28000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 28000
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 181794 3454 182414 28000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 7954 186914 28000
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 12454 191414 28000
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 28000
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 28000
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7954 222914 28000
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 12454 227414 28000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 16954 231914 28000
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 25954 240914 28000
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 7954 258914 28000
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 12454 263414 28000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 28000
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 25954 276914 28000
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 289794 3454 290414 28000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 28000
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 28000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 28000
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 28000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 25954 312914 28000
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 325794 3454 326414 28000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 7954 330914 28000
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 12454 335414 28000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 28000
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 28000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 25954 348914 28000
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 361794 3454 362414 28000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 7954 366914 28000
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 12454 371414 28000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 16954 375914 28000
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 21454 380414 28000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 25954 384914 28000
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 7954 402914 28000
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 12454 407414 28000
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 16954 411914 28000
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 21454 416414 28000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 25954 420914 28000
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 433794 3454 434414 28000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 7954 438914 28000
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 12454 443414 28000
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 16954 447914 28000
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 25954 456914 28000
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 7954 474914 28000
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 12454 479414 28000
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 16954 483914 28000
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 25954 492914 28000
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 7954 510914 28000
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 12454 515414 28000
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 16954 519914 28000
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 21454 524414 28000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 25954 528914 28000
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 538814 10981 538874 31590
rect 539363 31588 539364 31590
rect 539428 31588 539429 31652
rect 539363 31587 539429 31588
rect 539547 31108 539613 31109
rect 539547 31044 539548 31108
rect 539612 31044 539613 31108
rect 539547 31043 539613 31044
rect 539363 30564 539429 30565
rect 539363 30500 539364 30564
rect 539428 30500 539429 30564
rect 539363 30499 539429 30500
rect 539366 26250 539426 30499
rect 539550 28933 539610 31043
rect 539547 28932 539613 28933
rect 539547 28868 539548 28932
rect 539612 28868 539613 28932
rect 539547 28867 539613 28868
rect 538998 26190 539426 26250
rect 538998 21997 539058 26190
rect 538995 21996 539061 21997
rect 538995 21932 538996 21996
rect 539060 21932 539061 21996
rect 538995 21931 539061 21932
rect 540102 21861 540162 159563
rect 541019 158540 541085 158541
rect 541019 158476 541020 158540
rect 541084 158476 541085 158540
rect 541019 158475 541085 158476
rect 541022 146981 541082 158475
rect 541019 146980 541085 146981
rect 541019 146916 541020 146980
rect 541084 146916 541085 146980
rect 541019 146915 541085 146916
rect 541019 135148 541085 135149
rect 541019 135084 541020 135148
rect 541084 135084 541085 135148
rect 541019 135083 541085 135084
rect 540283 75852 540349 75853
rect 540283 75788 540284 75852
rect 540348 75788 540349 75852
rect 540283 75787 540349 75788
rect 540099 21860 540165 21861
rect 540099 21796 540100 21860
rect 540164 21796 540165 21860
rect 540099 21795 540165 21796
rect 540286 14925 540346 75787
rect 540283 14924 540349 14925
rect 540283 14860 540284 14924
rect 540348 14860 540349 14924
rect 540283 14859 540349 14860
rect 541022 11797 541082 135083
rect 541206 70957 541266 175883
rect 541387 153916 541453 153917
rect 541387 153852 541388 153916
rect 541452 153852 541453 153916
rect 541387 153851 541453 153852
rect 541390 147933 541450 153851
rect 541794 152000 542414 182898
rect 542494 200070 542738 200130
rect 541571 151740 541637 151741
rect 541571 151676 541572 151740
rect 541636 151676 541637 151740
rect 541571 151675 541637 151676
rect 541387 147932 541453 147933
rect 541387 147868 541388 147932
rect 541452 147868 541453 147932
rect 541387 147867 541453 147868
rect 541387 141132 541453 141133
rect 541387 141068 541388 141132
rect 541452 141068 541453 141132
rect 541387 141067 541453 141068
rect 541390 129981 541450 141067
rect 541574 139501 541634 151675
rect 542123 149020 542189 149021
rect 542123 148956 542124 149020
rect 542188 148956 542189 149020
rect 542123 148955 542189 148956
rect 541939 147660 542005 147661
rect 541939 147596 541940 147660
rect 542004 147596 542005 147660
rect 541939 147595 542005 147596
rect 541755 139636 541821 139637
rect 541755 139572 541756 139636
rect 541820 139572 541821 139636
rect 541755 139571 541821 139572
rect 541571 139500 541637 139501
rect 541571 139436 541572 139500
rect 541636 139436 541637 139500
rect 541571 139435 541637 139436
rect 541571 130252 541637 130253
rect 541571 130188 541572 130252
rect 541636 130188 541637 130252
rect 541571 130187 541637 130188
rect 541387 129980 541453 129981
rect 541387 129916 541388 129980
rect 541452 129916 541453 129980
rect 541387 129915 541453 129916
rect 541387 89996 541453 89997
rect 541387 89932 541388 89996
rect 541452 89932 541453 89996
rect 541387 89931 541453 89932
rect 541203 70956 541269 70957
rect 541203 70892 541204 70956
rect 541268 70892 541269 70956
rect 541203 70891 541269 70892
rect 541390 16557 541450 89931
rect 541387 16556 541453 16557
rect 541387 16492 541388 16556
rect 541452 16492 541453 16556
rect 541387 16491 541453 16492
rect 541019 11796 541085 11797
rect 541019 11732 541020 11796
rect 541084 11732 541085 11796
rect 541019 11731 541085 11732
rect 538811 10980 538877 10981
rect 538811 10916 538812 10980
rect 538876 10916 538877 10980
rect 538811 10915 538877 10916
rect 541574 6629 541634 130187
rect 541758 130117 541818 139571
rect 541942 138141 542002 147595
rect 542126 141269 542186 148955
rect 542123 141268 542189 141269
rect 542123 141204 542124 141268
rect 542188 141204 542189 141268
rect 542123 141203 542189 141204
rect 542307 140860 542373 140861
rect 542307 140796 542308 140860
rect 542372 140796 542373 140860
rect 542307 140795 542373 140796
rect 541939 138140 542005 138141
rect 541939 138076 541940 138140
rect 542004 138076 542005 138140
rect 541939 138075 542005 138076
rect 541755 130116 541821 130117
rect 541755 130052 541756 130116
rect 541820 130052 541821 130116
rect 541755 130051 541821 130052
rect 541755 129844 541821 129845
rect 541755 129780 541756 129844
rect 541820 129780 541821 129844
rect 541755 129779 541821 129780
rect 541758 89861 541818 129779
rect 542310 113117 542370 140795
rect 542307 113116 542373 113117
rect 542307 113052 542308 113116
rect 542372 113052 542373 113116
rect 542307 113051 542373 113052
rect 542494 109717 542554 200070
rect 542675 167788 542741 167789
rect 542675 167724 542676 167788
rect 542740 167724 542741 167788
rect 542675 167723 542741 167724
rect 542491 109716 542557 109717
rect 542491 109652 542492 109716
rect 542556 109652 542557 109716
rect 542491 109651 542557 109652
rect 542678 104277 542738 167723
rect 543963 165204 544029 165205
rect 543963 165140 543964 165204
rect 544028 165140 544029 165204
rect 543963 165139 544029 165140
rect 542859 156908 542925 156909
rect 542859 156844 542860 156908
rect 542924 156844 542925 156908
rect 542859 156843 542925 156844
rect 542862 144805 542922 156843
rect 543043 155820 543109 155821
rect 543043 155756 543044 155820
rect 543108 155756 543109 155820
rect 543043 155755 543109 155756
rect 542859 144804 542925 144805
rect 542859 144740 542860 144804
rect 542924 144740 542925 144804
rect 542859 144739 542925 144740
rect 543046 141133 543106 155755
rect 543779 155412 543845 155413
rect 543779 155348 543780 155412
rect 543844 155348 543845 155412
rect 543779 155347 543845 155348
rect 543595 144804 543661 144805
rect 543595 144740 543596 144804
rect 543660 144740 543661 144804
rect 543595 144739 543661 144740
rect 543043 141132 543109 141133
rect 543043 141068 543044 141132
rect 543108 141068 543109 141132
rect 543043 141067 543109 141068
rect 543598 137325 543658 144739
rect 543595 137324 543661 137325
rect 543595 137260 543596 137324
rect 543660 137260 543661 137324
rect 543595 137259 543661 137260
rect 543411 134468 543477 134469
rect 543411 134404 543412 134468
rect 543476 134404 543477 134468
rect 543411 134403 543477 134404
rect 543414 125493 543474 134403
rect 543411 125492 543477 125493
rect 543411 125428 543412 125492
rect 543476 125428 543477 125492
rect 543411 125427 543477 125428
rect 542859 124132 542925 124133
rect 542859 124068 542860 124132
rect 542924 124068 542925 124132
rect 542859 124067 542925 124068
rect 542675 104276 542741 104277
rect 542675 104212 542676 104276
rect 542740 104212 542741 104276
rect 542675 104211 542741 104212
rect 541755 89860 541821 89861
rect 541755 89796 541756 89860
rect 541820 89796 541821 89860
rect 541755 89795 541821 89796
rect 541571 6628 541637 6629
rect 541571 6564 541572 6628
rect 541636 6564 541637 6628
rect 541571 6563 541637 6564
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 541794 3454 542414 28000
rect 542862 23221 542922 124067
rect 543043 110668 543109 110669
rect 543043 110604 543044 110668
rect 543108 110604 543109 110668
rect 543043 110603 543109 110604
rect 542859 23220 542925 23221
rect 542859 23156 542860 23220
rect 542924 23156 542925 23220
rect 542859 23155 542925 23156
rect 543046 20229 543106 110603
rect 543227 106180 543293 106181
rect 543227 106116 543228 106180
rect 543292 106116 543293 106180
rect 543227 106115 543293 106116
rect 543043 20228 543109 20229
rect 543043 20164 543044 20228
rect 543108 20164 543109 20228
rect 543043 20163 543109 20164
rect 543230 16421 543290 106115
rect 543782 87957 543842 155347
rect 543966 125629 544026 165139
rect 544331 155956 544397 155957
rect 544331 155892 544332 155956
rect 544396 155892 544397 155956
rect 544331 155891 544397 155892
rect 544147 151196 544213 151197
rect 544147 151132 544148 151196
rect 544212 151132 544213 151196
rect 544147 151131 544213 151132
rect 543963 125628 544029 125629
rect 543963 125564 543964 125628
rect 544028 125564 544029 125628
rect 543963 125563 544029 125564
rect 544150 117333 544210 151131
rect 544334 129437 544394 155891
rect 545070 137322 545130 238171
rect 545251 232932 545317 232933
rect 545251 232868 545252 232932
rect 545316 232868 545317 232932
rect 545251 232867 545317 232868
rect 545254 137461 545314 232867
rect 546294 223954 546914 238000
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 545435 158404 545501 158405
rect 545435 158340 545436 158404
rect 545500 158340 545501 158404
rect 545435 158339 545501 158340
rect 545438 137730 545498 158339
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 545619 150108 545685 150109
rect 545619 150044 545620 150108
rect 545684 150044 545685 150108
rect 545619 150043 545685 150044
rect 545622 138030 545682 150043
rect 545622 137970 545866 138030
rect 545438 137670 545682 137730
rect 545251 137460 545317 137461
rect 545251 137396 545252 137460
rect 545316 137396 545317 137460
rect 545251 137395 545317 137396
rect 545070 137262 545498 137322
rect 545067 137188 545133 137189
rect 545067 137124 545068 137188
rect 545132 137124 545133 137188
rect 545067 137123 545133 137124
rect 545070 135149 545130 137123
rect 545067 135148 545133 135149
rect 545067 135084 545068 135148
rect 545132 135084 545133 135148
rect 545067 135083 545133 135084
rect 545438 132970 545498 137262
rect 545070 132910 545498 132970
rect 544331 129436 544397 129437
rect 544331 129372 544332 129436
rect 544396 129372 544397 129436
rect 544331 129371 544397 129372
rect 544515 127668 544581 127669
rect 544515 127604 544516 127668
rect 544580 127604 544581 127668
rect 544515 127603 544581 127604
rect 544147 117332 544213 117333
rect 544147 117268 544148 117332
rect 544212 117268 544213 117332
rect 544147 117267 544213 117268
rect 544331 115156 544397 115157
rect 544331 115092 544332 115156
rect 544396 115092 544397 115156
rect 544331 115091 544397 115092
rect 543963 110532 544029 110533
rect 543963 110468 543964 110532
rect 544028 110468 544029 110532
rect 543963 110467 544029 110468
rect 543779 87956 543845 87957
rect 543779 87892 543780 87956
rect 543844 87892 543845 87956
rect 543779 87891 543845 87892
rect 543966 55997 544026 110467
rect 543963 55996 544029 55997
rect 543963 55932 543964 55996
rect 544028 55932 544029 55996
rect 543963 55931 544029 55932
rect 544334 21725 544394 115091
rect 544518 110669 544578 127603
rect 544883 126988 544949 126989
rect 544883 126924 544884 126988
rect 544948 126924 544949 126988
rect 544883 126923 544949 126924
rect 544515 110668 544581 110669
rect 544515 110604 544516 110668
rect 544580 110604 544581 110668
rect 544515 110603 544581 110604
rect 544886 109037 544946 126923
rect 544883 109036 544949 109037
rect 544883 108972 544884 109036
rect 544948 108972 544949 109036
rect 544883 108971 544949 108972
rect 544515 86868 544581 86869
rect 544515 86804 544516 86868
rect 544580 86804 544581 86868
rect 544515 86803 544581 86804
rect 544518 23085 544578 86803
rect 544515 23084 544581 23085
rect 544515 23020 544516 23084
rect 544580 23020 544581 23084
rect 544515 23019 544581 23020
rect 545070 22813 545130 132910
rect 545622 132290 545682 137670
rect 545438 132230 545682 132290
rect 545251 131068 545317 131069
rect 545251 131004 545252 131068
rect 545316 131004 545317 131068
rect 545251 131003 545317 131004
rect 545067 22812 545133 22813
rect 545067 22748 545068 22812
rect 545132 22748 545133 22812
rect 545067 22747 545133 22748
rect 544331 21724 544397 21725
rect 544331 21660 544332 21724
rect 544396 21660 544397 21724
rect 544331 21659 544397 21660
rect 543227 16420 543293 16421
rect 543227 16356 543228 16420
rect 543292 16356 543293 16420
rect 543227 16355 543293 16356
rect 545254 16149 545314 131003
rect 545438 72997 545498 132230
rect 545806 128370 545866 137970
rect 545622 128310 545866 128370
rect 545622 126989 545682 128310
rect 545619 126988 545685 126989
rect 545619 126924 545620 126988
rect 545684 126924 545685 126988
rect 545619 126923 545685 126924
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 545619 89044 545685 89045
rect 545619 88980 545620 89044
rect 545684 88980 545685 89044
rect 545619 88979 545685 88980
rect 545435 72996 545501 72997
rect 545435 72932 545436 72996
rect 545500 72932 545501 72996
rect 545435 72931 545501 72932
rect 545622 17509 545682 88979
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 545619 17508 545685 17509
rect 545619 17444 545620 17508
rect 545684 17444 545685 17508
rect 545619 17443 545685 17444
rect 545251 16148 545317 16149
rect 545251 16084 545252 16148
rect 545316 16084 545317 16148
rect 545251 16083 545317 16084
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 7954 546914 43398
rect 547094 21589 547154 239531
rect 547643 166428 547709 166429
rect 547643 166364 547644 166428
rect 547708 166364 547709 166428
rect 547643 166363 547709 166364
rect 547275 157996 547341 157997
rect 547275 157932 547276 157996
rect 547340 157932 547341 157996
rect 547275 157931 547341 157932
rect 547278 124677 547338 157931
rect 547646 138030 547706 166363
rect 548011 157044 548077 157045
rect 548011 156980 548012 157044
rect 548076 156980 548077 157044
rect 548011 156979 548077 156980
rect 547646 137970 547890 138030
rect 547643 133924 547709 133925
rect 547643 133860 547644 133924
rect 547708 133860 547709 133924
rect 547643 133859 547709 133860
rect 547459 126988 547525 126989
rect 547459 126924 547460 126988
rect 547524 126924 547525 126988
rect 547459 126923 547525 126924
rect 547275 124676 547341 124677
rect 547275 124612 547276 124676
rect 547340 124612 547341 124676
rect 547275 124611 547341 124612
rect 547462 82925 547522 126923
rect 547646 126309 547706 133859
rect 547830 128485 547890 137970
rect 548014 130253 548074 156979
rect 548195 151332 548261 151333
rect 548195 151268 548196 151332
rect 548260 151268 548261 151332
rect 548195 151267 548261 151268
rect 548011 130252 548077 130253
rect 548011 130188 548012 130252
rect 548076 130188 548077 130252
rect 548011 130187 548077 130188
rect 547827 128484 547893 128485
rect 547827 128420 547828 128484
rect 547892 128420 547893 128484
rect 547827 128419 547893 128420
rect 547643 126308 547709 126309
rect 547643 126244 547644 126308
rect 547708 126244 547709 126308
rect 547643 126243 547709 126244
rect 547643 126172 547709 126173
rect 547643 126108 547644 126172
rect 547708 126108 547709 126172
rect 547643 126107 547709 126108
rect 547459 82924 547525 82925
rect 547459 82860 547460 82924
rect 547524 82860 547525 82924
rect 547459 82859 547525 82860
rect 547275 72452 547341 72453
rect 547275 72388 547276 72452
rect 547340 72388 547341 72452
rect 547275 72387 547341 72388
rect 547091 21588 547157 21589
rect 547091 21524 547092 21588
rect 547156 21524 547157 21588
rect 547091 21523 547157 21524
rect 547278 15061 547338 72387
rect 547646 23357 547706 126107
rect 548011 118828 548077 118829
rect 548011 118764 548012 118828
rect 548076 118764 548077 118828
rect 548011 118763 548077 118764
rect 548014 27029 548074 118763
rect 548198 92581 548258 151267
rect 548195 92580 548261 92581
rect 548195 92516 548196 92580
rect 548260 92516 548261 92580
rect 548195 92515 548261 92516
rect 548011 27028 548077 27029
rect 548011 26964 548012 27028
rect 548076 26964 548077 27028
rect 548011 26963 548077 26964
rect 547643 23356 547709 23357
rect 547643 23292 547644 23356
rect 547708 23292 547709 23356
rect 547643 23291 547709 23292
rect 548382 15877 548442 239667
rect 549483 238372 549549 238373
rect 549483 238308 549484 238372
rect 549548 238308 549549 238372
rect 549483 238307 549549 238308
rect 549486 18733 549546 238307
rect 549667 149156 549733 149157
rect 549667 149092 549668 149156
rect 549732 149092 549733 149156
rect 549667 149091 549733 149092
rect 549670 27437 549730 149091
rect 549667 27436 549733 27437
rect 549667 27372 549668 27436
rect 549732 27372 549733 27436
rect 549667 27371 549733 27372
rect 549483 18732 549549 18733
rect 549483 18668 549484 18732
rect 549548 18668 549549 18732
rect 549483 18667 549549 18668
rect 548379 15876 548445 15877
rect 548379 15812 548380 15876
rect 548444 15812 548445 15876
rect 548379 15811 548445 15812
rect 547275 15060 547341 15061
rect 547275 14996 547276 15060
rect 547340 14996 547341 15060
rect 547275 14995 547341 14996
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 550222 4861 550282 336635
rect 550403 262580 550469 262581
rect 550403 262516 550404 262580
rect 550468 262516 550469 262580
rect 550403 262515 550469 262516
rect 550406 29205 550466 262515
rect 550774 244290 550834 569875
rect 551507 441420 551573 441421
rect 551507 441356 551508 441420
rect 551572 441356 551573 441420
rect 551507 441355 551573 441356
rect 550590 244230 550834 244290
rect 550403 29204 550469 29205
rect 550403 29140 550404 29204
rect 550468 29140 550469 29204
rect 550403 29139 550469 29140
rect 550590 6357 550650 244230
rect 551510 238645 551570 441355
rect 551507 238644 551573 238645
rect 551507 238580 551508 238644
rect 551572 238580 551573 238644
rect 551507 238579 551573 238580
rect 550794 228454 551414 238000
rect 551694 237149 551754 684931
rect 552062 673981 552122 685883
rect 552427 679692 552493 679693
rect 552427 679628 552428 679692
rect 552492 679628 552493 679692
rect 552427 679627 552493 679628
rect 552059 673980 552125 673981
rect 552059 673916 552060 673980
rect 552124 673916 552125 673980
rect 552059 673915 552125 673916
rect 552243 673436 552309 673437
rect 552243 673372 552244 673436
rect 552308 673372 552309 673436
rect 552243 673371 552309 673372
rect 552059 641340 552125 641341
rect 552059 641276 552060 641340
rect 552124 641276 552125 641340
rect 552059 641275 552125 641276
rect 551691 237148 551757 237149
rect 551691 237084 551692 237148
rect 551756 237084 551757 237148
rect 551691 237083 551757 237084
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 552062 180029 552122 641275
rect 552246 237285 552306 673371
rect 552430 520981 552490 679627
rect 555294 664954 555914 700398
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 560523 682276 560589 682277
rect 560523 682212 560524 682276
rect 560588 682212 560589 682276
rect 560523 682211 560589 682212
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 557579 668540 557645 668541
rect 557579 668476 557580 668540
rect 557644 668476 557645 668540
rect 557579 668475 557645 668476
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 553347 628420 553413 628421
rect 553347 628356 553348 628420
rect 553412 628356 553413 628420
rect 553347 628355 553413 628356
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 553350 592050 553410 628355
rect 553166 591990 553410 592050
rect 555294 592954 555914 628398
rect 556291 608020 556357 608021
rect 556291 607956 556292 608020
rect 556356 607956 556357 608020
rect 556291 607955 556357 607956
rect 556107 599180 556173 599181
rect 556107 599116 556108 599180
rect 556172 599116 556173 599180
rect 556107 599115 556173 599116
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 553166 572730 553226 591990
rect 553166 572670 553410 572730
rect 553350 524430 553410 572670
rect 553166 524370 553410 524430
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 552427 520980 552493 520981
rect 552427 520916 552428 520980
rect 552492 520916 552493 520980
rect 552427 520915 552493 520916
rect 553166 514770 553226 524370
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 553166 514710 553410 514770
rect 553350 466470 553410 514710
rect 554819 506020 554885 506021
rect 554819 505956 554820 506020
rect 554884 505956 554885 506020
rect 554819 505955 554885 505956
rect 553531 491740 553597 491741
rect 553531 491676 553532 491740
rect 553596 491676 553597 491740
rect 553531 491675 553597 491676
rect 553166 466410 553410 466470
rect 553166 456810 553226 466410
rect 553166 456750 553410 456810
rect 553350 263610 553410 456750
rect 553166 263550 553410 263610
rect 553166 253950 553226 263550
rect 553166 253890 553410 253950
rect 553350 244290 553410 253890
rect 553166 244230 553410 244290
rect 552243 237284 552309 237285
rect 552243 237220 552244 237284
rect 552308 237220 552309 237284
rect 552243 237219 552309 237220
rect 553166 234630 553226 244230
rect 553166 234570 553410 234630
rect 552059 180028 552125 180029
rect 552059 179964 552060 180028
rect 552124 179964 552125 180028
rect 552059 179963 552125 179964
rect 552059 163572 552125 163573
rect 552059 163508 552060 163572
rect 552124 163508 552125 163572
rect 552059 163507 552125 163508
rect 551507 163436 551573 163437
rect 551507 163372 551508 163436
rect 551572 163372 551573 163436
rect 551507 163371 551573 163372
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 551510 51101 551570 163371
rect 551507 51100 551573 51101
rect 551507 51036 551508 51100
rect 551572 51036 551573 51100
rect 551507 51035 551573 51036
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 552062 29613 552122 163507
rect 552611 160988 552677 160989
rect 552611 160924 552612 160988
rect 552676 160924 552677 160988
rect 552611 160923 552677 160924
rect 552243 160716 552309 160717
rect 552243 160652 552244 160716
rect 552308 160652 552309 160716
rect 552243 160651 552309 160652
rect 552246 30837 552306 160651
rect 552427 153780 552493 153781
rect 552427 153716 552428 153780
rect 552492 153716 552493 153780
rect 552427 153715 552493 153716
rect 552243 30836 552309 30837
rect 552243 30772 552244 30836
rect 552308 30772 552309 30836
rect 552243 30771 552309 30772
rect 552059 29612 552125 29613
rect 552059 29548 552060 29612
rect 552124 29548 552125 29612
rect 552059 29547 552125 29548
rect 552430 27981 552490 153715
rect 552614 84693 552674 160923
rect 553350 138030 553410 234570
rect 553166 137970 553410 138030
rect 553166 128370 553226 137970
rect 553166 128310 553410 128370
rect 552611 84692 552677 84693
rect 552611 84628 552612 84692
rect 552676 84628 552677 84692
rect 552611 84627 552677 84628
rect 552427 27980 552493 27981
rect 552427 27916 552428 27980
rect 552492 27916 552493 27980
rect 552427 27915 552493 27916
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 553350 11933 553410 128310
rect 553534 22677 553594 491675
rect 553715 315620 553781 315621
rect 553715 315556 553716 315620
rect 553780 315556 553781 315620
rect 553715 315555 553781 315556
rect 553531 22676 553597 22677
rect 553531 22612 553532 22676
rect 553596 22612 553597 22676
rect 553531 22611 553597 22612
rect 553718 21317 553778 315555
rect 553899 158268 553965 158269
rect 553899 158204 553900 158268
rect 553964 158204 553965 158268
rect 553899 158203 553965 158204
rect 553902 22541 553962 158203
rect 553899 22540 553965 22541
rect 553899 22476 553900 22540
rect 553964 22476 553965 22540
rect 553899 22475 553965 22476
rect 553715 21316 553781 21317
rect 553715 21252 553716 21316
rect 553780 21252 553781 21316
rect 553715 21251 553781 21252
rect 554822 19005 554882 505955
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555003 404700 555069 404701
rect 555003 404636 555004 404700
rect 555068 404636 555069 404700
rect 555003 404635 555069 404636
rect 554819 19004 554885 19005
rect 554819 18940 554820 19004
rect 554884 18940 554885 19004
rect 554819 18939 554885 18940
rect 550587 6356 550653 6357
rect 550587 6292 550588 6356
rect 550652 6292 550653 6356
rect 550587 6291 550653 6292
rect 550219 4860 550285 4861
rect 550219 4796 550220 4860
rect 550284 4796 550285 4860
rect 550219 4795 550285 4796
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 -2266 551414 11898
rect 553347 11932 553413 11933
rect 553347 11868 553348 11932
rect 553412 11868 553413 11932
rect 553347 11867 553413 11868
rect 555006 7581 555066 404635
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555003 7580 555069 7581
rect 555003 7516 555004 7580
rect 555068 7516 555069 7580
rect 555003 7515 555069 7516
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 -3226 555914 16398
rect 556110 11661 556170 599115
rect 556294 19821 556354 607955
rect 556475 534580 556541 534581
rect 556475 534516 556476 534580
rect 556540 534516 556541 534580
rect 556475 534515 556541 534516
rect 556291 19820 556357 19821
rect 556291 19756 556292 19820
rect 556356 19756 556357 19820
rect 556291 19755 556357 19756
rect 556478 17237 556538 534515
rect 556659 494460 556725 494461
rect 556659 494396 556660 494460
rect 556724 494396 556725 494460
rect 556659 494395 556725 494396
rect 556475 17236 556541 17237
rect 556475 17172 556476 17236
rect 556540 17172 556541 17236
rect 556475 17171 556541 17172
rect 556107 11660 556173 11661
rect 556107 11596 556108 11660
rect 556172 11596 556173 11660
rect 556107 11595 556173 11596
rect 556662 10301 556722 494395
rect 557582 18461 557642 668475
rect 558867 649500 558933 649501
rect 558867 649436 558868 649500
rect 558932 649436 558933 649500
rect 558867 649435 558933 649436
rect 557763 633860 557829 633861
rect 557763 633796 557764 633860
rect 557828 633796 557829 633860
rect 557763 633795 557829 633796
rect 557579 18460 557645 18461
rect 557579 18396 557580 18460
rect 557644 18396 557645 18460
rect 557579 18395 557645 18396
rect 557766 12069 557826 633795
rect 557947 531860 558013 531861
rect 557947 531796 557948 531860
rect 558012 531796 558013 531860
rect 557947 531795 558013 531796
rect 557950 14517 558010 531795
rect 558131 497180 558197 497181
rect 558131 497116 558132 497180
rect 558196 497116 558197 497180
rect 558131 497115 558197 497116
rect 558134 16013 558194 497115
rect 558131 16012 558197 16013
rect 558131 15948 558132 16012
rect 558196 15948 558197 16012
rect 558131 15947 558197 15948
rect 557947 14516 558013 14517
rect 557947 14452 557948 14516
rect 558012 14452 558013 14516
rect 557947 14451 558013 14452
rect 557763 12068 557829 12069
rect 557763 12004 557764 12068
rect 557828 12004 557829 12068
rect 557763 12003 557829 12004
rect 556659 10300 556725 10301
rect 556659 10236 556660 10300
rect 556724 10236 556725 10300
rect 556659 10235 556725 10236
rect 558870 4997 558930 649435
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559051 612100 559117 612101
rect 559051 612036 559052 612100
rect 559116 612036 559117 612100
rect 559051 612035 559117 612036
rect 559054 6221 559114 612035
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559235 479500 559301 479501
rect 559235 479436 559236 479500
rect 559300 479436 559301 479500
rect 559235 479435 559301 479436
rect 559238 19957 559298 479435
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 560526 22949 560586 682211
rect 564294 673954 564914 709082
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 566043 700364 566109 700365
rect 566043 700300 566044 700364
rect 566108 700300 566109 700364
rect 566043 700299 566109 700300
rect 565123 679556 565189 679557
rect 565123 679492 565124 679556
rect 565188 679492 565189 679556
rect 565123 679491 565189 679492
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 563099 667860 563165 667861
rect 563099 667796 563100 667860
rect 563164 667796 563165 667860
rect 563099 667795 563165 667796
rect 561627 650860 561693 650861
rect 561627 650796 561628 650860
rect 561692 650796 561693 650860
rect 561627 650795 561693 650796
rect 560707 599860 560773 599861
rect 560707 599796 560708 599860
rect 560772 599796 560773 599860
rect 560707 599795 560773 599796
rect 560710 198661 560770 599795
rect 560891 546820 560957 546821
rect 560891 546756 560892 546820
rect 560956 546756 560957 546820
rect 560891 546755 560957 546756
rect 560707 198660 560773 198661
rect 560707 198596 560708 198660
rect 560772 198596 560773 198660
rect 560707 198595 560773 198596
rect 560894 197301 560954 546755
rect 561075 235244 561141 235245
rect 561075 235180 561076 235244
rect 561140 235180 561141 235244
rect 561075 235179 561141 235180
rect 560891 197300 560957 197301
rect 560891 197236 560892 197300
rect 560956 197236 560957 197300
rect 560891 197235 560957 197236
rect 560707 166292 560773 166293
rect 560707 166228 560708 166292
rect 560772 166228 560773 166292
rect 560707 166227 560773 166228
rect 560710 28525 560770 166227
rect 560707 28524 560773 28525
rect 560707 28460 560708 28524
rect 560772 28460 560773 28524
rect 560707 28459 560773 28460
rect 560523 22948 560589 22949
rect 560523 22884 560524 22948
rect 560588 22884 560589 22948
rect 560523 22883 560589 22884
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559235 19956 559301 19957
rect 559235 19892 559236 19956
rect 559300 19892 559301 19956
rect 559235 19891 559301 19892
rect 559051 6220 559117 6221
rect 559051 6156 559052 6220
rect 559116 6156 559117 6220
rect 559051 6155 559117 6156
rect 558867 4996 558933 4997
rect 558867 4932 558868 4996
rect 558932 4932 558933 4996
rect 558867 4931 558933 4932
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 -4186 560414 20898
rect 561078 20093 561138 235179
rect 561443 197436 561509 197437
rect 561443 197372 561444 197436
rect 561508 197372 561509 197436
rect 561443 197371 561509 197372
rect 561446 20909 561506 197371
rect 561630 29885 561690 650795
rect 561811 576740 561877 576741
rect 561811 576676 561812 576740
rect 561876 576676 561877 576740
rect 561811 576675 561877 576676
rect 561627 29884 561693 29885
rect 561627 29820 561628 29884
rect 561692 29820 561693 29884
rect 561627 29819 561693 29820
rect 561814 29341 561874 576675
rect 561995 552940 562061 552941
rect 561995 552876 561996 552940
rect 562060 552876 562061 552940
rect 561995 552875 562061 552876
rect 561811 29340 561877 29341
rect 561811 29276 561812 29340
rect 561876 29276 561877 29340
rect 561811 29275 561877 29276
rect 561998 28661 562058 552875
rect 562179 232660 562245 232661
rect 562179 232596 562180 232660
rect 562244 232596 562245 232660
rect 562179 232595 562245 232596
rect 562182 124133 562242 232595
rect 562179 124132 562245 124133
rect 562179 124068 562180 124132
rect 562244 124068 562245 124132
rect 562179 124067 562245 124068
rect 563102 28797 563162 667795
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 563283 602580 563349 602581
rect 563283 602516 563284 602580
rect 563348 602516 563349 602580
rect 563283 602515 563349 602516
rect 563099 28796 563165 28797
rect 563099 28732 563100 28796
rect 563164 28732 563165 28796
rect 563099 28731 563165 28732
rect 561995 28660 562061 28661
rect 561995 28596 561996 28660
rect 562060 28596 562061 28660
rect 561995 28595 562061 28596
rect 563286 24581 563346 602515
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 563467 159764 563533 159765
rect 563467 159700 563468 159764
rect 563532 159700 563533 159764
rect 563467 159699 563533 159700
rect 563283 24580 563349 24581
rect 563283 24516 563284 24580
rect 563348 24516 563349 24580
rect 563283 24515 563349 24516
rect 561443 20908 561509 20909
rect 561443 20844 561444 20908
rect 561508 20844 561509 20908
rect 561443 20843 561509 20844
rect 561075 20092 561141 20093
rect 561075 20028 561076 20092
rect 561140 20028 561141 20092
rect 561075 20027 561141 20028
rect 563470 6493 563530 159699
rect 563651 152556 563717 152557
rect 563651 152492 563652 152556
rect 563716 152492 563717 152556
rect 563651 152491 563717 152492
rect 563654 21181 563714 152491
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 565126 27301 565186 679491
rect 565307 663780 565373 663781
rect 565307 663716 565308 663780
rect 565372 663716 565373 663780
rect 565307 663715 565373 663716
rect 565123 27300 565189 27301
rect 565123 27236 565124 27300
rect 565188 27236 565189 27300
rect 565123 27235 565189 27236
rect 565310 27165 565370 663715
rect 565859 552124 565925 552125
rect 565859 552060 565860 552124
rect 565924 552060 565925 552124
rect 565859 552059 565925 552060
rect 565491 472700 565557 472701
rect 565491 472636 565492 472700
rect 565556 472636 565557 472700
rect 565491 472635 565557 472636
rect 565307 27164 565373 27165
rect 565307 27100 565308 27164
rect 565372 27100 565373 27164
rect 565307 27099 565373 27100
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 563651 21180 563717 21181
rect 563651 21116 563652 21180
rect 563716 21116 563717 21180
rect 563651 21115 563717 21116
rect 563467 6492 563533 6493
rect 563467 6428 563468 6492
rect 563532 6428 563533 6492
rect 563467 6427 563533 6428
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 -5146 564914 25398
rect 565494 24717 565554 472635
rect 565491 24716 565557 24717
rect 565491 24652 565492 24716
rect 565556 24652 565557 24716
rect 565491 24651 565557 24652
rect 565862 24037 565922 552059
rect 566046 249661 566106 700299
rect 566963 682412 567029 682413
rect 566963 682348 566964 682412
rect 567028 682348 567029 682412
rect 566963 682347 567029 682348
rect 566227 293180 566293 293181
rect 566227 293116 566228 293180
rect 566292 293116 566293 293180
rect 566227 293115 566293 293116
rect 566043 249660 566109 249661
rect 566043 249596 566044 249660
rect 566108 249596 566109 249660
rect 566043 249595 566109 249596
rect 566043 155276 566109 155277
rect 566043 155212 566044 155276
rect 566108 155212 566109 155276
rect 566043 155211 566109 155212
rect 566046 67693 566106 155211
rect 566043 67692 566109 67693
rect 566043 67628 566044 67692
rect 566108 67628 566109 67692
rect 566043 67627 566109 67628
rect 565859 24036 565925 24037
rect 565859 23972 565860 24036
rect 565924 23972 565925 24036
rect 565859 23971 565925 23972
rect 566230 3909 566290 293115
rect 566411 151468 566477 151469
rect 566411 151404 566412 151468
rect 566476 151404 566477 151468
rect 566411 151403 566477 151404
rect 566414 112437 566474 151403
rect 566411 112436 566477 112437
rect 566411 112372 566412 112436
rect 566476 112372 566477 112436
rect 566411 112371 566477 112372
rect 566966 25669 567026 682347
rect 568794 678454 569414 710042
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 569907 684860 569973 684861
rect 569907 684796 569908 684860
rect 569972 684796 569973 684860
rect 569907 684795 569973 684796
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 567331 586260 567397 586261
rect 567331 586196 567332 586260
rect 567396 586196 567397 586260
rect 567331 586195 567397 586196
rect 566963 25668 567029 25669
rect 566963 25604 566964 25668
rect 567028 25604 567029 25668
rect 566963 25603 567029 25604
rect 567334 24445 567394 586195
rect 567515 580820 567581 580821
rect 567515 580756 567516 580820
rect 567580 580756 567581 580820
rect 567515 580755 567581 580756
rect 567331 24444 567397 24445
rect 567331 24380 567332 24444
rect 567396 24380 567397 24444
rect 567331 24379 567397 24380
rect 567518 24309 567578 580755
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568619 566540 568685 566541
rect 568619 566476 568620 566540
rect 568684 566476 568685 566540
rect 568619 566475 568685 566476
rect 567699 286380 567765 286381
rect 567699 286316 567700 286380
rect 567764 286316 567765 286380
rect 567699 286315 567765 286316
rect 567515 24308 567581 24309
rect 567515 24244 567516 24308
rect 567580 24244 567581 24308
rect 567515 24243 567581 24244
rect 567702 21453 567762 286315
rect 568622 24173 568682 566475
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568619 24172 568685 24173
rect 568619 24108 568620 24172
rect 568684 24108 568685 24172
rect 568619 24107 568685 24108
rect 567699 21452 567765 21453
rect 567699 21388 567700 21452
rect 567764 21388 567765 21452
rect 567699 21387 567765 21388
rect 566227 3908 566293 3909
rect 566227 3844 566228 3908
rect 566292 3844 566293 3908
rect 566227 3843 566293 3844
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 -6106 569414 29898
rect 569910 14789 569970 684795
rect 573294 682954 573914 711002
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 575427 685268 575493 685269
rect 575427 685204 575428 685268
rect 575492 685204 575493 685268
rect 575427 685203 575493 685204
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 570091 681188 570157 681189
rect 570091 681124 570092 681188
rect 570156 681124 570157 681188
rect 570091 681123 570157 681124
rect 570094 17373 570154 681123
rect 570275 666500 570341 666501
rect 570275 666436 570276 666500
rect 570340 666436 570341 666500
rect 570275 666435 570341 666436
rect 570278 20909 570338 666435
rect 573294 646954 573914 682398
rect 574139 682004 574205 682005
rect 574139 681940 574140 682004
rect 574204 681940 574205 682004
rect 574139 681939 574205 681940
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 572667 625292 572733 625293
rect 572667 625228 572668 625292
rect 572732 625228 572733 625292
rect 572667 625227 572733 625228
rect 571379 601900 571445 601901
rect 571379 601836 571380 601900
rect 571444 601836 571445 601900
rect 571379 601835 571445 601836
rect 570275 20908 570341 20909
rect 570275 20844 570276 20908
rect 570340 20844 570341 20908
rect 570275 20843 570341 20844
rect 570091 17372 570157 17373
rect 570091 17308 570092 17372
rect 570156 17308 570157 17372
rect 570091 17307 570157 17308
rect 569907 14788 569973 14789
rect 569907 14724 569908 14788
rect 569972 14724 569973 14788
rect 569907 14723 569973 14724
rect 571382 3365 571442 601835
rect 571563 582180 571629 582181
rect 571563 582116 571564 582180
rect 571628 582116 571629 582180
rect 571563 582115 571629 582116
rect 571566 20773 571626 582115
rect 571563 20772 571629 20773
rect 571563 20708 571564 20772
rect 571628 20708 571629 20772
rect 571563 20707 571629 20708
rect 572670 19141 572730 625227
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 572667 19140 572733 19141
rect 572667 19076 572668 19140
rect 572732 19076 572733 19140
rect 572667 19075 572733 19076
rect 571379 3364 571445 3365
rect 571379 3300 571380 3364
rect 571444 3300 571445 3364
rect 571379 3299 571445 3300
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 -7066 573914 34398
rect 574142 18869 574202 681939
rect 574323 544780 574389 544781
rect 574323 544716 574324 544780
rect 574388 544716 574389 544780
rect 574323 544715 574389 544716
rect 574139 18868 574205 18869
rect 574139 18804 574140 18868
rect 574204 18804 574205 18868
rect 574139 18803 574205 18804
rect 574326 3773 574386 544715
rect 574323 3772 574389 3773
rect 574323 3708 574324 3772
rect 574388 3708 574389 3772
rect 574323 3707 574389 3708
rect 575430 3637 575490 685203
rect 577794 651454 578414 686898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 579659 685132 579725 685133
rect 579659 685068 579660 685132
rect 579724 685068 579725 685132
rect 579659 685067 579725 685068
rect 578555 680508 578621 680509
rect 578555 680444 578556 680508
rect 578620 680444 578621 680508
rect 578555 680443 578621 680444
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 576899 627060 576965 627061
rect 576899 626996 576900 627060
rect 576964 626996 576965 627060
rect 576899 626995 576965 626996
rect 575611 612780 575677 612781
rect 575611 612716 575612 612780
rect 575676 612716 575677 612780
rect 575611 612715 575677 612716
rect 575614 25805 575674 612715
rect 575611 25804 575677 25805
rect 575611 25740 575612 25804
rect 575676 25740 575677 25804
rect 575611 25739 575677 25740
rect 576902 18597 576962 626995
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 576899 18596 576965 18597
rect 576899 18532 576900 18596
rect 576964 18532 576965 18596
rect 576899 18531 576965 18532
rect 575427 3636 575493 3637
rect 575427 3572 575428 3636
rect 575492 3572 575493 3636
rect 575427 3571 575493 3572
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 3454 578414 38898
rect 578558 23765 578618 680443
rect 578739 646100 578805 646101
rect 578739 646036 578740 646100
rect 578804 646036 578805 646100
rect 578739 646035 578805 646036
rect 578742 24037 578802 646035
rect 578739 24036 578805 24037
rect 578739 23972 578740 24036
rect 578804 23972 578805 24036
rect 578739 23971 578805 23972
rect 578555 23764 578621 23765
rect 578555 23700 578556 23764
rect 578620 23700 578621 23764
rect 578555 23699 578621 23700
rect 579662 14653 579722 685067
rect 580947 669900 581013 669901
rect 580947 669836 580948 669900
rect 581012 669836 581013 669900
rect 580947 669835 581013 669836
rect 579843 435980 579909 435981
rect 579843 435916 579844 435980
rect 579908 435916 579909 435980
rect 579843 435915 579909 435916
rect 579846 17781 579906 435915
rect 579843 17780 579909 17781
rect 579843 17716 579844 17780
rect 579908 17716 579909 17780
rect 579843 17715 579909 17716
rect 580950 17645 581010 669835
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 580947 17644 581013 17645
rect 580947 17580 580948 17644
rect 581012 17580 581013 17644
rect 580947 17579 581013 17580
rect 579659 14652 579725 14653
rect 579659 14588 579660 14652
rect 579724 14588 579725 14652
rect 579659 14587 579725 14588
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 34328 655718 34564 655954
rect 34328 655398 34564 655634
rect 170056 655718 170292 655954
rect 170056 655398 170292 655634
rect 35008 651218 35244 651454
rect 35008 650898 35244 651134
rect 169376 651218 169612 651454
rect 169376 650898 169612 651134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 34328 619718 34564 619954
rect 34328 619398 34564 619634
rect 170056 619718 170292 619954
rect 170056 619398 170292 619634
rect 35008 615218 35244 615454
rect 35008 614898 35244 615134
rect 169376 615218 169612 615454
rect 169376 614898 169612 615134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 206328 655718 206564 655954
rect 206328 655398 206564 655634
rect 342056 655718 342292 655954
rect 342056 655398 342292 655634
rect 207008 651218 207244 651454
rect 207008 650898 207244 651134
rect 341376 651218 341612 651454
rect 341376 650898 341612 651134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 206328 619718 206564 619954
rect 206328 619398 206564 619634
rect 342056 619718 342292 619954
rect 342056 619398 342292 619634
rect 207008 615218 207244 615454
rect 207008 614898 207244 615134
rect 341376 615218 341612 615454
rect 341376 614898 341612 615134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 67610 547718 67846 547954
rect 67610 547398 67846 547634
rect 98330 547718 98566 547954
rect 98330 547398 98566 547634
rect 129050 547718 129286 547954
rect 129050 547398 129286 547634
rect 159770 547718 160006 547954
rect 159770 547398 160006 547634
rect 190490 547718 190726 547954
rect 190490 547398 190726 547634
rect 221210 547718 221446 547954
rect 221210 547398 221446 547634
rect 251930 547718 252166 547954
rect 251930 547398 252166 547634
rect 282650 547718 282886 547954
rect 282650 547398 282886 547634
rect 313370 547718 313606 547954
rect 313370 547398 313606 547634
rect 344090 547718 344326 547954
rect 344090 547398 344326 547634
rect 52250 543218 52486 543454
rect 52250 542898 52486 543134
rect 82970 543218 83206 543454
rect 82970 542898 83206 543134
rect 113690 543218 113926 543454
rect 113690 542898 113926 543134
rect 144410 543218 144646 543454
rect 144410 542898 144646 543134
rect 175130 543218 175366 543454
rect 175130 542898 175366 543134
rect 205850 543218 206086 543454
rect 205850 542898 206086 543134
rect 236570 543218 236806 543454
rect 236570 542898 236806 543134
rect 267290 543218 267526 543454
rect 267290 542898 267526 543134
rect 298010 543218 298246 543454
rect 298010 542898 298246 543134
rect 328730 543218 328966 543454
rect 328730 542898 328966 543134
rect 67610 511718 67846 511954
rect 67610 511398 67846 511634
rect 98330 511718 98566 511954
rect 98330 511398 98566 511634
rect 129050 511718 129286 511954
rect 129050 511398 129286 511634
rect 159770 511718 160006 511954
rect 159770 511398 160006 511634
rect 190490 511718 190726 511954
rect 190490 511398 190726 511634
rect 221210 511718 221446 511954
rect 221210 511398 221446 511634
rect 251930 511718 252166 511954
rect 251930 511398 252166 511634
rect 282650 511718 282886 511954
rect 282650 511398 282886 511634
rect 313370 511718 313606 511954
rect 313370 511398 313606 511634
rect 344090 511718 344326 511954
rect 344090 511398 344326 511634
rect 52250 507218 52486 507454
rect 52250 506898 52486 507134
rect 82970 507218 83206 507454
rect 82970 506898 83206 507134
rect 113690 507218 113926 507454
rect 113690 506898 113926 507134
rect 144410 507218 144646 507454
rect 144410 506898 144646 507134
rect 175130 507218 175366 507454
rect 175130 506898 175366 507134
rect 205850 507218 206086 507454
rect 205850 506898 206086 507134
rect 236570 507218 236806 507454
rect 236570 506898 236806 507134
rect 267290 507218 267526 507454
rect 267290 506898 267526 507134
rect 298010 507218 298246 507454
rect 298010 506898 298246 507134
rect 328730 507218 328966 507454
rect 328730 506898 328966 507134
rect 67610 475718 67846 475954
rect 67610 475398 67846 475634
rect 98330 475718 98566 475954
rect 98330 475398 98566 475634
rect 129050 475718 129286 475954
rect 129050 475398 129286 475634
rect 159770 475718 160006 475954
rect 159770 475398 160006 475634
rect 190490 475718 190726 475954
rect 190490 475398 190726 475634
rect 221210 475718 221446 475954
rect 221210 475398 221446 475634
rect 251930 475718 252166 475954
rect 251930 475398 252166 475634
rect 282650 475718 282886 475954
rect 282650 475398 282886 475634
rect 313370 475718 313606 475954
rect 313370 475398 313606 475634
rect 344090 475718 344326 475954
rect 344090 475398 344326 475634
rect 52250 471218 52486 471454
rect 52250 470898 52486 471134
rect 82970 471218 83206 471454
rect 82970 470898 83206 471134
rect 113690 471218 113926 471454
rect 113690 470898 113926 471134
rect 144410 471218 144646 471454
rect 144410 470898 144646 471134
rect 175130 471218 175366 471454
rect 175130 470898 175366 471134
rect 205850 471218 206086 471454
rect 205850 470898 206086 471134
rect 236570 471218 236806 471454
rect 236570 470898 236806 471134
rect 267290 471218 267526 471454
rect 267290 470898 267526 471134
rect 298010 471218 298246 471454
rect 298010 470898 298246 471134
rect 328730 471218 328966 471454
rect 328730 470898 328966 471134
rect 67610 439718 67846 439954
rect 67610 439398 67846 439634
rect 98330 439718 98566 439954
rect 98330 439398 98566 439634
rect 129050 439718 129286 439954
rect 129050 439398 129286 439634
rect 159770 439718 160006 439954
rect 159770 439398 160006 439634
rect 190490 439718 190726 439954
rect 190490 439398 190726 439634
rect 221210 439718 221446 439954
rect 221210 439398 221446 439634
rect 251930 439718 252166 439954
rect 251930 439398 252166 439634
rect 282650 439718 282886 439954
rect 282650 439398 282886 439634
rect 313370 439718 313606 439954
rect 313370 439398 313606 439634
rect 344090 439718 344326 439954
rect 344090 439398 344326 439634
rect 52250 435218 52486 435454
rect 52250 434898 52486 435134
rect 82970 435218 83206 435454
rect 82970 434898 83206 435134
rect 113690 435218 113926 435454
rect 113690 434898 113926 435134
rect 144410 435218 144646 435454
rect 144410 434898 144646 435134
rect 175130 435218 175366 435454
rect 175130 434898 175366 435134
rect 205850 435218 206086 435454
rect 205850 434898 206086 435134
rect 236570 435218 236806 435454
rect 236570 434898 236806 435134
rect 267290 435218 267526 435454
rect 267290 434898 267526 435134
rect 298010 435218 298246 435454
rect 298010 434898 298246 435134
rect 328730 435218 328966 435454
rect 328730 434898 328966 435134
rect 67610 403718 67846 403954
rect 67610 403398 67846 403634
rect 98330 403718 98566 403954
rect 98330 403398 98566 403634
rect 129050 403718 129286 403954
rect 129050 403398 129286 403634
rect 159770 403718 160006 403954
rect 159770 403398 160006 403634
rect 190490 403718 190726 403954
rect 190490 403398 190726 403634
rect 221210 403718 221446 403954
rect 221210 403398 221446 403634
rect 251930 403718 252166 403954
rect 251930 403398 252166 403634
rect 282650 403718 282886 403954
rect 282650 403398 282886 403634
rect 313370 403718 313606 403954
rect 313370 403398 313606 403634
rect 344090 403718 344326 403954
rect 344090 403398 344326 403634
rect 52250 399218 52486 399454
rect 52250 398898 52486 399134
rect 82970 399218 83206 399454
rect 82970 398898 83206 399134
rect 113690 399218 113926 399454
rect 113690 398898 113926 399134
rect 144410 399218 144646 399454
rect 144410 398898 144646 399134
rect 175130 399218 175366 399454
rect 175130 398898 175366 399134
rect 205850 399218 206086 399454
rect 205850 398898 206086 399134
rect 236570 399218 236806 399454
rect 236570 398898 236806 399134
rect 267290 399218 267526 399454
rect 267290 398898 267526 399134
rect 298010 399218 298246 399454
rect 298010 398898 298246 399134
rect 328730 399218 328966 399454
rect 328730 398898 328966 399134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 67610 367718 67846 367954
rect 67610 367398 67846 367634
rect 98330 367718 98566 367954
rect 98330 367398 98566 367634
rect 129050 367718 129286 367954
rect 129050 367398 129286 367634
rect 159770 367718 160006 367954
rect 159770 367398 160006 367634
rect 190490 367718 190726 367954
rect 190490 367398 190726 367634
rect 221210 367718 221446 367954
rect 221210 367398 221446 367634
rect 251930 367718 252166 367954
rect 251930 367398 252166 367634
rect 282650 367718 282886 367954
rect 282650 367398 282886 367634
rect 313370 367718 313606 367954
rect 313370 367398 313606 367634
rect 344090 367718 344326 367954
rect 344090 367398 344326 367634
rect 52250 363218 52486 363454
rect 52250 362898 52486 363134
rect 82970 363218 83206 363454
rect 82970 362898 83206 363134
rect 113690 363218 113926 363454
rect 113690 362898 113926 363134
rect 144410 363218 144646 363454
rect 144410 362898 144646 363134
rect 175130 363218 175366 363454
rect 175130 362898 175366 363134
rect 205850 363218 206086 363454
rect 205850 362898 206086 363134
rect 236570 363218 236806 363454
rect 236570 362898 236806 363134
rect 267290 363218 267526 363454
rect 267290 362898 267526 363134
rect 298010 363218 298246 363454
rect 298010 362898 298246 363134
rect 328730 363218 328966 363454
rect 328730 362898 328966 363134
rect 67610 331718 67846 331954
rect 67610 331398 67846 331634
rect 98330 331718 98566 331954
rect 98330 331398 98566 331634
rect 129050 331718 129286 331954
rect 129050 331398 129286 331634
rect 159770 331718 160006 331954
rect 159770 331398 160006 331634
rect 190490 331718 190726 331954
rect 190490 331398 190726 331634
rect 221210 331718 221446 331954
rect 221210 331398 221446 331634
rect 251930 331718 252166 331954
rect 251930 331398 252166 331634
rect 282650 331718 282886 331954
rect 282650 331398 282886 331634
rect 313370 331718 313606 331954
rect 313370 331398 313606 331634
rect 344090 331718 344326 331954
rect 344090 331398 344326 331634
rect 52250 327218 52486 327454
rect 52250 326898 52486 327134
rect 82970 327218 83206 327454
rect 82970 326898 83206 327134
rect 113690 327218 113926 327454
rect 113690 326898 113926 327134
rect 144410 327218 144646 327454
rect 144410 326898 144646 327134
rect 175130 327218 175366 327454
rect 175130 326898 175366 327134
rect 205850 327218 206086 327454
rect 205850 326898 206086 327134
rect 236570 327218 236806 327454
rect 236570 326898 236806 327134
rect 267290 327218 267526 327454
rect 267290 326898 267526 327134
rect 298010 327218 298246 327454
rect 298010 326898 298246 327134
rect 328730 327218 328966 327454
rect 328730 326898 328966 327134
rect 67610 295718 67846 295954
rect 67610 295398 67846 295634
rect 98330 295718 98566 295954
rect 98330 295398 98566 295634
rect 129050 295718 129286 295954
rect 129050 295398 129286 295634
rect 159770 295718 160006 295954
rect 159770 295398 160006 295634
rect 190490 295718 190726 295954
rect 190490 295398 190726 295634
rect 221210 295718 221446 295954
rect 221210 295398 221446 295634
rect 251930 295718 252166 295954
rect 251930 295398 252166 295634
rect 282650 295718 282886 295954
rect 282650 295398 282886 295634
rect 313370 295718 313606 295954
rect 313370 295398 313606 295634
rect 344090 295718 344326 295954
rect 344090 295398 344326 295634
rect 52250 291218 52486 291454
rect 52250 290898 52486 291134
rect 82970 291218 83206 291454
rect 82970 290898 83206 291134
rect 113690 291218 113926 291454
rect 113690 290898 113926 291134
rect 144410 291218 144646 291454
rect 144410 290898 144646 291134
rect 175130 291218 175366 291454
rect 175130 290898 175366 291134
rect 205850 291218 206086 291454
rect 205850 290898 206086 291134
rect 236570 291218 236806 291454
rect 236570 290898 236806 291134
rect 267290 291218 267526 291454
rect 267290 290898 267526 291134
rect 298010 291218 298246 291454
rect 298010 290898 298246 291134
rect 328730 291218 328966 291454
rect 328730 290898 328966 291134
rect 67610 259718 67846 259954
rect 67610 259398 67846 259634
rect 98330 259718 98566 259954
rect 98330 259398 98566 259634
rect 129050 259718 129286 259954
rect 129050 259398 129286 259634
rect 159770 259718 160006 259954
rect 159770 259398 160006 259634
rect 190490 259718 190726 259954
rect 190490 259398 190726 259634
rect 221210 259718 221446 259954
rect 221210 259398 221446 259634
rect 251930 259718 252166 259954
rect 251930 259398 252166 259634
rect 282650 259718 282886 259954
rect 282650 259398 282886 259634
rect 313370 259718 313606 259954
rect 313370 259398 313606 259634
rect 344090 259718 344326 259954
rect 344090 259398 344326 259634
rect 52250 255218 52486 255454
rect 52250 254898 52486 255134
rect 82970 255218 83206 255454
rect 82970 254898 83206 255134
rect 113690 255218 113926 255454
rect 113690 254898 113926 255134
rect 144410 255218 144646 255454
rect 144410 254898 144646 255134
rect 175130 255218 175366 255454
rect 175130 254898 175366 255134
rect 205850 255218 206086 255454
rect 205850 254898 206086 255134
rect 236570 255218 236806 255454
rect 236570 254898 236806 255134
rect 267290 255218 267526 255454
rect 267290 254898 267526 255134
rect 298010 255218 298246 255454
rect 298010 254898 298246 255134
rect 328730 255218 328966 255454
rect 328730 254898 328966 255134
rect 67610 223718 67846 223954
rect 67610 223398 67846 223634
rect 98330 223718 98566 223954
rect 98330 223398 98566 223634
rect 129050 223718 129286 223954
rect 129050 223398 129286 223634
rect 159770 223718 160006 223954
rect 159770 223398 160006 223634
rect 190490 223718 190726 223954
rect 190490 223398 190726 223634
rect 221210 223718 221446 223954
rect 221210 223398 221446 223634
rect 251930 223718 252166 223954
rect 251930 223398 252166 223634
rect 282650 223718 282886 223954
rect 282650 223398 282886 223634
rect 313370 223718 313606 223954
rect 313370 223398 313606 223634
rect 344090 223718 344326 223954
rect 344090 223398 344326 223634
rect 52250 219218 52486 219454
rect 52250 218898 52486 219134
rect 82970 219218 83206 219454
rect 82970 218898 83206 219134
rect 113690 219218 113926 219454
rect 113690 218898 113926 219134
rect 144410 219218 144646 219454
rect 144410 218898 144646 219134
rect 175130 219218 175366 219454
rect 175130 218898 175366 219134
rect 205850 219218 206086 219454
rect 205850 218898 206086 219134
rect 236570 219218 236806 219454
rect 236570 218898 236806 219134
rect 267290 219218 267526 219454
rect 267290 218898 267526 219134
rect 298010 219218 298246 219454
rect 298010 218898 298246 219134
rect 328730 219218 328966 219454
rect 328730 218898 328966 219134
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 429610 655718 429846 655954
rect 429610 655398 429846 655634
rect 460330 655718 460566 655954
rect 460330 655398 460566 655634
rect 491050 655718 491286 655954
rect 491050 655398 491286 655634
rect 521770 655718 522006 655954
rect 521770 655398 522006 655634
rect 414250 651218 414486 651454
rect 414250 650898 414486 651134
rect 444970 651218 445206 651454
rect 444970 650898 445206 651134
rect 475690 651218 475926 651454
rect 475690 650898 475926 651134
rect 506410 651218 506646 651454
rect 506410 650898 506646 651134
rect 537130 651218 537366 651454
rect 537130 650898 537366 651134
rect 429610 619718 429846 619954
rect 429610 619398 429846 619634
rect 460330 619718 460566 619954
rect 460330 619398 460566 619634
rect 491050 619718 491286 619954
rect 491050 619398 491286 619634
rect 521770 619718 522006 619954
rect 521770 619398 522006 619634
rect 414250 615218 414486 615454
rect 414250 614898 414486 615134
rect 444970 615218 445206 615454
rect 444970 614898 445206 615134
rect 475690 615218 475926 615454
rect 475690 614898 475926 615134
rect 506410 615218 506646 615454
rect 506410 614898 506646 615134
rect 537130 615218 537366 615454
rect 537130 614898 537366 615134
rect 429610 583718 429846 583954
rect 429610 583398 429846 583634
rect 460330 583718 460566 583954
rect 460330 583398 460566 583634
rect 491050 583718 491286 583954
rect 491050 583398 491286 583634
rect 521770 583718 522006 583954
rect 521770 583398 522006 583634
rect 414250 579218 414486 579454
rect 414250 578898 414486 579134
rect 444970 579218 445206 579454
rect 444970 578898 445206 579134
rect 475690 579218 475926 579454
rect 475690 578898 475926 579134
rect 506410 579218 506646 579454
rect 506410 578898 506646 579134
rect 537130 579218 537366 579454
rect 537130 578898 537366 579134
rect 429610 547718 429846 547954
rect 429610 547398 429846 547634
rect 460330 547718 460566 547954
rect 460330 547398 460566 547634
rect 491050 547718 491286 547954
rect 491050 547398 491286 547634
rect 521770 547718 522006 547954
rect 521770 547398 522006 547634
rect 414250 543218 414486 543454
rect 414250 542898 414486 543134
rect 444970 543218 445206 543454
rect 444970 542898 445206 543134
rect 475690 543218 475926 543454
rect 475690 542898 475926 543134
rect 506410 543218 506646 543454
rect 506410 542898 506646 543134
rect 537130 543218 537366 543454
rect 537130 542898 537366 543134
rect 429610 511718 429846 511954
rect 429610 511398 429846 511634
rect 460330 511718 460566 511954
rect 460330 511398 460566 511634
rect 491050 511718 491286 511954
rect 491050 511398 491286 511634
rect 521770 511718 522006 511954
rect 521770 511398 522006 511634
rect 414250 507218 414486 507454
rect 414250 506898 414486 507134
rect 444970 507218 445206 507454
rect 444970 506898 445206 507134
rect 475690 507218 475926 507454
rect 475690 506898 475926 507134
rect 506410 507218 506646 507454
rect 506410 506898 506646 507134
rect 537130 507218 537366 507454
rect 537130 506898 537366 507134
rect 429610 475718 429846 475954
rect 429610 475398 429846 475634
rect 460330 475718 460566 475954
rect 460330 475398 460566 475634
rect 491050 475718 491286 475954
rect 491050 475398 491286 475634
rect 521770 475718 522006 475954
rect 521770 475398 522006 475634
rect 414250 471218 414486 471454
rect 414250 470898 414486 471134
rect 444970 471218 445206 471454
rect 444970 470898 445206 471134
rect 475690 471218 475926 471454
rect 475690 470898 475926 471134
rect 506410 471218 506646 471454
rect 506410 470898 506646 471134
rect 537130 471218 537366 471454
rect 537130 470898 537366 471134
rect 429610 439718 429846 439954
rect 429610 439398 429846 439634
rect 460330 439718 460566 439954
rect 460330 439398 460566 439634
rect 491050 439718 491286 439954
rect 491050 439398 491286 439634
rect 521770 439718 522006 439954
rect 521770 439398 522006 439634
rect 414250 435218 414486 435454
rect 414250 434898 414486 435134
rect 444970 435218 445206 435454
rect 444970 434898 445206 435134
rect 475690 435218 475926 435454
rect 475690 434898 475926 435134
rect 506410 435218 506646 435454
rect 506410 434898 506646 435134
rect 537130 435218 537366 435454
rect 537130 434898 537366 435134
rect 429610 403718 429846 403954
rect 429610 403398 429846 403634
rect 460330 403718 460566 403954
rect 460330 403398 460566 403634
rect 491050 403718 491286 403954
rect 491050 403398 491286 403634
rect 521770 403718 522006 403954
rect 521770 403398 522006 403634
rect 414250 399218 414486 399454
rect 414250 398898 414486 399134
rect 444970 399218 445206 399454
rect 444970 398898 445206 399134
rect 475690 399218 475926 399454
rect 475690 398898 475926 399134
rect 506410 399218 506646 399454
rect 506410 398898 506646 399134
rect 537130 399218 537366 399454
rect 537130 398898 537366 399134
rect 429610 367718 429846 367954
rect 429610 367398 429846 367634
rect 460330 367718 460566 367954
rect 460330 367398 460566 367634
rect 491050 367718 491286 367954
rect 491050 367398 491286 367634
rect 521770 367718 522006 367954
rect 521770 367398 522006 367634
rect 414250 363218 414486 363454
rect 414250 362898 414486 363134
rect 444970 363218 445206 363454
rect 444970 362898 445206 363134
rect 475690 363218 475926 363454
rect 475690 362898 475926 363134
rect 506410 363218 506646 363454
rect 506410 362898 506646 363134
rect 537130 363218 537366 363454
rect 537130 362898 537366 363134
rect 429610 331718 429846 331954
rect 429610 331398 429846 331634
rect 460330 331718 460566 331954
rect 460330 331398 460566 331634
rect 491050 331718 491286 331954
rect 491050 331398 491286 331634
rect 521770 331718 522006 331954
rect 521770 331398 522006 331634
rect 414250 327218 414486 327454
rect 414250 326898 414486 327134
rect 444970 327218 445206 327454
rect 444970 326898 445206 327134
rect 475690 327218 475926 327454
rect 475690 326898 475926 327134
rect 506410 327218 506646 327454
rect 506410 326898 506646 327134
rect 537130 327218 537366 327454
rect 537130 326898 537366 327134
rect 429610 295718 429846 295954
rect 429610 295398 429846 295634
rect 460330 295718 460566 295954
rect 460330 295398 460566 295634
rect 491050 295718 491286 295954
rect 491050 295398 491286 295634
rect 521770 295718 522006 295954
rect 521770 295398 522006 295634
rect 414250 291218 414486 291454
rect 414250 290898 414486 291134
rect 444970 291218 445206 291454
rect 444970 290898 445206 291134
rect 475690 291218 475926 291454
rect 475690 290898 475926 291134
rect 506410 291218 506646 291454
rect 506410 290898 506646 291134
rect 537130 291218 537366 291454
rect 537130 290898 537366 291134
rect 429610 259718 429846 259954
rect 429610 259398 429846 259634
rect 460330 259718 460566 259954
rect 460330 259398 460566 259634
rect 491050 259718 491286 259954
rect 491050 259398 491286 259634
rect 521770 259718 522006 259954
rect 521770 259398 522006 259634
rect 414250 255218 414486 255454
rect 414250 254898 414486 255134
rect 444970 255218 445206 255454
rect 444970 254898 445206 255134
rect 475690 255218 475926 255454
rect 475690 254898 475926 255134
rect 506410 255218 506646 255454
rect 506410 254898 506646 255134
rect 537130 255218 537366 255454
rect 537130 254898 537366 255134
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 248570 147218 248806 147454
rect 248570 146898 248806 147134
rect 279290 147218 279526 147454
rect 279290 146898 279526 147134
rect 310010 147218 310246 147454
rect 310010 146898 310246 147134
rect 340730 147218 340966 147454
rect 340730 146898 340966 147134
rect 371450 147218 371686 147454
rect 371450 146898 371686 147134
rect 402170 147218 402406 147454
rect 402170 146898 402406 147134
rect 432890 147218 433126 147454
rect 432890 146898 433126 147134
rect 463610 147218 463846 147454
rect 463610 146898 463846 147134
rect 494330 147218 494566 147454
rect 494330 146898 494566 147134
rect 525050 147218 525286 147454
rect 525050 146898 525286 147134
rect 79610 115718 79846 115954
rect 79610 115398 79846 115634
rect 110330 115718 110566 115954
rect 110330 115398 110566 115634
rect 141050 115718 141286 115954
rect 141050 115398 141286 115634
rect 171770 115718 172006 115954
rect 171770 115398 172006 115634
rect 202490 115718 202726 115954
rect 202490 115398 202726 115634
rect 233210 115718 233446 115954
rect 233210 115398 233446 115634
rect 263930 115718 264166 115954
rect 263930 115398 264166 115634
rect 294650 115718 294886 115954
rect 294650 115398 294886 115634
rect 325370 115718 325606 115954
rect 325370 115398 325606 115634
rect 356090 115718 356326 115954
rect 356090 115398 356326 115634
rect 386810 115718 387046 115954
rect 386810 115398 387046 115634
rect 417530 115718 417766 115954
rect 417530 115398 417766 115634
rect 448250 115718 448486 115954
rect 448250 115398 448486 115634
rect 478970 115718 479206 115954
rect 478970 115398 479206 115634
rect 509690 115718 509926 115954
rect 509690 115398 509926 115634
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 248570 111218 248806 111454
rect 248570 110898 248806 111134
rect 279290 111218 279526 111454
rect 279290 110898 279526 111134
rect 310010 111218 310246 111454
rect 310010 110898 310246 111134
rect 340730 111218 340966 111454
rect 340730 110898 340966 111134
rect 371450 111218 371686 111454
rect 371450 110898 371686 111134
rect 402170 111218 402406 111454
rect 402170 110898 402406 111134
rect 432890 111218 433126 111454
rect 432890 110898 433126 111134
rect 463610 111218 463846 111454
rect 463610 110898 463846 111134
rect 494330 111218 494566 111454
rect 494330 110898 494566 111134
rect 525050 111218 525286 111454
rect 525050 110898 525286 111134
rect 79610 79718 79846 79954
rect 79610 79398 79846 79634
rect 110330 79718 110566 79954
rect 110330 79398 110566 79634
rect 141050 79718 141286 79954
rect 141050 79398 141286 79634
rect 171770 79718 172006 79954
rect 171770 79398 172006 79634
rect 202490 79718 202726 79954
rect 202490 79398 202726 79634
rect 233210 79718 233446 79954
rect 233210 79398 233446 79634
rect 263930 79718 264166 79954
rect 263930 79398 264166 79634
rect 294650 79718 294886 79954
rect 294650 79398 294886 79634
rect 325370 79718 325606 79954
rect 325370 79398 325606 79634
rect 356090 79718 356326 79954
rect 356090 79398 356326 79634
rect 386810 79718 387046 79954
rect 386810 79398 387046 79634
rect 417530 79718 417766 79954
rect 417530 79398 417766 79634
rect 448250 79718 448486 79954
rect 448250 79398 448486 79634
rect 478970 79718 479206 79954
rect 478970 79398 479206 79634
rect 509690 79718 509926 79954
rect 509690 79398 509926 79634
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 248570 75218 248806 75454
rect 248570 74898 248806 75134
rect 279290 75218 279526 75454
rect 279290 74898 279526 75134
rect 310010 75218 310246 75454
rect 310010 74898 310246 75134
rect 340730 75218 340966 75454
rect 340730 74898 340966 75134
rect 371450 75218 371686 75454
rect 371450 74898 371686 75134
rect 402170 75218 402406 75454
rect 402170 74898 402406 75134
rect 432890 75218 433126 75454
rect 432890 74898 433126 75134
rect 463610 75218 463846 75454
rect 463610 74898 463846 75134
rect 494330 75218 494566 75454
rect 494330 74898 494566 75134
rect 525050 75218 525286 75454
rect 525050 74898 525286 75134
rect 79610 43718 79846 43954
rect 79610 43398 79846 43634
rect 110330 43718 110566 43954
rect 110330 43398 110566 43634
rect 141050 43718 141286 43954
rect 141050 43398 141286 43634
rect 171770 43718 172006 43954
rect 171770 43398 172006 43634
rect 202490 43718 202726 43954
rect 202490 43398 202726 43634
rect 233210 43718 233446 43954
rect 233210 43398 233446 43634
rect 263930 43718 264166 43954
rect 263930 43398 264166 43634
rect 294650 43718 294886 43954
rect 294650 43398 294886 43634
rect 325370 43718 325606 43954
rect 325370 43398 325606 43634
rect 356090 43718 356326 43954
rect 356090 43398 356326 43634
rect 386810 43718 387046 43954
rect 386810 43398 387046 43634
rect 417530 43718 417766 43954
rect 417530 43398 417766 43634
rect 448250 43718 448486 43954
rect 448250 43398 448486 43634
rect 478970 43718 479206 43954
rect 478970 43398 479206 43634
rect 509690 43718 509926 43954
rect 509690 43398 509926 43634
rect 64250 39218 64486 39454
rect 64250 38898 64486 39134
rect 94970 39218 95206 39454
rect 94970 38898 95206 39134
rect 125690 39218 125926 39454
rect 125690 38898 125926 39134
rect 156410 39218 156646 39454
rect 156410 38898 156646 39134
rect 187130 39218 187366 39454
rect 187130 38898 187366 39134
rect 217850 39218 218086 39454
rect 217850 38898 218086 39134
rect 248570 39218 248806 39454
rect 248570 38898 248806 39134
rect 279290 39218 279526 39454
rect 279290 38898 279526 39134
rect 310010 39218 310246 39454
rect 310010 38898 310246 39134
rect 340730 39218 340966 39454
rect 340730 38898 340966 39134
rect 371450 39218 371686 39454
rect 371450 38898 371686 39134
rect 402170 39218 402406 39454
rect 402170 38898 402406 39134
rect 432890 39218 433126 39454
rect 432890 38898 433126 39134
rect 463610 39218 463846 39454
rect 463610 38898 463846 39134
rect 494330 39218 494566 39454
rect 494330 38898 494566 39134
rect 525050 39218 525286 39454
rect 525050 38898 525286 39134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 34328 655954
rect 34564 655718 170056 655954
rect 170292 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 206328 655954
rect 206564 655718 342056 655954
rect 342292 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 429610 655954
rect 429846 655718 460330 655954
rect 460566 655718 491050 655954
rect 491286 655718 521770 655954
rect 522006 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 34328 655634
rect 34564 655398 170056 655634
rect 170292 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 206328 655634
rect 206564 655398 342056 655634
rect 342292 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 429610 655634
rect 429846 655398 460330 655634
rect 460566 655398 491050 655634
rect 491286 655398 521770 655634
rect 522006 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 35008 651454
rect 35244 651218 169376 651454
rect 169612 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 207008 651454
rect 207244 651218 341376 651454
rect 341612 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 414250 651454
rect 414486 651218 444970 651454
rect 445206 651218 475690 651454
rect 475926 651218 506410 651454
rect 506646 651218 537130 651454
rect 537366 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 35008 651134
rect 35244 650898 169376 651134
rect 169612 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 207008 651134
rect 207244 650898 341376 651134
rect 341612 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 414250 651134
rect 414486 650898 444970 651134
rect 445206 650898 475690 651134
rect 475926 650898 506410 651134
rect 506646 650898 537130 651134
rect 537366 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 34328 619954
rect 34564 619718 170056 619954
rect 170292 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 206328 619954
rect 206564 619718 342056 619954
rect 342292 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 429610 619954
rect 429846 619718 460330 619954
rect 460566 619718 491050 619954
rect 491286 619718 521770 619954
rect 522006 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 34328 619634
rect 34564 619398 170056 619634
rect 170292 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 206328 619634
rect 206564 619398 342056 619634
rect 342292 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 429610 619634
rect 429846 619398 460330 619634
rect 460566 619398 491050 619634
rect 491286 619398 521770 619634
rect 522006 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 35008 615454
rect 35244 615218 169376 615454
rect 169612 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 207008 615454
rect 207244 615218 341376 615454
rect 341612 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 414250 615454
rect 414486 615218 444970 615454
rect 445206 615218 475690 615454
rect 475926 615218 506410 615454
rect 506646 615218 537130 615454
rect 537366 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 35008 615134
rect 35244 614898 169376 615134
rect 169612 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 207008 615134
rect 207244 614898 341376 615134
rect 341612 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 414250 615134
rect 414486 614898 444970 615134
rect 445206 614898 475690 615134
rect 475926 614898 506410 615134
rect 506646 614898 537130 615134
rect 537366 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 429610 583954
rect 429846 583718 460330 583954
rect 460566 583718 491050 583954
rect 491286 583718 521770 583954
rect 522006 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 429610 583634
rect 429846 583398 460330 583634
rect 460566 583398 491050 583634
rect 491286 583398 521770 583634
rect 522006 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 414250 579454
rect 414486 579218 444970 579454
rect 445206 579218 475690 579454
rect 475926 579218 506410 579454
rect 506646 579218 537130 579454
rect 537366 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 414250 579134
rect 414486 578898 444970 579134
rect 445206 578898 475690 579134
rect 475926 578898 506410 579134
rect 506646 578898 537130 579134
rect 537366 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 67610 547954
rect 67846 547718 98330 547954
rect 98566 547718 129050 547954
rect 129286 547718 159770 547954
rect 160006 547718 190490 547954
rect 190726 547718 221210 547954
rect 221446 547718 251930 547954
rect 252166 547718 282650 547954
rect 282886 547718 313370 547954
rect 313606 547718 344090 547954
rect 344326 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 429610 547954
rect 429846 547718 460330 547954
rect 460566 547718 491050 547954
rect 491286 547718 521770 547954
rect 522006 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 67610 547634
rect 67846 547398 98330 547634
rect 98566 547398 129050 547634
rect 129286 547398 159770 547634
rect 160006 547398 190490 547634
rect 190726 547398 221210 547634
rect 221446 547398 251930 547634
rect 252166 547398 282650 547634
rect 282886 547398 313370 547634
rect 313606 547398 344090 547634
rect 344326 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 429610 547634
rect 429846 547398 460330 547634
rect 460566 547398 491050 547634
rect 491286 547398 521770 547634
rect 522006 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 52250 543454
rect 52486 543218 82970 543454
rect 83206 543218 113690 543454
rect 113926 543218 144410 543454
rect 144646 543218 175130 543454
rect 175366 543218 205850 543454
rect 206086 543218 236570 543454
rect 236806 543218 267290 543454
rect 267526 543218 298010 543454
rect 298246 543218 328730 543454
rect 328966 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 414250 543454
rect 414486 543218 444970 543454
rect 445206 543218 475690 543454
rect 475926 543218 506410 543454
rect 506646 543218 537130 543454
rect 537366 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 52250 543134
rect 52486 542898 82970 543134
rect 83206 542898 113690 543134
rect 113926 542898 144410 543134
rect 144646 542898 175130 543134
rect 175366 542898 205850 543134
rect 206086 542898 236570 543134
rect 236806 542898 267290 543134
rect 267526 542898 298010 543134
rect 298246 542898 328730 543134
rect 328966 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 414250 543134
rect 414486 542898 444970 543134
rect 445206 542898 475690 543134
rect 475926 542898 506410 543134
rect 506646 542898 537130 543134
rect 537366 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 67610 511954
rect 67846 511718 98330 511954
rect 98566 511718 129050 511954
rect 129286 511718 159770 511954
rect 160006 511718 190490 511954
rect 190726 511718 221210 511954
rect 221446 511718 251930 511954
rect 252166 511718 282650 511954
rect 282886 511718 313370 511954
rect 313606 511718 344090 511954
rect 344326 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 429610 511954
rect 429846 511718 460330 511954
rect 460566 511718 491050 511954
rect 491286 511718 521770 511954
rect 522006 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 67610 511634
rect 67846 511398 98330 511634
rect 98566 511398 129050 511634
rect 129286 511398 159770 511634
rect 160006 511398 190490 511634
rect 190726 511398 221210 511634
rect 221446 511398 251930 511634
rect 252166 511398 282650 511634
rect 282886 511398 313370 511634
rect 313606 511398 344090 511634
rect 344326 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 429610 511634
rect 429846 511398 460330 511634
rect 460566 511398 491050 511634
rect 491286 511398 521770 511634
rect 522006 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 52250 507454
rect 52486 507218 82970 507454
rect 83206 507218 113690 507454
rect 113926 507218 144410 507454
rect 144646 507218 175130 507454
rect 175366 507218 205850 507454
rect 206086 507218 236570 507454
rect 236806 507218 267290 507454
rect 267526 507218 298010 507454
rect 298246 507218 328730 507454
rect 328966 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 414250 507454
rect 414486 507218 444970 507454
rect 445206 507218 475690 507454
rect 475926 507218 506410 507454
rect 506646 507218 537130 507454
rect 537366 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 52250 507134
rect 52486 506898 82970 507134
rect 83206 506898 113690 507134
rect 113926 506898 144410 507134
rect 144646 506898 175130 507134
rect 175366 506898 205850 507134
rect 206086 506898 236570 507134
rect 236806 506898 267290 507134
rect 267526 506898 298010 507134
rect 298246 506898 328730 507134
rect 328966 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 414250 507134
rect 414486 506898 444970 507134
rect 445206 506898 475690 507134
rect 475926 506898 506410 507134
rect 506646 506898 537130 507134
rect 537366 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 67610 475954
rect 67846 475718 98330 475954
rect 98566 475718 129050 475954
rect 129286 475718 159770 475954
rect 160006 475718 190490 475954
rect 190726 475718 221210 475954
rect 221446 475718 251930 475954
rect 252166 475718 282650 475954
rect 282886 475718 313370 475954
rect 313606 475718 344090 475954
rect 344326 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 429610 475954
rect 429846 475718 460330 475954
rect 460566 475718 491050 475954
rect 491286 475718 521770 475954
rect 522006 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 67610 475634
rect 67846 475398 98330 475634
rect 98566 475398 129050 475634
rect 129286 475398 159770 475634
rect 160006 475398 190490 475634
rect 190726 475398 221210 475634
rect 221446 475398 251930 475634
rect 252166 475398 282650 475634
rect 282886 475398 313370 475634
rect 313606 475398 344090 475634
rect 344326 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 429610 475634
rect 429846 475398 460330 475634
rect 460566 475398 491050 475634
rect 491286 475398 521770 475634
rect 522006 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 52250 471454
rect 52486 471218 82970 471454
rect 83206 471218 113690 471454
rect 113926 471218 144410 471454
rect 144646 471218 175130 471454
rect 175366 471218 205850 471454
rect 206086 471218 236570 471454
rect 236806 471218 267290 471454
rect 267526 471218 298010 471454
rect 298246 471218 328730 471454
rect 328966 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 414250 471454
rect 414486 471218 444970 471454
rect 445206 471218 475690 471454
rect 475926 471218 506410 471454
rect 506646 471218 537130 471454
rect 537366 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 52250 471134
rect 52486 470898 82970 471134
rect 83206 470898 113690 471134
rect 113926 470898 144410 471134
rect 144646 470898 175130 471134
rect 175366 470898 205850 471134
rect 206086 470898 236570 471134
rect 236806 470898 267290 471134
rect 267526 470898 298010 471134
rect 298246 470898 328730 471134
rect 328966 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 414250 471134
rect 414486 470898 444970 471134
rect 445206 470898 475690 471134
rect 475926 470898 506410 471134
rect 506646 470898 537130 471134
rect 537366 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 67610 439954
rect 67846 439718 98330 439954
rect 98566 439718 129050 439954
rect 129286 439718 159770 439954
rect 160006 439718 190490 439954
rect 190726 439718 221210 439954
rect 221446 439718 251930 439954
rect 252166 439718 282650 439954
rect 282886 439718 313370 439954
rect 313606 439718 344090 439954
rect 344326 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 429610 439954
rect 429846 439718 460330 439954
rect 460566 439718 491050 439954
rect 491286 439718 521770 439954
rect 522006 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 67610 439634
rect 67846 439398 98330 439634
rect 98566 439398 129050 439634
rect 129286 439398 159770 439634
rect 160006 439398 190490 439634
rect 190726 439398 221210 439634
rect 221446 439398 251930 439634
rect 252166 439398 282650 439634
rect 282886 439398 313370 439634
rect 313606 439398 344090 439634
rect 344326 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 429610 439634
rect 429846 439398 460330 439634
rect 460566 439398 491050 439634
rect 491286 439398 521770 439634
rect 522006 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 52250 435454
rect 52486 435218 82970 435454
rect 83206 435218 113690 435454
rect 113926 435218 144410 435454
rect 144646 435218 175130 435454
rect 175366 435218 205850 435454
rect 206086 435218 236570 435454
rect 236806 435218 267290 435454
rect 267526 435218 298010 435454
rect 298246 435218 328730 435454
rect 328966 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 414250 435454
rect 414486 435218 444970 435454
rect 445206 435218 475690 435454
rect 475926 435218 506410 435454
rect 506646 435218 537130 435454
rect 537366 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 52250 435134
rect 52486 434898 82970 435134
rect 83206 434898 113690 435134
rect 113926 434898 144410 435134
rect 144646 434898 175130 435134
rect 175366 434898 205850 435134
rect 206086 434898 236570 435134
rect 236806 434898 267290 435134
rect 267526 434898 298010 435134
rect 298246 434898 328730 435134
rect 328966 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 414250 435134
rect 414486 434898 444970 435134
rect 445206 434898 475690 435134
rect 475926 434898 506410 435134
rect 506646 434898 537130 435134
rect 537366 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 67610 403954
rect 67846 403718 98330 403954
rect 98566 403718 129050 403954
rect 129286 403718 159770 403954
rect 160006 403718 190490 403954
rect 190726 403718 221210 403954
rect 221446 403718 251930 403954
rect 252166 403718 282650 403954
rect 282886 403718 313370 403954
rect 313606 403718 344090 403954
rect 344326 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 429610 403954
rect 429846 403718 460330 403954
rect 460566 403718 491050 403954
rect 491286 403718 521770 403954
rect 522006 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 67610 403634
rect 67846 403398 98330 403634
rect 98566 403398 129050 403634
rect 129286 403398 159770 403634
rect 160006 403398 190490 403634
rect 190726 403398 221210 403634
rect 221446 403398 251930 403634
rect 252166 403398 282650 403634
rect 282886 403398 313370 403634
rect 313606 403398 344090 403634
rect 344326 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 429610 403634
rect 429846 403398 460330 403634
rect 460566 403398 491050 403634
rect 491286 403398 521770 403634
rect 522006 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 52250 399454
rect 52486 399218 82970 399454
rect 83206 399218 113690 399454
rect 113926 399218 144410 399454
rect 144646 399218 175130 399454
rect 175366 399218 205850 399454
rect 206086 399218 236570 399454
rect 236806 399218 267290 399454
rect 267526 399218 298010 399454
rect 298246 399218 328730 399454
rect 328966 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 414250 399454
rect 414486 399218 444970 399454
rect 445206 399218 475690 399454
rect 475926 399218 506410 399454
rect 506646 399218 537130 399454
rect 537366 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 52250 399134
rect 52486 398898 82970 399134
rect 83206 398898 113690 399134
rect 113926 398898 144410 399134
rect 144646 398898 175130 399134
rect 175366 398898 205850 399134
rect 206086 398898 236570 399134
rect 236806 398898 267290 399134
rect 267526 398898 298010 399134
rect 298246 398898 328730 399134
rect 328966 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 414250 399134
rect 414486 398898 444970 399134
rect 445206 398898 475690 399134
rect 475926 398898 506410 399134
rect 506646 398898 537130 399134
rect 537366 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 67610 367954
rect 67846 367718 98330 367954
rect 98566 367718 129050 367954
rect 129286 367718 159770 367954
rect 160006 367718 190490 367954
rect 190726 367718 221210 367954
rect 221446 367718 251930 367954
rect 252166 367718 282650 367954
rect 282886 367718 313370 367954
rect 313606 367718 344090 367954
rect 344326 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 429610 367954
rect 429846 367718 460330 367954
rect 460566 367718 491050 367954
rect 491286 367718 521770 367954
rect 522006 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 67610 367634
rect 67846 367398 98330 367634
rect 98566 367398 129050 367634
rect 129286 367398 159770 367634
rect 160006 367398 190490 367634
rect 190726 367398 221210 367634
rect 221446 367398 251930 367634
rect 252166 367398 282650 367634
rect 282886 367398 313370 367634
rect 313606 367398 344090 367634
rect 344326 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 429610 367634
rect 429846 367398 460330 367634
rect 460566 367398 491050 367634
rect 491286 367398 521770 367634
rect 522006 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 52250 363454
rect 52486 363218 82970 363454
rect 83206 363218 113690 363454
rect 113926 363218 144410 363454
rect 144646 363218 175130 363454
rect 175366 363218 205850 363454
rect 206086 363218 236570 363454
rect 236806 363218 267290 363454
rect 267526 363218 298010 363454
rect 298246 363218 328730 363454
rect 328966 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 414250 363454
rect 414486 363218 444970 363454
rect 445206 363218 475690 363454
rect 475926 363218 506410 363454
rect 506646 363218 537130 363454
rect 537366 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 52250 363134
rect 52486 362898 82970 363134
rect 83206 362898 113690 363134
rect 113926 362898 144410 363134
rect 144646 362898 175130 363134
rect 175366 362898 205850 363134
rect 206086 362898 236570 363134
rect 236806 362898 267290 363134
rect 267526 362898 298010 363134
rect 298246 362898 328730 363134
rect 328966 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 414250 363134
rect 414486 362898 444970 363134
rect 445206 362898 475690 363134
rect 475926 362898 506410 363134
rect 506646 362898 537130 363134
rect 537366 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 67610 331954
rect 67846 331718 98330 331954
rect 98566 331718 129050 331954
rect 129286 331718 159770 331954
rect 160006 331718 190490 331954
rect 190726 331718 221210 331954
rect 221446 331718 251930 331954
rect 252166 331718 282650 331954
rect 282886 331718 313370 331954
rect 313606 331718 344090 331954
rect 344326 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 429610 331954
rect 429846 331718 460330 331954
rect 460566 331718 491050 331954
rect 491286 331718 521770 331954
rect 522006 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 67610 331634
rect 67846 331398 98330 331634
rect 98566 331398 129050 331634
rect 129286 331398 159770 331634
rect 160006 331398 190490 331634
rect 190726 331398 221210 331634
rect 221446 331398 251930 331634
rect 252166 331398 282650 331634
rect 282886 331398 313370 331634
rect 313606 331398 344090 331634
rect 344326 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 429610 331634
rect 429846 331398 460330 331634
rect 460566 331398 491050 331634
rect 491286 331398 521770 331634
rect 522006 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 52250 327454
rect 52486 327218 82970 327454
rect 83206 327218 113690 327454
rect 113926 327218 144410 327454
rect 144646 327218 175130 327454
rect 175366 327218 205850 327454
rect 206086 327218 236570 327454
rect 236806 327218 267290 327454
rect 267526 327218 298010 327454
rect 298246 327218 328730 327454
rect 328966 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 414250 327454
rect 414486 327218 444970 327454
rect 445206 327218 475690 327454
rect 475926 327218 506410 327454
rect 506646 327218 537130 327454
rect 537366 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 52250 327134
rect 52486 326898 82970 327134
rect 83206 326898 113690 327134
rect 113926 326898 144410 327134
rect 144646 326898 175130 327134
rect 175366 326898 205850 327134
rect 206086 326898 236570 327134
rect 236806 326898 267290 327134
rect 267526 326898 298010 327134
rect 298246 326898 328730 327134
rect 328966 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 414250 327134
rect 414486 326898 444970 327134
rect 445206 326898 475690 327134
rect 475926 326898 506410 327134
rect 506646 326898 537130 327134
rect 537366 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 67610 295954
rect 67846 295718 98330 295954
rect 98566 295718 129050 295954
rect 129286 295718 159770 295954
rect 160006 295718 190490 295954
rect 190726 295718 221210 295954
rect 221446 295718 251930 295954
rect 252166 295718 282650 295954
rect 282886 295718 313370 295954
rect 313606 295718 344090 295954
rect 344326 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 429610 295954
rect 429846 295718 460330 295954
rect 460566 295718 491050 295954
rect 491286 295718 521770 295954
rect 522006 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 67610 295634
rect 67846 295398 98330 295634
rect 98566 295398 129050 295634
rect 129286 295398 159770 295634
rect 160006 295398 190490 295634
rect 190726 295398 221210 295634
rect 221446 295398 251930 295634
rect 252166 295398 282650 295634
rect 282886 295398 313370 295634
rect 313606 295398 344090 295634
rect 344326 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 429610 295634
rect 429846 295398 460330 295634
rect 460566 295398 491050 295634
rect 491286 295398 521770 295634
rect 522006 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 52250 291454
rect 52486 291218 82970 291454
rect 83206 291218 113690 291454
rect 113926 291218 144410 291454
rect 144646 291218 175130 291454
rect 175366 291218 205850 291454
rect 206086 291218 236570 291454
rect 236806 291218 267290 291454
rect 267526 291218 298010 291454
rect 298246 291218 328730 291454
rect 328966 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 414250 291454
rect 414486 291218 444970 291454
rect 445206 291218 475690 291454
rect 475926 291218 506410 291454
rect 506646 291218 537130 291454
rect 537366 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 52250 291134
rect 52486 290898 82970 291134
rect 83206 290898 113690 291134
rect 113926 290898 144410 291134
rect 144646 290898 175130 291134
rect 175366 290898 205850 291134
rect 206086 290898 236570 291134
rect 236806 290898 267290 291134
rect 267526 290898 298010 291134
rect 298246 290898 328730 291134
rect 328966 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 414250 291134
rect 414486 290898 444970 291134
rect 445206 290898 475690 291134
rect 475926 290898 506410 291134
rect 506646 290898 537130 291134
rect 537366 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 67610 259954
rect 67846 259718 98330 259954
rect 98566 259718 129050 259954
rect 129286 259718 159770 259954
rect 160006 259718 190490 259954
rect 190726 259718 221210 259954
rect 221446 259718 251930 259954
rect 252166 259718 282650 259954
rect 282886 259718 313370 259954
rect 313606 259718 344090 259954
rect 344326 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 429610 259954
rect 429846 259718 460330 259954
rect 460566 259718 491050 259954
rect 491286 259718 521770 259954
rect 522006 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 67610 259634
rect 67846 259398 98330 259634
rect 98566 259398 129050 259634
rect 129286 259398 159770 259634
rect 160006 259398 190490 259634
rect 190726 259398 221210 259634
rect 221446 259398 251930 259634
rect 252166 259398 282650 259634
rect 282886 259398 313370 259634
rect 313606 259398 344090 259634
rect 344326 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 429610 259634
rect 429846 259398 460330 259634
rect 460566 259398 491050 259634
rect 491286 259398 521770 259634
rect 522006 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 52250 255454
rect 52486 255218 82970 255454
rect 83206 255218 113690 255454
rect 113926 255218 144410 255454
rect 144646 255218 175130 255454
rect 175366 255218 205850 255454
rect 206086 255218 236570 255454
rect 236806 255218 267290 255454
rect 267526 255218 298010 255454
rect 298246 255218 328730 255454
rect 328966 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 414250 255454
rect 414486 255218 444970 255454
rect 445206 255218 475690 255454
rect 475926 255218 506410 255454
rect 506646 255218 537130 255454
rect 537366 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 52250 255134
rect 52486 254898 82970 255134
rect 83206 254898 113690 255134
rect 113926 254898 144410 255134
rect 144646 254898 175130 255134
rect 175366 254898 205850 255134
rect 206086 254898 236570 255134
rect 236806 254898 267290 255134
rect 267526 254898 298010 255134
rect 298246 254898 328730 255134
rect 328966 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 414250 255134
rect 414486 254898 444970 255134
rect 445206 254898 475690 255134
rect 475926 254898 506410 255134
rect 506646 254898 537130 255134
rect 537366 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 67610 223954
rect 67846 223718 98330 223954
rect 98566 223718 129050 223954
rect 129286 223718 159770 223954
rect 160006 223718 190490 223954
rect 190726 223718 221210 223954
rect 221446 223718 251930 223954
rect 252166 223718 282650 223954
rect 282886 223718 313370 223954
rect 313606 223718 344090 223954
rect 344326 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 67610 223634
rect 67846 223398 98330 223634
rect 98566 223398 129050 223634
rect 129286 223398 159770 223634
rect 160006 223398 190490 223634
rect 190726 223398 221210 223634
rect 221446 223398 251930 223634
rect 252166 223398 282650 223634
rect 282886 223398 313370 223634
rect 313606 223398 344090 223634
rect 344326 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 52250 219454
rect 52486 219218 82970 219454
rect 83206 219218 113690 219454
rect 113926 219218 144410 219454
rect 144646 219218 175130 219454
rect 175366 219218 205850 219454
rect 206086 219218 236570 219454
rect 236806 219218 267290 219454
rect 267526 219218 298010 219454
rect 298246 219218 328730 219454
rect 328966 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 52250 219134
rect 52486 218898 82970 219134
rect 83206 218898 113690 219134
rect 113926 218898 144410 219134
rect 144646 218898 175130 219134
rect 175366 218898 205850 219134
rect 206086 218898 236570 219134
rect 236806 218898 267290 219134
rect 267526 218898 298010 219134
rect 298246 218898 328730 219134
rect 328966 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 248570 147454
rect 248806 147218 279290 147454
rect 279526 147218 310010 147454
rect 310246 147218 340730 147454
rect 340966 147218 371450 147454
rect 371686 147218 402170 147454
rect 402406 147218 432890 147454
rect 433126 147218 463610 147454
rect 463846 147218 494330 147454
rect 494566 147218 525050 147454
rect 525286 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 248570 147134
rect 248806 146898 279290 147134
rect 279526 146898 310010 147134
rect 310246 146898 340730 147134
rect 340966 146898 371450 147134
rect 371686 146898 402170 147134
rect 402406 146898 432890 147134
rect 433126 146898 463610 147134
rect 463846 146898 494330 147134
rect 494566 146898 525050 147134
rect 525286 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 79610 115954
rect 79846 115718 110330 115954
rect 110566 115718 141050 115954
rect 141286 115718 171770 115954
rect 172006 115718 202490 115954
rect 202726 115718 233210 115954
rect 233446 115718 263930 115954
rect 264166 115718 294650 115954
rect 294886 115718 325370 115954
rect 325606 115718 356090 115954
rect 356326 115718 386810 115954
rect 387046 115718 417530 115954
rect 417766 115718 448250 115954
rect 448486 115718 478970 115954
rect 479206 115718 509690 115954
rect 509926 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 79610 115634
rect 79846 115398 110330 115634
rect 110566 115398 141050 115634
rect 141286 115398 171770 115634
rect 172006 115398 202490 115634
rect 202726 115398 233210 115634
rect 233446 115398 263930 115634
rect 264166 115398 294650 115634
rect 294886 115398 325370 115634
rect 325606 115398 356090 115634
rect 356326 115398 386810 115634
rect 387046 115398 417530 115634
rect 417766 115398 448250 115634
rect 448486 115398 478970 115634
rect 479206 115398 509690 115634
rect 509926 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 248570 111454
rect 248806 111218 279290 111454
rect 279526 111218 310010 111454
rect 310246 111218 340730 111454
rect 340966 111218 371450 111454
rect 371686 111218 402170 111454
rect 402406 111218 432890 111454
rect 433126 111218 463610 111454
rect 463846 111218 494330 111454
rect 494566 111218 525050 111454
rect 525286 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 248570 111134
rect 248806 110898 279290 111134
rect 279526 110898 310010 111134
rect 310246 110898 340730 111134
rect 340966 110898 371450 111134
rect 371686 110898 402170 111134
rect 402406 110898 432890 111134
rect 433126 110898 463610 111134
rect 463846 110898 494330 111134
rect 494566 110898 525050 111134
rect 525286 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 79610 79954
rect 79846 79718 110330 79954
rect 110566 79718 141050 79954
rect 141286 79718 171770 79954
rect 172006 79718 202490 79954
rect 202726 79718 233210 79954
rect 233446 79718 263930 79954
rect 264166 79718 294650 79954
rect 294886 79718 325370 79954
rect 325606 79718 356090 79954
rect 356326 79718 386810 79954
rect 387046 79718 417530 79954
rect 417766 79718 448250 79954
rect 448486 79718 478970 79954
rect 479206 79718 509690 79954
rect 509926 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 79610 79634
rect 79846 79398 110330 79634
rect 110566 79398 141050 79634
rect 141286 79398 171770 79634
rect 172006 79398 202490 79634
rect 202726 79398 233210 79634
rect 233446 79398 263930 79634
rect 264166 79398 294650 79634
rect 294886 79398 325370 79634
rect 325606 79398 356090 79634
rect 356326 79398 386810 79634
rect 387046 79398 417530 79634
rect 417766 79398 448250 79634
rect 448486 79398 478970 79634
rect 479206 79398 509690 79634
rect 509926 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 248570 75454
rect 248806 75218 279290 75454
rect 279526 75218 310010 75454
rect 310246 75218 340730 75454
rect 340966 75218 371450 75454
rect 371686 75218 402170 75454
rect 402406 75218 432890 75454
rect 433126 75218 463610 75454
rect 463846 75218 494330 75454
rect 494566 75218 525050 75454
rect 525286 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 248570 75134
rect 248806 74898 279290 75134
rect 279526 74898 310010 75134
rect 310246 74898 340730 75134
rect 340966 74898 371450 75134
rect 371686 74898 402170 75134
rect 402406 74898 432890 75134
rect 433126 74898 463610 75134
rect 463846 74898 494330 75134
rect 494566 74898 525050 75134
rect 525286 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 79610 43954
rect 79846 43718 110330 43954
rect 110566 43718 141050 43954
rect 141286 43718 171770 43954
rect 172006 43718 202490 43954
rect 202726 43718 233210 43954
rect 233446 43718 263930 43954
rect 264166 43718 294650 43954
rect 294886 43718 325370 43954
rect 325606 43718 356090 43954
rect 356326 43718 386810 43954
rect 387046 43718 417530 43954
rect 417766 43718 448250 43954
rect 448486 43718 478970 43954
rect 479206 43718 509690 43954
rect 509926 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 79610 43634
rect 79846 43398 110330 43634
rect 110566 43398 141050 43634
rect 141286 43398 171770 43634
rect 172006 43398 202490 43634
rect 202726 43398 233210 43634
rect 233446 43398 263930 43634
rect 264166 43398 294650 43634
rect 294886 43398 325370 43634
rect 325606 43398 356090 43634
rect 356326 43398 386810 43634
rect 387046 43398 417530 43634
rect 417766 43398 448250 43634
rect 448486 43398 478970 43634
rect 479206 43398 509690 43634
rect 509926 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 64250 39454
rect 64486 39218 94970 39454
rect 95206 39218 125690 39454
rect 125926 39218 156410 39454
rect 156646 39218 187130 39454
rect 187366 39218 217850 39454
rect 218086 39218 248570 39454
rect 248806 39218 279290 39454
rect 279526 39218 310010 39454
rect 310246 39218 340730 39454
rect 340966 39218 371450 39454
rect 371686 39218 402170 39454
rect 402406 39218 432890 39454
rect 433126 39218 463610 39454
rect 463846 39218 494330 39454
rect 494566 39218 525050 39454
rect 525286 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 64250 39134
rect 64486 38898 94970 39134
rect 95206 38898 125690 39134
rect 125926 38898 156410 39134
rect 156646 38898 187130 39134
rect 187366 38898 217850 39134
rect 218086 38898 248570 39134
rect 248806 38898 279290 39134
rect 279526 38898 310010 39134
rect 310246 38898 340730 39134
rect 340966 38898 371450 39134
rect 371686 38898 402170 39134
rect 402406 38898 432890 39134
rect 433126 38898 463610 39134
rect 463846 38898 494330 39134
rect 494566 38898 525050 39134
rect 525286 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use axi_node_intf_wrap  axi_interconnect_i
timestamp 0
transform 1 0 60000 0 1 30000
box 0 0 480000 120000
use mba_core_region  core_region_i
timestamp 0
transform 1 0 48000 0 1 200000
box 0 0 300000 360000
use sky130_sram_2kbyte_1rw1r_32x512_8  data_ram
timestamp 0
transform 1 0 206000 0 1 592000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_ram
timestamp 0
transform 1 0 34000 0 1 592000
box 0 0 136620 83308
use peripherals  peripherals_i
timestamp 0
transform 1 0 410000 0 1 240000
box 0 0 140000 440000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 590000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 677308 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 677308 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 677308 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 677308 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 562000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 677308 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 677308 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 677308 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 677308 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 152000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 152000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 152000 434414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 682000 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 152000 470414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 682000 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 152000 506414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 682000 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 28000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 152000 542414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 682000 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 677308 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 152000 83414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 677308 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 152000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 677308 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 152000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 677308 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 152000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 562000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 152000 227414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 677308 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 152000 263414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 677308 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 152000 299414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 677308 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 152000 335414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 677308 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 152000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 152000 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 152000 443414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 682000 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 152000 479414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 682000 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 28000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 152000 515414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 682000 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 682000 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 198000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 562000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 152000 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 152000 416414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 152000 452414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 152000 488414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 28000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 152000 524414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 677308 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 677308 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 677308 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 562000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 677308 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 677308 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 677308 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 677308 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 152000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 152000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 152000 425414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 152000 461414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 152000 497414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 152000 533414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 562000 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 152000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 152000 420914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 152000 456914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 152000 492914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 28000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 152000 528914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 590000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 677308 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 677308 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 677308 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 677308 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 562000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 677308 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 677308 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 677308 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 677308 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 152000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 152000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 152000 429914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 682000 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 152000 465914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 682000 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 152000 501914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 682000 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 152000 537914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 682000 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 590000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 677308 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 677308 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 677308 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 677308 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 562000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 677308 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 677308 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 677308 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 677308 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 152000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 152000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 152000 438914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 682000 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 152000 474914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 682000 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 28000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 152000 510914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 682000 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 682000 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 677308 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 152000 87914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 677308 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 152000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 677308 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 152000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 677308 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 152000 195914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 562000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 152000 231914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 677308 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 152000 267914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 677308 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 152000 303914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 677308 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 152000 339914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 677308 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 152000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 152000 411914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 682000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 152000 447914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 682000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 152000 483914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 682000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 28000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 152000 519914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 682000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
