magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< dnwell >>
rect -122 84 1072 7440
<< nwell >>
rect -202 7150 1152 7520
rect -202 168 168 7150
rect 782 168 1152 7150
rect -202 0 1152 168
<< pwell >>
rect 228 228 722 7090
<< mvnmos >>
rect 415 5956 535 6956
rect 415 4835 535 5835
rect 415 3714 535 4714
rect 415 2604 535 3604
rect 415 1483 535 2483
rect 415 362 535 1362
<< mvndiff >>
rect 362 6944 415 6956
rect 362 6910 370 6944
rect 404 6910 415 6944
rect 362 6876 415 6910
rect 362 6842 370 6876
rect 404 6842 415 6876
rect 362 6808 415 6842
rect 362 6774 370 6808
rect 404 6774 415 6808
rect 362 6740 415 6774
rect 362 6706 370 6740
rect 404 6706 415 6740
rect 362 6672 415 6706
rect 362 6638 370 6672
rect 404 6638 415 6672
rect 362 6604 415 6638
rect 362 6570 370 6604
rect 404 6570 415 6604
rect 362 6536 415 6570
rect 362 6502 370 6536
rect 404 6502 415 6536
rect 362 6468 415 6502
rect 362 6434 370 6468
rect 404 6434 415 6468
rect 362 6400 415 6434
rect 362 6366 370 6400
rect 404 6366 415 6400
rect 362 6332 415 6366
rect 362 6298 370 6332
rect 404 6298 415 6332
rect 362 6264 415 6298
rect 362 6230 370 6264
rect 404 6230 415 6264
rect 362 6196 415 6230
rect 362 6162 370 6196
rect 404 6162 415 6196
rect 362 6128 415 6162
rect 362 6094 370 6128
rect 404 6094 415 6128
rect 362 6060 415 6094
rect 362 6026 370 6060
rect 404 6026 415 6060
rect 362 5956 415 6026
rect 535 6944 588 6956
rect 535 6910 546 6944
rect 580 6910 588 6944
rect 535 6876 588 6910
rect 535 6842 546 6876
rect 580 6842 588 6876
rect 535 6808 588 6842
rect 535 6774 546 6808
rect 580 6774 588 6808
rect 535 6740 588 6774
rect 535 6706 546 6740
rect 580 6706 588 6740
rect 535 6672 588 6706
rect 535 6638 546 6672
rect 580 6638 588 6672
rect 535 6604 588 6638
rect 535 6570 546 6604
rect 580 6570 588 6604
rect 535 6536 588 6570
rect 535 6502 546 6536
rect 580 6502 588 6536
rect 535 6468 588 6502
rect 535 6434 546 6468
rect 580 6434 588 6468
rect 535 6400 588 6434
rect 535 6366 546 6400
rect 580 6366 588 6400
rect 535 6332 588 6366
rect 535 6298 546 6332
rect 580 6298 588 6332
rect 535 6264 588 6298
rect 535 6230 546 6264
rect 580 6230 588 6264
rect 535 6196 588 6230
rect 535 6162 546 6196
rect 580 6162 588 6196
rect 535 6128 588 6162
rect 535 6094 546 6128
rect 580 6094 588 6128
rect 535 6060 588 6094
rect 535 6026 546 6060
rect 580 6026 588 6060
rect 535 5956 588 6026
rect 362 5823 415 5835
rect 362 5789 370 5823
rect 404 5789 415 5823
rect 362 5755 415 5789
rect 362 5721 370 5755
rect 404 5721 415 5755
rect 362 5687 415 5721
rect 362 5653 370 5687
rect 404 5653 415 5687
rect 362 5619 415 5653
rect 362 5585 370 5619
rect 404 5585 415 5619
rect 362 5551 415 5585
rect 362 5517 370 5551
rect 404 5517 415 5551
rect 362 5483 415 5517
rect 362 5449 370 5483
rect 404 5449 415 5483
rect 362 5415 415 5449
rect 362 5381 370 5415
rect 404 5381 415 5415
rect 362 5347 415 5381
rect 362 5313 370 5347
rect 404 5313 415 5347
rect 362 5279 415 5313
rect 362 5245 370 5279
rect 404 5245 415 5279
rect 362 5211 415 5245
rect 362 5177 370 5211
rect 404 5177 415 5211
rect 362 5143 415 5177
rect 362 5109 370 5143
rect 404 5109 415 5143
rect 362 5075 415 5109
rect 362 5041 370 5075
rect 404 5041 415 5075
rect 362 5007 415 5041
rect 362 4973 370 5007
rect 404 4973 415 5007
rect 362 4939 415 4973
rect 362 4905 370 4939
rect 404 4905 415 4939
rect 362 4835 415 4905
rect 535 5823 588 5835
rect 535 5789 546 5823
rect 580 5789 588 5823
rect 535 5755 588 5789
rect 535 5721 546 5755
rect 580 5721 588 5755
rect 535 5687 588 5721
rect 535 5653 546 5687
rect 580 5653 588 5687
rect 535 5619 588 5653
rect 535 5585 546 5619
rect 580 5585 588 5619
rect 535 5551 588 5585
rect 535 5517 546 5551
rect 580 5517 588 5551
rect 535 5483 588 5517
rect 535 5449 546 5483
rect 580 5449 588 5483
rect 535 5415 588 5449
rect 535 5381 546 5415
rect 580 5381 588 5415
rect 535 5347 588 5381
rect 535 5313 546 5347
rect 580 5313 588 5347
rect 535 5279 588 5313
rect 535 5245 546 5279
rect 580 5245 588 5279
rect 535 5211 588 5245
rect 535 5177 546 5211
rect 580 5177 588 5211
rect 535 5143 588 5177
rect 535 5109 546 5143
rect 580 5109 588 5143
rect 535 5075 588 5109
rect 535 5041 546 5075
rect 580 5041 588 5075
rect 535 5007 588 5041
rect 535 4973 546 5007
rect 580 4973 588 5007
rect 535 4939 588 4973
rect 535 4905 546 4939
rect 580 4905 588 4939
rect 535 4835 588 4905
rect 362 4702 415 4714
rect 362 4668 370 4702
rect 404 4668 415 4702
rect 362 4634 415 4668
rect 362 4600 370 4634
rect 404 4600 415 4634
rect 362 4566 415 4600
rect 362 4532 370 4566
rect 404 4532 415 4566
rect 362 4498 415 4532
rect 362 4464 370 4498
rect 404 4464 415 4498
rect 362 4430 415 4464
rect 362 4396 370 4430
rect 404 4396 415 4430
rect 362 4362 415 4396
rect 362 4328 370 4362
rect 404 4328 415 4362
rect 362 4294 415 4328
rect 362 4260 370 4294
rect 404 4260 415 4294
rect 362 4226 415 4260
rect 362 4192 370 4226
rect 404 4192 415 4226
rect 362 4158 415 4192
rect 362 4124 370 4158
rect 404 4124 415 4158
rect 362 4090 415 4124
rect 362 4056 370 4090
rect 404 4056 415 4090
rect 362 4022 415 4056
rect 362 3988 370 4022
rect 404 3988 415 4022
rect 362 3954 415 3988
rect 362 3920 370 3954
rect 404 3920 415 3954
rect 362 3886 415 3920
rect 362 3852 370 3886
rect 404 3852 415 3886
rect 362 3818 415 3852
rect 362 3784 370 3818
rect 404 3784 415 3818
rect 362 3714 415 3784
rect 535 4702 588 4714
rect 535 4668 546 4702
rect 580 4668 588 4702
rect 535 4634 588 4668
rect 535 4600 546 4634
rect 580 4600 588 4634
rect 535 4566 588 4600
rect 535 4532 546 4566
rect 580 4532 588 4566
rect 535 4498 588 4532
rect 535 4464 546 4498
rect 580 4464 588 4498
rect 535 4430 588 4464
rect 535 4396 546 4430
rect 580 4396 588 4430
rect 535 4362 588 4396
rect 535 4328 546 4362
rect 580 4328 588 4362
rect 535 4294 588 4328
rect 535 4260 546 4294
rect 580 4260 588 4294
rect 535 4226 588 4260
rect 535 4192 546 4226
rect 580 4192 588 4226
rect 535 4158 588 4192
rect 535 4124 546 4158
rect 580 4124 588 4158
rect 535 4090 588 4124
rect 535 4056 546 4090
rect 580 4056 588 4090
rect 535 4022 588 4056
rect 535 3988 546 4022
rect 580 3988 588 4022
rect 535 3954 588 3988
rect 535 3920 546 3954
rect 580 3920 588 3954
rect 535 3886 588 3920
rect 535 3852 546 3886
rect 580 3852 588 3886
rect 535 3818 588 3852
rect 535 3784 546 3818
rect 580 3784 588 3818
rect 535 3714 588 3784
rect 362 3534 415 3604
rect 362 3500 370 3534
rect 404 3500 415 3534
rect 362 3466 415 3500
rect 362 3432 370 3466
rect 404 3432 415 3466
rect 362 3398 415 3432
rect 362 3364 370 3398
rect 404 3364 415 3398
rect 362 3330 415 3364
rect 362 3296 370 3330
rect 404 3296 415 3330
rect 362 3262 415 3296
rect 362 3228 370 3262
rect 404 3228 415 3262
rect 362 3194 415 3228
rect 362 3160 370 3194
rect 404 3160 415 3194
rect 362 3126 415 3160
rect 362 3092 370 3126
rect 404 3092 415 3126
rect 362 3058 415 3092
rect 362 3024 370 3058
rect 404 3024 415 3058
rect 362 2990 415 3024
rect 362 2956 370 2990
rect 404 2956 415 2990
rect 362 2922 415 2956
rect 362 2888 370 2922
rect 404 2888 415 2922
rect 362 2854 415 2888
rect 362 2820 370 2854
rect 404 2820 415 2854
rect 362 2786 415 2820
rect 362 2752 370 2786
rect 404 2752 415 2786
rect 362 2718 415 2752
rect 362 2684 370 2718
rect 404 2684 415 2718
rect 362 2650 415 2684
rect 362 2616 370 2650
rect 404 2616 415 2650
rect 362 2604 415 2616
rect 535 3534 588 3604
rect 535 3500 546 3534
rect 580 3500 588 3534
rect 535 3466 588 3500
rect 535 3432 546 3466
rect 580 3432 588 3466
rect 535 3398 588 3432
rect 535 3364 546 3398
rect 580 3364 588 3398
rect 535 3330 588 3364
rect 535 3296 546 3330
rect 580 3296 588 3330
rect 535 3262 588 3296
rect 535 3228 546 3262
rect 580 3228 588 3262
rect 535 3194 588 3228
rect 535 3160 546 3194
rect 580 3160 588 3194
rect 535 3126 588 3160
rect 535 3092 546 3126
rect 580 3092 588 3126
rect 535 3058 588 3092
rect 535 3024 546 3058
rect 580 3024 588 3058
rect 535 2990 588 3024
rect 535 2956 546 2990
rect 580 2956 588 2990
rect 535 2922 588 2956
rect 535 2888 546 2922
rect 580 2888 588 2922
rect 535 2854 588 2888
rect 535 2820 546 2854
rect 580 2820 588 2854
rect 535 2786 588 2820
rect 535 2752 546 2786
rect 580 2752 588 2786
rect 535 2718 588 2752
rect 535 2684 546 2718
rect 580 2684 588 2718
rect 535 2650 588 2684
rect 535 2616 546 2650
rect 580 2616 588 2650
rect 535 2604 588 2616
rect 362 2413 415 2483
rect 362 2379 370 2413
rect 404 2379 415 2413
rect 362 2345 415 2379
rect 362 2311 370 2345
rect 404 2311 415 2345
rect 362 2277 415 2311
rect 362 2243 370 2277
rect 404 2243 415 2277
rect 362 2209 415 2243
rect 362 2175 370 2209
rect 404 2175 415 2209
rect 362 2141 415 2175
rect 362 2107 370 2141
rect 404 2107 415 2141
rect 362 2073 415 2107
rect 362 2039 370 2073
rect 404 2039 415 2073
rect 362 2005 415 2039
rect 362 1971 370 2005
rect 404 1971 415 2005
rect 362 1937 415 1971
rect 362 1903 370 1937
rect 404 1903 415 1937
rect 362 1869 415 1903
rect 362 1835 370 1869
rect 404 1835 415 1869
rect 362 1801 415 1835
rect 362 1767 370 1801
rect 404 1767 415 1801
rect 362 1733 415 1767
rect 362 1699 370 1733
rect 404 1699 415 1733
rect 362 1665 415 1699
rect 362 1631 370 1665
rect 404 1631 415 1665
rect 362 1597 415 1631
rect 362 1563 370 1597
rect 404 1563 415 1597
rect 362 1529 415 1563
rect 362 1495 370 1529
rect 404 1495 415 1529
rect 362 1483 415 1495
rect 535 2413 588 2483
rect 535 2379 546 2413
rect 580 2379 588 2413
rect 535 2345 588 2379
rect 535 2311 546 2345
rect 580 2311 588 2345
rect 535 2277 588 2311
rect 535 2243 546 2277
rect 580 2243 588 2277
rect 535 2209 588 2243
rect 535 2175 546 2209
rect 580 2175 588 2209
rect 535 2141 588 2175
rect 535 2107 546 2141
rect 580 2107 588 2141
rect 535 2073 588 2107
rect 535 2039 546 2073
rect 580 2039 588 2073
rect 535 2005 588 2039
rect 535 1971 546 2005
rect 580 1971 588 2005
rect 535 1937 588 1971
rect 535 1903 546 1937
rect 580 1903 588 1937
rect 535 1869 588 1903
rect 535 1835 546 1869
rect 580 1835 588 1869
rect 535 1801 588 1835
rect 535 1767 546 1801
rect 580 1767 588 1801
rect 535 1733 588 1767
rect 535 1699 546 1733
rect 580 1699 588 1733
rect 535 1665 588 1699
rect 535 1631 546 1665
rect 580 1631 588 1665
rect 535 1597 588 1631
rect 535 1563 546 1597
rect 580 1563 588 1597
rect 535 1529 588 1563
rect 535 1495 546 1529
rect 580 1495 588 1529
rect 535 1483 588 1495
rect 362 1292 415 1362
rect 362 1258 370 1292
rect 404 1258 415 1292
rect 362 1224 415 1258
rect 362 1190 370 1224
rect 404 1190 415 1224
rect 362 1156 415 1190
rect 362 1122 370 1156
rect 404 1122 415 1156
rect 362 1088 415 1122
rect 362 1054 370 1088
rect 404 1054 415 1088
rect 362 1020 415 1054
rect 362 986 370 1020
rect 404 986 415 1020
rect 362 952 415 986
rect 362 918 370 952
rect 404 918 415 952
rect 362 884 415 918
rect 362 850 370 884
rect 404 850 415 884
rect 362 816 415 850
rect 362 782 370 816
rect 404 782 415 816
rect 362 748 415 782
rect 362 714 370 748
rect 404 714 415 748
rect 362 680 415 714
rect 362 646 370 680
rect 404 646 415 680
rect 362 612 415 646
rect 362 578 370 612
rect 404 578 415 612
rect 362 544 415 578
rect 362 510 370 544
rect 404 510 415 544
rect 362 476 415 510
rect 362 442 370 476
rect 404 442 415 476
rect 362 408 415 442
rect 362 374 370 408
rect 404 374 415 408
rect 362 362 415 374
rect 535 1292 588 1362
rect 535 1258 546 1292
rect 580 1258 588 1292
rect 535 1224 588 1258
rect 535 1190 546 1224
rect 580 1190 588 1224
rect 535 1156 588 1190
rect 535 1122 546 1156
rect 580 1122 588 1156
rect 535 1088 588 1122
rect 535 1054 546 1088
rect 580 1054 588 1088
rect 535 1020 588 1054
rect 535 986 546 1020
rect 580 986 588 1020
rect 535 952 588 986
rect 535 918 546 952
rect 580 918 588 952
rect 535 884 588 918
rect 535 850 546 884
rect 580 850 588 884
rect 535 816 588 850
rect 535 782 546 816
rect 580 782 588 816
rect 535 748 588 782
rect 535 714 546 748
rect 580 714 588 748
rect 535 680 588 714
rect 535 646 546 680
rect 580 646 588 680
rect 535 612 588 646
rect 535 578 546 612
rect 580 578 588 612
rect 535 544 588 578
rect 535 510 546 544
rect 580 510 588 544
rect 535 476 588 510
rect 535 442 546 476
rect 580 442 588 476
rect 535 408 588 442
rect 535 374 546 408
rect 580 374 588 408
rect 535 362 588 374
<< mvndiffc >>
rect 370 6910 404 6944
rect 370 6842 404 6876
rect 370 6774 404 6808
rect 370 6706 404 6740
rect 370 6638 404 6672
rect 370 6570 404 6604
rect 370 6502 404 6536
rect 370 6434 404 6468
rect 370 6366 404 6400
rect 370 6298 404 6332
rect 370 6230 404 6264
rect 370 6162 404 6196
rect 370 6094 404 6128
rect 370 6026 404 6060
rect 546 6910 580 6944
rect 546 6842 580 6876
rect 546 6774 580 6808
rect 546 6706 580 6740
rect 546 6638 580 6672
rect 546 6570 580 6604
rect 546 6502 580 6536
rect 546 6434 580 6468
rect 546 6366 580 6400
rect 546 6298 580 6332
rect 546 6230 580 6264
rect 546 6162 580 6196
rect 546 6094 580 6128
rect 546 6026 580 6060
rect 370 5789 404 5823
rect 370 5721 404 5755
rect 370 5653 404 5687
rect 370 5585 404 5619
rect 370 5517 404 5551
rect 370 5449 404 5483
rect 370 5381 404 5415
rect 370 5313 404 5347
rect 370 5245 404 5279
rect 370 5177 404 5211
rect 370 5109 404 5143
rect 370 5041 404 5075
rect 370 4973 404 5007
rect 370 4905 404 4939
rect 546 5789 580 5823
rect 546 5721 580 5755
rect 546 5653 580 5687
rect 546 5585 580 5619
rect 546 5517 580 5551
rect 546 5449 580 5483
rect 546 5381 580 5415
rect 546 5313 580 5347
rect 546 5245 580 5279
rect 546 5177 580 5211
rect 546 5109 580 5143
rect 546 5041 580 5075
rect 546 4973 580 5007
rect 546 4905 580 4939
rect 370 4668 404 4702
rect 370 4600 404 4634
rect 370 4532 404 4566
rect 370 4464 404 4498
rect 370 4396 404 4430
rect 370 4328 404 4362
rect 370 4260 404 4294
rect 370 4192 404 4226
rect 370 4124 404 4158
rect 370 4056 404 4090
rect 370 3988 404 4022
rect 370 3920 404 3954
rect 370 3852 404 3886
rect 370 3784 404 3818
rect 546 4668 580 4702
rect 546 4600 580 4634
rect 546 4532 580 4566
rect 546 4464 580 4498
rect 546 4396 580 4430
rect 546 4328 580 4362
rect 546 4260 580 4294
rect 546 4192 580 4226
rect 546 4124 580 4158
rect 546 4056 580 4090
rect 546 3988 580 4022
rect 546 3920 580 3954
rect 546 3852 580 3886
rect 546 3784 580 3818
rect 370 3500 404 3534
rect 370 3432 404 3466
rect 370 3364 404 3398
rect 370 3296 404 3330
rect 370 3228 404 3262
rect 370 3160 404 3194
rect 370 3092 404 3126
rect 370 3024 404 3058
rect 370 2956 404 2990
rect 370 2888 404 2922
rect 370 2820 404 2854
rect 370 2752 404 2786
rect 370 2684 404 2718
rect 370 2616 404 2650
rect 546 3500 580 3534
rect 546 3432 580 3466
rect 546 3364 580 3398
rect 546 3296 580 3330
rect 546 3228 580 3262
rect 546 3160 580 3194
rect 546 3092 580 3126
rect 546 3024 580 3058
rect 546 2956 580 2990
rect 546 2888 580 2922
rect 546 2820 580 2854
rect 546 2752 580 2786
rect 546 2684 580 2718
rect 546 2616 580 2650
rect 370 2379 404 2413
rect 370 2311 404 2345
rect 370 2243 404 2277
rect 370 2175 404 2209
rect 370 2107 404 2141
rect 370 2039 404 2073
rect 370 1971 404 2005
rect 370 1903 404 1937
rect 370 1835 404 1869
rect 370 1767 404 1801
rect 370 1699 404 1733
rect 370 1631 404 1665
rect 370 1563 404 1597
rect 370 1495 404 1529
rect 546 2379 580 2413
rect 546 2311 580 2345
rect 546 2243 580 2277
rect 546 2175 580 2209
rect 546 2107 580 2141
rect 546 2039 580 2073
rect 546 1971 580 2005
rect 546 1903 580 1937
rect 546 1835 580 1869
rect 546 1767 580 1801
rect 546 1699 580 1733
rect 546 1631 580 1665
rect 546 1563 580 1597
rect 546 1495 580 1529
rect 370 1258 404 1292
rect 370 1190 404 1224
rect 370 1122 404 1156
rect 370 1054 404 1088
rect 370 986 404 1020
rect 370 918 404 952
rect 370 850 404 884
rect 370 782 404 816
rect 370 714 404 748
rect 370 646 404 680
rect 370 578 404 612
rect 370 510 404 544
rect 370 442 404 476
rect 370 374 404 408
rect 546 1258 580 1292
rect 546 1190 580 1224
rect 546 1122 580 1156
rect 546 1054 580 1088
rect 546 986 580 1020
rect 546 918 580 952
rect 546 850 580 884
rect 546 782 580 816
rect 546 714 580 748
rect 546 646 580 680
rect 546 578 580 612
rect 546 510 580 544
rect 546 442 580 476
rect 546 374 580 408
<< mvpsubdiff >>
rect 254 7030 278 7064
rect 312 7030 391 7064
rect 425 7030 525 7064
rect 559 7040 696 7064
rect 559 7030 662 7040
rect 254 6972 288 7030
rect 662 6971 696 7006
rect 254 6904 288 6938
rect 254 6836 288 6870
rect 254 6768 288 6802
rect 254 6700 288 6734
rect 254 6632 288 6666
rect 254 6564 288 6598
rect 254 6496 288 6530
rect 254 6428 288 6462
rect 254 6360 288 6394
rect 254 6292 288 6326
rect 254 6224 288 6258
rect 254 6156 288 6190
rect 254 6088 288 6122
rect 254 6020 288 6054
rect 254 5952 288 5986
rect 662 6902 696 6937
rect 662 6833 696 6868
rect 662 6764 696 6799
rect 662 6695 696 6730
rect 662 6626 696 6661
rect 662 6557 696 6592
rect 662 6488 696 6523
rect 662 6419 696 6454
rect 662 6350 696 6385
rect 662 6281 696 6316
rect 662 6212 696 6247
rect 662 6143 696 6178
rect 662 6074 696 6109
rect 662 6005 696 6040
rect 254 5884 288 5918
rect 254 5816 288 5850
rect 662 5936 696 5971
rect 662 5867 696 5902
rect 254 5748 288 5782
rect 254 5680 288 5714
rect 254 5612 288 5646
rect 254 5544 288 5578
rect 254 5476 288 5510
rect 254 5408 288 5442
rect 254 5340 288 5374
rect 254 5272 288 5306
rect 254 5204 288 5238
rect 254 5136 288 5170
rect 254 5068 288 5102
rect 254 5000 288 5034
rect 254 4932 288 4966
rect 254 4864 288 4898
rect 662 5798 696 5833
rect 662 5729 696 5764
rect 662 5660 696 5695
rect 662 5591 696 5626
rect 662 5522 696 5557
rect 662 5453 696 5488
rect 662 5384 696 5419
rect 662 5315 696 5350
rect 662 5246 696 5281
rect 662 5177 696 5212
rect 662 5108 696 5143
rect 662 5039 696 5074
rect 662 4970 696 5005
rect 662 4901 696 4936
rect 254 4796 288 4830
rect 254 4728 288 4762
rect 662 4832 696 4867
rect 662 4763 696 4798
rect 254 4659 288 4694
rect 254 4590 288 4625
rect 254 4521 288 4556
rect 254 4452 288 4487
rect 254 4383 288 4418
rect 254 4314 288 4349
rect 254 4245 288 4280
rect 254 4176 288 4211
rect 254 4107 288 4142
rect 254 4038 288 4073
rect 254 3969 288 4004
rect 254 3900 288 3935
rect 254 3831 288 3866
rect 254 3762 288 3797
rect 254 3693 288 3728
rect 662 4694 696 4729
rect 662 4625 696 4660
rect 662 4556 696 4591
rect 662 4487 696 4522
rect 662 4418 696 4453
rect 662 4349 696 4384
rect 662 4280 696 4315
rect 662 4211 696 4246
rect 662 4142 696 4177
rect 662 4073 696 4108
rect 662 4004 696 4039
rect 662 3935 696 3970
rect 662 3866 696 3901
rect 662 3797 696 3832
rect 662 3728 696 3763
rect 254 3624 288 3659
rect 662 3659 696 3694
rect 254 3555 288 3590
rect 254 3486 288 3521
rect 254 3417 288 3452
rect 254 3348 288 3383
rect 254 3279 288 3314
rect 254 3210 288 3245
rect 254 3141 288 3176
rect 254 3072 288 3107
rect 254 3003 288 3038
rect 254 2934 288 2969
rect 254 2865 288 2900
rect 254 2796 288 2831
rect 254 2727 288 2762
rect 254 2658 288 2693
rect 254 2589 288 2624
rect 662 3590 696 3625
rect 662 3521 696 3556
rect 662 3452 696 3487
rect 662 3383 696 3418
rect 662 3314 696 3349
rect 662 3245 696 3280
rect 662 3176 696 3211
rect 662 3107 696 3142
rect 662 3038 696 3073
rect 662 2969 696 3004
rect 662 2900 696 2935
rect 662 2831 696 2866
rect 662 2762 696 2797
rect 662 2693 696 2728
rect 662 2624 696 2659
rect 254 2520 288 2555
rect 254 2451 288 2486
rect 662 2556 696 2590
rect 662 2488 696 2522
rect 254 2382 288 2417
rect 254 2313 288 2348
rect 254 2244 288 2279
rect 254 2175 288 2210
rect 254 2106 288 2141
rect 254 2037 288 2072
rect 254 1968 288 2003
rect 254 1899 288 1934
rect 254 1830 288 1865
rect 254 1761 288 1796
rect 254 1692 288 1727
rect 254 1623 288 1658
rect 254 1554 288 1589
rect 254 1485 288 1520
rect 662 2420 696 2454
rect 662 2352 696 2386
rect 662 2284 696 2318
rect 662 2216 696 2250
rect 662 2148 696 2182
rect 662 2080 696 2114
rect 662 2012 696 2046
rect 662 1944 696 1978
rect 662 1876 696 1910
rect 662 1808 696 1842
rect 662 1740 696 1774
rect 662 1672 696 1706
rect 662 1604 696 1638
rect 662 1536 696 1570
rect 254 1416 288 1451
rect 254 1347 288 1382
rect 662 1468 696 1502
rect 662 1400 696 1434
rect 254 1278 288 1313
rect 254 1209 288 1244
rect 254 1140 288 1175
rect 254 1071 288 1106
rect 254 1002 288 1037
rect 254 933 288 968
rect 254 864 288 899
rect 254 795 288 830
rect 254 726 288 761
rect 254 657 288 692
rect 254 588 288 623
rect 254 519 288 554
rect 254 450 288 485
rect 254 381 288 416
rect 662 1332 696 1366
rect 662 1264 696 1298
rect 662 1196 696 1230
rect 662 1128 696 1162
rect 662 1060 696 1094
rect 662 992 696 1026
rect 662 924 696 958
rect 662 856 696 890
rect 662 788 696 822
rect 662 720 696 754
rect 662 652 696 686
rect 662 584 696 618
rect 662 516 696 550
rect 662 448 696 482
rect 662 380 696 414
rect 254 312 288 347
rect 662 288 696 346
rect 288 278 352 288
rect 254 254 352 278
rect 386 254 423 288
rect 457 254 494 288
rect 528 254 566 288
rect 600 254 638 288
rect 672 254 696 288
<< mvnsubdiff >>
rect 68 7217 185 7251
rect 219 7217 261 7251
rect 295 7217 337 7251
rect 371 7217 413 7251
rect 447 7217 488 7251
rect 522 7217 563 7251
rect 597 7217 638 7251
rect 672 7217 713 7251
rect 747 7217 882 7251
rect 68 7101 102 7217
rect 68 7033 102 7067
rect 68 6965 102 6999
rect 68 6897 102 6931
rect 68 6829 102 6863
rect 68 6761 102 6795
rect 68 6693 102 6727
rect 68 6625 102 6659
rect 68 6557 102 6591
rect 68 6489 102 6523
rect 68 6421 102 6455
rect 68 6353 102 6387
rect 68 6285 102 6319
rect 68 6217 102 6251
rect 68 6149 102 6183
rect 68 6081 102 6115
rect 68 6013 102 6047
rect 68 5945 102 5979
rect 68 5877 102 5911
rect 68 5809 102 5843
rect 68 5741 102 5775
rect 68 5673 102 5707
rect 68 5605 102 5639
rect 68 5537 102 5571
rect 68 5469 102 5503
rect 68 5401 102 5435
rect 68 5333 102 5367
rect 68 5265 102 5299
rect 68 5197 102 5231
rect 68 5129 102 5163
rect 68 5061 102 5095
rect 68 4993 102 5027
rect 68 4925 102 4959
rect 68 4857 102 4891
rect 68 4789 102 4823
rect 68 4721 102 4755
rect 68 4653 102 4687
rect 68 4585 102 4619
rect 68 4517 102 4551
rect 68 4449 102 4483
rect 68 4381 102 4415
rect 68 4313 102 4347
rect 68 4245 102 4279
rect 68 4177 102 4211
rect 68 4109 102 4143
rect 68 4041 102 4075
rect 68 3973 102 4007
rect 68 3905 102 3939
rect 68 3837 102 3871
rect 68 3769 102 3803
rect 68 3701 102 3735
rect 68 3633 102 3667
rect 68 3565 102 3599
rect 68 3497 102 3531
rect 68 3429 102 3463
rect 68 3361 102 3395
rect 68 3293 102 3327
rect 68 3225 102 3259
rect 68 3157 102 3191
rect 68 3089 102 3123
rect 68 3021 102 3055
rect 68 2953 102 2987
rect 68 2885 102 2919
rect 68 2817 102 2851
rect 68 2749 102 2783
rect 68 2681 102 2715
rect 68 2613 102 2647
rect 68 2545 102 2579
rect 68 2477 102 2511
rect 68 2409 102 2443
rect 68 2341 102 2375
rect 68 2273 102 2307
rect 68 2205 102 2239
rect 68 2137 102 2171
rect 68 2069 102 2103
rect 68 2001 102 2035
rect 68 1933 102 1967
rect 68 1865 102 1899
rect 68 1797 102 1831
rect 68 1729 102 1763
rect 68 1661 102 1695
rect 68 1593 102 1627
rect 68 1525 102 1559
rect 68 1457 102 1491
rect 68 1389 102 1423
rect 68 1321 102 1355
rect 68 1253 102 1287
rect 68 1185 102 1219
rect 68 1117 102 1151
rect 68 1049 102 1083
rect 68 981 102 1015
rect 68 913 102 947
rect 68 845 102 879
rect 68 777 102 811
rect 68 709 102 743
rect 68 641 102 675
rect 68 573 102 607
rect 68 505 102 539
rect 68 437 102 471
rect 68 369 102 403
rect 68 300 102 335
rect 68 231 102 266
rect 68 101 102 197
rect 848 101 882 7217
rect 68 67 203 101
rect 237 67 273 101
rect 307 67 344 101
rect 378 67 415 101
rect 449 67 486 101
rect 520 67 557 101
rect 591 67 628 101
rect 662 67 699 101
rect 733 67 770 101
rect 804 67 882 101
<< mvpsubdiffcont >>
rect 278 7030 312 7064
rect 391 7030 425 7064
rect 525 7030 559 7064
rect 662 7006 696 7040
rect 254 6938 288 6972
rect 254 6870 288 6904
rect 254 6802 288 6836
rect 254 6734 288 6768
rect 254 6666 288 6700
rect 254 6598 288 6632
rect 254 6530 288 6564
rect 254 6462 288 6496
rect 254 6394 288 6428
rect 254 6326 288 6360
rect 254 6258 288 6292
rect 254 6190 288 6224
rect 254 6122 288 6156
rect 254 6054 288 6088
rect 254 5986 288 6020
rect 662 6937 696 6971
rect 662 6868 696 6902
rect 662 6799 696 6833
rect 662 6730 696 6764
rect 662 6661 696 6695
rect 662 6592 696 6626
rect 662 6523 696 6557
rect 662 6454 696 6488
rect 662 6385 696 6419
rect 662 6316 696 6350
rect 662 6247 696 6281
rect 662 6178 696 6212
rect 662 6109 696 6143
rect 662 6040 696 6074
rect 662 5971 696 6005
rect 254 5918 288 5952
rect 254 5850 288 5884
rect 662 5902 696 5936
rect 254 5782 288 5816
rect 254 5714 288 5748
rect 254 5646 288 5680
rect 254 5578 288 5612
rect 254 5510 288 5544
rect 254 5442 288 5476
rect 254 5374 288 5408
rect 254 5306 288 5340
rect 254 5238 288 5272
rect 254 5170 288 5204
rect 254 5102 288 5136
rect 254 5034 288 5068
rect 254 4966 288 5000
rect 254 4898 288 4932
rect 254 4830 288 4864
rect 662 5833 696 5867
rect 662 5764 696 5798
rect 662 5695 696 5729
rect 662 5626 696 5660
rect 662 5557 696 5591
rect 662 5488 696 5522
rect 662 5419 696 5453
rect 662 5350 696 5384
rect 662 5281 696 5315
rect 662 5212 696 5246
rect 662 5143 696 5177
rect 662 5074 696 5108
rect 662 5005 696 5039
rect 662 4936 696 4970
rect 662 4867 696 4901
rect 254 4762 288 4796
rect 254 4694 288 4728
rect 662 4798 696 4832
rect 662 4729 696 4763
rect 254 4625 288 4659
rect 254 4556 288 4590
rect 254 4487 288 4521
rect 254 4418 288 4452
rect 254 4349 288 4383
rect 254 4280 288 4314
rect 254 4211 288 4245
rect 254 4142 288 4176
rect 254 4073 288 4107
rect 254 4004 288 4038
rect 254 3935 288 3969
rect 254 3866 288 3900
rect 254 3797 288 3831
rect 254 3728 288 3762
rect 662 4660 696 4694
rect 662 4591 696 4625
rect 662 4522 696 4556
rect 662 4453 696 4487
rect 662 4384 696 4418
rect 662 4315 696 4349
rect 662 4246 696 4280
rect 662 4177 696 4211
rect 662 4108 696 4142
rect 662 4039 696 4073
rect 662 3970 696 4004
rect 662 3901 696 3935
rect 662 3832 696 3866
rect 662 3763 696 3797
rect 254 3659 288 3693
rect 254 3590 288 3624
rect 662 3694 696 3728
rect 662 3625 696 3659
rect 254 3521 288 3555
rect 254 3452 288 3486
rect 254 3383 288 3417
rect 254 3314 288 3348
rect 254 3245 288 3279
rect 254 3176 288 3210
rect 254 3107 288 3141
rect 254 3038 288 3072
rect 254 2969 288 3003
rect 254 2900 288 2934
rect 254 2831 288 2865
rect 254 2762 288 2796
rect 254 2693 288 2727
rect 254 2624 288 2658
rect 662 3556 696 3590
rect 662 3487 696 3521
rect 662 3418 696 3452
rect 662 3349 696 3383
rect 662 3280 696 3314
rect 662 3211 696 3245
rect 662 3142 696 3176
rect 662 3073 696 3107
rect 662 3004 696 3038
rect 662 2935 696 2969
rect 662 2866 696 2900
rect 662 2797 696 2831
rect 662 2728 696 2762
rect 662 2659 696 2693
rect 254 2555 288 2589
rect 254 2486 288 2520
rect 662 2590 696 2624
rect 662 2522 696 2556
rect 254 2417 288 2451
rect 254 2348 288 2382
rect 254 2279 288 2313
rect 254 2210 288 2244
rect 254 2141 288 2175
rect 254 2072 288 2106
rect 254 2003 288 2037
rect 254 1934 288 1968
rect 254 1865 288 1899
rect 254 1796 288 1830
rect 254 1727 288 1761
rect 254 1658 288 1692
rect 254 1589 288 1623
rect 254 1520 288 1554
rect 254 1451 288 1485
rect 662 2454 696 2488
rect 662 2386 696 2420
rect 662 2318 696 2352
rect 662 2250 696 2284
rect 662 2182 696 2216
rect 662 2114 696 2148
rect 662 2046 696 2080
rect 662 1978 696 2012
rect 662 1910 696 1944
rect 662 1842 696 1876
rect 662 1774 696 1808
rect 662 1706 696 1740
rect 662 1638 696 1672
rect 662 1570 696 1604
rect 662 1502 696 1536
rect 254 1382 288 1416
rect 662 1434 696 1468
rect 662 1366 696 1400
rect 254 1313 288 1347
rect 254 1244 288 1278
rect 254 1175 288 1209
rect 254 1106 288 1140
rect 254 1037 288 1071
rect 254 968 288 1002
rect 254 899 288 933
rect 254 830 288 864
rect 254 761 288 795
rect 254 692 288 726
rect 254 623 288 657
rect 254 554 288 588
rect 254 485 288 519
rect 254 416 288 450
rect 254 347 288 381
rect 662 1298 696 1332
rect 662 1230 696 1264
rect 662 1162 696 1196
rect 662 1094 696 1128
rect 662 1026 696 1060
rect 662 958 696 992
rect 662 890 696 924
rect 662 822 696 856
rect 662 754 696 788
rect 662 686 696 720
rect 662 618 696 652
rect 662 550 696 584
rect 662 482 696 516
rect 662 414 696 448
rect 662 346 696 380
rect 254 278 288 312
rect 352 254 386 288
rect 423 254 457 288
rect 494 254 528 288
rect 566 254 600 288
rect 638 254 672 288
<< mvnsubdiffcont >>
rect 185 7217 219 7251
rect 261 7217 295 7251
rect 337 7217 371 7251
rect 413 7217 447 7251
rect 488 7217 522 7251
rect 563 7217 597 7251
rect 638 7217 672 7251
rect 713 7217 747 7251
rect 68 7067 102 7101
rect 68 6999 102 7033
rect 68 6931 102 6965
rect 68 6863 102 6897
rect 68 6795 102 6829
rect 68 6727 102 6761
rect 68 6659 102 6693
rect 68 6591 102 6625
rect 68 6523 102 6557
rect 68 6455 102 6489
rect 68 6387 102 6421
rect 68 6319 102 6353
rect 68 6251 102 6285
rect 68 6183 102 6217
rect 68 6115 102 6149
rect 68 6047 102 6081
rect 68 5979 102 6013
rect 68 5911 102 5945
rect 68 5843 102 5877
rect 68 5775 102 5809
rect 68 5707 102 5741
rect 68 5639 102 5673
rect 68 5571 102 5605
rect 68 5503 102 5537
rect 68 5435 102 5469
rect 68 5367 102 5401
rect 68 5299 102 5333
rect 68 5231 102 5265
rect 68 5163 102 5197
rect 68 5095 102 5129
rect 68 5027 102 5061
rect 68 4959 102 4993
rect 68 4891 102 4925
rect 68 4823 102 4857
rect 68 4755 102 4789
rect 68 4687 102 4721
rect 68 4619 102 4653
rect 68 4551 102 4585
rect 68 4483 102 4517
rect 68 4415 102 4449
rect 68 4347 102 4381
rect 68 4279 102 4313
rect 68 4211 102 4245
rect 68 4143 102 4177
rect 68 4075 102 4109
rect 68 4007 102 4041
rect 68 3939 102 3973
rect 68 3871 102 3905
rect 68 3803 102 3837
rect 68 3735 102 3769
rect 68 3667 102 3701
rect 68 3599 102 3633
rect 68 3531 102 3565
rect 68 3463 102 3497
rect 68 3395 102 3429
rect 68 3327 102 3361
rect 68 3259 102 3293
rect 68 3191 102 3225
rect 68 3123 102 3157
rect 68 3055 102 3089
rect 68 2987 102 3021
rect 68 2919 102 2953
rect 68 2851 102 2885
rect 68 2783 102 2817
rect 68 2715 102 2749
rect 68 2647 102 2681
rect 68 2579 102 2613
rect 68 2511 102 2545
rect 68 2443 102 2477
rect 68 2375 102 2409
rect 68 2307 102 2341
rect 68 2239 102 2273
rect 68 2171 102 2205
rect 68 2103 102 2137
rect 68 2035 102 2069
rect 68 1967 102 2001
rect 68 1899 102 1933
rect 68 1831 102 1865
rect 68 1763 102 1797
rect 68 1695 102 1729
rect 68 1627 102 1661
rect 68 1559 102 1593
rect 68 1491 102 1525
rect 68 1423 102 1457
rect 68 1355 102 1389
rect 68 1287 102 1321
rect 68 1219 102 1253
rect 68 1151 102 1185
rect 68 1083 102 1117
rect 68 1015 102 1049
rect 68 947 102 981
rect 68 879 102 913
rect 68 811 102 845
rect 68 743 102 777
rect 68 675 102 709
rect 68 607 102 641
rect 68 539 102 573
rect 68 471 102 505
rect 68 403 102 437
rect 68 335 102 369
rect 68 266 102 300
rect 68 197 102 231
rect 203 67 237 101
rect 273 67 307 101
rect 344 67 378 101
rect 415 67 449 101
rect 486 67 520 101
rect 557 67 591 101
rect 628 67 662 101
rect 699 67 733 101
rect 770 67 804 101
<< poly >>
rect 415 6956 535 6982
rect 415 5916 535 5956
rect 415 5882 472 5916
rect 506 5882 535 5916
rect 415 5835 535 5882
rect 415 4795 535 4835
rect 415 4761 472 4795
rect 506 4761 535 4795
rect 415 4714 535 4761
rect 415 3676 535 3714
rect 415 3642 472 3676
rect 506 3642 535 3676
rect 415 3604 535 3642
rect 415 2556 535 2604
rect 415 2522 472 2556
rect 506 2522 535 2556
rect 415 2483 535 2522
rect 415 1435 535 1483
rect 415 1401 472 1435
rect 506 1401 535 1435
rect 415 1362 535 1401
rect 415 336 535 362
<< polycont >>
rect 472 5882 506 5916
rect 472 4761 506 4795
rect 472 3642 506 3676
rect 472 2522 506 2556
rect 472 1401 506 1435
<< locali >>
rect -44 7217 24 7251
rect 58 7217 96 7251
rect 130 7217 168 7251
rect 219 7217 247 7251
rect 295 7217 326 7251
rect 371 7217 405 7251
rect 447 7217 483 7251
rect 522 7217 561 7251
rect 597 7217 638 7251
rect 673 7217 713 7251
rect 751 7217 795 7251
rect 829 7217 882 7251
rect -44 7215 102 7217
rect -28 7181 102 7215
rect -62 7143 102 7181
rect -28 7109 102 7143
rect -62 7101 102 7109
rect -62 7071 68 7101
rect -28 7067 68 7071
rect -28 7037 102 7067
rect -62 7033 102 7037
rect -62 6999 68 7033
rect -28 6965 102 6999
rect -62 6931 68 6965
rect -62 6927 102 6931
rect -28 6897 102 6927
rect -28 6893 68 6897
rect -62 6863 68 6893
rect -62 6855 102 6863
rect -28 6829 102 6855
rect -28 6821 68 6829
rect -62 6795 68 6821
rect -62 6783 102 6795
rect -28 6761 102 6783
rect -28 6749 68 6761
rect -62 6727 68 6749
rect -62 6711 102 6727
rect -28 6693 102 6711
rect -28 6677 68 6693
rect -62 6659 68 6677
rect -62 6639 102 6659
rect -28 6625 102 6639
rect -28 6605 68 6625
rect -62 6591 68 6605
rect -62 6567 102 6591
rect -28 6557 102 6567
rect -28 6533 68 6557
rect -62 6523 68 6533
rect -62 6495 102 6523
rect -28 6489 102 6495
rect -28 6461 68 6489
rect -62 6455 68 6461
rect -62 6423 102 6455
rect -28 6421 102 6423
rect -28 6389 68 6421
rect -62 6387 68 6389
rect -62 6353 102 6387
rect -62 6351 68 6353
rect -28 6319 68 6351
rect -28 6317 102 6319
rect -62 6285 102 6317
rect -62 6279 68 6285
rect -28 6251 68 6279
rect -28 6245 102 6251
rect -62 6217 102 6245
rect -62 6207 68 6217
rect -28 6183 68 6207
rect -28 6173 102 6183
rect -62 6149 102 6173
rect -62 6135 68 6149
rect -28 6115 68 6135
rect -28 6101 102 6115
rect -62 6081 102 6101
rect -62 6063 68 6081
rect -28 6047 68 6063
rect -28 6029 102 6047
rect -62 6013 102 6029
rect -62 5991 68 6013
rect -28 5979 68 5991
rect -28 5957 102 5979
rect -62 5945 102 5957
rect -62 5919 68 5945
rect -28 5911 68 5919
rect -28 5885 102 5911
rect -62 5877 102 5885
rect -62 5847 68 5877
rect -28 5843 68 5847
rect -28 5813 102 5843
rect -62 5809 102 5813
rect -62 5775 68 5809
rect -28 5741 102 5775
rect -62 5707 68 5741
rect -62 5703 102 5707
rect -28 5673 102 5703
rect -28 5669 68 5673
rect -62 5639 68 5669
rect -62 5631 102 5639
rect -28 5605 102 5631
rect -28 5597 68 5605
rect -62 5571 68 5597
rect -62 5559 102 5571
rect -28 5537 102 5559
rect -28 5525 68 5537
rect -62 5503 68 5525
rect -62 5487 102 5503
rect -28 5469 102 5487
rect -28 5453 68 5469
rect -62 5435 68 5453
rect -62 5415 102 5435
rect -28 5401 102 5415
rect -28 5381 68 5401
rect -62 5367 68 5381
rect -62 5343 102 5367
rect -28 5333 102 5343
rect -28 5309 68 5333
rect -62 5299 68 5309
rect -62 5271 102 5299
rect -28 5265 102 5271
rect -28 5237 68 5265
rect -62 5231 68 5237
rect -62 5199 102 5231
rect -28 5197 102 5199
rect -28 5165 68 5197
rect -62 5163 68 5165
rect -62 5129 102 5163
rect -62 5127 68 5129
rect -28 5095 68 5127
rect -28 5093 102 5095
rect -62 5061 102 5093
rect -62 5055 68 5061
rect -28 5027 68 5055
rect -28 5021 102 5027
rect -62 4993 102 5021
rect -62 4983 68 4993
rect -28 4959 68 4983
rect -28 4949 102 4959
rect -62 4925 102 4949
rect -62 4911 68 4925
rect -28 4891 68 4911
rect -28 4877 102 4891
rect -62 4857 102 4877
rect -62 4839 68 4857
rect -28 4823 68 4839
rect -28 4805 102 4823
rect -62 4789 102 4805
rect -62 4767 68 4789
rect -28 4755 68 4767
rect -28 4733 102 4755
rect -62 4721 102 4733
rect -62 4695 68 4721
rect -28 4687 68 4695
rect -28 4661 102 4687
rect -62 4653 102 4661
rect -62 4623 68 4653
rect -28 4619 68 4623
rect -28 4589 102 4619
rect -62 4585 102 4589
rect -62 4551 68 4585
rect -28 4517 102 4551
rect -62 4483 68 4517
rect -62 4479 102 4483
rect -28 4449 102 4479
rect -28 4445 68 4449
rect -62 4415 68 4445
rect -62 4407 102 4415
rect -28 4381 102 4407
rect -28 4373 68 4381
rect -62 4347 68 4373
rect -62 4335 102 4347
rect -28 4313 102 4335
rect -28 4301 68 4313
rect -62 4279 68 4301
rect -62 4263 102 4279
rect -28 4245 102 4263
rect -28 4229 68 4245
rect -62 4211 68 4229
rect -62 4191 102 4211
rect -28 4177 102 4191
rect -28 4157 68 4177
rect -62 4143 68 4157
rect -62 4119 102 4143
rect -28 4109 102 4119
rect -28 4085 68 4109
rect -62 4075 68 4085
rect -62 4047 102 4075
rect -28 4041 102 4047
rect -28 4013 68 4041
rect -62 4007 68 4013
rect -62 3975 102 4007
rect -28 3973 102 3975
rect -28 3941 68 3973
rect -62 3939 68 3941
rect -62 3905 102 3939
rect -62 3903 68 3905
rect -28 3871 68 3903
rect -28 3869 102 3871
rect -62 3837 102 3869
rect -62 3831 68 3837
rect -28 3803 68 3831
rect -28 3797 102 3803
rect -62 3769 102 3797
rect -62 3759 68 3769
rect -28 3735 68 3759
rect -28 3725 102 3735
rect -62 3701 102 3725
rect -62 3687 68 3701
rect -28 3667 68 3687
rect -28 3653 102 3667
rect -62 3633 102 3653
rect -62 3615 68 3633
rect -28 3599 68 3615
rect -28 3581 102 3599
rect -62 3565 102 3581
rect -62 3543 68 3565
rect -28 3531 68 3543
rect -28 3509 102 3531
rect -62 3497 102 3509
rect -62 3471 68 3497
rect -28 3463 68 3471
rect -28 3437 102 3463
rect -62 3436 102 3437
rect -62 3399 -28 3436
rect -62 3327 -28 3365
rect -62 3262 -28 3293
rect 24 3429 102 3436
rect 24 3395 68 3429
rect 24 3361 102 3395
rect 24 3327 68 3361
rect 24 3293 102 3327
rect 24 3262 68 3293
rect -62 3259 68 3262
rect -62 3255 102 3259
rect -28 3225 102 3255
rect -28 3221 68 3225
rect -62 3191 68 3221
rect -62 3183 102 3191
rect -28 3157 102 3183
rect -28 3149 68 3157
rect -62 3123 68 3149
rect -62 3111 102 3123
rect -28 3089 102 3111
rect -28 3077 68 3089
rect -62 3055 68 3077
rect -62 3039 102 3055
rect -28 3021 102 3039
rect -28 3005 68 3021
rect -62 2987 68 3005
rect -62 2967 102 2987
rect -28 2953 102 2967
rect -28 2933 68 2953
rect -62 2919 68 2933
rect -62 2895 102 2919
rect -28 2885 102 2895
rect -28 2861 68 2885
rect -62 2851 68 2861
rect -62 2823 102 2851
rect -28 2817 102 2823
rect -28 2789 68 2817
rect -62 2783 68 2789
rect -62 2751 102 2783
rect -28 2749 102 2751
rect -28 2717 68 2749
rect -62 2715 68 2717
rect -62 2681 102 2715
rect -62 2679 68 2681
rect -28 2647 68 2679
rect -28 2645 102 2647
rect -62 2613 102 2645
rect -62 2607 68 2613
rect -28 2579 68 2607
rect -28 2573 102 2579
rect -62 2545 102 2573
rect -62 2535 68 2545
rect -28 2511 68 2535
rect -28 2501 102 2511
rect -62 2477 102 2501
rect -62 2463 68 2477
rect -28 2443 68 2463
rect -28 2429 102 2443
rect -62 2409 102 2429
rect -62 2391 68 2409
rect -28 2375 68 2391
rect -28 2357 102 2375
rect -62 2341 102 2357
rect -62 2319 68 2341
rect -28 2307 68 2319
rect -28 2285 102 2307
rect -62 2273 102 2285
rect -62 2247 68 2273
rect -28 2239 68 2247
rect -28 2213 102 2239
rect -62 2205 102 2213
rect -62 2175 68 2205
rect -28 2171 68 2175
rect -28 2141 102 2171
rect -62 2137 102 2141
rect -62 2103 68 2137
rect -28 2069 102 2103
rect -62 2035 68 2069
rect -62 2031 102 2035
rect -28 2001 102 2031
rect -28 1997 68 2001
rect -62 1967 68 1997
rect -62 1959 102 1967
rect -28 1933 102 1959
rect -28 1925 68 1933
rect -62 1899 68 1925
rect -62 1887 102 1899
rect -28 1865 102 1887
rect -28 1853 68 1865
rect -62 1831 68 1853
rect -62 1815 102 1831
rect -28 1797 102 1815
rect -28 1781 68 1797
rect -62 1763 68 1781
rect -62 1743 102 1763
rect -28 1729 102 1743
rect -28 1709 68 1729
rect -62 1695 68 1709
rect -62 1670 102 1695
rect -28 1661 102 1670
rect -28 1636 68 1661
rect -62 1627 68 1636
rect -62 1597 102 1627
rect -28 1593 102 1597
rect -28 1563 68 1593
rect -62 1559 68 1563
rect -62 1525 102 1559
rect -62 1524 68 1525
rect -28 1491 68 1524
rect -28 1490 102 1491
rect -62 1457 102 1490
rect -62 1451 68 1457
rect -28 1423 68 1451
rect -28 1417 102 1423
rect -62 1389 102 1417
rect -62 1378 68 1389
rect -28 1355 68 1378
rect -28 1344 102 1355
rect -62 1321 102 1344
rect -62 1305 68 1321
rect -28 1287 68 1305
rect -28 1271 102 1287
rect -62 1253 102 1271
rect -62 1232 68 1253
rect -28 1219 68 1232
rect -28 1198 102 1219
rect -62 1185 102 1198
rect -62 1159 68 1185
rect -28 1151 68 1159
rect -28 1125 102 1151
rect -62 1117 102 1125
rect -62 1086 68 1117
rect -28 1083 68 1086
rect -28 1052 102 1083
rect -62 1049 102 1052
rect -62 1015 68 1049
rect -62 1013 102 1015
rect -28 981 102 1013
rect -28 979 68 981
rect -62 947 68 979
rect -62 940 102 947
rect -28 913 102 940
rect -28 906 68 913
rect -62 879 68 906
rect -62 867 102 879
rect -28 845 102 867
rect -28 833 68 845
rect -62 811 68 833
rect -62 794 102 811
rect -28 777 102 794
rect -28 760 68 777
rect -62 743 68 760
rect -62 721 102 743
rect -28 709 102 721
rect -28 687 68 709
rect -62 675 68 687
rect -62 648 102 675
rect -28 641 102 648
rect -28 614 68 641
rect -62 607 68 614
rect -62 575 102 607
rect -28 573 102 575
rect -28 541 68 573
rect -62 539 68 541
rect -62 505 102 539
rect -62 502 68 505
rect -28 471 68 502
rect -28 468 102 471
rect -62 437 102 468
rect -62 429 68 437
rect -28 403 68 429
rect -28 395 102 403
rect -62 369 102 395
rect -62 356 68 369
rect -28 335 68 356
rect -28 322 102 335
rect -62 300 102 322
rect -62 283 68 300
rect -28 266 68 283
rect -28 249 102 266
rect -62 231 102 249
rect -62 210 68 231
rect -28 197 68 210
rect -28 176 102 197
rect -62 137 102 176
rect 154 7064 796 7165
rect 154 7055 278 7064
rect 312 7055 391 7064
rect 425 7055 525 7064
rect 559 7055 796 7064
rect 154 7021 225 7055
rect 259 7030 278 7055
rect 259 7021 305 7030
rect 339 7021 385 7055
rect 425 7030 465 7055
rect 419 7021 465 7030
rect 499 7030 525 7055
rect 580 7040 796 7055
rect 499 7021 546 7030
rect 580 7021 662 7040
rect 154 7006 662 7021
rect 696 7006 796 7040
rect 154 7000 796 7006
rect 154 6982 318 7000
rect 154 6948 225 6982
rect 259 6972 318 6982
rect 154 6938 254 6948
rect 288 6938 318 6972
rect 523 6982 796 7000
rect 154 6909 318 6938
rect 154 6875 225 6909
rect 259 6904 318 6909
rect 154 6870 254 6875
rect 288 6870 318 6904
rect 154 6836 318 6870
rect 154 6802 225 6836
rect 288 6802 318 6836
rect 154 6768 318 6802
rect 154 6763 254 6768
rect 154 6729 225 6763
rect 288 6734 318 6768
rect 259 6729 318 6734
rect 154 6700 318 6729
rect 154 6690 254 6700
rect 154 6656 225 6690
rect 288 6666 318 6700
rect 259 6656 318 6666
rect 154 6632 318 6656
rect 154 6617 254 6632
rect 154 6583 225 6617
rect 288 6598 318 6632
rect 259 6583 318 6598
rect 154 6564 318 6583
rect 154 6544 254 6564
rect 154 6510 225 6544
rect 288 6530 318 6564
rect 259 6510 318 6530
rect 154 6496 318 6510
rect 154 6471 254 6496
rect 154 6437 225 6471
rect 288 6462 318 6496
rect 259 6437 318 6462
rect 154 6428 318 6437
rect 154 6398 254 6428
rect 154 6364 225 6398
rect 288 6394 318 6428
rect 259 6364 318 6394
rect 154 6360 318 6364
rect 154 6326 254 6360
rect 288 6326 318 6360
rect 154 6325 318 6326
rect 154 6291 225 6325
rect 259 6292 318 6325
rect 154 6258 254 6291
rect 288 6258 318 6292
rect 154 6252 318 6258
rect 154 6218 225 6252
rect 259 6224 318 6252
rect 154 6190 254 6218
rect 288 6190 318 6224
rect 154 6179 318 6190
rect 154 6145 225 6179
rect 259 6156 318 6179
rect 154 6122 254 6145
rect 288 6122 318 6156
rect 154 6106 318 6122
rect 154 6072 225 6106
rect 259 6088 318 6106
rect 154 6054 254 6072
rect 288 6054 318 6088
rect 154 6033 318 6054
rect 154 5999 225 6033
rect 259 6020 318 6033
rect 154 5986 254 5999
rect 288 5986 318 6020
rect 154 5960 318 5986
rect 154 5926 225 5960
rect 259 5952 318 5960
rect 154 5918 254 5926
rect 288 5918 318 5952
rect 154 5887 318 5918
rect 154 5853 225 5887
rect 259 5884 318 5887
rect 154 5850 254 5853
rect 288 5850 318 5884
rect 154 5816 318 5850
rect 154 5814 254 5816
rect 154 5780 225 5814
rect 288 5782 318 5816
rect 259 5780 318 5782
rect 154 5748 318 5780
rect 154 5741 254 5748
rect 154 5707 225 5741
rect 288 5714 318 5748
rect 259 5707 318 5714
rect 154 5680 318 5707
rect 154 5668 254 5680
rect 154 5634 225 5668
rect 288 5646 318 5680
rect 259 5634 318 5646
rect 154 5612 318 5634
rect 154 5595 254 5612
rect 154 5561 225 5595
rect 288 5578 318 5612
rect 259 5561 318 5578
rect 154 5544 318 5561
rect 154 5522 254 5544
rect 154 5488 225 5522
rect 288 5510 318 5544
rect 259 5488 318 5510
rect 154 5476 318 5488
rect 154 5449 254 5476
rect 154 5415 225 5449
rect 288 5442 318 5476
rect 259 5415 318 5442
rect 154 5408 318 5415
rect 154 5376 254 5408
rect 154 5342 225 5376
rect 288 5374 318 5408
rect 259 5342 318 5374
rect 154 5340 318 5342
rect 154 5306 254 5340
rect 288 5306 318 5340
rect 154 5303 318 5306
rect 154 5269 225 5303
rect 259 5272 318 5303
rect 154 5238 254 5269
rect 288 5238 318 5272
rect 154 5230 318 5238
rect 154 5196 225 5230
rect 259 5204 318 5230
rect 154 5170 254 5196
rect 288 5170 318 5204
rect 154 5157 318 5170
rect 154 5123 225 5157
rect 259 5136 318 5157
rect 154 5102 254 5123
rect 288 5102 318 5136
rect 154 5084 318 5102
rect 154 5050 225 5084
rect 259 5068 318 5084
rect 154 5034 254 5050
rect 288 5034 318 5068
rect 154 5011 318 5034
rect 154 4977 225 5011
rect 259 5000 318 5011
rect 154 4966 254 4977
rect 288 4966 318 5000
rect 154 4938 318 4966
rect 154 4904 225 4938
rect 259 4932 318 4938
rect 154 4898 254 4904
rect 288 4898 318 4932
rect 154 4865 318 4898
rect 154 4831 225 4865
rect 259 4864 318 4865
rect 154 4830 254 4831
rect 288 4830 318 4864
rect 154 4796 318 4830
rect 154 4792 254 4796
rect 154 4758 225 4792
rect 288 4762 318 4796
rect 259 4758 318 4762
rect 154 4728 318 4758
rect 154 4719 254 4728
rect 154 4685 225 4719
rect 288 4694 318 4728
rect 259 4685 318 4694
rect 154 4659 318 4685
rect 154 4646 254 4659
rect 154 4612 225 4646
rect 288 4625 318 4659
rect 259 4612 318 4625
rect 154 4590 318 4612
rect 154 4573 254 4590
rect 154 4539 225 4573
rect 288 4556 318 4590
rect 259 4539 318 4556
rect 154 4521 318 4539
rect 154 4500 254 4521
rect 154 4466 225 4500
rect 288 4487 318 4521
rect 259 4466 318 4487
rect 154 4452 318 4466
rect 154 4427 254 4452
rect 154 4393 225 4427
rect 288 4418 318 4452
rect 259 4393 318 4418
rect 154 4383 318 4393
rect 154 4354 254 4383
rect 154 4320 225 4354
rect 288 4349 318 4383
rect 259 4320 318 4349
rect 154 4314 318 4320
rect 154 4281 254 4314
rect 154 4247 225 4281
rect 288 4280 318 4314
rect 259 4247 318 4280
rect 154 4245 318 4247
rect 154 4211 254 4245
rect 288 4211 318 4245
rect 154 4208 318 4211
rect 154 4174 225 4208
rect 259 4176 318 4208
rect 154 4142 254 4174
rect 288 4142 318 4176
rect 154 4135 318 4142
rect 154 4101 225 4135
rect 259 4107 318 4135
rect 154 4073 254 4101
rect 288 4073 318 4107
rect 154 4062 318 4073
rect 154 4028 225 4062
rect 259 4038 318 4062
rect 154 4004 254 4028
rect 288 4004 318 4038
rect 154 3989 318 4004
rect 154 3955 225 3989
rect 259 3969 318 3989
rect 154 3935 254 3955
rect 288 3935 318 3969
rect 154 3916 318 3935
rect 154 3882 225 3916
rect 259 3900 318 3916
rect 154 3866 254 3882
rect 288 3866 318 3900
rect 154 3843 318 3866
rect 154 3809 225 3843
rect 259 3831 318 3843
rect 154 3797 254 3809
rect 288 3797 318 3831
rect 154 3770 318 3797
rect 154 3736 225 3770
rect 259 3762 318 3770
rect 154 3728 254 3736
rect 288 3728 318 3762
rect 154 3697 318 3728
rect 154 3663 225 3697
rect 259 3693 318 3697
rect 154 3659 254 3663
rect 288 3659 318 3693
rect 154 3624 318 3659
rect 154 3590 225 3624
rect 288 3590 318 3624
rect 154 3555 318 3590
rect 154 3551 254 3555
rect 154 3517 225 3551
rect 288 3521 318 3555
rect 259 3517 318 3521
rect 154 3486 318 3517
rect 154 3478 254 3486
rect 154 3444 225 3478
rect 288 3452 318 3486
rect 259 3444 318 3452
rect 154 3417 318 3444
rect 154 3405 254 3417
rect 154 3371 225 3405
rect 288 3383 318 3417
rect 259 3371 318 3383
rect 154 3348 318 3371
rect 154 3332 254 3348
rect 154 3298 225 3332
rect 288 3314 318 3348
rect 259 3298 318 3314
rect 154 3279 318 3298
rect 154 3260 254 3279
rect 154 3226 225 3260
rect 288 3245 318 3279
rect 259 3226 318 3245
rect 154 3210 318 3226
rect 154 3188 254 3210
rect 154 3154 225 3188
rect 288 3176 318 3210
rect 259 3154 318 3176
rect 154 3141 318 3154
rect 154 3116 254 3141
rect 154 3082 225 3116
rect 288 3107 318 3141
rect 259 3082 318 3107
rect 154 3072 318 3082
rect 154 3044 254 3072
rect 154 3010 225 3044
rect 288 3038 318 3072
rect 259 3010 318 3038
rect 154 3003 318 3010
rect 154 2972 254 3003
rect 154 2938 225 2972
rect 288 2969 318 3003
rect 259 2938 318 2969
rect 154 2934 318 2938
rect 154 2900 254 2934
rect 288 2900 318 2934
rect 154 2866 225 2900
rect 259 2866 318 2900
rect 154 2865 318 2866
rect 154 2831 254 2865
rect 288 2831 318 2865
rect 154 2828 318 2831
rect 154 2794 225 2828
rect 259 2796 318 2828
rect 154 2762 254 2794
rect 288 2762 318 2796
rect 154 2756 318 2762
rect 154 2722 225 2756
rect 259 2727 318 2756
rect 154 2693 254 2722
rect 288 2693 318 2727
rect 154 2684 318 2693
rect 154 2650 225 2684
rect 259 2658 318 2684
rect 154 2624 254 2650
rect 288 2624 318 2658
rect 154 2612 318 2624
rect 154 2578 225 2612
rect 259 2589 318 2612
rect 154 2555 254 2578
rect 288 2555 318 2589
rect 154 2540 318 2555
rect 154 2506 225 2540
rect 259 2520 318 2540
rect 154 2486 254 2506
rect 288 2486 318 2520
rect 154 2468 318 2486
rect 154 2434 225 2468
rect 259 2451 318 2468
rect 154 2417 254 2434
rect 288 2417 318 2451
rect 154 2396 318 2417
rect 154 2362 225 2396
rect 259 2382 318 2396
rect 154 2348 254 2362
rect 288 2348 318 2382
rect 154 2324 318 2348
rect 154 2290 225 2324
rect 259 2313 318 2324
rect 154 2279 254 2290
rect 288 2279 318 2313
rect 154 2252 318 2279
rect 154 2218 225 2252
rect 259 2244 318 2252
rect 154 2210 254 2218
rect 288 2210 318 2244
rect 154 2180 318 2210
rect 154 2146 225 2180
rect 259 2175 318 2180
rect 154 2141 254 2146
rect 288 2141 318 2175
rect 154 2108 318 2141
rect 154 2074 225 2108
rect 259 2106 318 2108
rect 154 2072 254 2074
rect 288 2072 318 2106
rect 154 2037 318 2072
rect 154 2036 254 2037
rect 154 2002 225 2036
rect 288 2003 318 2037
rect 259 2002 318 2003
rect 154 1968 318 2002
rect 154 1964 254 1968
rect 154 1930 225 1964
rect 288 1934 318 1968
rect 259 1930 318 1934
rect 154 1899 318 1930
rect 154 1892 254 1899
rect 154 1858 225 1892
rect 288 1865 318 1899
rect 259 1858 318 1865
rect 154 1830 318 1858
rect 154 1820 254 1830
rect 154 1786 225 1820
rect 288 1796 318 1830
rect 259 1786 318 1796
rect 154 1761 318 1786
rect 154 1748 254 1761
rect 154 1714 225 1748
rect 288 1727 318 1761
rect 259 1714 318 1727
rect 154 1692 318 1714
rect 154 1676 254 1692
rect 154 1642 225 1676
rect 288 1658 318 1692
rect 259 1642 318 1658
rect 154 1623 318 1642
rect 154 1604 254 1623
rect 154 1570 225 1604
rect 288 1589 318 1623
rect 259 1570 318 1589
rect 154 1554 318 1570
rect 154 1532 254 1554
rect 154 1498 225 1532
rect 288 1520 318 1554
rect 259 1498 318 1520
rect 154 1485 318 1498
rect 154 1460 254 1485
rect 154 1426 225 1460
rect 288 1451 318 1485
rect 259 1426 318 1451
rect 154 1416 318 1426
rect 154 1388 254 1416
rect 154 1354 225 1388
rect 288 1382 318 1416
rect 259 1354 318 1382
rect 154 1347 318 1354
rect 154 1316 254 1347
rect 154 1282 225 1316
rect 288 1313 318 1347
rect 259 1282 318 1313
rect 154 1278 318 1282
rect 154 1244 254 1278
rect 288 1244 318 1278
rect 154 1210 225 1244
rect 259 1210 318 1244
rect 154 1209 318 1210
rect 154 1175 254 1209
rect 288 1175 318 1209
rect 154 1172 318 1175
rect 154 1138 225 1172
rect 259 1140 318 1172
rect 154 1106 254 1138
rect 288 1106 318 1140
rect 154 1100 318 1106
rect 154 1066 225 1100
rect 259 1071 318 1100
rect 154 1037 254 1066
rect 288 1037 318 1071
rect 154 1028 318 1037
rect 154 994 225 1028
rect 259 1002 318 1028
rect 154 968 254 994
rect 288 968 318 1002
rect 154 956 318 968
rect 154 922 225 956
rect 259 933 318 956
rect 154 899 254 922
rect 288 899 318 933
rect 154 884 318 899
rect 154 850 225 884
rect 259 864 318 884
rect 154 830 254 850
rect 288 830 318 864
rect 154 812 318 830
rect 154 778 225 812
rect 259 795 318 812
rect 154 761 254 778
rect 288 761 318 795
rect 154 740 318 761
rect 154 706 225 740
rect 259 726 318 740
rect 154 692 254 706
rect 288 692 318 726
rect 154 668 318 692
rect 154 634 225 668
rect 259 657 318 668
rect 154 623 254 634
rect 288 623 318 657
rect 154 596 318 623
rect 154 562 225 596
rect 259 588 318 596
rect 154 554 254 562
rect 288 554 318 588
rect 154 524 318 554
rect 154 490 225 524
rect 259 519 318 524
rect 154 485 254 490
rect 288 485 318 519
rect 154 452 318 485
rect 154 418 225 452
rect 259 450 318 452
rect 154 416 254 418
rect 288 416 318 450
rect 154 381 318 416
rect 154 380 254 381
rect 154 346 225 380
rect 288 347 318 381
rect 370 6944 471 6960
rect 404 6910 471 6944
rect 370 6892 471 6910
rect 404 6842 471 6892
rect 370 6819 471 6842
rect 404 6774 471 6819
rect 370 6746 471 6774
rect 404 6706 471 6746
rect 370 6673 471 6706
rect 404 6638 471 6673
rect 370 6604 471 6638
rect 404 6566 471 6604
rect 370 6536 471 6566
rect 404 6493 471 6536
rect 370 6468 471 6493
rect 404 6420 471 6468
rect 370 6400 471 6420
rect 404 6347 471 6400
rect 370 6332 471 6347
rect 404 6274 471 6332
rect 370 6264 471 6274
rect 404 6201 471 6264
rect 370 6196 471 6201
rect 404 6094 471 6196
rect 370 6089 471 6094
rect 404 6026 471 6089
rect 370 6016 471 6026
rect 404 5982 471 6016
rect 370 5966 471 5982
rect 523 6948 546 6982
rect 580 6971 796 6982
rect 580 6948 662 6971
rect 523 6944 662 6948
rect 523 6910 546 6944
rect 580 6937 662 6944
rect 696 6937 796 6971
rect 580 6910 796 6937
rect 523 6909 796 6910
rect 523 6842 546 6909
rect 580 6902 796 6909
rect 580 6868 662 6902
rect 696 6868 796 6902
rect 580 6842 796 6868
rect 523 6836 796 6842
rect 523 6774 546 6836
rect 580 6833 796 6836
rect 580 6799 662 6833
rect 696 6799 796 6833
rect 580 6774 796 6799
rect 523 6764 796 6774
rect 523 6763 662 6764
rect 523 6706 546 6763
rect 580 6730 662 6763
rect 696 6730 796 6764
rect 580 6706 796 6730
rect 523 6695 796 6706
rect 523 6690 662 6695
rect 523 6638 546 6690
rect 580 6661 662 6690
rect 696 6661 796 6695
rect 580 6638 796 6661
rect 523 6626 796 6638
rect 523 6617 662 6626
rect 523 6570 546 6617
rect 580 6592 662 6617
rect 696 6592 796 6626
rect 580 6570 796 6592
rect 523 6557 796 6570
rect 523 6544 662 6557
rect 523 6502 546 6544
rect 580 6523 662 6544
rect 696 6523 796 6557
rect 580 6502 796 6523
rect 523 6488 796 6502
rect 523 6471 662 6488
rect 523 6434 546 6471
rect 580 6454 662 6471
rect 696 6454 796 6488
rect 580 6434 796 6454
rect 523 6419 796 6434
rect 523 6400 662 6419
rect 523 6364 546 6400
rect 580 6385 662 6400
rect 696 6385 796 6419
rect 580 6364 796 6385
rect 523 6350 796 6364
rect 523 6332 662 6350
rect 523 6291 546 6332
rect 580 6316 662 6332
rect 696 6316 796 6350
rect 580 6291 796 6316
rect 523 6281 796 6291
rect 523 6264 662 6281
rect 523 6218 546 6264
rect 580 6247 662 6264
rect 696 6247 796 6281
rect 580 6218 796 6247
rect 523 6212 796 6218
rect 523 6196 662 6212
rect 523 6145 546 6196
rect 580 6178 662 6196
rect 696 6178 796 6212
rect 580 6145 796 6178
rect 523 6143 796 6145
rect 523 6128 662 6143
rect 523 6072 546 6128
rect 580 6109 662 6128
rect 696 6109 796 6143
rect 580 6074 796 6109
rect 580 6072 662 6074
rect 523 6060 662 6072
rect 523 5999 546 6060
rect 580 6040 662 6060
rect 696 6040 796 6074
rect 580 6005 796 6040
rect 580 5999 662 6005
rect 523 5971 662 5999
rect 696 5971 796 6005
rect 523 5966 796 5971
rect 370 5943 438 5966
rect 404 5909 438 5943
rect 546 5960 796 5966
rect 370 5870 438 5909
rect 404 5836 438 5870
rect 370 5823 438 5836
rect 404 5763 438 5823
rect 370 5755 438 5763
rect 404 5690 438 5755
rect 370 5687 438 5690
rect 404 5653 438 5687
rect 370 5651 438 5653
rect 404 5585 438 5651
rect 370 5578 438 5585
rect 404 5517 438 5578
rect 370 5505 438 5517
rect 404 5449 438 5505
rect 370 5432 438 5449
rect 404 5381 438 5432
rect 370 5359 438 5381
rect 404 5313 438 5359
rect 370 5286 438 5313
rect 404 5245 438 5286
rect 370 5213 438 5245
rect 404 5177 438 5213
rect 370 5143 438 5177
rect 404 5106 438 5143
rect 370 5075 438 5106
rect 404 5033 438 5075
rect 370 5007 438 5033
rect 404 4960 438 5007
rect 370 4939 438 4960
rect 404 4887 438 4939
rect 370 4848 438 4887
rect 404 4814 438 4848
rect 370 4775 438 4814
rect 404 4741 438 4775
rect 370 4702 438 4741
rect 404 4668 438 4702
rect 370 4634 438 4668
rect 404 4595 438 4634
rect 370 4566 438 4595
rect 404 4522 438 4566
rect 370 4498 438 4522
rect 404 4449 438 4498
rect 370 4430 438 4449
rect 404 4376 438 4430
rect 370 4362 438 4376
rect 404 4303 438 4362
rect 370 4294 438 4303
rect 404 4230 438 4294
rect 370 4226 438 4230
rect 404 4192 438 4226
rect 370 4191 438 4192
rect 404 4124 438 4191
rect 370 4118 438 4124
rect 404 4056 438 4118
rect 370 4045 438 4056
rect 404 3988 438 4045
rect 370 3972 438 3988
rect 404 3920 438 3972
rect 370 3899 438 3920
rect 404 3852 438 3899
rect 370 3826 438 3852
rect 404 3784 438 3826
rect 370 3753 438 3784
rect 404 3719 438 3753
rect 370 3680 438 3719
rect 404 3646 438 3680
rect 370 3607 438 3646
rect 404 3573 438 3607
rect 370 3534 438 3573
rect 404 3500 438 3534
rect 370 3466 438 3500
rect 404 3427 438 3466
rect 370 3398 438 3427
rect 404 3354 438 3398
rect 370 3330 438 3354
rect 404 3281 438 3330
rect 370 3262 438 3281
rect 404 3207 438 3262
rect 370 3194 438 3207
rect 404 3129 438 3194
rect 370 3126 438 3129
rect 404 3092 438 3126
rect 370 3090 438 3092
rect 404 3024 438 3090
rect 370 3018 438 3024
rect 404 2956 438 3018
rect 370 2946 438 2956
rect 404 2888 438 2946
rect 370 2874 438 2888
rect 404 2820 438 2874
rect 370 2802 438 2820
rect 404 2752 438 2802
rect 370 2730 438 2752
rect 404 2684 438 2730
rect 370 2658 438 2684
rect 404 2616 438 2658
rect 370 2586 438 2616
rect 404 2552 438 2586
rect 370 2514 438 2552
rect 404 2480 438 2514
rect 370 2442 438 2480
rect 404 2379 438 2442
rect 370 2370 438 2379
rect 404 2311 438 2370
rect 370 2298 438 2311
rect 404 2243 438 2298
rect 370 2226 438 2243
rect 404 2175 438 2226
rect 370 2154 438 2175
rect 404 2107 438 2154
rect 370 2082 438 2107
rect 404 2039 438 2082
rect 370 2010 438 2039
rect 404 1971 438 2010
rect 370 1938 438 1971
rect 404 1903 438 1938
rect 370 1869 438 1903
rect 404 1832 438 1869
rect 370 1801 438 1832
rect 404 1760 438 1801
rect 370 1733 438 1760
rect 404 1688 438 1733
rect 370 1665 438 1688
rect 404 1616 438 1665
rect 370 1597 438 1616
rect 404 1544 438 1597
rect 370 1529 438 1544
rect 404 1472 438 1529
rect 370 1434 438 1472
rect 404 1400 438 1434
rect 370 1362 438 1400
rect 472 5922 506 5932
rect 472 5849 506 5882
rect 472 5776 506 5815
rect 472 5703 506 5742
rect 472 5630 506 5669
rect 472 5557 506 5596
rect 472 5484 506 5523
rect 472 5411 506 5450
rect 472 5338 506 5377
rect 472 5265 506 5304
rect 472 5192 506 5231
rect 472 5119 506 5158
rect 472 5046 506 5085
rect 472 4973 506 5012
rect 472 4900 506 4939
rect 472 4827 506 4866
rect 472 4754 506 4761
rect 472 4681 506 4720
rect 472 4608 506 4647
rect 472 4535 506 4574
rect 472 4461 506 4501
rect 472 4387 506 4427
rect 472 4313 506 4353
rect 472 4239 506 4279
rect 472 4165 506 4205
rect 472 4091 506 4131
rect 472 4017 506 4057
rect 472 3943 506 3983
rect 472 3869 506 3909
rect 472 3795 506 3835
rect 472 3721 506 3761
rect 472 3676 506 3687
rect 472 3572 506 3613
rect 472 3498 506 3538
rect 472 3424 506 3464
rect 472 3350 506 3390
rect 472 3276 506 3316
rect 472 3202 506 3242
rect 472 3128 506 3168
rect 472 3054 506 3094
rect 472 2980 506 3020
rect 472 2906 506 2946
rect 472 2832 506 2872
rect 472 2758 506 2798
rect 472 2684 506 2724
rect 472 2610 506 2650
rect 472 2556 506 2576
rect 472 2462 506 2502
rect 472 2388 506 2428
rect 472 2314 506 2354
rect 472 2241 506 2280
rect 472 2168 506 2207
rect 472 2095 506 2134
rect 472 2022 506 2061
rect 472 1949 506 1988
rect 472 1876 506 1915
rect 472 1803 506 1842
rect 472 1730 506 1769
rect 472 1657 506 1696
rect 472 1584 506 1623
rect 472 1511 506 1550
rect 472 1435 506 1477
rect 472 1385 506 1401
rect 580 5936 796 5960
rect 580 5926 662 5936
rect 546 5902 662 5926
rect 696 5902 796 5936
rect 546 5887 796 5902
rect 580 5867 796 5887
rect 580 5853 662 5867
rect 546 5833 662 5853
rect 696 5833 796 5867
rect 546 5823 796 5833
rect 580 5798 796 5823
rect 580 5780 662 5798
rect 546 5764 662 5780
rect 696 5764 796 5798
rect 546 5755 796 5764
rect 580 5729 796 5755
rect 580 5707 662 5729
rect 546 5695 662 5707
rect 696 5695 796 5729
rect 546 5687 796 5695
rect 580 5660 796 5687
rect 580 5634 662 5660
rect 546 5626 662 5634
rect 696 5626 796 5660
rect 546 5619 796 5626
rect 580 5591 796 5619
rect 580 5561 662 5591
rect 546 5557 662 5561
rect 696 5557 796 5591
rect 546 5551 796 5557
rect 580 5522 796 5551
rect 580 5488 662 5522
rect 696 5488 796 5522
rect 546 5483 796 5488
rect 580 5453 796 5483
rect 580 5419 662 5453
rect 696 5419 796 5453
rect 580 5384 796 5419
rect 580 5381 662 5384
rect 546 5376 662 5381
rect 580 5350 662 5376
rect 696 5350 796 5384
rect 580 5315 796 5350
rect 580 5313 662 5315
rect 546 5303 662 5313
rect 580 5281 662 5303
rect 696 5281 796 5315
rect 580 5246 796 5281
rect 580 5245 662 5246
rect 546 5230 662 5245
rect 580 5212 662 5230
rect 696 5212 796 5246
rect 580 5177 796 5212
rect 546 5157 662 5177
rect 580 5143 662 5157
rect 696 5143 796 5177
rect 580 5109 796 5143
rect 546 5108 796 5109
rect 546 5084 662 5108
rect 580 5074 662 5084
rect 696 5074 796 5108
rect 580 5041 796 5074
rect 546 5039 796 5041
rect 546 5011 662 5039
rect 580 5005 662 5011
rect 696 5005 796 5039
rect 580 4973 796 5005
rect 546 4970 796 4973
rect 546 4939 662 4970
rect 580 4936 662 4939
rect 696 4936 796 4970
rect 580 4904 796 4936
rect 546 4901 796 4904
rect 546 4867 662 4901
rect 696 4867 796 4901
rect 546 4865 796 4867
rect 580 4832 796 4865
rect 580 4831 662 4832
rect 546 4798 662 4831
rect 696 4798 796 4832
rect 546 4792 796 4798
rect 580 4763 796 4792
rect 580 4758 662 4763
rect 546 4729 662 4758
rect 696 4729 796 4763
rect 546 4719 796 4729
rect 580 4694 796 4719
rect 580 4668 662 4694
rect 546 4660 662 4668
rect 696 4660 796 4694
rect 546 4646 796 4660
rect 580 4625 796 4646
rect 580 4600 662 4625
rect 546 4591 662 4600
rect 696 4591 796 4625
rect 546 4573 796 4591
rect 580 4556 796 4573
rect 580 4532 662 4556
rect 546 4522 662 4532
rect 696 4522 796 4556
rect 546 4500 796 4522
rect 580 4487 796 4500
rect 580 4464 662 4487
rect 546 4453 662 4464
rect 696 4453 796 4487
rect 546 4430 796 4453
rect 580 4418 796 4430
rect 580 4392 662 4418
rect 546 4384 662 4392
rect 696 4384 796 4418
rect 546 4362 796 4384
rect 580 4349 796 4362
rect 580 4318 662 4349
rect 546 4315 662 4318
rect 696 4315 796 4349
rect 546 4294 796 4315
rect 580 4280 796 4294
rect 580 4246 662 4280
rect 696 4246 796 4280
rect 580 4244 796 4246
rect 546 4226 796 4244
rect 580 4211 796 4226
rect 580 4177 662 4211
rect 696 4177 796 4211
rect 580 4170 796 4177
rect 546 4158 796 4170
rect 580 4142 796 4158
rect 580 4108 662 4142
rect 696 4108 796 4142
rect 580 4096 796 4108
rect 546 4090 796 4096
rect 580 4073 796 4090
rect 580 4039 662 4073
rect 696 4039 796 4073
rect 580 4004 796 4039
rect 580 3988 662 4004
rect 546 3982 662 3988
rect 580 3970 662 3982
rect 696 3970 796 4004
rect 580 3935 796 3970
rect 580 3920 662 3935
rect 546 3908 662 3920
rect 580 3901 662 3908
rect 696 3901 796 3935
rect 580 3866 796 3901
rect 580 3852 662 3866
rect 546 3834 662 3852
rect 580 3832 662 3834
rect 696 3832 796 3866
rect 580 3797 796 3832
rect 580 3784 662 3797
rect 546 3763 662 3784
rect 696 3763 796 3797
rect 546 3760 796 3763
rect 580 3728 796 3760
rect 580 3726 662 3728
rect 546 3694 662 3726
rect 696 3694 796 3728
rect 546 3670 796 3694
rect 580 3659 796 3670
rect 580 3636 662 3659
rect 546 3625 662 3636
rect 696 3625 796 3659
rect 546 3597 796 3625
rect 580 3590 796 3597
rect 580 3563 662 3590
rect 546 3556 662 3563
rect 696 3556 796 3590
rect 546 3534 796 3556
rect 580 3521 796 3534
rect 580 3490 662 3521
rect 546 3487 662 3490
rect 696 3487 796 3521
rect 546 3466 796 3487
rect 580 3452 796 3466
rect 580 3418 662 3452
rect 696 3418 796 3452
rect 580 3417 796 3418
rect 546 3398 796 3417
rect 580 3383 796 3398
rect 580 3349 662 3383
rect 696 3349 796 3383
rect 580 3344 796 3349
rect 546 3330 796 3344
rect 580 3314 796 3330
rect 580 3280 662 3314
rect 696 3280 796 3314
rect 580 3271 796 3280
rect 546 3262 796 3271
rect 580 3245 796 3262
rect 580 3211 662 3245
rect 696 3211 796 3245
rect 580 3198 796 3211
rect 546 3194 796 3198
rect 580 3176 796 3194
rect 580 3160 662 3176
rect 546 3159 662 3160
rect 580 3142 662 3159
rect 696 3142 796 3176
rect 580 3107 796 3142
rect 580 3092 662 3107
rect 546 3086 662 3092
rect 580 3073 662 3086
rect 696 3073 796 3107
rect 580 3038 796 3073
rect 580 3024 662 3038
rect 546 3013 662 3024
rect 580 3004 662 3013
rect 696 3004 796 3038
rect 580 2969 796 3004
rect 580 2956 662 2969
rect 546 2940 662 2956
rect 580 2935 662 2940
rect 696 2935 796 2969
rect 580 2900 796 2935
rect 580 2888 662 2900
rect 546 2867 662 2888
rect 580 2866 662 2867
rect 696 2866 796 2900
rect 580 2831 796 2866
rect 580 2820 662 2831
rect 546 2797 662 2820
rect 696 2797 796 2831
rect 546 2794 796 2797
rect 580 2762 796 2794
rect 580 2752 662 2762
rect 546 2728 662 2752
rect 696 2728 796 2762
rect 546 2721 796 2728
rect 580 2693 796 2721
rect 580 2684 662 2693
rect 546 2659 662 2684
rect 696 2659 796 2693
rect 546 2650 796 2659
rect 580 2624 796 2650
rect 580 2614 662 2624
rect 546 2590 662 2614
rect 696 2590 796 2624
rect 546 2575 796 2590
rect 580 2556 796 2575
rect 580 2541 662 2556
rect 546 2522 662 2541
rect 696 2522 796 2556
rect 546 2502 796 2522
rect 580 2488 796 2502
rect 580 2468 662 2488
rect 546 2454 662 2468
rect 696 2454 796 2488
rect 546 2429 796 2454
rect 580 2420 796 2429
rect 580 2386 662 2420
rect 696 2386 796 2420
rect 580 2379 796 2386
rect 546 2356 796 2379
rect 580 2352 796 2356
rect 580 2318 662 2352
rect 696 2318 796 2352
rect 580 2311 796 2318
rect 546 2284 796 2311
rect 546 2283 662 2284
rect 580 2250 662 2283
rect 696 2250 796 2284
rect 580 2243 796 2250
rect 546 2216 796 2243
rect 546 2210 662 2216
rect 580 2182 662 2210
rect 696 2182 796 2216
rect 580 2175 796 2182
rect 546 2148 796 2175
rect 546 2141 662 2148
rect 580 2114 662 2141
rect 696 2114 796 2148
rect 580 2103 796 2114
rect 546 2080 796 2103
rect 546 2073 662 2080
rect 580 2046 662 2073
rect 696 2046 796 2080
rect 580 2030 796 2046
rect 546 2012 796 2030
rect 546 2005 662 2012
rect 580 1978 662 2005
rect 696 1978 796 2012
rect 580 1957 796 1978
rect 546 1944 796 1957
rect 546 1937 662 1944
rect 580 1910 662 1937
rect 696 1910 796 1944
rect 580 1884 796 1910
rect 546 1876 796 1884
rect 546 1869 662 1876
rect 580 1842 662 1869
rect 696 1842 796 1876
rect 580 1811 796 1842
rect 546 1808 796 1811
rect 546 1801 662 1808
rect 580 1774 662 1801
rect 696 1774 796 1808
rect 580 1740 796 1774
rect 580 1738 662 1740
rect 546 1733 662 1738
rect 580 1706 662 1733
rect 696 1706 796 1740
rect 580 1672 796 1706
rect 580 1638 662 1672
rect 696 1638 796 1672
rect 580 1631 796 1638
rect 546 1626 796 1631
rect 580 1604 796 1626
rect 580 1570 662 1604
rect 696 1570 796 1604
rect 580 1563 796 1570
rect 546 1553 796 1563
rect 580 1536 796 1553
rect 580 1502 662 1536
rect 696 1502 796 1536
rect 580 1495 796 1502
rect 546 1480 796 1495
rect 580 1468 796 1480
rect 580 1446 662 1468
rect 546 1434 662 1446
rect 696 1434 796 1468
rect 546 1407 796 1434
rect 404 1351 438 1362
rect 580 1400 796 1407
rect 580 1373 662 1400
rect 546 1366 662 1373
rect 696 1366 796 1400
rect 546 1351 796 1366
rect 404 1328 471 1351
rect 370 1292 471 1328
rect 404 1256 471 1292
rect 370 1224 471 1256
rect 404 1184 471 1224
rect 370 1156 471 1184
rect 404 1112 471 1156
rect 370 1088 471 1112
rect 404 1040 471 1088
rect 370 1020 471 1040
rect 404 968 471 1020
rect 370 952 471 968
rect 404 896 471 952
rect 370 884 471 896
rect 404 824 471 884
rect 370 816 471 824
rect 404 752 471 816
rect 370 748 471 752
rect 404 646 471 748
rect 370 642 471 646
rect 404 578 471 642
rect 370 570 471 578
rect 404 510 471 570
rect 370 498 471 510
rect 404 442 471 498
rect 370 426 471 442
rect 404 374 471 426
rect 370 358 471 374
rect 523 1334 796 1351
rect 523 1300 546 1334
rect 580 1332 796 1334
rect 580 1300 662 1332
rect 523 1298 662 1300
rect 696 1298 796 1332
rect 523 1292 796 1298
rect 523 1227 546 1292
rect 580 1264 796 1292
rect 580 1230 662 1264
rect 696 1230 796 1264
rect 580 1227 796 1230
rect 523 1224 796 1227
rect 523 1190 546 1224
rect 580 1196 796 1224
rect 580 1190 662 1196
rect 523 1188 662 1190
rect 523 1122 546 1188
rect 580 1162 662 1188
rect 696 1162 796 1196
rect 580 1128 796 1162
rect 580 1122 662 1128
rect 523 1115 662 1122
rect 523 1054 546 1115
rect 580 1094 662 1115
rect 696 1094 796 1128
rect 580 1060 796 1094
rect 580 1054 662 1060
rect 523 1042 662 1054
rect 523 986 546 1042
rect 580 1026 662 1042
rect 696 1026 796 1060
rect 580 992 796 1026
rect 580 986 662 992
rect 523 969 662 986
rect 523 918 546 969
rect 580 958 662 969
rect 696 958 796 992
rect 580 924 796 958
rect 580 918 662 924
rect 523 896 662 918
rect 523 850 546 896
rect 580 890 662 896
rect 696 890 796 924
rect 580 856 796 890
rect 580 850 662 856
rect 523 823 662 850
rect 523 782 546 823
rect 580 822 662 823
rect 696 822 796 856
rect 580 788 796 822
rect 580 782 662 788
rect 523 754 662 782
rect 696 754 796 788
rect 523 750 796 754
rect 523 714 546 750
rect 580 720 796 750
rect 580 714 662 720
rect 523 686 662 714
rect 696 686 796 720
rect 523 680 796 686
rect 523 643 546 680
rect 580 652 796 680
rect 580 643 662 652
rect 523 618 662 643
rect 696 618 796 652
rect 523 612 796 618
rect 523 570 546 612
rect 580 584 796 612
rect 580 570 662 584
rect 523 550 662 570
rect 696 550 796 584
rect 523 544 796 550
rect 523 496 546 544
rect 580 516 796 544
rect 580 496 662 516
rect 523 482 662 496
rect 696 482 796 516
rect 523 476 796 482
rect 523 422 546 476
rect 580 448 796 476
rect 580 422 662 448
rect 523 414 662 422
rect 696 414 796 448
rect 523 408 796 414
rect 259 346 318 347
rect 154 318 318 346
rect 523 348 546 408
rect 580 380 796 408
rect 580 348 662 380
rect 523 346 662 348
rect 696 346 796 380
rect 523 318 796 346
rect 154 312 796 318
rect 154 308 254 312
rect 288 308 796 312
rect 154 274 225 308
rect 288 278 306 308
rect 259 274 306 278
rect 340 288 386 308
rect 340 274 352 288
rect 154 254 352 274
rect 420 288 466 308
rect 500 288 546 308
rect 580 288 796 308
rect 420 274 423 288
rect 386 254 423 274
rect 457 274 466 288
rect 528 274 546 288
rect 457 254 494 274
rect 528 254 566 274
rect 600 254 638 288
rect 672 254 796 288
rect 154 153 796 254
rect -28 103 102 137
rect -44 101 102 103
rect 848 101 882 7217
rect -44 67 28 101
rect 62 67 106 101
rect 140 67 184 101
rect 237 67 262 101
rect 307 67 340 101
rect 378 67 415 101
rect 452 67 486 101
rect 530 67 557 101
rect 608 67 628 101
rect 686 67 699 101
rect 764 67 770 101
rect 804 67 808 101
rect 842 67 882 101
<< viali >>
rect 24 7217 58 7251
rect 96 7217 130 7251
rect 168 7217 185 7251
rect 185 7217 202 7251
rect 247 7217 261 7251
rect 261 7217 281 7251
rect 326 7217 337 7251
rect 337 7217 360 7251
rect 405 7217 413 7251
rect 413 7217 439 7251
rect 483 7217 488 7251
rect 488 7217 517 7251
rect 561 7217 563 7251
rect 563 7217 595 7251
rect 639 7217 672 7251
rect 672 7217 673 7251
rect 717 7217 747 7251
rect 747 7217 751 7251
rect 795 7217 829 7251
rect -62 7181 -28 7215
rect -62 7109 -28 7143
rect -62 7037 -28 7071
rect -62 6965 -28 6999
rect -62 6893 -28 6927
rect -62 6821 -28 6855
rect -62 6749 -28 6783
rect -62 6677 -28 6711
rect -62 6605 -28 6639
rect -62 6533 -28 6567
rect -62 6461 -28 6495
rect -62 6389 -28 6423
rect -62 6317 -28 6351
rect -62 6245 -28 6279
rect -62 6173 -28 6207
rect -62 6101 -28 6135
rect -62 6029 -28 6063
rect -62 5957 -28 5991
rect -62 5885 -28 5919
rect -62 5813 -28 5847
rect -62 5741 -28 5775
rect -62 5669 -28 5703
rect -62 5597 -28 5631
rect -62 5525 -28 5559
rect -62 5453 -28 5487
rect -62 5381 -28 5415
rect -62 5309 -28 5343
rect -62 5237 -28 5271
rect -62 5165 -28 5199
rect -62 5093 -28 5127
rect -62 5021 -28 5055
rect -62 4949 -28 4983
rect -62 4877 -28 4911
rect -62 4805 -28 4839
rect -62 4733 -28 4767
rect -62 4661 -28 4695
rect -62 4589 -28 4623
rect -62 4517 -28 4551
rect -62 4445 -28 4479
rect -62 4373 -28 4407
rect -62 4301 -28 4335
rect -62 4229 -28 4263
rect -62 4157 -28 4191
rect -62 4085 -28 4119
rect -62 4013 -28 4047
rect -62 3941 -28 3975
rect -62 3869 -28 3903
rect -62 3797 -28 3831
rect -62 3725 -28 3759
rect -62 3653 -28 3687
rect -62 3581 -28 3615
rect -62 3509 -28 3543
rect -62 3437 -28 3471
rect -62 3365 -28 3399
rect -62 3293 -28 3327
rect -62 3221 -28 3255
rect -62 3149 -28 3183
rect -62 3077 -28 3111
rect -62 3005 -28 3039
rect -62 2933 -28 2967
rect -62 2861 -28 2895
rect -62 2789 -28 2823
rect -62 2717 -28 2751
rect -62 2645 -28 2679
rect -62 2573 -28 2607
rect -62 2501 -28 2535
rect -62 2429 -28 2463
rect -62 2357 -28 2391
rect -62 2285 -28 2319
rect -62 2213 -28 2247
rect -62 2141 -28 2175
rect -62 2069 -28 2103
rect -62 1997 -28 2031
rect -62 1925 -28 1959
rect -62 1853 -28 1887
rect -62 1781 -28 1815
rect -62 1709 -28 1743
rect -62 1636 -28 1670
rect -62 1563 -28 1597
rect -62 1490 -28 1524
rect -62 1417 -28 1451
rect -62 1344 -28 1378
rect -62 1271 -28 1305
rect -62 1198 -28 1232
rect -62 1125 -28 1159
rect -62 1052 -28 1086
rect -62 979 -28 1013
rect -62 906 -28 940
rect -62 833 -28 867
rect -62 760 -28 794
rect -62 687 -28 721
rect -62 614 -28 648
rect -62 541 -28 575
rect -62 468 -28 502
rect -62 395 -28 429
rect -62 322 -28 356
rect -62 249 -28 283
rect -62 176 -28 210
rect 225 7021 259 7055
rect 305 7030 312 7055
rect 312 7030 339 7055
rect 305 7021 339 7030
rect 385 7030 391 7055
rect 391 7030 419 7055
rect 385 7021 419 7030
rect 465 7021 499 7055
rect 546 7030 559 7055
rect 559 7030 580 7055
rect 546 7021 580 7030
rect 225 6972 259 6982
rect 225 6948 254 6972
rect 254 6948 259 6972
rect 225 6904 259 6909
rect 225 6875 254 6904
rect 254 6875 259 6904
rect 225 6802 254 6836
rect 254 6802 259 6836
rect 225 6734 254 6763
rect 254 6734 259 6763
rect 225 6729 259 6734
rect 225 6666 254 6690
rect 254 6666 259 6690
rect 225 6656 259 6666
rect 225 6598 254 6617
rect 254 6598 259 6617
rect 225 6583 259 6598
rect 225 6530 254 6544
rect 254 6530 259 6544
rect 225 6510 259 6530
rect 225 6462 254 6471
rect 254 6462 259 6471
rect 225 6437 259 6462
rect 225 6394 254 6398
rect 254 6394 259 6398
rect 225 6364 259 6394
rect 225 6292 259 6325
rect 225 6291 254 6292
rect 254 6291 259 6292
rect 225 6224 259 6252
rect 225 6218 254 6224
rect 254 6218 259 6224
rect 225 6156 259 6179
rect 225 6145 254 6156
rect 254 6145 259 6156
rect 225 6088 259 6106
rect 225 6072 254 6088
rect 254 6072 259 6088
rect 225 6020 259 6033
rect 225 5999 254 6020
rect 254 5999 259 6020
rect 225 5952 259 5960
rect 225 5926 254 5952
rect 254 5926 259 5952
rect 225 5884 259 5887
rect 225 5853 254 5884
rect 254 5853 259 5884
rect 225 5782 254 5814
rect 254 5782 259 5814
rect 225 5780 259 5782
rect 225 5714 254 5741
rect 254 5714 259 5741
rect 225 5707 259 5714
rect 225 5646 254 5668
rect 254 5646 259 5668
rect 225 5634 259 5646
rect 225 5578 254 5595
rect 254 5578 259 5595
rect 225 5561 259 5578
rect 225 5510 254 5522
rect 254 5510 259 5522
rect 225 5488 259 5510
rect 225 5442 254 5449
rect 254 5442 259 5449
rect 225 5415 259 5442
rect 225 5374 254 5376
rect 254 5374 259 5376
rect 225 5342 259 5374
rect 225 5272 259 5303
rect 225 5269 254 5272
rect 254 5269 259 5272
rect 225 5204 259 5230
rect 225 5196 254 5204
rect 254 5196 259 5204
rect 225 5136 259 5157
rect 225 5123 254 5136
rect 254 5123 259 5136
rect 225 5068 259 5084
rect 225 5050 254 5068
rect 254 5050 259 5068
rect 225 5000 259 5011
rect 225 4977 254 5000
rect 254 4977 259 5000
rect 225 4932 259 4938
rect 225 4904 254 4932
rect 254 4904 259 4932
rect 225 4864 259 4865
rect 225 4831 254 4864
rect 254 4831 259 4864
rect 225 4762 254 4792
rect 254 4762 259 4792
rect 225 4758 259 4762
rect 225 4694 254 4719
rect 254 4694 259 4719
rect 225 4685 259 4694
rect 225 4625 254 4646
rect 254 4625 259 4646
rect 225 4612 259 4625
rect 225 4556 254 4573
rect 254 4556 259 4573
rect 225 4539 259 4556
rect 225 4487 254 4500
rect 254 4487 259 4500
rect 225 4466 259 4487
rect 225 4418 254 4427
rect 254 4418 259 4427
rect 225 4393 259 4418
rect 225 4349 254 4354
rect 254 4349 259 4354
rect 225 4320 259 4349
rect 225 4280 254 4281
rect 254 4280 259 4281
rect 225 4247 259 4280
rect 225 4176 259 4208
rect 225 4174 254 4176
rect 254 4174 259 4176
rect 225 4107 259 4135
rect 225 4101 254 4107
rect 254 4101 259 4107
rect 225 4038 259 4062
rect 225 4028 254 4038
rect 254 4028 259 4038
rect 225 3969 259 3989
rect 225 3955 254 3969
rect 254 3955 259 3969
rect 225 3900 259 3916
rect 225 3882 254 3900
rect 254 3882 259 3900
rect 225 3831 259 3843
rect 225 3809 254 3831
rect 254 3809 259 3831
rect 225 3762 259 3770
rect 225 3736 254 3762
rect 254 3736 259 3762
rect 225 3693 259 3697
rect 225 3663 254 3693
rect 254 3663 259 3693
rect 225 3590 254 3624
rect 254 3590 259 3624
rect 225 3521 254 3551
rect 254 3521 259 3551
rect 225 3517 259 3521
rect 225 3452 254 3478
rect 254 3452 259 3478
rect 225 3444 259 3452
rect 225 3383 254 3405
rect 254 3383 259 3405
rect 225 3371 259 3383
rect 225 3314 254 3332
rect 254 3314 259 3332
rect 225 3298 259 3314
rect 225 3245 254 3260
rect 254 3245 259 3260
rect 225 3226 259 3245
rect 225 3176 254 3188
rect 254 3176 259 3188
rect 225 3154 259 3176
rect 225 3107 254 3116
rect 254 3107 259 3116
rect 225 3082 259 3107
rect 225 3038 254 3044
rect 254 3038 259 3044
rect 225 3010 259 3038
rect 225 2969 254 2972
rect 254 2969 259 2972
rect 225 2938 259 2969
rect 225 2866 259 2900
rect 225 2796 259 2828
rect 225 2794 254 2796
rect 254 2794 259 2796
rect 225 2727 259 2756
rect 225 2722 254 2727
rect 254 2722 259 2727
rect 225 2658 259 2684
rect 225 2650 254 2658
rect 254 2650 259 2658
rect 225 2589 259 2612
rect 225 2578 254 2589
rect 254 2578 259 2589
rect 225 2520 259 2540
rect 225 2506 254 2520
rect 254 2506 259 2520
rect 225 2451 259 2468
rect 225 2434 254 2451
rect 254 2434 259 2451
rect 225 2382 259 2396
rect 225 2362 254 2382
rect 254 2362 259 2382
rect 225 2313 259 2324
rect 225 2290 254 2313
rect 254 2290 259 2313
rect 225 2244 259 2252
rect 225 2218 254 2244
rect 254 2218 259 2244
rect 225 2175 259 2180
rect 225 2146 254 2175
rect 254 2146 259 2175
rect 225 2106 259 2108
rect 225 2074 254 2106
rect 254 2074 259 2106
rect 225 2003 254 2036
rect 254 2003 259 2036
rect 225 2002 259 2003
rect 225 1934 254 1964
rect 254 1934 259 1964
rect 225 1930 259 1934
rect 225 1865 254 1892
rect 254 1865 259 1892
rect 225 1858 259 1865
rect 225 1796 254 1820
rect 254 1796 259 1820
rect 225 1786 259 1796
rect 225 1727 254 1748
rect 254 1727 259 1748
rect 225 1714 259 1727
rect 225 1658 254 1676
rect 254 1658 259 1676
rect 225 1642 259 1658
rect 225 1589 254 1604
rect 254 1589 259 1604
rect 225 1570 259 1589
rect 225 1520 254 1532
rect 254 1520 259 1532
rect 225 1498 259 1520
rect 225 1451 254 1460
rect 254 1451 259 1460
rect 225 1426 259 1451
rect 225 1382 254 1388
rect 254 1382 259 1388
rect 225 1354 259 1382
rect 225 1313 254 1316
rect 254 1313 259 1316
rect 225 1282 259 1313
rect 225 1210 259 1244
rect 225 1140 259 1172
rect 225 1138 254 1140
rect 254 1138 259 1140
rect 225 1071 259 1100
rect 225 1066 254 1071
rect 254 1066 259 1071
rect 225 1002 259 1028
rect 225 994 254 1002
rect 254 994 259 1002
rect 225 933 259 956
rect 225 922 254 933
rect 254 922 259 933
rect 225 864 259 884
rect 225 850 254 864
rect 254 850 259 864
rect 225 795 259 812
rect 225 778 254 795
rect 254 778 259 795
rect 225 726 259 740
rect 225 706 254 726
rect 254 706 259 726
rect 225 657 259 668
rect 225 634 254 657
rect 254 634 259 657
rect 225 588 259 596
rect 225 562 254 588
rect 254 562 259 588
rect 225 519 259 524
rect 225 490 254 519
rect 254 490 259 519
rect 225 450 259 452
rect 225 418 254 450
rect 254 418 259 450
rect 225 347 254 380
rect 254 347 259 380
rect 370 6876 404 6892
rect 370 6858 404 6876
rect 370 6808 404 6819
rect 370 6785 404 6808
rect 370 6740 404 6746
rect 370 6712 404 6740
rect 370 6672 404 6673
rect 370 6639 404 6672
rect 370 6570 404 6600
rect 370 6566 404 6570
rect 370 6502 404 6527
rect 370 6493 404 6502
rect 370 6434 404 6454
rect 370 6420 404 6434
rect 370 6366 404 6381
rect 370 6347 404 6366
rect 370 6298 404 6308
rect 370 6274 404 6298
rect 370 6230 404 6235
rect 370 6201 404 6230
rect 370 6128 404 6162
rect 370 6060 404 6089
rect 370 6055 404 6060
rect 370 5982 404 6016
rect 546 6948 580 6982
rect 546 6876 580 6909
rect 546 6875 580 6876
rect 546 6808 580 6836
rect 546 6802 580 6808
rect 546 6740 580 6763
rect 546 6729 580 6740
rect 546 6672 580 6690
rect 546 6656 580 6672
rect 546 6604 580 6617
rect 546 6583 580 6604
rect 546 6536 580 6544
rect 546 6510 580 6536
rect 546 6468 580 6471
rect 546 6437 580 6468
rect 546 6366 580 6398
rect 546 6364 580 6366
rect 546 6298 580 6325
rect 546 6291 580 6298
rect 546 6230 580 6252
rect 546 6218 580 6230
rect 546 6162 580 6179
rect 546 6145 580 6162
rect 546 6094 580 6106
rect 546 6072 580 6094
rect 546 6026 580 6033
rect 546 5999 580 6026
rect 370 5909 404 5943
rect 370 5836 404 5870
rect 370 5789 404 5797
rect 370 5763 404 5789
rect 370 5721 404 5724
rect 370 5690 404 5721
rect 370 5619 404 5651
rect 370 5617 404 5619
rect 370 5551 404 5578
rect 370 5544 404 5551
rect 370 5483 404 5505
rect 370 5471 404 5483
rect 370 5415 404 5432
rect 370 5398 404 5415
rect 370 5347 404 5359
rect 370 5325 404 5347
rect 370 5279 404 5286
rect 370 5252 404 5279
rect 370 5211 404 5213
rect 370 5179 404 5211
rect 370 5109 404 5140
rect 370 5106 404 5109
rect 370 5041 404 5067
rect 370 5033 404 5041
rect 370 4973 404 4994
rect 370 4960 404 4973
rect 370 4905 404 4921
rect 370 4887 404 4905
rect 370 4814 404 4848
rect 370 4741 404 4775
rect 370 4668 404 4702
rect 370 4600 404 4629
rect 370 4595 404 4600
rect 370 4532 404 4556
rect 370 4522 404 4532
rect 370 4464 404 4483
rect 370 4449 404 4464
rect 370 4396 404 4410
rect 370 4376 404 4396
rect 370 4328 404 4337
rect 370 4303 404 4328
rect 370 4260 404 4264
rect 370 4230 404 4260
rect 370 4158 404 4191
rect 370 4157 404 4158
rect 370 4090 404 4118
rect 370 4084 404 4090
rect 370 4022 404 4045
rect 370 4011 404 4022
rect 370 3954 404 3972
rect 370 3938 404 3954
rect 370 3886 404 3899
rect 370 3865 404 3886
rect 370 3818 404 3826
rect 370 3792 404 3818
rect 370 3719 404 3753
rect 370 3646 404 3680
rect 370 3573 404 3607
rect 370 3500 404 3534
rect 370 3432 404 3461
rect 370 3427 404 3432
rect 370 3364 404 3388
rect 370 3354 404 3364
rect 370 3296 404 3315
rect 370 3281 404 3296
rect 370 3228 404 3241
rect 370 3207 404 3228
rect 370 3160 404 3163
rect 370 3129 404 3160
rect 370 3058 404 3090
rect 370 3056 404 3058
rect 370 2990 404 3018
rect 370 2984 404 2990
rect 370 2922 404 2946
rect 370 2912 404 2922
rect 370 2854 404 2874
rect 370 2840 404 2854
rect 370 2786 404 2802
rect 370 2768 404 2786
rect 370 2718 404 2730
rect 370 2696 404 2718
rect 370 2650 404 2658
rect 370 2624 404 2650
rect 370 2552 404 2586
rect 370 2480 404 2514
rect 370 2413 404 2442
rect 370 2408 404 2413
rect 370 2345 404 2370
rect 370 2336 404 2345
rect 370 2277 404 2298
rect 370 2264 404 2277
rect 370 2209 404 2226
rect 370 2192 404 2209
rect 370 2141 404 2154
rect 370 2120 404 2141
rect 370 2073 404 2082
rect 370 2048 404 2073
rect 370 2005 404 2010
rect 370 1976 404 2005
rect 370 1937 404 1938
rect 370 1904 404 1937
rect 370 1835 404 1866
rect 370 1832 404 1835
rect 370 1767 404 1794
rect 370 1760 404 1767
rect 370 1699 404 1722
rect 370 1688 404 1699
rect 370 1631 404 1650
rect 370 1616 404 1631
rect 370 1563 404 1578
rect 370 1544 404 1563
rect 370 1495 404 1506
rect 370 1472 404 1495
rect 370 1400 404 1434
rect 472 5916 506 5922
rect 472 5888 506 5916
rect 472 5815 506 5849
rect 472 5742 506 5776
rect 472 5669 506 5703
rect 472 5596 506 5630
rect 472 5523 506 5557
rect 472 5450 506 5484
rect 472 5377 506 5411
rect 472 5304 506 5338
rect 472 5231 506 5265
rect 472 5158 506 5192
rect 472 5085 506 5119
rect 472 5012 506 5046
rect 472 4939 506 4973
rect 472 4866 506 4900
rect 472 4795 506 4827
rect 472 4793 506 4795
rect 472 4720 506 4754
rect 472 4647 506 4681
rect 472 4574 506 4608
rect 472 4501 506 4535
rect 472 4427 506 4461
rect 472 4353 506 4387
rect 472 4279 506 4313
rect 472 4205 506 4239
rect 472 4131 506 4165
rect 472 4057 506 4091
rect 472 3983 506 4017
rect 472 3909 506 3943
rect 472 3835 506 3869
rect 472 3761 506 3795
rect 472 3687 506 3721
rect 472 3642 506 3647
rect 472 3613 506 3642
rect 472 3538 506 3572
rect 472 3464 506 3498
rect 472 3390 506 3424
rect 472 3316 506 3350
rect 472 3242 506 3276
rect 472 3168 506 3202
rect 472 3094 506 3128
rect 472 3020 506 3054
rect 472 2946 506 2980
rect 472 2872 506 2906
rect 472 2798 506 2832
rect 472 2724 506 2758
rect 472 2650 506 2684
rect 472 2576 506 2610
rect 472 2522 506 2536
rect 472 2502 506 2522
rect 472 2428 506 2462
rect 472 2354 506 2388
rect 472 2280 506 2314
rect 472 2207 506 2241
rect 472 2134 506 2168
rect 472 2061 506 2095
rect 472 1988 506 2022
rect 472 1915 506 1949
rect 472 1842 506 1876
rect 472 1769 506 1803
rect 472 1696 506 1730
rect 472 1623 506 1657
rect 472 1550 506 1584
rect 472 1477 506 1511
rect 546 5926 580 5960
rect 546 5853 580 5887
rect 546 5789 580 5814
rect 546 5780 580 5789
rect 546 5721 580 5741
rect 546 5707 580 5721
rect 546 5653 580 5668
rect 546 5634 580 5653
rect 546 5585 580 5595
rect 546 5561 580 5585
rect 546 5517 580 5522
rect 546 5488 580 5517
rect 546 5415 580 5449
rect 546 5347 580 5376
rect 546 5342 580 5347
rect 546 5279 580 5303
rect 546 5269 580 5279
rect 546 5211 580 5230
rect 546 5196 580 5211
rect 546 5143 580 5157
rect 546 5123 580 5143
rect 546 5075 580 5084
rect 546 5050 580 5075
rect 546 5007 580 5011
rect 546 4977 580 5007
rect 546 4905 580 4938
rect 546 4904 580 4905
rect 546 4831 580 4865
rect 546 4758 580 4792
rect 546 4702 580 4719
rect 546 4685 580 4702
rect 546 4634 580 4646
rect 546 4612 580 4634
rect 546 4566 580 4573
rect 546 4539 580 4566
rect 546 4498 580 4500
rect 546 4466 580 4498
rect 546 4396 580 4426
rect 546 4392 580 4396
rect 546 4328 580 4352
rect 546 4318 580 4328
rect 546 4260 580 4278
rect 546 4244 580 4260
rect 546 4192 580 4204
rect 546 4170 580 4192
rect 546 4124 580 4130
rect 546 4096 580 4124
rect 546 4022 580 4056
rect 546 3954 580 3982
rect 546 3948 580 3954
rect 546 3886 580 3908
rect 546 3874 580 3886
rect 546 3818 580 3834
rect 546 3800 580 3818
rect 546 3726 580 3760
rect 546 3636 580 3670
rect 546 3563 580 3597
rect 546 3500 580 3524
rect 546 3490 580 3500
rect 546 3432 580 3451
rect 546 3417 580 3432
rect 546 3364 580 3378
rect 546 3344 580 3364
rect 546 3296 580 3305
rect 546 3271 580 3296
rect 546 3228 580 3232
rect 546 3198 580 3228
rect 546 3126 580 3159
rect 546 3125 580 3126
rect 546 3058 580 3086
rect 546 3052 580 3058
rect 546 2990 580 3013
rect 546 2979 580 2990
rect 546 2922 580 2940
rect 546 2906 580 2922
rect 546 2854 580 2867
rect 546 2833 580 2854
rect 546 2786 580 2794
rect 546 2760 580 2786
rect 546 2718 580 2721
rect 546 2687 580 2718
rect 546 2616 580 2648
rect 546 2614 580 2616
rect 546 2541 580 2575
rect 546 2468 580 2502
rect 546 2413 580 2429
rect 546 2395 580 2413
rect 546 2345 580 2356
rect 546 2322 580 2345
rect 546 2277 580 2283
rect 546 2249 580 2277
rect 546 2209 580 2210
rect 546 2176 580 2209
rect 546 2107 580 2137
rect 546 2103 580 2107
rect 546 2039 580 2064
rect 546 2030 580 2039
rect 546 1971 580 1991
rect 546 1957 580 1971
rect 546 1903 580 1918
rect 546 1884 580 1903
rect 546 1835 580 1845
rect 546 1811 580 1835
rect 546 1767 580 1772
rect 546 1738 580 1767
rect 546 1665 580 1699
rect 546 1597 580 1626
rect 546 1592 580 1597
rect 546 1529 580 1553
rect 546 1519 580 1529
rect 546 1446 580 1480
rect 370 1328 404 1362
rect 546 1373 580 1407
rect 370 1258 404 1290
rect 370 1256 404 1258
rect 370 1190 404 1218
rect 370 1184 404 1190
rect 370 1122 404 1146
rect 370 1112 404 1122
rect 370 1054 404 1074
rect 370 1040 404 1054
rect 370 986 404 1002
rect 370 968 404 986
rect 370 918 404 930
rect 370 896 404 918
rect 370 850 404 858
rect 370 824 404 850
rect 370 782 404 786
rect 370 752 404 782
rect 370 680 404 714
rect 370 612 404 642
rect 370 608 404 612
rect 370 544 404 570
rect 370 536 404 544
rect 370 476 404 498
rect 370 464 404 476
rect 370 408 404 426
rect 370 392 404 408
rect 546 1300 580 1334
rect 546 1258 580 1261
rect 546 1227 580 1258
rect 546 1156 580 1188
rect 546 1154 580 1156
rect 546 1088 580 1115
rect 546 1081 580 1088
rect 546 1020 580 1042
rect 546 1008 580 1020
rect 546 952 580 969
rect 546 935 580 952
rect 546 884 580 896
rect 546 862 580 884
rect 546 816 580 823
rect 546 789 580 816
rect 546 748 580 750
rect 546 716 580 748
rect 546 646 580 677
rect 546 643 580 646
rect 546 578 580 604
rect 546 570 580 578
rect 546 510 580 530
rect 546 496 580 510
rect 546 442 580 456
rect 546 422 580 442
rect 225 346 259 347
rect 546 374 580 382
rect 546 348 580 374
rect 225 278 254 308
rect 254 278 259 308
rect 225 274 259 278
rect 306 274 340 308
rect 386 274 420 308
rect 466 288 500 308
rect 546 288 580 308
rect 466 274 494 288
rect 494 274 500 288
rect 546 274 566 288
rect 566 274 580 288
rect -62 103 -28 137
rect 28 67 62 101
rect 106 67 140 101
rect 184 67 203 101
rect 203 67 218 101
rect 262 67 273 101
rect 273 67 296 101
rect 340 67 344 101
rect 344 67 374 101
rect 418 67 449 101
rect 449 67 452 101
rect 496 67 520 101
rect 520 67 530 101
rect 574 67 591 101
rect 591 67 608 101
rect 652 67 662 101
rect 662 67 686 101
rect 730 67 733 101
rect 733 67 764 101
rect 808 67 842 101
<< metal1 >>
tri 798 7257 886 7345 se
rect 12 7251 886 7257
rect -68 7215 -22 7227
rect -68 7181 -62 7215
rect -28 7181 -22 7215
rect 12 7217 24 7251
rect 58 7217 96 7251
rect 130 7217 168 7251
rect 202 7217 247 7251
rect 281 7217 326 7251
rect 360 7217 405 7251
rect 439 7217 483 7251
rect 517 7217 561 7251
rect 595 7217 639 7251
rect 673 7217 717 7251
rect 751 7217 795 7251
rect 829 7217 886 7251
rect 12 7211 886 7217
rect -68 7143 -22 7181
rect -68 7109 -62 7143
rect -28 7109 -22 7143
tri -22 7137 52 7211 nw
tri 806 7137 880 7211 ne
rect 880 7137 886 7211
tri 880 7131 886 7137 ne
rect -68 7071 -22 7109
rect -68 7037 -62 7071
rect -28 7037 -22 7071
rect -68 6999 -22 7037
rect -68 6965 -62 6999
rect -28 6965 -22 6999
rect -68 6927 -22 6965
rect -68 6893 -62 6927
rect -28 6893 -22 6927
rect -68 6855 -22 6893
rect 195 7055 604 7123
rect 195 7021 225 7055
rect 259 7021 305 7055
rect 339 7021 385 7055
rect 419 7021 465 7055
rect 499 7021 546 7055
rect 580 7021 604 7055
rect 195 7015 604 7021
rect 195 7008 299 7015
tri 299 7008 306 7015 nw
tri 500 7009 506 7015 ne
rect 506 7009 604 7015
tri 506 7008 507 7009 ne
rect 507 7008 604 7009
rect 195 7001 292 7008
tri 292 7001 299 7008 nw
tri 507 7003 512 7008 ne
rect 512 7003 604 7008
tri 512 7001 514 7003 ne
rect 514 7001 604 7003
rect 195 6995 286 7001
tri 286 6995 292 7001 nw
tri 514 6997 518 7001 ne
rect 518 6997 604 7001
tri 518 6995 520 6997 ne
rect 520 6995 604 6997
rect 195 6988 279 6995
tri 279 6988 286 6995 nw
tri 520 6993 522 6995 ne
rect 522 6993 604 6995
tri 522 6988 527 6993 ne
rect 527 6988 604 6993
rect 195 6982 273 6988
tri 273 6982 279 6988 nw
tri 527 6987 528 6988 ne
rect 528 6987 604 6988
tri 528 6982 533 6987 ne
rect 533 6982 604 6987
rect 195 6948 225 6982
rect 259 6981 272 6982
tri 272 6981 273 6982 nw
tri 533 6981 534 6982 ne
rect 534 6981 546 6982
rect 259 6975 266 6981
tri 266 6975 272 6981 nw
tri 534 6975 540 6981 ne
rect 259 6948 265 6975
tri 265 6974 266 6975 nw
rect 195 6909 265 6948
rect 195 6882 225 6909
tri 195 6875 202 6882 ne
rect 202 6875 225 6882
rect 259 6875 265 6909
rect 540 6948 546 6981
rect 580 6948 604 6982
rect 540 6909 604 6948
tri 202 6864 213 6875 ne
rect 213 6864 265 6875
tri 213 6858 219 6864 ne
rect -68 6821 -62 6855
rect -28 6821 -22 6855
rect -68 6783 -22 6821
rect -68 6749 -62 6783
rect -28 6749 -22 6783
rect -68 6711 -22 6749
rect -68 6677 -62 6711
rect -28 6677 -22 6711
rect -68 6639 -22 6677
rect -68 6605 -62 6639
rect -28 6605 -22 6639
rect -68 6567 -22 6605
rect -68 6533 -62 6567
rect -28 6533 -22 6567
rect -68 6495 -22 6533
rect -68 6461 -62 6495
rect -28 6461 -22 6495
rect -68 6423 -22 6461
rect -68 6389 -62 6423
rect -28 6389 -22 6423
rect -68 6351 -22 6389
rect -68 6317 -62 6351
rect -28 6317 -22 6351
rect -68 6279 -22 6317
rect -68 6245 -62 6279
rect -28 6245 -22 6279
rect -68 6207 -22 6245
rect -68 6173 -62 6207
rect -28 6173 -22 6207
rect -68 6135 -22 6173
rect -68 6101 -62 6135
rect -28 6101 -22 6135
rect -68 6063 -22 6101
rect -68 6029 -62 6063
rect -28 6029 -22 6063
rect 219 6836 265 6864
rect 219 6802 225 6836
rect 259 6802 265 6836
rect 219 6763 265 6802
rect 219 6729 225 6763
rect 259 6729 265 6763
rect 219 6690 265 6729
rect 219 6656 225 6690
rect 259 6656 265 6690
rect 219 6617 265 6656
rect 219 6583 225 6617
rect 259 6583 265 6617
rect 219 6544 265 6583
rect 219 6510 225 6544
rect 259 6510 265 6544
rect 219 6471 265 6510
rect 219 6437 225 6471
rect 259 6437 265 6471
rect 219 6398 265 6437
rect 219 6364 225 6398
rect 259 6364 265 6398
rect 219 6325 265 6364
rect 219 6291 225 6325
rect 259 6291 265 6325
rect 219 6252 265 6291
rect 219 6218 225 6252
rect 259 6218 265 6252
rect 219 6179 265 6218
rect 219 6145 225 6179
rect 259 6145 265 6179
rect 219 6106 265 6145
rect 219 6072 225 6106
rect 259 6072 265 6106
tri 218 6055 219 6056 se
rect 219 6055 265 6072
rect -68 5991 -22 6029
rect -68 5957 -62 5991
rect -28 5957 -22 5991
rect -68 5919 -22 5957
rect -68 5885 -62 5919
rect -28 5885 -22 5919
rect -68 5847 -22 5885
rect -68 5813 -62 5847
rect -28 5813 -22 5847
rect -68 5775 -22 5813
rect -68 5741 -62 5775
rect -28 5741 -22 5775
rect -68 5703 -22 5741
tri 213 6050 218 6055 se
rect 218 6050 265 6055
rect 213 6044 265 6050
rect 213 5962 265 5992
rect 213 5887 265 5910
rect 213 5880 225 5887
rect 259 5880 265 5887
rect 213 5814 265 5828
rect 213 5798 225 5814
rect 259 5798 265 5814
rect 213 5741 265 5746
rect 213 5740 225 5741
tri 213 5734 219 5740 ne
rect -68 5669 -62 5703
rect -28 5669 -22 5703
rect -68 5631 -22 5669
rect -68 5597 -62 5631
rect -28 5597 -22 5631
rect -68 5559 -22 5597
rect -68 5525 -62 5559
rect -28 5525 -22 5559
rect -68 5487 -22 5525
rect -68 5453 -62 5487
rect -28 5453 -22 5487
rect -68 5415 -22 5453
rect -68 5381 -62 5415
rect -28 5381 -22 5415
rect -68 5343 -22 5381
rect -68 5309 -62 5343
rect -28 5309 -22 5343
rect -68 5271 -22 5309
rect -68 5237 -62 5271
rect -28 5237 -22 5271
rect -68 5199 -22 5237
rect -68 5165 -62 5199
rect -28 5165 -22 5199
rect -68 5127 -22 5165
rect -68 5093 -62 5127
rect -28 5093 -22 5127
rect -68 5055 -22 5093
rect -68 5021 -62 5055
rect -28 5021 -22 5055
rect -68 4983 -22 5021
rect -68 4949 -62 4983
rect -28 4949 -22 4983
rect -68 4911 -22 4949
rect -68 4877 -62 4911
rect -28 4877 -22 4911
rect -68 4839 -22 4877
rect -68 4805 -62 4839
rect -28 4805 -22 4839
rect -68 4767 -22 4805
rect -68 4733 -62 4767
rect -28 4733 -22 4767
rect -68 4695 -22 4733
rect -68 4661 -62 4695
rect -28 4661 -22 4695
rect -68 4623 -22 4661
rect -68 4589 -62 4623
rect -28 4589 -22 4623
rect -68 4551 -22 4589
rect -68 4517 -62 4551
rect -28 4517 -22 4551
rect -68 4479 -22 4517
rect -68 4445 -62 4479
rect -28 4445 -22 4479
rect -68 4407 -22 4445
rect -68 4373 -62 4407
rect -28 4373 -22 4407
rect -68 4335 -22 4373
rect -68 4301 -62 4335
rect -28 4301 -22 4335
rect -68 4263 -22 4301
rect -68 4229 -62 4263
rect -28 4229 -22 4263
rect -68 4191 -22 4229
rect -68 4157 -62 4191
rect -28 4157 -22 4191
rect -68 4119 -22 4157
rect -68 4085 -62 4119
rect -28 4085 -22 4119
rect -68 4047 -22 4085
rect -68 4013 -62 4047
rect -28 4013 -22 4047
rect 219 5707 225 5740
rect 259 5707 265 5741
rect 219 5668 265 5707
rect 219 5634 225 5668
rect 259 5634 265 5668
rect 219 5595 265 5634
rect 219 5561 225 5595
rect 259 5561 265 5595
rect 219 5522 265 5561
rect 219 5488 225 5522
rect 259 5488 265 5522
rect 219 5449 265 5488
rect 219 5415 225 5449
rect 259 5415 265 5449
rect 219 5376 265 5415
rect 219 5342 225 5376
rect 259 5342 265 5376
rect 219 5303 265 5342
rect 219 5269 225 5303
rect 259 5269 265 5303
rect 219 5230 265 5269
rect 219 5196 225 5230
rect 259 5196 265 5230
rect 219 5157 265 5196
rect 219 5123 225 5157
rect 259 5123 265 5157
rect 219 5084 265 5123
rect 219 5050 225 5084
rect 259 5050 265 5084
rect 219 5011 265 5050
rect 219 4977 225 5011
rect 259 4977 265 5011
rect 219 4938 265 4977
rect 219 4904 225 4938
rect 259 4904 265 4938
rect 219 4865 265 4904
rect 219 4831 225 4865
rect 259 4831 265 4865
rect 219 4792 265 4831
rect 219 4758 225 4792
rect 259 4758 265 4792
rect 219 4719 265 4758
rect 219 4685 225 4719
rect 259 4685 265 4719
rect 219 4646 265 4685
rect 219 4612 225 4646
rect 259 4612 265 4646
rect 219 4573 265 4612
rect 219 4539 225 4573
rect 259 4539 265 4573
rect 219 4500 265 4539
rect 219 4466 225 4500
rect 259 4466 265 4500
rect 219 4427 265 4466
rect 219 4393 225 4427
rect 259 4393 265 4427
rect 219 4354 265 4393
rect 219 4320 225 4354
rect 259 4320 265 4354
rect 219 4281 265 4320
rect 219 4247 225 4281
rect 259 4247 265 4281
rect 219 4208 265 4247
rect 219 4174 225 4208
rect 259 4174 265 4208
rect 219 4135 265 4174
rect 219 4101 225 4135
rect 259 4101 265 4135
rect 219 4062 265 4101
tri 217 4028 219 4030 se
rect 219 4028 225 4062
rect 259 4028 265 4062
rect -68 3975 -22 4013
rect -68 3941 -62 3975
rect -28 3941 -22 3975
rect -68 3903 -22 3941
rect -68 3869 -62 3903
rect -28 3869 -22 3903
rect -68 3831 -22 3869
rect -68 3797 -62 3831
rect -28 3797 -22 3831
rect -68 3759 -22 3797
rect -68 3725 -62 3759
rect -28 3725 -22 3759
rect -68 3687 -22 3725
tri 213 4024 217 4028 se
rect 217 4024 265 4028
rect 213 4018 265 4024
rect 213 3955 225 3966
rect 259 3955 265 3966
rect 213 3936 265 3955
rect 213 3882 225 3884
rect 259 3882 265 3884
rect 213 3854 265 3882
rect 213 3772 265 3802
rect 213 3714 265 3720
tri 213 3708 219 3714 ne
rect -68 3653 -62 3687
rect -28 3653 -22 3687
rect -68 3615 -22 3653
rect -68 3581 -62 3615
rect -28 3581 -22 3615
rect -68 3543 -22 3581
rect -68 3509 -62 3543
rect -28 3509 -22 3543
rect -68 3471 -22 3509
rect -68 3437 -62 3471
rect -28 3437 -22 3471
rect -68 3399 -22 3437
rect -68 3365 -62 3399
rect -28 3365 -22 3399
rect -68 3327 -22 3365
rect -68 3293 -62 3327
rect -28 3293 -22 3327
rect -68 3255 -22 3293
rect -68 3221 -62 3255
rect -28 3221 -22 3255
rect -68 3183 -22 3221
rect -68 3149 -62 3183
rect -28 3149 -22 3183
rect -68 3111 -22 3149
rect -68 3077 -62 3111
rect -28 3077 -22 3111
rect -68 3039 -22 3077
rect -68 3005 -62 3039
rect -28 3005 -22 3039
rect -68 2967 -22 3005
rect -68 2933 -62 2967
rect -28 2933 -22 2967
rect -68 2895 -22 2933
rect -68 2861 -62 2895
rect -28 2861 -22 2895
rect -68 2823 -22 2861
rect -68 2789 -62 2823
rect -28 2789 -22 2823
rect -68 2751 -22 2789
rect -68 2717 -62 2751
rect -28 2717 -22 2751
rect -68 2679 -22 2717
rect -68 2645 -62 2679
rect -28 2645 -22 2679
rect -68 2607 -22 2645
rect -68 2573 -62 2607
rect -28 2573 -22 2607
rect -68 2535 -22 2573
rect -68 2501 -62 2535
rect -28 2501 -22 2535
rect -68 2463 -22 2501
rect -68 2429 -62 2463
rect -28 2429 -22 2463
rect -68 2391 -22 2429
rect -68 2357 -62 2391
rect -28 2357 -22 2391
rect -68 2319 -22 2357
rect -68 2285 -62 2319
rect -28 2285 -22 2319
rect -68 2247 -22 2285
rect -68 2213 -62 2247
rect -28 2213 -22 2247
rect -68 2175 -22 2213
rect -68 2141 -62 2175
rect -28 2141 -22 2175
rect -68 2103 -22 2141
rect -68 2069 -62 2103
rect -28 2069 -22 2103
rect -68 2031 -22 2069
rect -68 1997 -62 2031
rect -28 1997 -22 2031
rect -68 1959 -22 1997
rect -68 1925 -62 1959
rect -28 1925 -22 1959
rect -68 1887 -22 1925
rect -68 1853 -62 1887
rect -28 1853 -22 1887
rect -68 1815 -22 1853
rect -68 1781 -62 1815
rect -28 1781 -22 1815
rect -68 1743 -22 1781
rect -68 1709 -62 1743
rect -28 1709 -22 1743
rect -68 1670 -22 1709
rect -68 1636 -62 1670
rect -28 1636 -22 1670
rect -68 1597 -22 1636
rect -68 1563 -62 1597
rect -28 1563 -22 1597
rect -68 1524 -22 1563
rect -68 1490 -62 1524
rect -28 1490 -22 1524
rect -68 1451 -22 1490
rect -68 1417 -62 1451
rect -28 1417 -22 1451
rect -68 1378 -22 1417
rect -68 1344 -62 1378
rect -28 1344 -22 1378
rect 219 3697 265 3714
rect 219 3663 225 3697
rect 259 3663 265 3697
rect 219 3624 265 3663
rect 219 3590 225 3624
rect 259 3590 265 3624
rect 219 3551 265 3590
rect 219 3517 225 3551
rect 259 3517 265 3551
rect 219 3478 265 3517
rect 219 3444 225 3478
rect 259 3444 265 3478
rect 219 3405 265 3444
rect 219 3371 225 3405
rect 259 3371 265 3405
rect 219 3332 265 3371
rect 219 3298 225 3332
rect 259 3298 265 3332
rect 219 3260 265 3298
rect 219 3226 225 3260
rect 259 3226 265 3260
rect 219 3188 265 3226
rect 219 3154 225 3188
rect 259 3154 265 3188
rect 219 3116 265 3154
rect 219 3082 225 3116
rect 259 3082 265 3116
rect 219 3044 265 3082
rect 219 3010 225 3044
rect 259 3010 265 3044
rect 219 2972 265 3010
rect 219 2938 225 2972
rect 259 2938 265 2972
rect 219 2900 265 2938
rect 219 2866 225 2900
rect 259 2866 265 2900
rect 219 2828 265 2866
rect 219 2794 225 2828
rect 259 2794 265 2828
rect 219 2756 265 2794
rect 219 2722 225 2756
rect 259 2722 265 2756
rect 219 2684 265 2722
rect 219 2650 225 2684
rect 259 2650 265 2684
rect 219 2612 265 2650
rect 219 2578 225 2612
rect 259 2578 265 2612
rect 219 2540 265 2578
rect 219 2506 225 2540
rect 259 2506 265 2540
rect 219 2468 265 2506
rect 219 2434 225 2468
rect 259 2434 265 2468
rect 219 2396 265 2434
rect 219 2362 225 2396
rect 259 2362 265 2396
rect 219 2324 265 2362
rect 219 2290 225 2324
rect 259 2290 265 2324
rect 219 2252 265 2290
rect 219 2218 225 2252
rect 259 2218 265 2252
rect 219 2180 265 2218
rect 219 2146 225 2180
rect 259 2146 265 2180
rect 219 2108 265 2146
rect 219 2074 225 2108
rect 259 2074 265 2108
rect 219 2036 265 2074
rect 219 2002 225 2036
rect 259 2002 265 2036
rect 219 1964 265 2002
rect 219 1930 225 1964
rect 259 1930 265 1964
rect 219 1892 265 1930
rect 219 1858 225 1892
rect 259 1858 265 1892
rect 219 1820 265 1858
rect 219 1786 225 1820
rect 259 1786 265 1820
rect 219 1748 265 1786
rect 219 1714 225 1748
rect 259 1714 265 1748
rect 219 1676 265 1714
rect 219 1642 225 1676
rect 259 1642 265 1676
rect 219 1604 265 1642
rect 219 1570 225 1604
rect 259 1570 265 1604
rect 219 1532 265 1570
rect 219 1498 225 1532
rect 259 1498 265 1532
rect 219 1460 265 1498
rect 219 1426 225 1460
rect 259 1426 265 1460
rect 219 1388 265 1426
rect -68 1305 -22 1344
rect -68 1271 -62 1305
rect -28 1271 -22 1305
rect -68 1232 -22 1271
rect -68 1198 -62 1232
rect -28 1198 -22 1232
rect -68 1159 -22 1198
rect -68 1125 -62 1159
rect -28 1125 -22 1159
rect -68 1086 -22 1125
rect -68 1052 -62 1086
rect -28 1052 -22 1086
rect -68 1013 -22 1052
tri 213 1359 219 1365 se
rect 219 1359 225 1388
rect 213 1354 225 1359
rect 259 1354 265 1388
rect 213 1353 265 1354
rect 213 1282 225 1301
rect 259 1282 265 1301
rect 213 1271 265 1282
rect 213 1210 225 1219
rect 259 1210 265 1219
rect 213 1189 265 1210
rect 213 1107 265 1137
rect 213 1049 265 1055
tri 213 1043 219 1049 ne
rect -68 979 -62 1013
rect -28 979 -22 1013
rect -68 940 -22 979
rect -68 906 -62 940
rect -28 906 -22 940
rect -68 867 -22 906
rect -68 833 -62 867
rect -28 833 -22 867
rect -68 794 -22 833
rect -68 760 -62 794
rect -28 760 -22 794
rect -68 721 -22 760
rect -68 687 -62 721
rect -28 687 -22 721
rect -68 648 -22 687
rect -68 614 -62 648
rect -28 614 -22 648
rect -68 575 -22 614
rect -68 541 -62 575
rect -28 541 -22 575
rect -68 502 -22 541
rect -68 468 -62 502
rect -28 468 -22 502
rect 219 1028 265 1049
rect 219 994 225 1028
rect 259 994 265 1028
rect 219 956 265 994
rect 219 922 225 956
rect 259 922 265 956
rect 219 884 265 922
rect 219 850 225 884
rect 259 850 265 884
rect 219 812 265 850
rect 219 778 225 812
rect 259 778 265 812
rect 219 740 265 778
rect 219 706 225 740
rect 259 706 265 740
rect 219 668 265 706
rect 219 634 225 668
rect 259 634 265 668
rect 219 596 265 634
rect 219 562 225 596
rect 259 562 265 596
rect 219 524 265 562
rect 219 490 225 524
rect 259 490 265 524
tri 213 478 219 484 se
rect 219 478 265 490
rect -68 429 -22 468
tri 199 464 213 478 se
rect 213 464 265 478
rect -68 395 -62 429
rect -28 395 -22 429
rect -68 356 -22 395
rect -68 322 -62 356
rect -28 322 -22 356
rect -68 283 -22 322
rect -68 249 -62 283
rect -28 249 -22 283
rect -68 210 -22 249
tri 195 460 199 464 se
rect 199 460 265 464
rect 195 452 265 460
rect 195 418 225 452
rect 259 418 265 452
rect 195 380 265 418
rect 364 6892 410 6904
rect 364 6858 370 6892
rect 404 6858 410 6892
rect 364 6819 410 6858
rect 364 6785 370 6819
rect 404 6785 410 6819
rect 364 6746 410 6785
rect 364 6712 370 6746
rect 404 6712 410 6746
rect 364 6673 410 6712
rect 364 6639 370 6673
rect 404 6639 410 6673
rect 364 6600 410 6639
rect 364 6566 370 6600
rect 404 6566 410 6600
rect 364 6527 410 6566
rect 364 6493 370 6527
rect 404 6493 410 6527
rect 364 6454 410 6493
rect 364 6420 370 6454
rect 404 6420 410 6454
rect 364 6381 410 6420
rect 364 6347 370 6381
rect 404 6347 410 6381
rect 364 6308 410 6347
rect 364 6274 370 6308
rect 404 6274 410 6308
rect 364 6235 410 6274
rect 364 6201 370 6235
rect 404 6201 410 6235
rect 364 6162 410 6201
rect 364 6128 370 6162
rect 404 6128 410 6162
rect 364 6089 410 6128
rect 364 6055 370 6089
rect 404 6055 410 6089
rect 364 6016 410 6055
rect 364 5982 370 6016
rect 404 5982 410 6016
rect 364 5943 410 5982
rect 364 5909 370 5943
rect 404 5909 410 5943
rect 540 6875 546 6909
rect 580 6882 604 6909
rect 580 6875 586 6882
rect 540 6836 586 6875
tri 586 6864 604 6882 nw
rect 540 6802 546 6836
rect 580 6802 586 6836
rect 540 6763 586 6802
rect 540 6729 546 6763
rect 580 6729 586 6763
rect 540 6690 586 6729
rect 540 6656 546 6690
rect 580 6656 586 6690
rect 540 6617 586 6656
rect 540 6583 546 6617
rect 580 6583 586 6617
rect 540 6544 586 6583
rect 540 6510 546 6544
rect 580 6510 586 6544
rect 540 6471 586 6510
rect 540 6437 546 6471
rect 580 6437 586 6471
rect 540 6398 586 6437
rect 540 6364 546 6398
rect 580 6364 586 6398
rect 540 6325 586 6364
rect 540 6291 546 6325
rect 580 6291 586 6325
rect 540 6252 586 6291
rect 540 6218 546 6252
rect 580 6218 586 6252
rect 540 6179 586 6218
rect 540 6145 546 6179
rect 580 6145 586 6179
rect 540 6106 586 6145
rect 540 6072 546 6106
rect 580 6072 586 6106
rect 540 6050 586 6072
tri 586 6050 592 6056 sw
rect 540 6044 592 6050
rect 540 5962 592 5992
rect 364 5870 410 5909
rect 364 5836 370 5870
rect 404 5836 410 5870
rect 364 5797 410 5836
rect 364 5763 370 5797
rect 404 5763 410 5797
rect 364 5724 410 5763
rect 364 5690 370 5724
rect 404 5690 410 5724
rect 364 5651 410 5690
rect 364 5617 370 5651
rect 404 5617 410 5651
rect 364 5578 410 5617
rect 364 5544 370 5578
rect 404 5544 410 5578
rect 364 5505 410 5544
rect 364 5471 370 5505
rect 404 5471 410 5505
rect 364 5432 410 5471
rect 364 5398 370 5432
rect 404 5398 410 5432
rect 364 5359 410 5398
rect 364 5325 370 5359
rect 404 5325 410 5359
rect 364 5286 410 5325
rect 364 5252 370 5286
rect 404 5252 410 5286
rect 364 5213 410 5252
rect 364 5179 370 5213
rect 404 5179 410 5213
rect 364 5140 410 5179
rect 364 5106 370 5140
rect 404 5106 410 5140
rect 364 5067 410 5106
rect 364 5033 370 5067
rect 404 5033 410 5067
rect 364 4994 410 5033
rect 364 4960 370 4994
rect 404 4960 410 4994
rect 364 4921 410 4960
rect 364 4887 370 4921
rect 404 4887 410 4921
rect 364 4848 410 4887
rect 364 4814 370 4848
rect 404 4814 410 4848
rect 364 4775 410 4814
rect 364 4741 370 4775
rect 404 4741 410 4775
rect 364 4702 410 4741
rect 364 4668 370 4702
rect 404 4668 410 4702
rect 364 4629 410 4668
rect 364 4595 370 4629
rect 404 4595 410 4629
rect 364 4556 410 4595
rect 364 4522 370 4556
rect 404 4522 410 4556
rect 364 4483 410 4522
rect 364 4449 370 4483
rect 404 4449 410 4483
rect 364 4410 410 4449
rect 364 4376 370 4410
rect 404 4376 410 4410
rect 364 4337 410 4376
rect 364 4303 370 4337
rect 404 4303 410 4337
rect 364 4264 410 4303
rect 364 4230 370 4264
rect 404 4230 410 4264
rect 364 4191 410 4230
rect 364 4157 370 4191
rect 404 4157 410 4191
rect 364 4118 410 4157
rect 364 4084 370 4118
rect 404 4084 410 4118
rect 364 4045 410 4084
rect 364 4011 370 4045
rect 404 4011 410 4045
rect 364 3972 410 4011
rect 364 3938 370 3972
rect 404 3938 410 3972
rect 364 3899 410 3938
rect 364 3865 370 3899
rect 404 3865 410 3899
rect 364 3826 410 3865
rect 364 3792 370 3826
rect 404 3792 410 3826
rect 364 3753 410 3792
rect 364 3719 370 3753
rect 404 3719 410 3753
rect 364 3680 410 3719
rect 364 3646 370 3680
rect 404 3646 410 3680
rect 364 3607 410 3646
rect 364 3573 370 3607
rect 404 3573 410 3607
rect 364 3534 410 3573
rect 364 3500 370 3534
rect 404 3500 410 3534
rect 364 3461 410 3500
rect 364 3427 370 3461
rect 404 3427 410 3461
rect 364 3388 410 3427
rect 364 3354 370 3388
rect 404 3354 410 3388
rect 364 3315 410 3354
rect 364 3281 370 3315
rect 404 3281 410 3315
rect 364 3241 410 3281
rect 364 3207 370 3241
rect 404 3207 410 3241
rect 364 3163 410 3207
rect 364 3129 370 3163
rect 404 3129 410 3163
rect 364 3090 410 3129
rect 364 3056 370 3090
rect 404 3056 410 3090
rect 364 3018 410 3056
rect 364 2984 370 3018
rect 404 2984 410 3018
rect 364 2946 410 2984
rect 364 2912 370 2946
rect 404 2912 410 2946
rect 364 2874 410 2912
rect 364 2840 370 2874
rect 404 2840 410 2874
rect 364 2802 410 2840
rect 364 2768 370 2802
rect 404 2768 410 2802
rect 364 2730 410 2768
rect 364 2696 370 2730
rect 404 2696 410 2730
rect 364 2658 410 2696
rect 364 2624 370 2658
rect 404 2624 410 2658
rect 364 2586 410 2624
rect 364 2552 370 2586
rect 404 2552 410 2586
rect 364 2514 410 2552
rect 364 2480 370 2514
rect 404 2480 410 2514
rect 364 2442 410 2480
rect 364 2408 370 2442
rect 404 2408 410 2442
rect 364 2370 410 2408
rect 364 2336 370 2370
rect 404 2336 410 2370
rect 364 2298 410 2336
rect 364 2264 370 2298
rect 404 2264 410 2298
rect 364 2226 410 2264
rect 364 2192 370 2226
rect 404 2192 410 2226
rect 364 2154 410 2192
rect 364 2120 370 2154
rect 404 2120 410 2154
rect 364 2082 410 2120
rect 364 2048 370 2082
rect 404 2048 410 2082
rect 364 2010 410 2048
rect 364 1976 370 2010
rect 404 1976 410 2010
rect 364 1938 410 1976
rect 364 1904 370 1938
rect 404 1904 410 1938
rect 364 1866 410 1904
rect 364 1832 370 1866
rect 404 1832 410 1866
rect 364 1794 410 1832
rect 364 1760 370 1794
rect 404 1760 410 1794
rect 364 1722 410 1760
rect 364 1688 370 1722
rect 404 1688 410 1722
rect 364 1650 410 1688
rect 364 1616 370 1650
rect 404 1616 410 1650
rect 364 1578 410 1616
rect 364 1544 370 1578
rect 404 1544 410 1578
rect 364 1506 410 1544
rect 364 1472 370 1506
rect 404 1472 410 1506
rect 364 1434 410 1472
rect 466 5922 512 5934
rect 466 5888 472 5922
rect 506 5888 512 5922
rect 466 5849 512 5888
rect 466 5815 472 5849
rect 506 5815 512 5849
rect 466 5776 512 5815
rect 466 5742 472 5776
rect 506 5742 512 5776
rect 466 5703 512 5742
rect 466 5669 472 5703
rect 506 5669 512 5703
rect 466 5630 512 5669
rect 466 5596 472 5630
rect 506 5596 512 5630
rect 466 5557 512 5596
rect 466 5523 472 5557
rect 506 5523 512 5557
rect 466 5484 512 5523
rect 466 5450 472 5484
rect 506 5450 512 5484
rect 466 5411 512 5450
rect 466 5377 472 5411
rect 506 5377 512 5411
rect 466 5338 512 5377
rect 466 5304 472 5338
rect 506 5304 512 5338
rect 466 5265 512 5304
rect 466 5231 472 5265
rect 506 5231 512 5265
rect 466 5192 512 5231
rect 466 5158 472 5192
rect 506 5158 512 5192
rect 466 5119 512 5158
rect 466 5085 472 5119
rect 506 5085 512 5119
rect 466 5046 512 5085
rect 466 5012 472 5046
rect 506 5012 512 5046
rect 466 4973 512 5012
rect 466 4939 472 4973
rect 506 4939 512 4973
rect 466 4900 512 4939
rect 466 4866 472 4900
rect 506 4866 512 4900
rect 466 4827 512 4866
rect 466 4793 472 4827
rect 506 4793 512 4827
rect 466 4754 512 4793
rect 466 4720 472 4754
rect 506 4720 512 4754
rect 466 4681 512 4720
rect 466 4647 472 4681
rect 506 4647 512 4681
rect 466 4608 512 4647
rect 466 4574 472 4608
rect 506 4574 512 4608
rect 466 4535 512 4574
rect 466 4501 472 4535
rect 506 4501 512 4535
rect 466 4461 512 4501
rect 466 4427 472 4461
rect 506 4427 512 4461
rect 466 4387 512 4427
rect 466 4353 472 4387
rect 506 4353 512 4387
rect 466 4313 512 4353
rect 466 4279 472 4313
rect 506 4279 512 4313
rect 466 4239 512 4279
rect 466 4205 472 4239
rect 506 4205 512 4239
rect 466 4165 512 4205
rect 466 4131 472 4165
rect 506 4131 512 4165
rect 466 4091 512 4131
rect 466 4057 472 4091
rect 506 4057 512 4091
rect 466 4017 512 4057
rect 466 3983 472 4017
rect 506 3983 512 4017
rect 466 3943 512 3983
rect 466 3909 472 3943
rect 506 3909 512 3943
rect 466 3869 512 3909
rect 466 3835 472 3869
rect 506 3835 512 3869
rect 466 3795 512 3835
rect 466 3761 472 3795
rect 506 3761 512 3795
rect 466 3721 512 3761
rect 466 3687 472 3721
rect 506 3687 512 3721
rect 466 3647 512 3687
rect 466 3613 472 3647
rect 506 3613 512 3647
rect 466 3572 512 3613
rect 466 3538 472 3572
rect 506 3538 512 3572
rect 466 3498 512 3538
rect 466 3464 472 3498
rect 506 3464 512 3498
rect 466 3424 512 3464
rect 466 3390 472 3424
rect 506 3390 512 3424
rect 466 3350 512 3390
rect 466 3316 472 3350
rect 506 3316 512 3350
rect 466 3276 512 3316
rect 466 3242 472 3276
rect 506 3242 512 3276
rect 466 3202 512 3242
rect 466 3168 472 3202
rect 506 3168 512 3202
rect 466 3128 512 3168
rect 466 3094 472 3128
rect 506 3094 512 3128
rect 466 3054 512 3094
rect 466 3020 472 3054
rect 506 3020 512 3054
rect 466 2980 512 3020
rect 466 2946 472 2980
rect 506 2946 512 2980
rect 466 2906 512 2946
rect 466 2872 472 2906
rect 506 2872 512 2906
rect 466 2832 512 2872
rect 466 2798 472 2832
rect 506 2798 512 2832
rect 466 2758 512 2798
rect 466 2724 472 2758
rect 506 2724 512 2758
rect 466 2684 512 2724
rect 466 2650 472 2684
rect 506 2650 512 2684
rect 466 2610 512 2650
rect 466 2576 472 2610
rect 506 2576 512 2610
rect 466 2536 512 2576
rect 466 2502 472 2536
rect 506 2502 512 2536
rect 466 2462 512 2502
rect 466 2428 472 2462
rect 506 2428 512 2462
rect 466 2388 512 2428
rect 466 2354 472 2388
rect 506 2354 512 2388
rect 466 2314 512 2354
rect 466 2280 472 2314
rect 506 2280 512 2314
rect 466 2241 512 2280
rect 466 2207 472 2241
rect 506 2207 512 2241
rect 466 2168 512 2207
rect 466 2134 472 2168
rect 506 2134 512 2168
rect 466 2095 512 2134
rect 466 2061 472 2095
rect 506 2061 512 2095
rect 466 2022 512 2061
rect 466 1988 472 2022
rect 506 1988 512 2022
rect 466 1949 512 1988
rect 466 1915 472 1949
rect 506 1915 512 1949
rect 466 1876 512 1915
rect 466 1842 472 1876
rect 506 1842 512 1876
rect 466 1803 512 1842
rect 466 1769 472 1803
rect 506 1769 512 1803
rect 466 1730 512 1769
rect 466 1696 472 1730
rect 506 1696 512 1730
rect 466 1657 512 1696
rect 466 1623 472 1657
rect 506 1623 512 1657
rect 466 1584 512 1623
rect 466 1550 472 1584
rect 506 1550 512 1584
rect 466 1511 512 1550
rect 466 1477 472 1511
rect 506 1477 512 1511
rect 466 1465 512 1477
rect 540 5887 592 5910
rect 540 5880 546 5887
rect 580 5880 592 5887
rect 540 5814 592 5828
rect 540 5798 546 5814
rect 580 5798 592 5814
rect 540 5741 592 5746
rect 540 5707 546 5741
rect 580 5740 592 5741
rect 580 5707 586 5740
tri 586 5734 592 5740 nw
rect 540 5668 586 5707
rect 540 5634 546 5668
rect 580 5634 586 5668
rect 540 5595 586 5634
rect 540 5561 546 5595
rect 580 5561 586 5595
rect 540 5522 586 5561
rect 540 5488 546 5522
rect 580 5488 586 5522
rect 540 5449 586 5488
rect 540 5415 546 5449
rect 580 5415 586 5449
rect 540 5376 586 5415
rect 540 5342 546 5376
rect 580 5342 586 5376
rect 540 5303 586 5342
rect 540 5269 546 5303
rect 580 5269 586 5303
rect 540 5230 586 5269
rect 540 5196 546 5230
rect 580 5196 586 5230
rect 540 5157 586 5196
rect 540 5123 546 5157
rect 580 5123 586 5157
rect 540 5084 586 5123
rect 540 5050 546 5084
rect 580 5050 586 5084
rect 540 5011 586 5050
rect 540 4977 546 5011
rect 580 4977 586 5011
rect 540 4938 586 4977
rect 540 4904 546 4938
rect 580 4904 586 4938
rect 540 4865 586 4904
rect 540 4831 546 4865
rect 580 4831 586 4865
rect 540 4792 586 4831
rect 540 4758 546 4792
rect 580 4758 586 4792
rect 540 4719 586 4758
rect 540 4685 546 4719
rect 580 4685 586 4719
rect 540 4646 586 4685
rect 540 4612 546 4646
rect 580 4612 586 4646
rect 540 4573 586 4612
rect 540 4539 546 4573
rect 580 4539 586 4573
rect 540 4500 586 4539
rect 540 4466 546 4500
rect 580 4466 586 4500
rect 540 4426 586 4466
rect 540 4392 546 4426
rect 580 4392 586 4426
rect 540 4352 586 4392
rect 540 4318 546 4352
rect 580 4318 586 4352
rect 540 4278 586 4318
rect 540 4244 546 4278
rect 580 4244 586 4278
rect 540 4204 586 4244
rect 540 4170 546 4204
rect 580 4170 586 4204
rect 540 4130 586 4170
rect 540 4096 546 4130
rect 580 4096 586 4130
rect 540 4056 586 4096
rect 540 4022 546 4056
rect 580 4024 586 4056
tri 586 4024 592 4030 sw
rect 580 4022 592 4024
rect 540 4018 592 4022
rect 540 3948 546 3966
rect 580 3948 592 3966
rect 540 3936 592 3948
rect 540 3874 546 3884
rect 580 3874 592 3884
rect 540 3854 592 3874
rect 540 3800 546 3802
rect 580 3800 592 3802
rect 540 3772 592 3800
rect 540 3714 592 3720
rect 540 3670 586 3714
tri 586 3708 592 3714 nw
rect 540 3636 546 3670
rect 580 3636 586 3670
rect 540 3597 586 3636
rect 540 3563 546 3597
rect 580 3563 586 3597
rect 540 3524 586 3563
rect 540 3490 546 3524
rect 580 3490 586 3524
rect 540 3451 586 3490
rect 540 3417 546 3451
rect 580 3417 586 3451
rect 540 3378 586 3417
rect 540 3344 546 3378
rect 580 3344 586 3378
rect 540 3305 586 3344
rect 540 3271 546 3305
rect 580 3271 586 3305
rect 540 3232 586 3271
rect 540 3198 546 3232
rect 580 3198 586 3232
rect 540 3159 586 3198
rect 540 3125 546 3159
rect 580 3125 586 3159
rect 540 3086 586 3125
rect 540 3052 546 3086
rect 580 3052 586 3086
rect 540 3013 586 3052
rect 540 2979 546 3013
rect 580 2979 586 3013
rect 540 2940 586 2979
rect 540 2906 546 2940
rect 580 2906 586 2940
rect 540 2867 586 2906
rect 540 2833 546 2867
rect 580 2833 586 2867
rect 540 2794 586 2833
rect 540 2760 546 2794
rect 580 2760 586 2794
rect 540 2721 586 2760
rect 540 2687 546 2721
rect 580 2687 586 2721
rect 540 2648 586 2687
rect 540 2614 546 2648
rect 580 2614 586 2648
rect 540 2575 586 2614
rect 540 2541 546 2575
rect 580 2541 586 2575
rect 540 2502 586 2541
rect 540 2468 546 2502
rect 580 2468 586 2502
rect 540 2429 586 2468
rect 540 2395 546 2429
rect 580 2395 586 2429
rect 540 2356 586 2395
rect 540 2322 546 2356
rect 580 2322 586 2356
rect 540 2283 586 2322
rect 540 2249 546 2283
rect 580 2249 586 2283
rect 540 2210 586 2249
rect 540 2176 546 2210
rect 580 2176 586 2210
rect 540 2137 586 2176
rect 540 2103 546 2137
rect 580 2103 586 2137
rect 540 2064 586 2103
rect 540 2030 546 2064
rect 580 2030 586 2064
rect 540 1991 586 2030
rect 540 1957 546 1991
rect 580 1957 586 1991
rect 540 1918 586 1957
rect 540 1884 546 1918
rect 580 1884 586 1918
rect 540 1845 586 1884
rect 540 1811 546 1845
rect 580 1811 586 1845
rect 540 1772 586 1811
rect 540 1738 546 1772
rect 580 1738 586 1772
rect 540 1699 586 1738
rect 540 1665 546 1699
rect 580 1665 586 1699
rect 540 1626 586 1665
rect 540 1592 546 1626
rect 580 1592 586 1626
rect 540 1553 586 1592
rect 540 1519 546 1553
rect 580 1519 586 1553
rect 540 1480 586 1519
rect 364 1400 370 1434
rect 404 1400 410 1434
rect 364 1362 410 1400
rect 364 1328 370 1362
rect 404 1328 410 1362
rect 364 1290 410 1328
rect 364 1256 370 1290
rect 404 1256 410 1290
rect 364 1218 410 1256
rect 364 1184 370 1218
rect 404 1184 410 1218
rect 364 1146 410 1184
rect 364 1112 370 1146
rect 404 1112 410 1146
rect 364 1074 410 1112
rect 364 1040 370 1074
rect 404 1040 410 1074
rect 364 1002 410 1040
rect 364 968 370 1002
rect 404 968 410 1002
rect 364 930 410 968
rect 364 896 370 930
rect 404 896 410 930
rect 364 858 410 896
rect 364 824 370 858
rect 404 824 410 858
rect 364 786 410 824
rect 364 752 370 786
rect 404 752 410 786
rect 364 714 410 752
rect 364 680 370 714
rect 404 680 410 714
rect 364 642 410 680
rect 364 608 370 642
rect 404 608 410 642
rect 364 570 410 608
rect 364 536 370 570
rect 404 536 410 570
rect 364 498 410 536
rect 364 464 370 498
rect 404 464 410 498
rect 364 426 410 464
rect 364 392 370 426
rect 404 392 410 426
rect 364 380 410 392
rect 540 1446 546 1480
rect 580 1446 586 1480
rect 540 1407 586 1446
rect 540 1373 546 1407
rect 580 1373 586 1407
rect 540 1359 586 1373
tri 586 1359 592 1365 sw
rect 540 1353 592 1359
rect 540 1300 546 1301
rect 580 1300 592 1301
rect 540 1271 592 1300
rect 540 1189 592 1219
rect 540 1115 592 1137
rect 540 1107 546 1115
rect 580 1107 592 1115
rect 540 1049 592 1055
rect 540 1042 586 1049
tri 586 1043 592 1049 nw
rect 540 1008 546 1042
rect 580 1008 586 1042
rect 540 969 586 1008
rect 540 935 546 969
rect 580 935 586 969
rect 540 896 586 935
rect 540 862 546 896
rect 580 862 586 896
rect 540 823 586 862
rect 540 789 546 823
rect 580 789 586 823
rect 540 750 586 789
rect 540 716 546 750
rect 580 716 586 750
rect 540 677 586 716
rect 540 643 546 677
rect 580 643 586 677
rect 540 604 586 643
rect 540 570 546 604
rect 580 570 586 604
rect 540 530 586 570
rect 540 496 546 530
rect 580 496 586 530
rect 540 460 586 496
tri 586 460 604 478 sw
rect 540 456 604 460
rect 540 422 546 456
rect 580 422 604 456
rect 540 382 604 422
rect 195 346 225 380
rect 259 367 265 380
tri 265 367 266 368 sw
rect 259 348 266 367
tri 266 348 285 367 sw
tri 521 348 540 367 se
rect 540 348 546 382
rect 580 348 604 382
rect 259 346 285 348
rect 195 327 285 346
tri 285 327 306 348 sw
tri 506 333 521 348 se
rect 521 333 604 348
tri 500 327 506 333 se
rect 506 327 604 333
rect 195 308 604 327
rect 195 274 225 308
rect 259 274 306 308
rect 340 274 386 308
rect 420 274 466 308
rect 500 274 546 308
rect 580 274 604 308
rect 195 219 604 274
rect -68 176 -62 210
rect -28 176 -22 210
rect -68 137 -22 176
tri 845 144 908 207 se
rect 908 144 936 207
rect -68 103 -62 137
rect -28 107 -22 137
tri -22 107 15 144 sw
tri 808 107 845 144 se
rect 845 107 936 144
rect -28 103 15 107
rect -68 61 15 103
rect 16 101 936 107
rect 16 67 28 101
rect 62 67 106 101
rect 140 67 184 101
rect 218 67 262 101
rect 296 67 340 101
rect 374 67 418 101
rect 452 67 496 101
rect 530 67 574 101
rect 608 67 652 101
rect 686 67 730 101
rect 764 67 808 101
rect 842 67 936 101
rect 16 61 936 67
<< via1 >>
rect 213 6033 265 6044
rect 213 5999 225 6033
rect 225 5999 259 6033
rect 259 5999 265 6033
rect 213 5992 265 5999
rect 213 5960 265 5962
rect 213 5926 225 5960
rect 225 5926 259 5960
rect 259 5926 265 5960
rect 213 5910 265 5926
rect 213 5853 225 5880
rect 225 5853 259 5880
rect 259 5853 265 5880
rect 213 5828 265 5853
rect 213 5780 225 5798
rect 225 5780 259 5798
rect 259 5780 265 5798
rect 213 5746 265 5780
rect 213 3989 265 4018
rect 213 3966 225 3989
rect 225 3966 259 3989
rect 259 3966 265 3989
rect 213 3916 265 3936
rect 213 3884 225 3916
rect 225 3884 259 3916
rect 259 3884 265 3916
rect 213 3843 265 3854
rect 213 3809 225 3843
rect 225 3809 259 3843
rect 259 3809 265 3843
rect 213 3802 265 3809
rect 213 3770 265 3772
rect 213 3736 225 3770
rect 225 3736 259 3770
rect 259 3736 265 3770
rect 213 3720 265 3736
rect 213 1316 265 1353
rect 213 1301 225 1316
rect 225 1301 259 1316
rect 259 1301 265 1316
rect 213 1244 265 1271
rect 213 1219 225 1244
rect 225 1219 259 1244
rect 259 1219 265 1244
rect 213 1172 265 1189
rect 213 1138 225 1172
rect 225 1138 259 1172
rect 259 1138 265 1172
rect 213 1137 265 1138
rect 213 1100 265 1107
rect 213 1066 225 1100
rect 225 1066 259 1100
rect 259 1066 265 1100
rect 213 1055 265 1066
rect 540 6033 592 6044
rect 540 5999 546 6033
rect 546 5999 580 6033
rect 580 5999 592 6033
rect 540 5992 592 5999
rect 540 5960 592 5962
rect 540 5926 546 5960
rect 546 5926 580 5960
rect 580 5926 592 5960
rect 540 5910 592 5926
rect 540 5853 546 5880
rect 546 5853 580 5880
rect 580 5853 592 5880
rect 540 5828 592 5853
rect 540 5780 546 5798
rect 546 5780 580 5798
rect 580 5780 592 5798
rect 540 5746 592 5780
rect 540 3982 592 4018
rect 540 3966 546 3982
rect 546 3966 580 3982
rect 580 3966 592 3982
rect 540 3908 592 3936
rect 540 3884 546 3908
rect 546 3884 580 3908
rect 580 3884 592 3908
rect 540 3834 592 3854
rect 540 3802 546 3834
rect 546 3802 580 3834
rect 580 3802 592 3834
rect 540 3760 592 3772
rect 540 3726 546 3760
rect 546 3726 580 3760
rect 580 3726 592 3760
rect 540 3720 592 3726
rect 540 1334 592 1353
rect 540 1301 546 1334
rect 546 1301 580 1334
rect 580 1301 592 1334
rect 540 1261 592 1271
rect 540 1227 546 1261
rect 546 1227 580 1261
rect 580 1227 592 1261
rect 540 1219 592 1227
rect 540 1188 592 1189
rect 540 1154 546 1188
rect 546 1154 580 1188
rect 580 1154 592 1188
rect 540 1137 592 1154
rect 540 1081 546 1107
rect 546 1081 580 1107
rect 580 1081 592 1107
rect 540 1055 592 1081
<< metal2 >>
rect 213 6044 592 6050
rect 265 5992 540 6044
rect 213 5962 592 5992
rect 265 5910 540 5962
rect 213 5880 592 5910
rect 265 5828 540 5880
rect 213 5798 592 5828
rect 265 5746 540 5798
rect 213 5740 592 5746
rect 213 4018 592 4024
rect 265 3966 540 4018
rect 213 3936 592 3966
rect 265 3884 540 3936
rect 213 3854 592 3884
rect 265 3802 540 3854
rect 213 3772 592 3802
rect 265 3720 540 3772
rect 213 3714 592 3720
rect 213 1353 592 1359
rect 265 1301 540 1353
rect 213 1271 592 1301
rect 265 1219 540 1271
rect 213 1189 592 1219
rect 265 1137 540 1189
rect 213 1107 592 1137
rect 265 1055 540 1107
rect 213 1049 592 1055
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_0
timestamp 1649977179
transform 1 0 415 0 -1 5835
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_1
timestamp 1649977179
transform 1 0 415 0 -1 6956
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_2
timestamp 1649977179
transform 1 0 415 0 1 1483
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_3
timestamp 1649977179
transform 1 0 415 0 1 362
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_4
timestamp 1649977179
transform 1 0 415 0 -1 4714
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_5
timestamp 1649977179
transform 1 0 415 0 1 2604
box -28 0 148 471
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1649977179
transform 1 0 456 0 1 1385
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1649977179
transform 1 0 456 0 1 3626
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_2
timestamp 1649977179
transform 1 0 456 0 1 5866
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_3
timestamp 1649977179
transform 1 0 456 0 1 4745
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_4
timestamp 1649977179
transform 1 0 456 0 1 2506
box 0 0 1 1
<< labels >>
flabel metal1 s 466 3284 512 3414 0 FreeSans 200 0 0 0 PD_H
port 1 nsew
flabel metal1 s 367 2854 410 2984 0 FreeSans 200 0 0 0 PAD
port 2 nsew
flabel metal1 s 365 4748 408 4878 0 FreeSans 200 0 0 0 PAD
port 2 nsew
flabel metal1 s 466 4318 512 4448 0 FreeSans 200 0 0 0 PD_H
port 1 nsew
<< properties >>
string GDS_END 5603770
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 5542226
<< end >>
