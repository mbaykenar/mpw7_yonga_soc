magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -42 416 913 1116
<< pwell >>
rect 40 118 846 310
<< mvnmos >>
rect 119 144 239 284
rect 295 144 415 284
rect 471 144 591 284
rect 647 144 767 284
<< mvpmos >>
rect 119 750 239 950
rect 295 750 415 950
rect 471 750 591 950
rect 647 750 767 950
rect 119 482 239 682
rect 295 482 415 682
rect 471 482 591 682
rect 647 482 767 682
<< mvndiff >>
rect 66 272 119 284
rect 66 238 74 272
rect 108 238 119 272
rect 66 204 119 238
rect 66 170 74 204
rect 108 170 119 204
rect 66 144 119 170
rect 239 272 295 284
rect 239 238 250 272
rect 284 238 295 272
rect 239 204 295 238
rect 239 170 250 204
rect 284 170 295 204
rect 239 144 295 170
rect 415 272 471 284
rect 415 238 426 272
rect 460 238 471 272
rect 415 204 471 238
rect 415 170 426 204
rect 460 170 471 204
rect 415 144 471 170
rect 591 272 647 284
rect 591 238 602 272
rect 636 238 647 272
rect 591 204 647 238
rect 591 170 602 204
rect 636 170 647 204
rect 591 144 647 170
rect 767 272 820 284
rect 767 238 778 272
rect 812 238 820 272
rect 767 204 820 238
rect 767 170 778 204
rect 812 170 820 204
rect 767 144 820 170
<< mvpdiff >>
rect 66 932 119 950
rect 66 898 74 932
rect 108 898 119 932
rect 66 864 119 898
rect 66 830 74 864
rect 108 830 119 864
rect 66 796 119 830
rect 66 762 74 796
rect 108 762 119 796
rect 66 750 119 762
rect 239 932 295 950
rect 239 898 250 932
rect 284 898 295 932
rect 239 864 295 898
rect 239 830 250 864
rect 284 830 295 864
rect 239 796 295 830
rect 239 762 250 796
rect 284 762 295 796
rect 239 750 295 762
rect 415 932 471 950
rect 415 898 426 932
rect 460 898 471 932
rect 415 864 471 898
rect 415 830 426 864
rect 460 830 471 864
rect 415 796 471 830
rect 415 762 426 796
rect 460 762 471 796
rect 415 750 471 762
rect 591 932 647 950
rect 591 898 602 932
rect 636 898 647 932
rect 591 864 647 898
rect 591 830 602 864
rect 636 830 647 864
rect 591 796 647 830
rect 591 762 602 796
rect 636 762 647 796
rect 591 750 647 762
rect 767 932 820 950
rect 767 898 778 932
rect 812 898 820 932
rect 767 864 820 898
rect 767 830 778 864
rect 812 830 820 864
rect 767 796 820 830
rect 767 762 778 796
rect 812 762 820 796
rect 767 750 820 762
rect 66 670 119 682
rect 66 636 74 670
rect 108 636 119 670
rect 66 602 119 636
rect 66 568 74 602
rect 108 568 119 602
rect 66 534 119 568
rect 66 500 74 534
rect 108 500 119 534
rect 66 482 119 500
rect 239 670 295 682
rect 239 636 250 670
rect 284 636 295 670
rect 239 602 295 636
rect 239 568 250 602
rect 284 568 295 602
rect 239 534 295 568
rect 239 500 250 534
rect 284 500 295 534
rect 239 482 295 500
rect 415 670 471 682
rect 415 636 426 670
rect 460 636 471 670
rect 415 602 471 636
rect 415 568 426 602
rect 460 568 471 602
rect 415 534 471 568
rect 415 500 426 534
rect 460 500 471 534
rect 415 482 471 500
rect 591 670 647 682
rect 591 636 602 670
rect 636 636 647 670
rect 591 602 647 636
rect 591 568 602 602
rect 636 568 647 602
rect 591 534 647 568
rect 591 500 602 534
rect 636 500 647 534
rect 591 482 647 500
rect 767 670 820 682
rect 767 636 778 670
rect 812 636 820 670
rect 767 602 820 636
rect 767 568 778 602
rect 812 568 820 602
rect 767 534 820 568
rect 767 500 778 534
rect 812 500 820 534
rect 767 482 820 500
<< mvndiffc >>
rect 74 238 108 272
rect 74 170 108 204
rect 250 238 284 272
rect 250 170 284 204
rect 426 238 460 272
rect 426 170 460 204
rect 602 238 636 272
rect 602 170 636 204
rect 778 238 812 272
rect 778 170 812 204
<< mvpdiffc >>
rect 74 898 108 932
rect 74 830 108 864
rect 74 762 108 796
rect 250 898 284 932
rect 250 830 284 864
rect 250 762 284 796
rect 426 898 460 932
rect 426 830 460 864
rect 426 762 460 796
rect 602 898 636 932
rect 602 830 636 864
rect 602 762 636 796
rect 778 898 812 932
rect 778 830 812 864
rect 778 762 812 796
rect 74 636 108 670
rect 74 568 108 602
rect 74 500 108 534
rect 250 636 284 670
rect 250 568 284 602
rect 250 500 284 534
rect 426 636 460 670
rect 426 568 460 602
rect 426 500 460 534
rect 602 636 636 670
rect 602 568 636 602
rect 602 500 636 534
rect 778 636 812 670
rect 778 568 812 602
rect 778 500 812 534
<< poly >>
rect 119 950 239 976
rect 295 950 415 976
rect 471 950 591 976
rect 647 950 767 976
rect 119 682 239 750
rect 295 682 415 750
rect 471 682 591 750
rect 647 682 767 750
rect 119 434 239 482
rect 119 400 165 434
rect 199 400 239 434
rect 119 366 239 400
rect 119 332 165 366
rect 199 332 239 366
rect 119 284 239 332
rect 295 407 415 482
rect 471 407 591 482
rect 295 391 591 407
rect 295 357 318 391
rect 352 357 386 391
rect 420 357 454 391
rect 488 357 522 391
rect 556 357 591 391
rect 295 341 591 357
rect 295 284 415 341
rect 471 284 591 341
rect 647 434 767 482
rect 647 400 687 434
rect 721 400 767 434
rect 647 366 767 400
rect 647 332 687 366
rect 721 332 767 366
rect 647 284 767 332
rect 119 118 239 144
rect 295 118 415 144
rect 471 118 591 144
rect 647 118 767 144
<< polycont >>
rect 165 400 199 434
rect 165 332 199 366
rect 318 357 352 391
rect 386 357 420 391
rect 454 357 488 391
rect 522 357 556 391
rect 687 400 721 434
rect 687 332 721 366
<< locali >>
rect 74 932 108 944
rect 74 864 108 872
rect 74 796 108 830
rect 74 670 108 762
rect 74 602 108 636
rect 74 534 108 568
rect 250 932 284 950
rect 250 864 284 898
rect 250 796 284 830
rect 250 670 284 762
rect 250 602 284 636
rect 250 534 284 568
rect 74 484 108 500
rect 249 500 250 519
rect 426 932 460 944
rect 426 864 460 872
rect 426 796 460 830
rect 426 670 460 762
rect 426 602 460 636
rect 426 534 460 568
rect 284 500 287 519
rect 249 485 287 500
rect 602 932 636 950
rect 602 864 636 898
rect 602 796 636 830
rect 602 670 636 762
rect 602 602 636 636
rect 602 534 636 568
rect 149 433 165 434
rect 199 433 215 434
rect 144 400 165 433
rect 144 399 182 400
rect 149 366 215 399
rect 149 332 165 366
rect 199 332 215 366
rect 74 272 108 288
rect 74 227 108 238
rect 74 155 108 170
rect 250 272 284 485
rect 426 484 460 500
rect 600 500 602 519
rect 778 932 812 944
rect 778 864 812 872
rect 778 796 812 830
rect 778 670 812 762
rect 778 602 812 636
rect 778 534 812 568
rect 636 500 638 519
rect 600 485 638 500
rect 318 399 319 407
rect 353 399 421 433
rect 455 399 522 433
rect 318 391 556 399
rect 352 357 386 391
rect 420 357 454 391
rect 488 357 522 391
rect 318 341 556 357
rect 250 204 284 238
rect 250 154 284 170
rect 426 272 460 288
rect 426 227 460 238
rect 426 155 460 170
rect 602 272 636 485
rect 778 484 812 500
rect 671 400 687 434
rect 723 400 737 434
rect 671 366 737 400
rect 671 332 687 366
rect 721 362 737 366
rect 723 332 737 362
rect 602 204 636 238
rect 602 154 636 170
rect 778 272 812 288
rect 778 227 812 238
rect 778 155 812 170
<< viali >>
rect 74 944 108 978
rect 74 898 108 906
rect 74 872 108 898
rect 215 485 249 519
rect 426 944 460 978
rect 426 898 460 906
rect 426 872 460 898
rect 287 485 321 519
rect 110 399 144 433
rect 182 400 199 433
rect 199 400 216 433
rect 182 399 216 400
rect 74 204 108 227
rect 74 193 108 204
rect 74 121 108 155
rect 566 485 600 519
rect 778 944 812 978
rect 778 898 812 906
rect 778 872 812 898
rect 638 485 672 519
rect 319 399 353 433
rect 421 399 455 433
rect 522 399 556 433
rect 426 204 460 227
rect 426 193 460 204
rect 426 121 460 155
rect 689 400 721 434
rect 721 400 723 434
rect 689 332 721 362
rect 721 332 723 362
rect 689 328 723 332
rect 778 204 812 227
rect 778 193 812 204
rect 778 121 812 155
<< metal1 >>
rect 24 978 847 1062
rect 24 944 74 978
rect 108 944 426 978
rect 460 944 778 978
rect 812 944 847 978
rect 24 906 847 944
rect 24 872 74 906
rect 108 872 426 906
rect 460 872 778 906
rect 812 872 847 906
rect 24 859 847 872
rect 203 519 684 525
rect 203 485 215 519
rect 249 485 287 519
rect 321 485 566 519
rect 600 485 638 519
rect 672 485 684 519
rect 203 479 684 485
tri 676 439 683 446 se
rect 683 439 729 446
rect 98 434 729 439
rect 98 433 689 434
rect 98 399 110 433
rect 144 399 182 433
rect 216 399 319 433
rect 353 399 421 433
rect 455 399 522 433
rect 556 400 689 433
rect 723 400 729 434
rect 556 399 729 400
rect 98 393 729 399
tri 649 362 680 393 ne
rect 680 362 729 393
tri 680 359 683 362 ne
rect 683 328 689 362
rect 723 328 729 362
rect 683 316 729 328
rect 24 227 847 239
rect 24 193 74 227
rect 108 193 426 227
rect 460 193 778 227
rect 812 193 847 227
rect 24 155 847 193
rect 24 121 74 155
rect 108 121 426 155
rect 460 121 778 155
rect 812 121 847 155
rect 24 24 847 121
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808615  sky130_fd_pr__model__nfet_highvoltage__example_55959141808615_0
timestamp 1649977179
transform 1 0 119 0 -1 284
box -28 0 676 63
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808616  sky130_fd_pr__model__pfet_highvoltage__example_55959141808616_0
timestamp 1649977179
transform 1 0 119 0 -1 682
box -28 0 676 97
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808616  sky130_fd_pr__model__pfet_highvoltage__example_55959141808616_1
timestamp 1649977179
transform 1 0 119 0 1 750
box -28 0 676 97
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1649977179
transform 0 -1 812 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1649977179
transform 0 -1 812 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1649977179
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1649977179
transform 0 -1 460 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1649977179
transform 0 -1 460 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1649977179
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1649977179
transform 0 -1 215 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1649977179
transform 0 -1 737 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808612  sky130_fd_pr__via_pol1__example_55959141808612_0
timestamp 1649977179
transform 1 0 302 0 1 341
box 0 0 1 1
<< labels >>
flabel metal1 s 149 396 200 437 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 s 352 488 401 522 0 FreeSans 200 0 0 0 OUT
port 2 nsew
<< properties >>
string GDS_END 7954714
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7950372
<< end >>
