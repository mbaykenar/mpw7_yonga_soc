magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 2 67 631 203
rect 2 21 443 67
rect 30 -17 64 21
<< locali >>
rect 96 213 184 255
rect 283 179 333 425
rect 582 255 625 393
rect 520 213 625 255
rect 107 145 341 179
rect 107 51 173 145
rect 275 51 341 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 331 81 493
rect 115 365 165 527
rect 199 459 425 493
rect 199 331 249 459
rect 17 289 249 331
rect 367 378 425 459
rect 367 289 418 378
rect 479 323 513 492
rect 555 429 605 527
rect 452 289 513 323
rect 452 249 486 289
rect 375 215 486 249
rect 443 179 486 215
rect 17 17 73 179
rect 207 17 241 111
rect 375 17 409 179
rect 443 145 513 179
rect 479 89 513 145
rect 555 17 606 169
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 520 213 625 255 6 A
port 1 nsew signal input
rlabel locali s 582 255 625 393 6 A
port 1 nsew signal input
rlabel locali s 96 213 184 255 6 SLEEP
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 2 21 443 67 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 2 67 631 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 275 51 341 145 6 X
port 7 nsew signal output
rlabel locali s 107 51 173 145 6 X
port 7 nsew signal output
rlabel locali s 107 145 341 179 6 X
port 7 nsew signal output
rlabel locali s 283 179 333 425 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2376910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2370968
<< end >>
