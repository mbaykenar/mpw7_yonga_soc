magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 367 47 397 177
rect 451 47 481 177
rect 535 47 565 177
<< scpmoshvt >>
rect 79 297 109 497
rect 151 297 181 497
rect 367 297 397 497
rect 451 297 481 497
rect 535 297 565 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 129 163 177
rect 109 95 119 129
rect 153 95 163 129
rect 109 47 163 95
rect 193 93 367 177
rect 193 59 203 93
rect 237 59 271 93
rect 305 59 367 93
rect 193 47 367 59
rect 397 129 451 177
rect 397 95 407 129
rect 441 95 451 129
rect 397 47 451 95
rect 481 47 535 177
rect 565 161 617 177
rect 565 127 575 161
rect 609 127 617 161
rect 565 93 617 127
rect 565 59 575 93
rect 609 59 617 93
rect 565 47 617 59
<< pdiff >>
rect 27 483 79 497
rect 27 449 35 483
rect 69 449 79 483
rect 27 415 79 449
rect 27 381 35 415
rect 69 381 79 415
rect 27 297 79 381
rect 109 297 151 497
rect 181 481 233 497
rect 181 447 191 481
rect 225 447 233 481
rect 181 413 233 447
rect 181 379 191 413
rect 225 379 233 413
rect 181 345 233 379
rect 181 311 191 345
rect 225 311 233 345
rect 181 297 233 311
rect 299 481 367 497
rect 299 447 307 481
rect 341 447 367 481
rect 299 413 367 447
rect 299 379 323 413
rect 357 379 367 413
rect 299 297 367 379
rect 397 481 451 497
rect 397 447 407 481
rect 441 447 451 481
rect 397 297 451 447
rect 481 489 535 497
rect 481 455 491 489
rect 525 455 535 489
rect 481 297 535 455
rect 565 477 617 497
rect 565 443 575 477
rect 609 443 617 477
rect 565 391 617 443
rect 565 357 575 391
rect 609 357 617 391
rect 565 297 617 357
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 95 153 129
rect 203 59 237 93
rect 271 59 305 93
rect 407 95 441 129
rect 575 127 609 161
rect 575 59 609 93
<< pdiffc >>
rect 35 449 69 483
rect 35 381 69 415
rect 191 447 225 481
rect 191 379 225 413
rect 191 311 225 345
rect 307 447 341 481
rect 323 379 357 413
rect 407 447 441 481
rect 491 455 525 489
rect 575 443 609 477
rect 575 357 609 391
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 367 497 397 523
rect 451 497 481 523
rect 535 497 565 523
rect 79 265 109 297
rect 55 249 109 265
rect 55 215 65 249
rect 99 215 109 249
rect 55 199 109 215
rect 151 265 181 297
rect 367 265 397 297
rect 451 265 481 297
rect 535 265 565 297
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 271 249 397 265
rect 271 215 282 249
rect 316 215 397 249
rect 271 199 397 215
rect 439 249 493 265
rect 439 215 449 249
rect 483 215 493 249
rect 439 199 493 215
rect 535 249 600 265
rect 535 215 556 249
rect 590 215 600 249
rect 535 199 600 215
rect 79 177 109 199
rect 163 177 193 199
rect 367 177 397 199
rect 451 177 481 199
rect 535 177 565 199
rect 79 21 109 47
rect 163 21 193 47
rect 367 21 397 47
rect 451 21 481 47
rect 535 21 565 47
<< polycont >>
rect 65 215 99 249
rect 161 215 195 249
rect 282 215 316 249
rect 449 215 483 249
rect 556 215 590 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 483 85 527
rect 19 449 35 483
rect 69 449 85 483
rect 19 415 85 449
rect 19 381 35 415
rect 69 381 85 415
rect 19 361 85 381
rect 175 481 241 493
rect 175 447 191 481
rect 225 447 241 481
rect 175 413 241 447
rect 175 379 191 413
rect 225 379 241 413
rect 175 345 241 379
rect 284 481 357 493
rect 284 447 307 481
rect 341 447 357 481
rect 391 481 457 493
rect 391 447 407 481
rect 441 447 457 481
rect 284 413 357 447
rect 284 379 323 413
rect 423 391 457 447
rect 491 489 541 527
rect 525 455 541 489
rect 491 427 541 455
rect 575 477 626 493
rect 609 443 626 477
rect 575 391 626 443
rect 357 379 389 391
rect 284 357 389 379
rect 423 357 575 391
rect 609 357 626 391
rect 30 249 104 323
rect 175 311 191 345
rect 225 323 241 345
rect 225 311 316 323
rect 175 289 316 311
rect 30 215 65 249
rect 99 215 104 249
rect 30 199 104 215
rect 145 249 248 255
rect 145 215 161 249
rect 195 215 248 249
rect 145 202 248 215
rect 282 249 316 289
rect 282 166 316 215
rect 19 161 85 165
rect 19 127 35 161
rect 69 127 85 161
rect 19 93 85 127
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 119 132 316 166
rect 355 165 389 357
rect 449 249 522 323
rect 483 215 522 249
rect 449 199 522 215
rect 556 249 614 323
rect 590 215 614 249
rect 556 199 614 215
rect 119 129 153 132
rect 355 129 441 165
rect 119 51 153 95
rect 187 93 321 98
rect 187 59 203 93
rect 237 59 271 93
rect 305 59 321 93
rect 187 17 321 59
rect 355 95 407 129
rect 355 51 441 95
rect 488 85 522 199
rect 559 161 625 165
rect 559 127 575 161
rect 609 127 625 161
rect 559 93 625 127
rect 559 59 575 93
rect 609 59 625 93
rect 559 17 625 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 304 425 338 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 304 357 338 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 396 85 430 119 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 488 85 522 119 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 488 153 522 187 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 488 221 522 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 488 289 522 323 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 580 221 614 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A2_N
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2bb2oi_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3915202
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3908354
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
