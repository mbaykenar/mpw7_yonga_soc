magic
tech sky130B
timestamp 1649977179
<< properties >>
string GDS_END 59022
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 58698
<< end >>
