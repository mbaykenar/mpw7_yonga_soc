magic
tech sky130B
magscale 12 1
timestamp 1598787041
<< metal5 >>
rect 0 90 45 105
rect 30 75 45 90
rect 0 60 45 75
rect 0 15 15 60
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
