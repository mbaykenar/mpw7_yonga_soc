magic
tech sky130A
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_0
timestamp 1649977179
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
flabel comment s -25 150 -25 150 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7185802
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7185028
<< end >>
