magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 4 21 367 203
rect 29 -17 63 21
<< locali >>
rect 19 337 74 491
rect 19 299 136 337
rect 19 135 67 265
rect 101 165 136 299
rect 170 199 253 265
rect 289 199 348 265
rect 101 129 167 165
rect 122 53 167 129
rect 207 75 253 199
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 108 405 174 491
rect 208 439 247 527
rect 283 405 349 491
rect 108 371 349 405
rect 170 305 349 371
rect 22 17 88 95
rect 289 17 349 163
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 207 75 253 199 6 A1
port 1 nsew signal input
rlabel locali s 170 199 253 265 6 A1
port 1 nsew signal input
rlabel locali s 289 199 348 265 6 A2
port 2 nsew signal input
rlabel locali s 19 135 67 265 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 4 21 367 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 122 53 167 129 6 Y
port 8 nsew signal output
rlabel locali s 101 129 167 165 6 Y
port 8 nsew signal output
rlabel locali s 101 165 136 299 6 Y
port 8 nsew signal output
rlabel locali s 19 299 136 337 6 Y
port 8 nsew signal output
rlabel locali s 19 337 74 491 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4042676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4038006
<< end >>
