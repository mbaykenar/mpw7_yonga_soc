magic
tech sky130B
magscale 12 1
timestamp 1598766739
<< metal5 >>
rect 0 90 15 105
rect 0 75 30 90
rect 45 75 60 105
rect 0 60 60 75
rect 0 0 15 60
rect 30 45 60 60
rect 45 0 60 45
<< properties >>
string FIXED_BBOX 0 -30 75 105
<< end >>
