magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< pwell >>
rect 10 10 462 230
<< nmoslvt >>
rect 92 36 122 204
rect 178 36 208 204
rect 264 36 294 204
rect 350 36 380 204
<< ndiff >>
rect 36 173 92 204
rect 36 139 47 173
rect 81 139 92 173
rect 36 101 92 139
rect 36 67 47 101
rect 81 67 92 101
rect 36 36 92 67
rect 122 173 178 204
rect 122 139 133 173
rect 167 139 178 173
rect 122 101 178 139
rect 122 67 133 101
rect 167 67 178 101
rect 122 36 178 67
rect 208 173 264 204
rect 208 139 219 173
rect 253 139 264 173
rect 208 101 264 139
rect 208 67 219 101
rect 253 67 264 101
rect 208 36 264 67
rect 294 173 350 204
rect 294 139 305 173
rect 339 139 350 173
rect 294 101 350 139
rect 294 67 305 101
rect 339 67 350 101
rect 294 36 350 67
rect 380 173 436 204
rect 380 139 391 173
rect 425 139 436 173
rect 380 101 436 139
rect 380 67 391 101
rect 425 67 436 101
rect 380 36 436 67
<< ndiffc >>
rect 47 139 81 173
rect 47 67 81 101
rect 133 139 167 173
rect 133 67 167 101
rect 219 139 253 173
rect 219 67 253 101
rect 305 139 339 173
rect 305 67 339 101
rect 391 139 425 173
rect 391 67 425 101
<< poly >>
rect 92 285 380 301
rect 92 251 117 285
rect 151 251 185 285
rect 219 251 253 285
rect 287 251 321 285
rect 355 251 380 285
rect 92 230 380 251
rect 92 204 122 230
rect 178 204 208 230
rect 264 204 294 230
rect 350 204 380 230
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
<< polycont >>
rect 117 251 151 285
rect 185 251 219 285
rect 253 251 287 285
rect 321 251 355 285
<< locali >>
rect 101 285 371 301
rect 101 251 111 285
rect 151 251 183 285
rect 219 251 253 285
rect 289 251 321 285
rect 361 251 371 285
rect 101 235 371 251
rect 47 173 81 189
rect 47 101 81 139
rect 47 51 81 67
rect 133 173 167 189
rect 133 101 167 139
rect 133 51 167 67
rect 219 173 253 189
rect 219 101 253 139
rect 219 51 253 67
rect 305 173 339 189
rect 305 101 339 139
rect 305 51 339 67
rect 391 173 425 189
rect 391 101 425 139
rect 391 51 425 67
<< viali >>
rect 111 251 117 285
rect 117 251 145 285
rect 183 251 185 285
rect 185 251 217 285
rect 255 251 287 285
rect 287 251 289 285
rect 327 251 355 285
rect 355 251 361 285
rect 47 139 81 173
rect 47 67 81 101
rect 133 139 167 173
rect 133 67 167 101
rect 219 139 253 173
rect 219 67 253 101
rect 305 139 339 173
rect 305 67 339 101
rect 391 139 425 173
rect 391 67 425 101
<< metal1 >>
rect 99 285 373 297
rect 99 251 111 285
rect 145 251 183 285
rect 217 251 255 285
rect 289 251 327 285
rect 361 251 373 285
rect 99 239 373 251
rect 41 173 87 189
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 124 175 176 189
rect 124 111 176 123
rect 124 51 176 59
rect 213 173 259 189
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 296 175 348 189
rect 296 111 348 123
rect 296 51 348 59
rect 385 173 431 189
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 41 -89 431 -29
<< via1 >>
rect 124 173 176 175
rect 124 139 133 173
rect 133 139 167 173
rect 167 139 176 173
rect 124 123 176 139
rect 124 101 176 111
rect 124 67 133 101
rect 133 67 167 101
rect 167 67 176 101
rect 124 59 176 67
rect 296 173 348 175
rect 296 139 305 173
rect 305 139 339 173
rect 339 139 348 173
rect 296 123 348 139
rect 296 101 348 111
rect 296 67 305 101
rect 305 67 339 101
rect 339 67 348 101
rect 296 59 348 67
<< metal2 >>
rect 117 186 183 195
rect 117 130 122 186
rect 178 130 183 186
rect 117 123 124 130
rect 176 123 183 130
rect 117 111 183 123
rect 117 106 124 111
rect 176 106 183 111
rect 117 50 122 106
rect 178 50 183 106
rect 117 41 183 50
rect 289 186 355 195
rect 289 130 294 186
rect 350 130 355 186
rect 289 123 296 130
rect 348 123 355 130
rect 289 111 355 123
rect 289 106 296 111
rect 348 106 355 111
rect 289 50 294 106
rect 350 50 355 106
rect 289 41 355 50
<< via2 >>
rect 122 175 178 186
rect 122 130 124 175
rect 124 130 176 175
rect 176 130 178 175
rect 122 59 124 106
rect 124 59 176 106
rect 176 59 178 106
rect 122 50 178 59
rect 294 175 350 186
rect 294 130 296 175
rect 296 130 348 175
rect 348 130 350 175
rect 294 59 296 106
rect 296 59 348 106
rect 348 59 350 106
rect 294 50 350 59
<< metal3 >>
rect 117 186 355 195
rect 117 130 122 186
rect 178 130 294 186
rect 350 130 355 186
rect 117 129 355 130
rect 117 106 183 129
rect 117 50 122 106
rect 178 50 183 106
rect 117 41 183 50
rect 289 106 355 129
rect 289 50 294 106
rect 350 50 355 106
rect 289 41 355 50
<< labels >>
flabel metal3 s 117 129 355 195 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 41 -89 431 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal1 s 99 239 373 297 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel pwell s 73 217 90 227 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 5864406
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5857248
string path 8.050 4.725 8.050 1.275 
<< end >>
