magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__dfl1sd__example_5595914180823  sky130_fd_pr__dfl1sd__example_5595914180823_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180823  sky130_fd_pr__dfl1sd__example_5595914180823_1
timestamp 1649977179
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 63 128 63 0 FreeSans 300 0 0 0 D
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7860112
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7859062
<< end >>
