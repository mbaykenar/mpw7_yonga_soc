magic
tech sky130B
magscale 1 2
timestamp 1662552612
<< obsli1 >>
rect 1104 2159 48852 27761
<< obsm1 >>
rect 14 2128 49666 27792
<< metal2 >>
rect 18 29200 74 30000
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 1950 29200 2006 30000
rect 2594 29200 2650 30000
rect 3238 29200 3294 30000
rect 3882 29200 3938 30000
rect 4526 29200 4582 30000
rect 5170 29200 5226 30000
rect 5814 29200 5870 30000
rect 6458 29200 6514 30000
rect 7102 29200 7158 30000
rect 7746 29200 7802 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 9678 29200 9734 30000
rect 10322 29200 10378 30000
rect 10966 29200 11022 30000
rect 11610 29200 11666 30000
rect 12254 29200 12310 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14186 29200 14242 30000
rect 14830 29200 14886 30000
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 16762 29200 16818 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 18694 29200 18750 30000
rect 19338 29200 19394 30000
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21270 29200 21326 30000
rect 21914 29200 21970 30000
rect 22558 29200 22614 30000
rect 23202 29200 23258 30000
rect 23846 29200 23902 30000
rect 24490 29200 24546 30000
rect 25134 29200 25190 30000
rect 25778 29200 25834 30000
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 27710 29200 27766 30000
rect 28354 29200 28410 30000
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 30286 29200 30342 30000
rect 30930 29200 30986 30000
rect 31574 29200 31630 30000
rect 32218 29200 32274 30000
rect 32862 29200 32918 30000
rect 33506 29200 33562 30000
rect 34150 29200 34206 30000
rect 34794 29200 34850 30000
rect 35438 29200 35494 30000
rect 36082 29200 36138 30000
rect 36726 29200 36782 30000
rect 37370 29200 37426 30000
rect 38014 29200 38070 30000
rect 38658 29200 38714 30000
rect 39302 29200 39358 30000
rect 39946 29200 40002 30000
rect 40590 29200 40646 30000
rect 41234 29200 41290 30000
rect 41878 29200 41934 30000
rect 42522 29200 42578 30000
rect 43166 29200 43222 30000
rect 43810 29200 43866 30000
rect 44454 29200 44510 30000
rect 45098 29200 45154 30000
rect 45742 29200 45798 30000
rect 46386 29200 46442 30000
rect 47030 29200 47086 30000
rect 47674 29200 47730 30000
rect 48318 29200 48374 30000
rect 48962 29200 49018 30000
rect 49606 29200 49662 30000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
<< obsm2 >>
rect 130 29144 606 29345
rect 774 29144 1250 29345
rect 1418 29144 1894 29345
rect 2062 29144 2538 29345
rect 2706 29144 3182 29345
rect 3350 29144 3826 29345
rect 3994 29144 4470 29345
rect 4638 29144 5114 29345
rect 5282 29144 5758 29345
rect 5926 29144 6402 29345
rect 6570 29144 7046 29345
rect 7214 29144 7690 29345
rect 7858 29144 8334 29345
rect 8502 29144 8978 29345
rect 9146 29144 9622 29345
rect 9790 29144 10266 29345
rect 10434 29144 10910 29345
rect 11078 29144 11554 29345
rect 11722 29144 12198 29345
rect 12366 29144 12842 29345
rect 13010 29144 13486 29345
rect 13654 29144 14130 29345
rect 14298 29144 14774 29345
rect 14942 29144 15418 29345
rect 15586 29144 16062 29345
rect 16230 29144 16706 29345
rect 16874 29144 17350 29345
rect 17518 29144 17994 29345
rect 18162 29144 18638 29345
rect 18806 29144 19282 29345
rect 19450 29144 19926 29345
rect 20094 29144 20570 29345
rect 20738 29144 21214 29345
rect 21382 29144 21858 29345
rect 22026 29144 22502 29345
rect 22670 29144 23146 29345
rect 23314 29144 23790 29345
rect 23958 29144 24434 29345
rect 24602 29144 25078 29345
rect 25246 29144 25722 29345
rect 25890 29144 26366 29345
rect 26534 29144 27010 29345
rect 27178 29144 27654 29345
rect 27822 29144 28298 29345
rect 28466 29144 28942 29345
rect 29110 29144 29586 29345
rect 29754 29144 30230 29345
rect 30398 29144 30874 29345
rect 31042 29144 31518 29345
rect 31686 29144 32162 29345
rect 32330 29144 32806 29345
rect 32974 29144 33450 29345
rect 33618 29144 34094 29345
rect 34262 29144 34738 29345
rect 34906 29144 35382 29345
rect 35550 29144 36026 29345
rect 36194 29144 36670 29345
rect 36838 29144 37314 29345
rect 37482 29144 37958 29345
rect 38126 29144 38602 29345
rect 38770 29144 39246 29345
rect 39414 29144 39890 29345
rect 40058 29144 40534 29345
rect 40702 29144 41178 29345
rect 41346 29144 41822 29345
rect 41990 29144 42466 29345
rect 42634 29144 43110 29345
rect 43278 29144 43754 29345
rect 43922 29144 44398 29345
rect 44566 29144 45042 29345
rect 45210 29144 45686 29345
rect 45854 29144 46330 29345
rect 46498 29144 46974 29345
rect 47142 29144 47618 29345
rect 47786 29144 48262 29345
rect 48430 29144 48906 29345
rect 49074 29144 49550 29345
rect 20 856 49660 29144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
rect 39414 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41178 856
rect 41346 31 41822 856
rect 41990 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45042 856
rect 45210 31 45686 856
rect 45854 31 46330 856
rect 46498 31 46974 856
rect 47142 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 49550 856
<< metal3 >>
rect 0 29248 800 29368
rect 49200 29248 50000 29368
rect 0 28568 800 28688
rect 49200 28568 50000 28688
rect 0 27888 800 28008
rect 49200 27888 50000 28008
rect 0 27208 800 27328
rect 49200 27208 50000 27328
rect 0 26528 800 26648
rect 49200 26528 50000 26648
rect 0 25848 800 25968
rect 49200 25848 50000 25968
rect 0 25168 800 25288
rect 49200 25168 50000 25288
rect 0 24488 800 24608
rect 49200 24488 50000 24608
rect 0 23808 800 23928
rect 49200 23808 50000 23928
rect 0 23128 800 23248
rect 49200 23128 50000 23248
rect 0 22448 800 22568
rect 49200 22448 50000 22568
rect 0 21768 800 21888
rect 49200 21768 50000 21888
rect 0 21088 800 21208
rect 49200 21088 50000 21208
rect 0 20408 800 20528
rect 49200 20408 50000 20528
rect 0 19728 800 19848
rect 49200 19728 50000 19848
rect 0 19048 800 19168
rect 49200 19048 50000 19168
rect 0 18368 800 18488
rect 49200 18368 50000 18488
rect 0 17688 800 17808
rect 49200 17688 50000 17808
rect 0 17008 800 17128
rect 49200 17008 50000 17128
rect 0 16328 800 16448
rect 49200 16328 50000 16448
rect 0 15648 800 15768
rect 49200 15648 50000 15768
rect 0 14968 800 15088
rect 49200 14968 50000 15088
rect 0 14288 800 14408
rect 49200 14288 50000 14408
rect 0 13608 800 13728
rect 49200 13608 50000 13728
rect 0 12928 800 13048
rect 49200 12928 50000 13048
rect 0 12248 800 12368
rect 49200 12248 50000 12368
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 0 10888 800 11008
rect 49200 10888 50000 11008
rect 0 10208 800 10328
rect 49200 10208 50000 10328
rect 0 9528 800 9648
rect 49200 9528 50000 9648
rect 0 8848 800 8968
rect 49200 8848 50000 8968
rect 0 8168 800 8288
rect 49200 8168 50000 8288
rect 0 7488 800 7608
rect 49200 7488 50000 7608
rect 0 6808 800 6928
rect 49200 6808 50000 6928
rect 0 6128 800 6248
rect 49200 6128 50000 6248
rect 0 5448 800 5568
rect 49200 5448 50000 5568
rect 0 4768 800 4888
rect 49200 4768 50000 4888
rect 0 4088 800 4208
rect 49200 4088 50000 4208
rect 0 3408 800 3528
rect 49200 3408 50000 3528
rect 0 2728 800 2848
rect 49200 2728 50000 2848
rect 0 2048 800 2168
rect 49200 2048 50000 2168
rect 0 1368 800 1488
rect 49200 1368 50000 1488
rect 0 688 800 808
rect 49200 688 50000 808
rect 0 8 800 128
rect 49200 8 50000 128
<< obsm3 >>
rect 880 29168 49120 29341
rect 800 28768 49200 29168
rect 880 28488 49120 28768
rect 800 28088 49200 28488
rect 880 27808 49120 28088
rect 800 27408 49200 27808
rect 880 27128 49120 27408
rect 800 26728 49200 27128
rect 880 26448 49120 26728
rect 800 26048 49200 26448
rect 880 25768 49120 26048
rect 800 25368 49200 25768
rect 880 25088 49120 25368
rect 800 24688 49200 25088
rect 880 24408 49120 24688
rect 800 24008 49200 24408
rect 880 23728 49120 24008
rect 800 23328 49200 23728
rect 880 23048 49120 23328
rect 800 22648 49200 23048
rect 880 22368 49120 22648
rect 800 21968 49200 22368
rect 880 21688 49120 21968
rect 800 21288 49200 21688
rect 880 21008 49120 21288
rect 800 20608 49200 21008
rect 880 20328 49120 20608
rect 800 19928 49200 20328
rect 880 19648 49120 19928
rect 800 19248 49200 19648
rect 880 18968 49120 19248
rect 800 18568 49200 18968
rect 880 18288 49120 18568
rect 800 17888 49200 18288
rect 880 17608 49120 17888
rect 800 17208 49200 17608
rect 880 16928 49120 17208
rect 800 16528 49200 16928
rect 880 16248 49120 16528
rect 800 15848 49200 16248
rect 880 15568 49120 15848
rect 800 15168 49200 15568
rect 880 14888 49120 15168
rect 800 14488 49200 14888
rect 880 14208 49120 14488
rect 800 13808 49200 14208
rect 880 13528 49120 13808
rect 800 13128 49200 13528
rect 880 12848 49120 13128
rect 800 12448 49200 12848
rect 880 12168 49120 12448
rect 800 11768 49200 12168
rect 880 11488 49120 11768
rect 800 11088 49200 11488
rect 880 10808 49120 11088
rect 800 10408 49200 10808
rect 880 10128 49120 10408
rect 800 9728 49200 10128
rect 880 9448 49120 9728
rect 800 9048 49200 9448
rect 880 8768 49120 9048
rect 800 8368 49200 8768
rect 880 8088 49120 8368
rect 800 7688 49200 8088
rect 880 7408 49120 7688
rect 800 7008 49200 7408
rect 880 6728 49120 7008
rect 800 6328 49200 6728
rect 880 6048 49120 6328
rect 800 5648 49200 6048
rect 880 5368 49120 5648
rect 800 4968 49200 5368
rect 880 4688 49120 4968
rect 800 4288 49200 4688
rect 880 4008 49120 4288
rect 800 3608 49200 4008
rect 880 3328 49120 3608
rect 800 2928 49200 3328
rect 880 2648 49120 2928
rect 800 2248 49200 2648
rect 880 1968 49120 2248
rect 800 1568 49200 1968
rect 880 1288 49120 1568
rect 800 888 49200 1288
rect 880 608 49120 888
rect 800 208 49200 608
rect 880 35 49120 208
<< metal4 >>
rect 6918 2128 7238 27792
rect 12892 2128 13212 27792
rect 18866 2128 19186 27792
rect 24840 2128 25160 27792
rect 30814 2128 31134 27792
rect 36788 2128 37108 27792
rect 42762 2128 43082 27792
<< labels >>
rlabel metal3 s 49200 14968 50000 15088 6 clk_i
port 1 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 clk_o
port 2 nsew signal output
rlabel metal2 s 4526 29200 4582 30000 6 clk_sel_i
port 3 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 clk_standalone_i
port 4 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 fll_ack_o
port 5 nsew signal output
rlabel metal3 s 49200 29248 50000 29368 6 fll_add_i[0]
port 6 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 fll_add_i[1]
port 7 nsew signal input
rlabel metal2 s 16762 29200 16818 30000 6 fll_data_i[0]
port 8 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 fll_data_i[10]
port 9 nsew signal input
rlabel metal2 s 3238 29200 3294 30000 6 fll_data_i[11]
port 10 nsew signal input
rlabel metal3 s 49200 21088 50000 21208 6 fll_data_i[12]
port 11 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 fll_data_i[13]
port 12 nsew signal input
rlabel metal2 s 32862 29200 32918 30000 6 fll_data_i[14]
port 13 nsew signal input
rlabel metal2 s 14186 29200 14242 30000 6 fll_data_i[15]
port 14 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 fll_data_i[16]
port 15 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 fll_data_i[17]
port 16 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 fll_data_i[18]
port 17 nsew signal input
rlabel metal2 s 31574 29200 31630 30000 6 fll_data_i[19]
port 18 nsew signal input
rlabel metal2 s 27066 29200 27122 30000 6 fll_data_i[1]
port 19 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 fll_data_i[20]
port 20 nsew signal input
rlabel metal3 s 49200 10208 50000 10328 6 fll_data_i[21]
port 21 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 fll_data_i[22]
port 22 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 fll_data_i[23]
port 23 nsew signal input
rlabel metal3 s 49200 10888 50000 11008 6 fll_data_i[24]
port 24 nsew signal input
rlabel metal2 s 39302 29200 39358 30000 6 fll_data_i[25]
port 25 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 fll_data_i[26]
port 26 nsew signal input
rlabel metal2 s 44454 29200 44510 30000 6 fll_data_i[27]
port 27 nsew signal input
rlabel metal2 s 2594 29200 2650 30000 6 fll_data_i[28]
port 28 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 fll_data_i[29]
port 29 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 fll_data_i[2]
port 30 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 fll_data_i[30]
port 31 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 fll_data_i[31]
port 32 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 fll_data_i[3]
port 33 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 fll_data_i[4]
port 34 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 fll_data_i[5]
port 35 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 fll_data_i[6]
port 36 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 fll_data_i[7]
port 37 nsew signal input
rlabel metal2 s 29642 29200 29698 30000 6 fll_data_i[8]
port 38 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 fll_data_i[9]
port 39 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 fll_lock_o
port 40 nsew signal output
rlabel metal3 s 49200 12248 50000 12368 6 fll_r_data_o[0]
port 41 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 fll_r_data_o[10]
port 42 nsew signal output
rlabel metal2 s 5170 29200 5226 30000 6 fll_r_data_o[11]
port 43 nsew signal output
rlabel metal2 s 30930 29200 30986 30000 6 fll_r_data_o[12]
port 44 nsew signal output
rlabel metal3 s 49200 4768 50000 4888 6 fll_r_data_o[13]
port 45 nsew signal output
rlabel metal3 s 49200 4088 50000 4208 6 fll_r_data_o[14]
port 46 nsew signal output
rlabel metal3 s 49200 15648 50000 15768 6 fll_r_data_o[15]
port 47 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 fll_r_data_o[16]
port 48 nsew signal output
rlabel metal2 s 46386 29200 46442 30000 6 fll_r_data_o[17]
port 49 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 fll_r_data_o[18]
port 50 nsew signal output
rlabel metal3 s 49200 17008 50000 17128 6 fll_r_data_o[19]
port 51 nsew signal output
rlabel metal2 s 26422 29200 26478 30000 6 fll_r_data_o[1]
port 52 nsew signal output
rlabel metal2 s 18694 29200 18750 30000 6 fll_r_data_o[20]
port 53 nsew signal output
rlabel metal2 s 6458 29200 6514 30000 6 fll_r_data_o[21]
port 54 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 fll_r_data_o[22]
port 55 nsew signal output
rlabel metal2 s 43166 29200 43222 30000 6 fll_r_data_o[23]
port 56 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 fll_r_data_o[24]
port 57 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 fll_r_data_o[25]
port 58 nsew signal output
rlabel metal3 s 49200 26528 50000 26648 6 fll_r_data_o[26]
port 59 nsew signal output
rlabel metal2 s 1950 29200 2006 30000 6 fll_r_data_o[27]
port 60 nsew signal output
rlabel metal2 s 41234 29200 41290 30000 6 fll_r_data_o[28]
port 61 nsew signal output
rlabel metal2 s 20626 29200 20682 30000 6 fll_r_data_o[29]
port 62 nsew signal output
rlabel metal3 s 49200 23808 50000 23928 6 fll_r_data_o[2]
port 63 nsew signal output
rlabel metal2 s 32218 29200 32274 30000 6 fll_r_data_o[30]
port 64 nsew signal output
rlabel metal3 s 49200 9528 50000 9648 6 fll_r_data_o[31]
port 65 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 fll_r_data_o[3]
port 66 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 fll_r_data_o[4]
port 67 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 fll_r_data_o[5]
port 68 nsew signal output
rlabel metal3 s 49200 20408 50000 20528 6 fll_r_data_o[6]
port 69 nsew signal output
rlabel metal2 s 10966 29200 11022 30000 6 fll_r_data_o[7]
port 70 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 fll_r_data_o[8]
port 71 nsew signal output
rlabel metal2 s 18050 29200 18106 30000 6 fll_r_data_o[9]
port 72 nsew signal output
rlabel metal2 s 42522 29200 42578 30000 6 fll_req_i
port 73 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 fll_wrn_i
port 74 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 io_oeb[0]
port 75 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 io_oeb[10]
port 76 nsew signal output
rlabel metal2 s 28998 29200 29054 30000 6 io_oeb[11]
port 77 nsew signal output
rlabel metal2 s 35438 29200 35494 30000 6 io_oeb[12]
port 78 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 io_oeb[13]
port 79 nsew signal output
rlabel metal2 s 34794 29200 34850 30000 6 io_oeb[14]
port 80 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_oeb[15]
port 81 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 io_oeb[16]
port 82 nsew signal output
rlabel metal2 s 40590 29200 40646 30000 6 io_oeb[17]
port 83 nsew signal output
rlabel metal2 s 1306 29200 1362 30000 6 io_oeb[18]
port 84 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 io_oeb[19]
port 85 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 io_oeb[1]
port 86 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 io_oeb[20]
port 87 nsew signal output
rlabel metal3 s 49200 25848 50000 25968 6 io_oeb[21]
port 88 nsew signal output
rlabel metal3 s 49200 2728 50000 2848 6 io_oeb[22]
port 89 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 io_oeb[23]
port 90 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 io_oeb[24]
port 91 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 io_oeb[25]
port 92 nsew signal output
rlabel metal2 s 21914 29200 21970 30000 6 io_oeb[26]
port 93 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 io_oeb[27]
port 94 nsew signal output
rlabel metal3 s 49200 11568 50000 11688 6 io_oeb[28]
port 95 nsew signal output
rlabel metal2 s 45742 29200 45798 30000 6 io_oeb[29]
port 96 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 io_oeb[2]
port 97 nsew signal output
rlabel metal3 s 49200 688 50000 808 6 io_oeb[30]
port 98 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_oeb[31]
port 99 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_oeb[32]
port 100 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 io_oeb[33]
port 101 nsew signal output
rlabel metal2 s 23202 29200 23258 30000 6 io_oeb[34]
port 102 nsew signal output
rlabel metal2 s 47674 29200 47730 30000 6 io_oeb[35]
port 103 nsew signal output
rlabel metal2 s 33506 29200 33562 30000 6 io_oeb[36]
port 104 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_oeb[37]
port 105 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 io_oeb[3]
port 106 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_oeb[4]
port 107 nsew signal output
rlabel metal2 s 7102 29200 7158 30000 6 io_oeb[5]
port 108 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_oeb[6]
port 109 nsew signal output
rlabel metal3 s 49200 6808 50000 6928 6 io_oeb[7]
port 110 nsew signal output
rlabel metal2 s 662 29200 718 30000 6 io_oeb[8]
port 111 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_oeb[9]
port 112 nsew signal output
rlabel metal2 s 11610 29200 11666 30000 6 io_out[0]
port 113 nsew signal output
rlabel metal2 s 27710 29200 27766 30000 6 io_out[10]
port 114 nsew signal output
rlabel metal3 s 49200 27208 50000 27328 6 io_out[11]
port 115 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[12]
port 116 nsew signal output
rlabel metal2 s 22558 29200 22614 30000 6 io_out[13]
port 117 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 io_out[14]
port 118 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 io_out[15]
port 119 nsew signal output
rlabel metal2 s 23846 29200 23902 30000 6 io_out[16]
port 120 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 io_out[17]
port 121 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 io_out[18]
port 122 nsew signal output
rlabel metal3 s 0 8 800 128 6 io_out[19]
port 123 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 io_out[1]
port 124 nsew signal output
rlabel metal3 s 49200 18368 50000 18488 6 io_out[20]
port 125 nsew signal output
rlabel metal2 s 28354 29200 28410 30000 6 io_out[21]
port 126 nsew signal output
rlabel metal2 s 49606 29200 49662 30000 6 io_out[22]
port 127 nsew signal output
rlabel metal2 s 9678 29200 9734 30000 6 io_out[23]
port 128 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 io_out[24]
port 129 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 io_out[25]
port 130 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 io_out[2]
port 131 nsew signal output
rlabel metal2 s 12898 29200 12954 30000 6 io_out[3]
port 132 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_out[4]
port 133 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_out[5]
port 134 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 io_out[6]
port 135 nsew signal output
rlabel metal2 s 12254 29200 12310 30000 6 io_out[7]
port 136 nsew signal output
rlabel metal2 s 47030 29200 47086 30000 6 io_out[8]
port 137 nsew signal output
rlabel metal2 s 48962 29200 49018 30000 6 io_out[9]
port 138 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[0]
port 139 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out[10]
port 140 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[11]
port 141 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 la_data_out[12]
port 142 nsew signal output
rlabel metal3 s 49200 28568 50000 28688 6 la_data_out[13]
port 143 nsew signal output
rlabel metal2 s 38658 29200 38714 30000 6 la_data_out[14]
port 144 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 la_data_out[15]
port 145 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 la_data_out[16]
port 146 nsew signal output
rlabel metal3 s 49200 3408 50000 3528 6 la_data_out[17]
port 147 nsew signal output
rlabel metal2 s 24490 29200 24546 30000 6 la_data_out[18]
port 148 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_data_out[19]
port 149 nsew signal output
rlabel metal3 s 49200 8 50000 128 6 la_data_out[1]
port 150 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_data_out[20]
port 151 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[21]
port 152 nsew signal output
rlabel metal3 s 49200 25168 50000 25288 6 la_data_out[22]
port 153 nsew signal output
rlabel metal3 s 49200 16328 50000 16448 6 la_data_out[23]
port 154 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 la_data_out[24]
port 155 nsew signal output
rlabel metal2 s 14830 29200 14886 30000 6 la_data_out[25]
port 156 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[26]
port 157 nsew signal output
rlabel metal2 s 36082 29200 36138 30000 6 la_data_out[27]
port 158 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out[28]
port 159 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 la_data_out[29]
port 160 nsew signal output
rlabel metal2 s 41878 29200 41934 30000 6 la_data_out[2]
port 161 nsew signal output
rlabel metal3 s 49200 1368 50000 1488 6 la_data_out[30]
port 162 nsew signal output
rlabel metal3 s 49200 14288 50000 14408 6 la_data_out[31]
port 163 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 la_data_out[32]
port 164 nsew signal output
rlabel metal3 s 49200 23128 50000 23248 6 la_data_out[33]
port 165 nsew signal output
rlabel metal2 s 5814 29200 5870 30000 6 la_data_out[34]
port 166 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 la_data_out[35]
port 167 nsew signal output
rlabel metal3 s 49200 24488 50000 24608 6 la_data_out[36]
port 168 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[37]
port 169 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 la_data_out[38]
port 170 nsew signal output
rlabel metal2 s 13542 29200 13598 30000 6 la_data_out[39]
port 171 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out[3]
port 172 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[40]
port 173 nsew signal output
rlabel metal2 s 38014 29200 38070 30000 6 la_data_out[41]
port 174 nsew signal output
rlabel metal3 s 49200 13608 50000 13728 6 la_data_out[42]
port 175 nsew signal output
rlabel metal2 s 19338 29200 19394 30000 6 la_data_out[43]
port 176 nsew signal output
rlabel metal2 s 21270 29200 21326 30000 6 la_data_out[44]
port 177 nsew signal output
rlabel metal2 s 19982 29200 20038 30000 6 la_data_out[45]
port 178 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 la_data_out[46]
port 179 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 la_data_out[47]
port 180 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 la_data_out[48]
port 181 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la_data_out[49]
port 182 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 la_data_out[4]
port 183 nsew signal output
rlabel metal2 s 7746 29200 7802 30000 6 la_data_out[50]
port 184 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 la_data_out[51]
port 185 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 la_data_out[52]
port 186 nsew signal output
rlabel metal3 s 49200 6128 50000 6248 6 la_data_out[53]
port 187 nsew signal output
rlabel metal3 s 49200 22448 50000 22568 6 la_data_out[54]
port 188 nsew signal output
rlabel metal2 s 9034 29200 9090 30000 6 la_data_out[55]
port 189 nsew signal output
rlabel metal3 s 49200 12928 50000 13048 6 la_data_out[56]
port 190 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[57]
port 191 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 la_data_out[58]
port 192 nsew signal output
rlabel metal3 s 49200 27888 50000 28008 6 la_data_out[59]
port 193 nsew signal output
rlabel metal2 s 30286 29200 30342 30000 6 la_data_out[5]
port 194 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 la_data_out[60]
port 195 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 la_data_out[61]
port 196 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 la_data_out[62]
port 197 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[63]
port 198 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_data_out[6]
port 199 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[7]
port 200 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 la_data_out[8]
port 201 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 la_data_out[9]
port 202 nsew signal output
rlabel metal3 s 49200 2048 50000 2168 6 rstn_i
port 203 nsew signal input
rlabel metal2 s 48318 29200 48374 30000 6 rstn_o
port 204 nsew signal output
rlabel metal3 s 49200 19728 50000 19848 6 scan_en_i
port 205 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 scan_i
port 206 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 scan_o
port 207 nsew signal output
rlabel metal3 s 49200 7488 50000 7608 6 testmode_i
port 208 nsew signal input
rlabel metal2 s 662 0 718 800 6 user_irq[0]
port 209 nsew signal output
rlabel metal3 s 49200 21768 50000 21888 6 user_irq[1]
port 210 nsew signal output
rlabel metal2 s 45098 29200 45154 30000 6 user_irq[2]
port 211 nsew signal output
rlabel metal4 s 6918 2128 7238 27792 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 18866 2128 19186 27792 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 30814 2128 31134 27792 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 42762 2128 43082 27792 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 12892 2128 13212 27792 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 24840 2128 25160 27792 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 36788 2128 37108 27792 6 vssd1
port 213 nsew ground bidirectional
rlabel metal2 s 41234 0 41290 800 6 wbs_ack_o
port 214 nsew signal output
rlabel metal2 s 43810 29200 43866 30000 6 wbs_dat_o[0]
port 215 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 wbs_dat_o[10]
port 216 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 wbs_dat_o[11]
port 217 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[12]
port 218 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[13]
port 219 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[14]
port 220 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_o[15]
port 221 nsew signal output
rlabel metal2 s 10322 29200 10378 30000 6 wbs_dat_o[16]
port 222 nsew signal output
rlabel metal2 s 25778 29200 25834 30000 6 wbs_dat_o[17]
port 223 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_o[18]
port 224 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_o[19]
port 225 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_o[1]
port 226 nsew signal output
rlabel metal2 s 34150 29200 34206 30000 6 wbs_dat_o[20]
port 227 nsew signal output
rlabel metal2 s 25134 29200 25190 30000 6 wbs_dat_o[21]
port 228 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[22]
port 229 nsew signal output
rlabel metal2 s 39946 29200 40002 30000 6 wbs_dat_o[23]
port 230 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_o[24]
port 231 nsew signal output
rlabel metal2 s 18 29200 74 30000 6 wbs_dat_o[25]
port 232 nsew signal output
rlabel metal3 s 49200 19048 50000 19168 6 wbs_dat_o[26]
port 233 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[27]
port 234 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[28]
port 235 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 wbs_dat_o[29]
port 236 nsew signal output
rlabel metal3 s 49200 17688 50000 17808 6 wbs_dat_o[2]
port 237 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[30]
port 238 nsew signal output
rlabel metal2 s 37370 29200 37426 30000 6 wbs_dat_o[31]
port 239 nsew signal output
rlabel metal2 s 36726 29200 36782 30000 6 wbs_dat_o[3]
port 240 nsew signal output
rlabel metal2 s 8390 29200 8446 30000 6 wbs_dat_o[4]
port 241 nsew signal output
rlabel metal2 s 15474 29200 15530 30000 6 wbs_dat_o[5]
port 242 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[6]
port 243 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 wbs_dat_o[7]
port 244 nsew signal output
rlabel metal2 s 3882 29200 3938 30000 6 wbs_dat_o[8]
port 245 nsew signal output
rlabel metal3 s 49200 8848 50000 8968 6 wbs_dat_o[9]
port 246 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 50000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 756922
string GDS_FILE /home/mbaykenar/Desktop/workspace/mpw7_yonga_soc/openlane/clk_rst_gen/runs/22_09_07_15_09/results/signoff/clk_rst_gen.magic.gds
string GDS_START 87268
<< end >>

