magic
tech sky130A
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1649977179
transform -1 0 -14 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_1
timestamp 1649977179
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
flabel comment s -42 97 -42 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7391320
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7390202
<< end >>
