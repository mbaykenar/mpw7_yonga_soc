magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -71 728 917 742
rect -71 10 919 728
rect 1114 -948 1386 -492
<< pwell >>
rect 1327 1915 1413 1936
rect -43 1911 43 1913
rect 698 1911 2065 1915
rect -43 1353 2065 1911
rect 4 1263 2065 1353
rect 4 1011 2049 1263
rect 4 964 464 1011
rect 1435 919 2049 1011
rect 980 55 1367 707
rect 1630 -1302 1950 -1050
<< nmos >>
rect 1712 -1276 1762 -1076
rect 1818 -1276 1868 -1076
<< mvnmos >>
rect 1514 1289 1634 1889
rect 1690 1289 1810 1889
rect 1866 1289 1986 1889
rect 86 990 206 1190
rect 262 990 382 1190
rect 1514 945 1714 1095
rect 1770 945 1970 1095
rect 1168 81 1288 681
<< mvpmos >>
rect 130 526 230 676
rect 130 207 230 357
rect 396 76 516 676
rect 572 76 692 676
<< mvnnmos >>
rect 181 1685 361 1885
rect 417 1685 597 1885
rect 777 1689 957 1889
rect 1013 1689 1193 1889
rect 181 1391 361 1591
rect 417 1391 597 1591
rect 777 1391 957 1591
rect 1013 1391 1193 1591
<< pmoshvt >>
rect 1150 -721 1350 -671
rect 1150 -827 1350 -777
<< nmoslvt >>
rect 648 1037 678 1237
rect 734 1037 764 1237
rect 820 1037 850 1237
rect 906 1037 936 1237
rect 992 1037 1022 1237
rect 1078 1037 1108 1237
rect 1164 1037 1194 1237
rect 1250 1037 1280 1237
<< ndiff >>
rect 592 1225 648 1237
rect 592 1191 603 1225
rect 637 1191 648 1225
rect 592 1157 648 1191
rect 592 1123 603 1157
rect 637 1123 648 1157
rect 592 1089 648 1123
rect 592 1055 603 1089
rect 637 1055 648 1089
rect 592 1037 648 1055
rect 678 1225 734 1237
rect 678 1191 689 1225
rect 723 1191 734 1225
rect 678 1157 734 1191
rect 678 1123 689 1157
rect 723 1123 734 1157
rect 678 1089 734 1123
rect 678 1055 689 1089
rect 723 1055 734 1089
rect 678 1037 734 1055
rect 764 1225 820 1237
rect 764 1191 775 1225
rect 809 1191 820 1225
rect 764 1157 820 1191
rect 764 1123 775 1157
rect 809 1123 820 1157
rect 764 1089 820 1123
rect 764 1055 775 1089
rect 809 1055 820 1089
rect 764 1037 820 1055
rect 850 1225 906 1237
rect 850 1191 861 1225
rect 895 1191 906 1225
rect 850 1157 906 1191
rect 850 1123 861 1157
rect 895 1123 906 1157
rect 850 1089 906 1123
rect 850 1055 861 1089
rect 895 1055 906 1089
rect 850 1037 906 1055
rect 936 1225 992 1237
rect 936 1191 947 1225
rect 981 1191 992 1225
rect 936 1157 992 1191
rect 936 1123 947 1157
rect 981 1123 992 1157
rect 936 1089 992 1123
rect 936 1055 947 1089
rect 981 1055 992 1089
rect 936 1037 992 1055
rect 1022 1225 1078 1237
rect 1022 1191 1033 1225
rect 1067 1191 1078 1225
rect 1022 1157 1078 1191
rect 1022 1123 1033 1157
rect 1067 1123 1078 1157
rect 1022 1089 1078 1123
rect 1022 1055 1033 1089
rect 1067 1055 1078 1089
rect 1022 1037 1078 1055
rect 1108 1225 1164 1237
rect 1108 1191 1119 1225
rect 1153 1191 1164 1225
rect 1108 1157 1164 1191
rect 1108 1123 1119 1157
rect 1153 1123 1164 1157
rect 1108 1089 1164 1123
rect 1108 1055 1119 1089
rect 1153 1055 1164 1089
rect 1108 1037 1164 1055
rect 1194 1225 1250 1237
rect 1194 1191 1205 1225
rect 1239 1191 1250 1225
rect 1194 1157 1250 1191
rect 1194 1123 1205 1157
rect 1239 1123 1250 1157
rect 1194 1089 1250 1123
rect 1194 1055 1205 1089
rect 1239 1055 1250 1089
rect 1194 1037 1250 1055
rect 1280 1225 1333 1237
rect 1280 1191 1291 1225
rect 1325 1191 1333 1225
rect 1280 1157 1333 1191
rect 1280 1123 1291 1157
rect 1325 1123 1333 1157
rect 1280 1089 1333 1123
rect 1280 1055 1291 1089
rect 1325 1055 1333 1089
rect 1280 1037 1333 1055
rect 1656 -1094 1712 -1076
rect 1656 -1128 1667 -1094
rect 1701 -1128 1712 -1094
rect 1656 -1162 1712 -1128
rect 1656 -1196 1667 -1162
rect 1701 -1196 1712 -1162
rect 1656 -1230 1712 -1196
rect 1656 -1264 1667 -1230
rect 1701 -1264 1712 -1230
rect 1656 -1276 1712 -1264
rect 1762 -1094 1818 -1076
rect 1762 -1128 1773 -1094
rect 1807 -1128 1818 -1094
rect 1762 -1162 1818 -1128
rect 1762 -1196 1773 -1162
rect 1807 -1196 1818 -1162
rect 1762 -1230 1818 -1196
rect 1762 -1264 1773 -1230
rect 1807 -1264 1818 -1230
rect 1762 -1276 1818 -1264
rect 1868 -1094 1924 -1076
rect 1868 -1128 1879 -1094
rect 1913 -1128 1924 -1094
rect 1868 -1162 1924 -1128
rect 1868 -1196 1879 -1162
rect 1913 -1196 1924 -1162
rect 1868 -1230 1924 -1196
rect 1868 -1264 1879 -1230
rect 1913 -1264 1924 -1230
rect 1868 -1276 1924 -1264
<< pdiff >>
rect 1150 -626 1350 -618
rect 1150 -660 1168 -626
rect 1202 -660 1236 -626
rect 1270 -660 1304 -626
rect 1338 -660 1350 -626
rect 1150 -671 1350 -660
rect 1150 -732 1350 -721
rect 1150 -766 1168 -732
rect 1202 -766 1236 -732
rect 1270 -766 1304 -732
rect 1338 -766 1350 -732
rect 1150 -777 1350 -766
rect 1150 -838 1350 -827
rect 1150 -872 1168 -838
rect 1202 -872 1236 -838
rect 1270 -872 1304 -838
rect 1338 -872 1350 -838
rect 1150 -880 1350 -872
<< mvndiff >>
rect 128 1867 181 1885
rect 128 1833 136 1867
rect 170 1833 181 1867
rect 128 1799 181 1833
rect 128 1765 136 1799
rect 170 1765 181 1799
rect 128 1731 181 1765
rect 128 1697 136 1731
rect 170 1697 181 1731
rect 128 1685 181 1697
rect 361 1867 417 1885
rect 361 1833 372 1867
rect 406 1833 417 1867
rect 361 1799 417 1833
rect 361 1765 372 1799
rect 406 1765 417 1799
rect 361 1731 417 1765
rect 361 1697 372 1731
rect 406 1697 417 1731
rect 361 1685 417 1697
rect 597 1867 650 1885
rect 597 1833 608 1867
rect 642 1833 650 1867
rect 597 1799 650 1833
rect 597 1765 608 1799
rect 642 1765 650 1799
rect 597 1731 650 1765
rect 597 1697 608 1731
rect 642 1697 650 1731
rect 597 1685 650 1697
rect 724 1877 777 1889
rect 724 1843 732 1877
rect 766 1843 777 1877
rect 724 1809 777 1843
rect 724 1775 732 1809
rect 766 1775 777 1809
rect 724 1741 777 1775
rect 724 1707 732 1741
rect 766 1707 777 1741
rect 724 1689 777 1707
rect 957 1877 1013 1889
rect 957 1843 968 1877
rect 1002 1843 1013 1877
rect 957 1809 1013 1843
rect 957 1775 968 1809
rect 1002 1775 1013 1809
rect 957 1741 1013 1775
rect 957 1707 968 1741
rect 1002 1707 1013 1741
rect 957 1689 1013 1707
rect 1193 1877 1246 1889
rect 1193 1843 1204 1877
rect 1238 1843 1246 1877
rect 1193 1809 1246 1843
rect 1193 1775 1204 1809
rect 1238 1775 1246 1809
rect 1193 1741 1246 1775
rect 1193 1707 1204 1741
rect 1238 1707 1246 1741
rect 1193 1689 1246 1707
rect 128 1573 181 1591
rect 128 1539 136 1573
rect 170 1539 181 1573
rect 128 1505 181 1539
rect 128 1471 136 1505
rect 170 1471 181 1505
rect 128 1437 181 1471
rect 128 1403 136 1437
rect 170 1403 181 1437
rect 128 1391 181 1403
rect 361 1573 417 1591
rect 361 1539 372 1573
rect 406 1539 417 1573
rect 361 1505 417 1539
rect 361 1471 372 1505
rect 406 1471 417 1505
rect 361 1437 417 1471
rect 361 1403 372 1437
rect 406 1403 417 1437
rect 361 1391 417 1403
rect 597 1573 650 1591
rect 597 1539 608 1573
rect 642 1539 650 1573
rect 597 1505 650 1539
rect 597 1471 608 1505
rect 642 1471 650 1505
rect 597 1437 650 1471
rect 597 1403 608 1437
rect 642 1403 650 1437
rect 597 1391 650 1403
rect 724 1573 777 1591
rect 724 1539 732 1573
rect 766 1539 777 1573
rect 724 1505 777 1539
rect 724 1471 732 1505
rect 766 1471 777 1505
rect 724 1437 777 1471
rect 724 1403 732 1437
rect 766 1403 777 1437
rect 724 1391 777 1403
rect 957 1573 1013 1591
rect 957 1539 968 1573
rect 1002 1539 1013 1573
rect 957 1505 1013 1539
rect 957 1471 968 1505
rect 1002 1471 1013 1505
rect 957 1437 1013 1471
rect 957 1403 968 1437
rect 1002 1403 1013 1437
rect 957 1391 1013 1403
rect 1193 1573 1246 1591
rect 1193 1539 1204 1573
rect 1238 1539 1246 1573
rect 1193 1505 1246 1539
rect 1193 1471 1204 1505
rect 1238 1471 1246 1505
rect 1193 1437 1246 1471
rect 1193 1403 1204 1437
rect 1238 1403 1246 1437
rect 1461 1811 1514 1889
rect 1461 1777 1469 1811
rect 1503 1777 1514 1811
rect 1461 1743 1514 1777
rect 1461 1709 1469 1743
rect 1503 1709 1514 1743
rect 1461 1675 1514 1709
rect 1461 1641 1469 1675
rect 1503 1641 1514 1675
rect 1461 1607 1514 1641
rect 1461 1573 1469 1607
rect 1503 1573 1514 1607
rect 1461 1539 1514 1573
rect 1461 1505 1469 1539
rect 1503 1505 1514 1539
rect 1461 1471 1514 1505
rect 1461 1437 1469 1471
rect 1503 1437 1514 1471
rect 1193 1391 1246 1403
rect 1461 1403 1514 1437
rect 1461 1369 1469 1403
rect 1503 1369 1514 1403
rect 1461 1335 1514 1369
rect 1461 1301 1469 1335
rect 1503 1301 1514 1335
rect 1461 1289 1514 1301
rect 1634 1811 1690 1889
rect 1634 1777 1645 1811
rect 1679 1777 1690 1811
rect 1634 1743 1690 1777
rect 1634 1709 1645 1743
rect 1679 1709 1690 1743
rect 1634 1675 1690 1709
rect 1634 1641 1645 1675
rect 1679 1641 1690 1675
rect 1634 1607 1690 1641
rect 1634 1573 1645 1607
rect 1679 1573 1690 1607
rect 1634 1539 1690 1573
rect 1634 1505 1645 1539
rect 1679 1505 1690 1539
rect 1634 1471 1690 1505
rect 1634 1437 1645 1471
rect 1679 1437 1690 1471
rect 1634 1403 1690 1437
rect 1634 1369 1645 1403
rect 1679 1369 1690 1403
rect 1634 1335 1690 1369
rect 1634 1301 1645 1335
rect 1679 1301 1690 1335
rect 1634 1289 1690 1301
rect 1810 1811 1866 1889
rect 1810 1777 1821 1811
rect 1855 1777 1866 1811
rect 1810 1743 1866 1777
rect 1810 1709 1821 1743
rect 1855 1709 1866 1743
rect 1810 1675 1866 1709
rect 1810 1641 1821 1675
rect 1855 1641 1866 1675
rect 1810 1607 1866 1641
rect 1810 1573 1821 1607
rect 1855 1573 1866 1607
rect 1810 1539 1866 1573
rect 1810 1505 1821 1539
rect 1855 1505 1866 1539
rect 1810 1471 1866 1505
rect 1810 1437 1821 1471
rect 1855 1437 1866 1471
rect 1810 1403 1866 1437
rect 1810 1369 1821 1403
rect 1855 1369 1866 1403
rect 1810 1335 1866 1369
rect 1810 1301 1821 1335
rect 1855 1301 1866 1335
rect 1810 1289 1866 1301
rect 1986 1811 2039 1889
rect 1986 1777 1997 1811
rect 2031 1777 2039 1811
rect 1986 1743 2039 1777
rect 1986 1709 1997 1743
rect 2031 1709 2039 1743
rect 1986 1675 2039 1709
rect 1986 1641 1997 1675
rect 2031 1641 2039 1675
rect 1986 1607 2039 1641
rect 1986 1573 1997 1607
rect 2031 1573 2039 1607
rect 1986 1539 2039 1573
rect 1986 1505 1997 1539
rect 2031 1505 2039 1539
rect 1986 1471 2039 1505
rect 1986 1437 1997 1471
rect 2031 1437 2039 1471
rect 1986 1403 2039 1437
rect 1986 1369 1997 1403
rect 2031 1369 2039 1403
rect 1986 1335 2039 1369
rect 1986 1301 1997 1335
rect 2031 1301 2039 1335
rect 1986 1289 2039 1301
rect 30 1178 86 1190
rect 30 1144 41 1178
rect 75 1144 86 1178
rect 30 1110 86 1144
rect 30 1076 41 1110
rect 75 1076 86 1110
rect 30 1042 86 1076
rect 30 1008 41 1042
rect 75 1008 86 1042
rect 30 990 86 1008
rect 206 1178 262 1190
rect 206 1144 217 1178
rect 251 1144 262 1178
rect 206 1110 262 1144
rect 206 1076 217 1110
rect 251 1076 262 1110
rect 206 1042 262 1076
rect 206 1008 217 1042
rect 251 1008 262 1042
rect 206 990 262 1008
rect 382 1178 438 1190
rect 382 1144 393 1178
rect 427 1144 438 1178
rect 382 1110 438 1144
rect 382 1076 393 1110
rect 427 1076 438 1110
rect 382 1042 438 1076
rect 382 1008 393 1042
rect 427 1008 438 1042
rect 1461 1083 1514 1095
rect 1461 1049 1469 1083
rect 1503 1049 1514 1083
rect 1461 1015 1514 1049
rect 382 990 438 1008
rect 1461 981 1469 1015
rect 1503 981 1514 1015
rect 1461 945 1514 981
rect 1714 1083 1770 1095
rect 1714 1049 1725 1083
rect 1759 1049 1770 1083
rect 1714 1015 1770 1049
rect 1714 981 1725 1015
rect 1759 981 1770 1015
rect 1714 945 1770 981
rect 1970 1083 2023 1095
rect 1970 1049 1981 1083
rect 2015 1049 2023 1083
rect 1970 1015 2023 1049
rect 1970 981 1981 1015
rect 2015 981 2023 1015
rect 1970 945 2023 981
rect 1115 669 1168 681
rect 1115 635 1123 669
rect 1157 635 1168 669
rect 1115 601 1168 635
rect 1115 567 1123 601
rect 1157 567 1168 601
rect 1115 533 1168 567
rect 1115 499 1123 533
rect 1157 499 1168 533
rect 1115 465 1168 499
rect 1115 431 1123 465
rect 1157 431 1168 465
rect 1115 397 1168 431
rect 1115 363 1123 397
rect 1157 363 1168 397
rect 1115 329 1168 363
rect 1115 295 1123 329
rect 1157 295 1168 329
rect 1115 261 1168 295
rect 1115 227 1123 261
rect 1157 227 1168 261
rect 1115 193 1168 227
rect 1115 159 1123 193
rect 1157 159 1168 193
rect 1115 81 1168 159
rect 1288 669 1341 681
rect 1288 635 1299 669
rect 1333 635 1341 669
rect 1288 601 1341 635
rect 1288 567 1299 601
rect 1333 567 1341 601
rect 1288 533 1341 567
rect 1288 499 1299 533
rect 1333 499 1341 533
rect 1288 465 1341 499
rect 1288 431 1299 465
rect 1333 431 1341 465
rect 1288 397 1341 431
rect 1288 363 1299 397
rect 1333 363 1341 397
rect 1288 329 1341 363
rect 1288 295 1299 329
rect 1333 295 1341 329
rect 1288 261 1341 295
rect 1288 227 1299 261
rect 1333 227 1341 261
rect 1288 193 1341 227
rect 1288 159 1299 193
rect 1333 159 1341 193
rect 1288 81 1341 159
<< mvpdiff >>
rect 77 664 130 676
rect 77 630 85 664
rect 119 630 130 664
rect 77 596 130 630
rect 77 562 85 596
rect 119 562 130 596
rect 77 526 130 562
rect 230 664 283 676
rect 230 630 241 664
rect 275 630 283 664
rect 230 596 283 630
rect 230 562 241 596
rect 275 562 283 596
rect 230 526 283 562
rect 343 664 396 676
rect 343 630 351 664
rect 385 630 396 664
rect 343 596 396 630
rect 343 562 351 596
rect 385 562 396 596
rect 343 528 396 562
rect 343 494 351 528
rect 385 494 396 528
rect 343 460 396 494
rect 343 426 351 460
rect 385 426 396 460
rect 343 392 396 426
rect 343 358 351 392
rect 385 358 396 392
rect 77 345 130 357
rect 77 311 85 345
rect 119 311 130 345
rect 77 277 130 311
rect 77 243 85 277
rect 119 243 130 277
rect 77 207 130 243
rect 230 345 283 357
rect 230 311 241 345
rect 275 311 283 345
rect 230 277 283 311
rect 230 243 241 277
rect 275 243 283 277
rect 230 207 283 243
rect 343 324 396 358
rect 343 290 351 324
rect 385 290 396 324
rect 343 256 396 290
rect 343 222 351 256
rect 385 222 396 256
rect 343 188 396 222
rect 343 154 351 188
rect 385 154 396 188
rect 343 76 396 154
rect 516 664 572 676
rect 516 630 527 664
rect 561 630 572 664
rect 516 596 572 630
rect 516 562 527 596
rect 561 562 572 596
rect 516 528 572 562
rect 516 494 527 528
rect 561 494 572 528
rect 516 460 572 494
rect 516 426 527 460
rect 561 426 572 460
rect 516 392 572 426
rect 516 358 527 392
rect 561 358 572 392
rect 516 324 572 358
rect 516 290 527 324
rect 561 290 572 324
rect 516 256 572 290
rect 516 222 527 256
rect 561 222 572 256
rect 516 188 572 222
rect 516 154 527 188
rect 561 154 572 188
rect 516 76 572 154
rect 692 664 745 676
rect 692 630 703 664
rect 737 630 745 664
rect 692 596 745 630
rect 692 562 703 596
rect 737 562 745 596
rect 692 528 745 562
rect 692 494 703 528
rect 737 494 745 528
rect 692 460 745 494
rect 692 426 703 460
rect 737 426 745 460
rect 692 392 745 426
rect 692 358 703 392
rect 737 358 745 392
rect 692 324 745 358
rect 692 290 703 324
rect 737 290 745 324
rect 692 256 745 290
rect 692 222 703 256
rect 737 222 745 256
rect 692 188 745 222
rect 692 154 703 188
rect 737 154 745 188
rect 692 76 745 154
<< ndiffc >>
rect 603 1191 637 1225
rect 603 1123 637 1157
rect 603 1055 637 1089
rect 689 1191 723 1225
rect 689 1123 723 1157
rect 689 1055 723 1089
rect 775 1191 809 1225
rect 775 1123 809 1157
rect 775 1055 809 1089
rect 861 1191 895 1225
rect 861 1123 895 1157
rect 861 1055 895 1089
rect 947 1191 981 1225
rect 947 1123 981 1157
rect 947 1055 981 1089
rect 1033 1191 1067 1225
rect 1033 1123 1067 1157
rect 1033 1055 1067 1089
rect 1119 1191 1153 1225
rect 1119 1123 1153 1157
rect 1119 1055 1153 1089
rect 1205 1191 1239 1225
rect 1205 1123 1239 1157
rect 1205 1055 1239 1089
rect 1291 1191 1325 1225
rect 1291 1123 1325 1157
rect 1291 1055 1325 1089
rect 1667 -1128 1701 -1094
rect 1667 -1196 1701 -1162
rect 1667 -1264 1701 -1230
rect 1773 -1128 1807 -1094
rect 1773 -1196 1807 -1162
rect 1773 -1264 1807 -1230
rect 1879 -1128 1913 -1094
rect 1879 -1196 1913 -1162
rect 1879 -1264 1913 -1230
<< pdiffc >>
rect 1168 -660 1202 -626
rect 1236 -660 1270 -626
rect 1304 -660 1338 -626
rect 1168 -766 1202 -732
rect 1236 -766 1270 -732
rect 1304 -766 1338 -732
rect 1168 -872 1202 -838
rect 1236 -872 1270 -838
rect 1304 -872 1338 -838
<< mvndiffc >>
rect 136 1833 170 1867
rect 136 1765 170 1799
rect 136 1697 170 1731
rect 372 1833 406 1867
rect 372 1765 406 1799
rect 372 1697 406 1731
rect 608 1833 642 1867
rect 608 1765 642 1799
rect 608 1697 642 1731
rect 732 1843 766 1877
rect 732 1775 766 1809
rect 732 1707 766 1741
rect 968 1843 1002 1877
rect 968 1775 1002 1809
rect 968 1707 1002 1741
rect 1204 1843 1238 1877
rect 1204 1775 1238 1809
rect 1204 1707 1238 1741
rect 136 1539 170 1573
rect 136 1471 170 1505
rect 136 1403 170 1437
rect 372 1539 406 1573
rect 372 1471 406 1505
rect 372 1403 406 1437
rect 608 1539 642 1573
rect 608 1471 642 1505
rect 608 1403 642 1437
rect 732 1539 766 1573
rect 732 1471 766 1505
rect 732 1403 766 1437
rect 968 1539 1002 1573
rect 968 1471 1002 1505
rect 968 1403 1002 1437
rect 1204 1539 1238 1573
rect 1204 1471 1238 1505
rect 1204 1403 1238 1437
rect 1469 1777 1503 1811
rect 1469 1709 1503 1743
rect 1469 1641 1503 1675
rect 1469 1573 1503 1607
rect 1469 1505 1503 1539
rect 1469 1437 1503 1471
rect 1469 1369 1503 1403
rect 1469 1301 1503 1335
rect 1645 1777 1679 1811
rect 1645 1709 1679 1743
rect 1645 1641 1679 1675
rect 1645 1573 1679 1607
rect 1645 1505 1679 1539
rect 1645 1437 1679 1471
rect 1645 1369 1679 1403
rect 1645 1301 1679 1335
rect 1821 1777 1855 1811
rect 1821 1709 1855 1743
rect 1821 1641 1855 1675
rect 1821 1573 1855 1607
rect 1821 1505 1855 1539
rect 1821 1437 1855 1471
rect 1821 1369 1855 1403
rect 1821 1301 1855 1335
rect 1997 1777 2031 1811
rect 1997 1709 2031 1743
rect 1997 1641 2031 1675
rect 1997 1573 2031 1607
rect 1997 1505 2031 1539
rect 1997 1437 2031 1471
rect 1997 1369 2031 1403
rect 1997 1301 2031 1335
rect 41 1144 75 1178
rect 41 1076 75 1110
rect 41 1008 75 1042
rect 217 1144 251 1178
rect 217 1076 251 1110
rect 217 1008 251 1042
rect 393 1144 427 1178
rect 393 1076 427 1110
rect 393 1008 427 1042
rect 1469 1049 1503 1083
rect 1469 981 1503 1015
rect 1725 1049 1759 1083
rect 1725 981 1759 1015
rect 1981 1049 2015 1083
rect 1981 981 2015 1015
rect 1123 635 1157 669
rect 1123 567 1157 601
rect 1123 499 1157 533
rect 1123 431 1157 465
rect 1123 363 1157 397
rect 1123 295 1157 329
rect 1123 227 1157 261
rect 1123 159 1157 193
rect 1299 635 1333 669
rect 1299 567 1333 601
rect 1299 499 1333 533
rect 1299 431 1333 465
rect 1299 363 1333 397
rect 1299 295 1333 329
rect 1299 227 1333 261
rect 1299 159 1333 193
<< mvpdiffc >>
rect 85 630 119 664
rect 85 562 119 596
rect 241 630 275 664
rect 241 562 275 596
rect 351 630 385 664
rect 351 562 385 596
rect 351 494 385 528
rect 351 426 385 460
rect 351 358 385 392
rect 85 311 119 345
rect 85 243 119 277
rect 241 311 275 345
rect 241 243 275 277
rect 351 290 385 324
rect 351 222 385 256
rect 351 154 385 188
rect 527 630 561 664
rect 527 562 561 596
rect 527 494 561 528
rect 527 426 561 460
rect 527 358 561 392
rect 527 290 561 324
rect 527 222 561 256
rect 527 154 561 188
rect 703 630 737 664
rect 703 562 737 596
rect 703 494 737 528
rect 703 426 737 460
rect 703 358 737 392
rect 703 290 737 324
rect 703 222 737 256
rect 703 154 737 188
<< nsubdiff >>
rect 1150 -562 1174 -528
rect 1208 -562 1292 -528
rect 1326 -562 1350 -528
<< mvpsubdiff >>
rect -17 1863 17 1887
rect -17 1792 17 1829
rect -17 1721 17 1758
rect -17 1650 17 1687
rect 1353 1886 1387 1910
rect 1353 1818 1387 1852
rect 1353 1750 1387 1784
rect -17 1579 17 1616
rect 1353 1682 1387 1716
rect 1353 1614 1387 1648
rect -17 1508 17 1545
rect -17 1437 17 1474
rect -17 1379 17 1403
rect 1353 1546 1387 1580
rect 1353 1429 1387 1512
rect 1006 657 1040 681
rect 1006 583 1040 623
rect 1006 509 1040 549
rect 1006 435 1040 475
rect 1006 361 1040 401
rect 1006 287 1040 327
rect 1006 213 1040 253
rect 1006 139 1040 179
rect 1006 81 1040 105
<< mvnsubdiff >>
rect 0 94 77 128
rect 111 94 145 128
rect 179 94 203 128
rect 819 638 853 662
rect 819 566 853 604
rect 819 494 853 532
rect 819 422 853 460
rect 819 350 853 388
rect 819 278 853 316
rect 819 206 853 244
rect 819 134 853 172
rect 819 76 853 100
<< nsubdiffcont >>
rect 1174 -562 1208 -528
rect 1292 -562 1326 -528
<< mvpsubdiffcont >>
rect -17 1829 17 1863
rect -17 1758 17 1792
rect -17 1687 17 1721
rect 1353 1852 1387 1886
rect 1353 1784 1387 1818
rect 1353 1716 1387 1750
rect -17 1616 17 1650
rect 1353 1648 1387 1682
rect -17 1545 17 1579
rect -17 1474 17 1508
rect -17 1403 17 1437
rect 1353 1580 1387 1614
rect 1353 1512 1387 1546
rect 1006 623 1040 657
rect 1006 549 1040 583
rect 1006 475 1040 509
rect 1006 401 1040 435
rect 1006 327 1040 361
rect 1006 253 1040 287
rect 1006 179 1040 213
rect 1006 105 1040 139
<< mvnsubdiffcont >>
rect 77 94 111 128
rect 145 94 179 128
rect 819 604 853 638
rect 819 532 853 566
rect 819 460 853 494
rect 819 388 853 422
rect 819 316 853 350
rect 819 244 853 278
rect 819 172 853 206
rect 819 100 853 134
<< poly >>
rect 181 1990 1200 2019
rect 181 1956 211 1990
rect 245 1956 279 1990
rect 313 1956 347 1990
rect 381 1956 415 1990
rect 449 1956 483 1990
rect 517 1956 551 1990
rect 585 1956 619 1990
rect 653 1956 687 1990
rect 721 1956 755 1990
rect 789 1956 823 1990
rect 857 1956 891 1990
rect 925 1956 959 1990
rect 993 1956 1027 1990
rect 1061 1956 1095 1990
rect 1129 1956 1200 1990
rect 181 1911 1200 1956
rect 1506 1971 1640 1987
rect 1506 1937 1522 1971
rect 1556 1937 1590 1971
rect 1624 1937 1640 1971
rect 1506 1921 1640 1937
rect 1683 1965 1817 1981
rect 1683 1931 1699 1965
rect 1733 1931 1767 1965
rect 1801 1931 1817 1965
rect 181 1885 361 1911
rect 417 1885 597 1911
rect 777 1889 957 1911
rect 1013 1889 1193 1911
rect 1514 1889 1634 1921
rect 1683 1915 1817 1931
rect 1866 1975 2005 1991
rect 1866 1941 1887 1975
rect 1921 1941 1955 1975
rect 1989 1941 2005 1975
rect 1866 1915 2005 1941
rect 1690 1889 1810 1915
rect 1866 1889 1986 1915
rect 181 1591 361 1685
rect 417 1591 597 1685
rect 777 1591 957 1689
rect 1013 1591 1193 1689
rect 181 1365 361 1391
rect 417 1365 597 1391
rect 777 1365 957 1391
rect 1013 1365 1193 1391
rect 181 1305 1200 1365
rect 1514 1263 1634 1289
rect 1690 1263 1810 1289
rect 1866 1263 1986 1289
rect 648 1237 678 1263
rect 734 1237 764 1263
rect 820 1237 850 1263
rect 906 1237 936 1263
rect 992 1237 1022 1263
rect 1078 1237 1108 1263
rect 1164 1237 1194 1263
rect 1250 1237 1280 1263
rect 86 1190 206 1216
rect 262 1190 382 1216
rect 1514 1179 1714 1201
rect 1514 1145 1569 1179
rect 1603 1145 1637 1179
rect 1671 1145 1714 1179
rect 1514 1095 1714 1145
rect 1770 1169 1970 1187
rect 1770 1135 1852 1169
rect 1886 1135 1920 1169
rect 1954 1135 1970 1169
rect 1770 1095 1970 1135
rect 648 1011 678 1037
rect 734 1011 764 1037
rect 820 1011 850 1037
rect 906 1011 936 1037
rect 992 1011 1022 1037
rect 1078 1011 1108 1037
rect 1164 1011 1194 1037
rect 1250 1011 1280 1037
rect 86 927 206 990
rect 65 911 206 927
rect 65 877 81 911
rect 115 877 149 911
rect 183 877 206 911
rect 65 861 206 877
rect 130 702 206 861
rect 262 897 382 990
rect 262 863 303 897
rect 337 863 382 897
rect 262 829 382 863
rect 634 907 949 1011
rect 992 988 1302 1011
rect 992 954 1039 988
rect 1073 954 1107 988
rect 1141 954 1175 988
rect 1209 954 1243 988
rect 1277 954 1302 988
rect 992 934 1302 954
rect 1514 919 1714 945
rect 1770 919 1970 945
rect 634 873 695 907
rect 729 873 763 907
rect 797 873 831 907
rect 865 873 899 907
rect 933 873 949 907
rect 634 829 949 873
rect 262 795 303 829
rect 337 828 382 829
rect 337 795 516 828
rect 262 762 516 795
rect 130 676 230 702
rect 396 676 516 762
rect 572 758 712 774
rect 572 724 588 758
rect 622 724 656 758
rect 690 724 712 758
rect 572 708 712 724
rect 1154 763 1336 779
rect 1154 729 1218 763
rect 1252 729 1286 763
rect 1320 729 1336 763
rect 572 676 692 708
rect 1154 707 1336 729
rect 1168 681 1288 707
rect 130 500 230 526
rect 130 439 297 455
rect 130 405 174 439
rect 208 405 242 439
rect 276 405 297 439
rect 130 389 297 405
rect 130 357 230 389
rect 130 181 230 207
rect 396 50 516 76
rect 572 24 692 76
rect 1168 55 1288 81
rect 1477 -671 1611 -655
rect 1124 -721 1150 -671
rect 1350 -705 1493 -671
rect 1527 -705 1561 -671
rect 1595 -705 1611 -671
rect 1350 -721 1611 -705
rect 1124 -827 1150 -777
rect 1350 -793 1611 -777
rect 1350 -827 1493 -793
rect 1527 -827 1561 -793
rect 1595 -827 1611 -793
rect 1477 -843 1611 -827
rect 1628 -1000 1762 -984
rect 1628 -1034 1644 -1000
rect 1678 -1034 1712 -1000
rect 1746 -1034 1762 -1000
rect 1628 -1050 1762 -1034
rect 1712 -1076 1762 -1050
rect 1818 -1000 1952 -984
rect 1818 -1034 1834 -1000
rect 1868 -1034 1902 -1000
rect 1936 -1034 1952 -1000
rect 1818 -1050 1952 -1034
rect 1818 -1076 1868 -1050
rect 1712 -1302 1762 -1276
rect 1818 -1302 1868 -1276
<< polycont >>
rect 211 1956 245 1990
rect 279 1956 313 1990
rect 347 1956 381 1990
rect 415 1956 449 1990
rect 483 1956 517 1990
rect 551 1956 585 1990
rect 619 1956 653 1990
rect 687 1956 721 1990
rect 755 1956 789 1990
rect 823 1956 857 1990
rect 891 1956 925 1990
rect 959 1956 993 1990
rect 1027 1956 1061 1990
rect 1095 1956 1129 1990
rect 1522 1937 1556 1971
rect 1590 1937 1624 1971
rect 1699 1931 1733 1965
rect 1767 1931 1801 1965
rect 1887 1941 1921 1975
rect 1955 1941 1989 1975
rect 1569 1145 1603 1179
rect 1637 1145 1671 1179
rect 1852 1135 1886 1169
rect 1920 1135 1954 1169
rect 81 877 115 911
rect 149 877 183 911
rect 303 863 337 897
rect 1039 954 1073 988
rect 1107 954 1141 988
rect 1175 954 1209 988
rect 1243 954 1277 988
rect 695 873 729 907
rect 763 873 797 907
rect 831 873 865 907
rect 899 873 933 907
rect 303 795 337 829
rect 588 724 622 758
rect 656 724 690 758
rect 1218 729 1252 763
rect 1286 729 1320 763
rect 174 405 208 439
rect 242 405 276 439
rect 1493 -705 1527 -671
rect 1561 -705 1595 -671
rect 1493 -827 1527 -793
rect 1561 -827 1595 -793
rect 1644 -1034 1678 -1000
rect 1712 -1034 1746 -1000
rect 1834 -1034 1868 -1000
rect 1902 -1034 1936 -1000
<< locali >>
rect 195 1956 211 1990
rect 245 1956 279 1990
rect 317 1956 347 1990
rect 389 1956 415 1990
rect 461 1956 483 1990
rect 533 1956 551 1990
rect 605 1956 619 1990
rect 677 1956 687 1990
rect 749 1956 755 1990
rect 821 1956 823 1990
rect 857 1956 859 1990
rect 925 1956 931 1990
rect 993 1956 1003 1990
rect 1061 1956 1075 1990
rect 1129 1956 1147 1990
rect 1506 1937 1522 1971
rect 1556 1937 1590 1971
rect 1624 1937 1640 1971
rect -17 1863 17 1887
rect -17 1792 17 1829
rect -17 1721 17 1758
rect -17 1650 17 1687
rect -17 1579 17 1584
rect -17 1508 17 1512
rect -17 1437 17 1440
rect -17 1402 17 1403
rect -17 1330 17 1368
rect 136 1867 170 1883
rect 136 1799 170 1833
rect 136 1731 170 1765
rect 136 1668 170 1697
rect 342 1867 448 1883
rect 342 1833 372 1867
rect 406 1833 448 1867
rect 342 1799 448 1833
rect 342 1765 372 1799
rect 406 1765 448 1799
rect 342 1731 448 1765
rect 342 1697 372 1731
rect 406 1697 448 1731
rect 342 1674 448 1697
rect 376 1640 414 1674
rect 608 1867 642 1883
rect 608 1799 642 1833
rect 608 1731 642 1765
rect 608 1691 642 1697
rect 136 1573 170 1634
rect 608 1610 642 1657
rect 136 1505 170 1528
rect 136 1456 170 1471
rect 136 1352 170 1403
rect 372 1582 406 1589
rect 372 1510 406 1539
rect 372 1438 406 1471
rect 372 1387 406 1403
rect 608 1573 642 1576
rect 608 1528 642 1539
rect 608 1437 642 1471
rect 608 1352 642 1403
rect 136 1275 642 1352
rect 732 1877 766 1893
rect 732 1841 766 1843
rect 931 1877 1037 1893
rect 931 1843 968 1877
rect 1002 1843 1037 1877
rect 732 1809 773 1841
rect 766 1775 773 1809
rect 732 1741 773 1775
rect 766 1707 773 1741
rect 732 1691 773 1707
rect 766 1657 773 1691
rect 931 1809 1037 1843
rect 931 1775 968 1809
rect 1002 1775 1037 1809
rect 931 1741 1037 1775
rect 931 1707 968 1741
rect 1002 1707 1037 1741
rect 931 1693 1037 1707
rect 965 1659 1003 1693
rect 1204 1877 1238 1893
rect 1204 1841 1238 1843
rect 1353 1886 1387 1910
rect 1517 1867 1639 1937
rect 1683 1931 1699 1965
rect 1733 1931 1767 1965
rect 1801 1931 1817 1965
rect 1871 1941 1887 1975
rect 1921 1941 1955 1975
rect 1989 1941 2005 1975
rect 1204 1809 1239 1841
rect 1238 1775 1239 1809
rect 1204 1741 1239 1775
rect 1238 1707 1239 1741
rect 732 1610 773 1657
rect 766 1576 773 1610
rect 732 1573 773 1576
rect 766 1539 773 1573
rect 732 1528 773 1539
rect 766 1471 773 1528
rect 732 1437 773 1471
rect 766 1403 773 1437
rect 732 1352 773 1403
rect 968 1532 1002 1539
rect 968 1437 1002 1471
rect 968 1387 1002 1403
rect 1204 1573 1239 1707
rect 1238 1539 1239 1573
rect 1204 1505 1239 1539
rect 1238 1471 1239 1505
rect 1204 1437 1239 1471
rect 1238 1403 1239 1437
rect 1353 1818 1387 1852
rect 1353 1750 1387 1784
rect 1353 1682 1387 1716
rect 1353 1614 1387 1648
rect 1353 1564 1387 1580
rect 1469 1811 1503 1827
rect 1469 1743 1503 1777
rect 1469 1691 1503 1709
rect 1469 1615 1503 1641
rect 1353 1546 1354 1564
rect 1387 1512 1388 1530
rect 1353 1483 1388 1512
rect 1353 1449 1354 1483
rect 1353 1429 1388 1449
rect 1204 1352 1239 1403
rect 732 1275 1239 1352
rect 1354 1402 1388 1429
rect 1354 1321 1388 1368
rect 1469 1539 1503 1573
rect 1469 1471 1503 1505
rect 1469 1403 1503 1437
rect 1469 1335 1503 1369
rect 1469 1285 1503 1301
rect 41 1178 75 1194
rect 41 1110 75 1144
rect 41 1042 75 1076
rect 41 999 75 1008
rect 217 1178 251 1200
rect 217 1110 251 1128
rect 217 1042 251 1076
rect 75 965 113 999
rect 217 992 251 1008
rect 388 1178 427 1194
rect 388 1144 393 1178
rect 388 1110 427 1144
rect 388 1076 393 1110
rect 485 1079 561 1275
rect 603 1234 637 1241
rect 603 1162 637 1191
rect 603 1089 637 1123
rect 388 1042 427 1076
rect 497 1045 535 1079
rect 388 1008 393 1042
rect 388 1006 427 1008
rect 65 877 81 911
rect 117 877 149 911
rect 189 877 206 911
rect 303 897 337 925
rect 303 829 337 863
rect 241 779 247 813
rect 281 795 303 813
rect 281 779 319 795
rect 85 664 119 680
rect 85 596 119 630
rect 85 345 119 562
rect 241 664 275 779
rect 388 680 447 1006
rect 485 999 561 1045
rect 603 1039 637 1055
rect 689 1225 723 1241
rect 689 1157 723 1191
rect 689 1089 723 1123
rect 689 999 723 1055
rect 775 1234 809 1241
rect 775 1162 809 1191
rect 775 1089 809 1123
rect 775 1039 809 1055
rect 861 1225 895 1241
rect 861 1157 895 1191
rect 861 1089 895 1123
rect 861 999 895 1055
rect 947 1234 981 1241
rect 947 1162 981 1191
rect 947 1089 981 1123
rect 947 1039 981 1055
rect 1033 1225 1067 1275
rect 1033 1157 1067 1191
rect 1033 1089 1067 1123
rect 1033 1039 1067 1055
rect 1119 1234 1153 1241
rect 1119 1162 1153 1191
rect 1119 1089 1153 1123
rect 1119 1039 1153 1055
rect 1205 1225 1239 1275
rect 1548 1251 1594 1867
rect 1205 1157 1239 1191
rect 1205 1089 1239 1123
rect 1205 1039 1239 1055
rect 1291 1234 1325 1241
rect 1291 1162 1325 1191
rect 1291 1089 1325 1123
rect 1291 1039 1325 1055
rect 1364 1217 1594 1251
rect 1645 1811 1679 1827
rect 1645 1743 1679 1777
rect 1645 1675 1679 1709
rect 1645 1607 1679 1641
rect 1645 1539 1679 1573
rect 1645 1493 1679 1505
rect 1645 1421 1679 1437
rect 1645 1335 1679 1369
rect 1713 1566 1787 1931
rect 1713 1532 1727 1566
rect 1761 1532 1787 1566
rect 1713 1490 1787 1532
rect 1713 1456 1727 1490
rect 1761 1456 1787 1490
rect 1713 1364 1787 1456
rect 1821 1811 1855 1827
rect 1821 1743 1855 1777
rect 1821 1675 1855 1709
rect 1821 1607 1855 1641
rect 1821 1539 1855 1573
rect 1821 1471 1855 1505
rect 1821 1403 1855 1437
rect 1889 1653 1963 1941
rect 1889 1619 1924 1653
rect 1958 1619 1963 1653
rect 1889 1577 1963 1619
rect 1889 1543 1924 1577
rect 1958 1543 1963 1577
rect 1889 1425 1963 1543
rect 1997 1811 2031 1857
rect 1997 1743 2031 1777
rect 1997 1675 2031 1709
rect 1997 1607 2031 1641
rect 1997 1539 2031 1573
rect 1997 1471 2031 1505
rect 1821 1335 1855 1369
rect 485 961 895 999
rect 1023 954 1033 988
rect 1073 954 1107 988
rect 1142 954 1175 988
rect 1217 954 1243 988
rect 1292 954 1293 988
rect 553 878 591 912
rect 572 758 625 878
rect 679 873 695 907
rect 729 873 763 907
rect 797 873 831 907
rect 865 873 899 907
rect 933 873 949 907
rect 572 724 588 758
rect 622 724 656 758
rect 690 724 712 758
rect 797 739 949 873
rect 1364 822 1415 1217
rect 1645 1179 1679 1301
rect 1725 1309 1821 1324
rect 1725 1203 1749 1309
rect 1997 1403 2031 1437
rect 1997 1335 2031 1369
rect 1553 1145 1569 1179
rect 1603 1145 1637 1179
rect 1671 1145 1687 1179
rect 1079 779 1117 813
rect 1151 779 1157 813
rect 241 596 275 630
rect 241 439 275 562
rect 351 664 363 680
rect 397 646 435 680
rect 527 664 561 680
rect 385 630 433 646
rect 351 596 433 630
rect 385 562 433 596
rect 351 528 433 562
rect 385 494 433 528
rect 351 460 433 494
rect 158 405 174 439
rect 208 405 242 439
rect 276 405 297 439
rect 385 426 433 460
rect 351 392 433 426
rect 85 277 119 280
rect 85 242 119 243
rect 85 170 119 208
rect 85 128 119 136
rect 241 345 314 361
rect 275 311 314 345
rect 241 277 314 311
rect 275 243 314 277
rect 0 94 77 128
rect 111 94 145 128
rect 179 94 203 128
rect 241 102 314 243
rect 385 358 433 392
rect 351 324 433 358
rect 385 290 433 324
rect 351 256 433 290
rect 385 222 433 256
rect 351 188 433 222
rect 385 154 433 188
rect 351 138 433 154
rect 527 596 561 630
rect 527 528 561 562
rect 527 460 561 494
rect 527 392 561 426
rect 527 324 561 358
rect 527 256 561 280
rect 527 188 561 208
rect 598 102 669 724
rect 797 705 817 739
rect 851 705 889 739
rect 923 705 949 739
rect 1109 681 1157 779
rect 1200 763 1415 822
rect 1456 1083 1505 1111
rect 1456 1049 1469 1083
rect 1503 1049 1505 1083
rect 1574 1065 1680 1145
rect 1725 1083 1796 1203
rect 1997 1169 2031 1301
rect 1836 1135 1852 1169
rect 1886 1135 1920 1169
rect 1954 1135 2031 1169
rect 1456 1015 1505 1049
rect 1456 981 1469 1015
rect 1503 981 1505 1015
rect 1759 1049 1796 1083
rect 1725 1015 1796 1049
rect 1456 819 1505 981
rect 1582 957 1620 991
rect 1759 981 1796 1015
rect 1725 965 1796 981
rect 1830 999 1864 1037
rect 1548 929 1654 957
rect 1548 858 1796 929
rect 1490 785 1528 819
rect 1658 769 1796 858
rect 1898 817 1947 1135
rect 1981 1083 2015 1099
rect 1981 1015 2015 1048
rect 1981 965 2015 976
rect 1932 783 1970 817
rect 1200 729 1218 763
rect 1252 729 1286 763
rect 1320 751 1415 763
rect 1320 732 1465 751
rect 1320 729 1381 732
rect 1367 698 1381 729
rect 1415 698 1465 732
rect 703 666 737 680
rect 703 596 737 630
rect 703 528 737 560
rect 703 460 737 494
rect 703 392 737 426
rect 703 324 737 358
rect 703 256 737 290
rect 703 188 737 222
rect 703 138 737 154
rect 819 638 853 662
rect 819 566 853 604
rect 819 494 853 532
rect 819 422 853 460
rect 819 350 853 388
rect 819 314 853 316
rect 819 278 853 280
rect 819 242 853 244
rect 819 206 853 208
rect 819 170 853 172
rect 241 49 669 102
rect 819 134 853 136
rect 819 76 853 100
rect 1006 657 1040 681
rect 1006 583 1040 610
rect 1006 509 1040 538
rect 1006 435 1040 475
rect 1006 361 1040 401
rect 1006 287 1040 327
rect 1006 213 1040 253
rect 1006 139 1040 179
rect 1109 647 1117 681
rect 1151 669 1157 681
rect 1109 635 1123 647
rect 1109 609 1157 635
rect 1109 575 1117 609
rect 1151 601 1157 609
rect 1109 567 1123 575
rect 1109 533 1157 567
rect 1109 499 1123 533
rect 1109 465 1157 499
rect 1109 431 1123 465
rect 1109 397 1157 431
rect 1109 363 1123 397
rect 1109 329 1157 363
rect 1109 295 1123 329
rect 1109 261 1157 295
rect 1109 227 1123 261
rect 1109 193 1157 227
rect 1109 159 1123 193
rect 1109 113 1157 159
rect 1299 620 1333 635
rect 1367 656 1465 698
rect 1367 622 1381 656
rect 1415 622 1465 656
rect 1299 533 1333 567
rect 1299 465 1333 499
rect 1299 397 1333 431
rect 1299 329 1333 363
rect 1299 261 1333 295
rect 1299 193 1333 227
rect 1299 143 1333 159
rect 1006 81 1040 105
rect 1090 -562 1147 -528
rect 1208 -562 1238 -528
rect 1272 -562 1292 -528
rect 1326 -562 1350 -528
rect 1153 -626 1317 -603
rect 1152 -660 1168 -626
rect 1202 -660 1236 -626
rect 1270 -660 1304 -626
rect 1351 -637 1389 -603
rect 1338 -660 1354 -637
rect 1404 -705 1493 -671
rect 1533 -705 1561 -671
rect 1605 -705 1611 -671
rect 1090 -766 1147 -732
rect 1202 -766 1236 -732
rect 1272 -766 1304 -732
rect 1338 -766 1354 -732
rect 1404 -838 1439 -705
rect 1477 -827 1493 -793
rect 1533 -827 1561 -793
rect 1605 -827 1611 -793
rect 1152 -872 1168 -838
rect 1202 -872 1236 -838
rect 1270 -872 1304 -838
rect 1338 -856 1439 -838
rect 1152 -890 1333 -872
rect 1367 -890 1405 -856
rect 1439 -890 1487 -864
rect 1152 -898 1487 -890
rect 1618 -1034 1644 -1000
rect 1690 -1034 1712 -1000
rect 1746 -1034 1762 -1000
rect 1818 -1034 1821 -1000
rect 1868 -1034 1893 -1000
rect 1936 -1034 1952 -1000
rect 1618 -1110 1656 -1076
rect 1690 -1094 1701 -1078
rect 1667 -1162 1701 -1128
rect 1667 -1230 1701 -1196
rect 1667 -1280 1701 -1264
rect 1773 -1094 1807 -1078
rect 1773 -1156 1807 -1128
rect 1773 -1228 1807 -1196
rect 1773 -1280 1807 -1264
rect 1879 -1082 1913 -1078
rect 1913 -1116 1951 -1082
rect 1879 -1162 1913 -1128
rect 1879 -1230 1913 -1196
rect 1879 -1280 1913 -1264
<< viali >>
rect 211 1956 245 1990
rect 283 1956 313 1990
rect 313 1956 317 1990
rect 355 1956 381 1990
rect 381 1956 389 1990
rect 427 1956 449 1990
rect 449 1956 461 1990
rect 499 1956 517 1990
rect 517 1956 533 1990
rect 571 1956 585 1990
rect 585 1956 605 1990
rect 643 1956 653 1990
rect 653 1956 677 1990
rect 715 1956 721 1990
rect 721 1956 749 1990
rect 787 1956 789 1990
rect 789 1956 821 1990
rect 859 1956 891 1990
rect 891 1956 893 1990
rect 931 1956 959 1990
rect 959 1956 965 1990
rect 1003 1956 1027 1990
rect 1027 1956 1037 1990
rect 1075 1956 1095 1990
rect 1095 1956 1109 1990
rect 1147 1956 1181 1990
rect -17 1616 17 1618
rect -17 1584 17 1616
rect -17 1545 17 1546
rect -17 1512 17 1545
rect -17 1440 17 1474
rect -17 1368 17 1402
rect -17 1296 17 1330
rect 136 1634 170 1668
rect 342 1640 376 1674
rect 414 1640 448 1674
rect 608 1657 642 1691
rect 136 1539 170 1562
rect 136 1528 170 1539
rect 136 1437 170 1456
rect 136 1422 170 1437
rect 372 1573 406 1582
rect 372 1548 406 1573
rect 372 1505 406 1510
rect 372 1476 406 1505
rect 372 1437 406 1438
rect 372 1404 406 1437
rect 608 1576 642 1610
rect 608 1505 642 1528
rect 608 1494 642 1505
rect 732 1657 766 1691
rect 931 1659 965 1693
rect 1003 1659 1037 1693
rect 732 1576 766 1610
rect 732 1505 766 1528
rect 732 1494 766 1505
rect 968 1573 1002 1604
rect 968 1570 1002 1573
rect 968 1505 1002 1532
rect 968 1498 1002 1505
rect 1469 1675 1503 1691
rect 1469 1657 1503 1675
rect 1469 1607 1503 1615
rect 1469 1581 1503 1607
rect 1354 1546 1388 1564
rect 1354 1530 1387 1546
rect 1387 1530 1388 1546
rect 1354 1449 1388 1483
rect 1354 1368 1388 1402
rect 1354 1287 1388 1321
rect 217 1200 251 1234
rect 217 1144 251 1162
rect 217 1128 251 1144
rect 41 965 75 999
rect 113 965 147 999
rect 603 1225 637 1234
rect 603 1200 637 1225
rect 603 1157 637 1162
rect 603 1128 637 1157
rect 463 1045 497 1079
rect 535 1045 569 1079
rect 83 877 115 911
rect 115 877 117 911
rect 155 877 183 911
rect 183 877 189 911
rect 247 779 281 813
rect 319 795 337 813
rect 337 795 353 813
rect 319 779 353 795
rect 775 1225 809 1234
rect 775 1200 809 1225
rect 775 1157 809 1162
rect 775 1128 809 1157
rect 947 1225 981 1234
rect 947 1200 981 1225
rect 947 1157 981 1162
rect 947 1128 981 1157
rect 1119 1225 1153 1234
rect 1119 1200 1153 1225
rect 1119 1157 1153 1162
rect 1119 1128 1153 1157
rect 1291 1225 1325 1234
rect 1291 1200 1325 1225
rect 1291 1157 1325 1162
rect 1291 1128 1325 1157
rect 1645 1471 1679 1493
rect 1645 1459 1679 1471
rect 1645 1403 1679 1421
rect 1645 1387 1679 1403
rect 1727 1532 1761 1566
rect 1727 1456 1761 1490
rect 1924 1619 1958 1653
rect 1924 1543 1958 1577
rect 1033 954 1039 988
rect 1039 954 1067 988
rect 1108 954 1141 988
rect 1141 954 1142 988
rect 1183 954 1209 988
rect 1209 954 1217 988
rect 1258 954 1277 988
rect 1277 954 1292 988
rect 519 878 553 912
rect 591 878 625 912
rect 1749 1301 1821 1309
rect 1821 1301 1855 1309
rect 1749 1203 1855 1301
rect 1045 779 1079 813
rect 1117 779 1151 813
rect 363 664 397 680
rect 363 646 385 664
rect 385 646 397 664
rect 435 646 469 680
rect 85 311 119 314
rect 85 280 119 311
rect 85 208 119 242
rect 85 136 119 170
rect 527 290 561 314
rect 527 280 561 290
rect 527 222 561 242
rect 527 208 561 222
rect 527 154 561 170
rect 527 136 561 154
rect 817 705 851 739
rect 889 705 923 739
rect 1548 957 1582 991
rect 1620 957 1654 991
rect 1830 1037 1864 1071
rect 1830 965 1864 999
rect 1456 785 1490 819
rect 1528 785 1562 819
rect 1981 1049 2015 1082
rect 1981 1048 2015 1049
rect 1981 981 2015 1010
rect 1981 976 2015 981
rect 1898 783 1932 817
rect 1970 783 2004 817
rect 1381 698 1415 732
rect 703 664 737 666
rect 703 632 737 664
rect 703 562 737 594
rect 703 560 737 562
rect 819 280 853 314
rect 819 208 853 242
rect 819 136 853 170
rect 1006 623 1040 644
rect 1006 610 1040 623
rect 1006 549 1040 572
rect 1006 538 1040 549
rect 1117 669 1151 681
rect 1117 647 1123 669
rect 1123 647 1151 669
rect 1117 601 1151 609
rect 1117 575 1123 601
rect 1123 575 1151 601
rect 1299 669 1333 692
rect 1299 658 1333 669
rect 1381 622 1415 656
rect 1299 601 1333 620
rect 1299 586 1333 601
rect 1056 -562 1090 -528
rect 1147 -562 1174 -528
rect 1174 -562 1181 -528
rect 1238 -562 1272 -528
rect 1317 -626 1351 -603
rect 1317 -637 1338 -626
rect 1338 -637 1351 -626
rect 1389 -637 1423 -603
rect 1499 -705 1527 -671
rect 1527 -705 1533 -671
rect 1571 -705 1595 -671
rect 1595 -705 1605 -671
rect 1056 -766 1090 -732
rect 1147 -766 1168 -732
rect 1168 -766 1181 -732
rect 1238 -766 1270 -732
rect 1270 -766 1272 -732
rect 1499 -827 1527 -793
rect 1527 -827 1533 -793
rect 1571 -827 1595 -793
rect 1595 -827 1605 -793
rect 1333 -872 1338 -856
rect 1338 -872 1367 -856
rect 1333 -890 1367 -872
rect 1405 -890 1439 -856
rect 1584 -1034 1618 -1000
rect 1656 -1034 1678 -1000
rect 1678 -1034 1690 -1000
rect 1821 -1034 1834 -1000
rect 1834 -1034 1855 -1000
rect 1893 -1034 1902 -1000
rect 1902 -1034 1927 -1000
rect 1584 -1110 1618 -1076
rect 1656 -1094 1690 -1076
rect 1656 -1110 1667 -1094
rect 1667 -1110 1690 -1094
rect 1773 -1162 1807 -1156
rect 1773 -1190 1807 -1162
rect 1773 -1230 1807 -1228
rect 1773 -1262 1807 -1230
rect 1879 -1094 1913 -1082
rect 1879 -1116 1913 -1094
rect 1951 -1116 1985 -1082
<< metal1 >>
rect -7 1990 2077 2019
rect -7 1956 211 1990
rect 245 1956 283 1990
rect 317 1956 355 1990
rect 389 1956 427 1990
rect 461 1956 499 1990
rect 533 1956 571 1990
rect 605 1956 643 1990
rect 677 1956 715 1990
rect 749 1956 787 1990
rect 821 1956 859 1990
rect 893 1956 931 1990
rect 965 1956 1003 1990
rect 1037 1956 1075 1990
rect 1109 1956 1147 1990
rect 1181 1956 2077 1990
rect -7 1818 2077 1956
rect 602 1691 648 1703
rect 127 1674 179 1680
rect -23 1618 23 1630
rect -23 1584 -17 1618
rect 17 1584 23 1618
rect -23 1546 23 1584
rect -23 1512 -17 1546
rect 17 1512 23 1546
rect -23 1474 23 1512
rect -23 1440 -17 1474
rect 17 1456 23 1474
rect 127 1606 179 1622
rect 330 1674 460 1680
rect 330 1640 342 1674
rect 376 1640 414 1674
rect 448 1640 460 1674
rect 330 1634 460 1640
rect 602 1657 608 1691
rect 642 1657 648 1691
tri 330 1619 345 1634 ne
rect 345 1619 433 1634
tri 433 1619 448 1634 nw
tri 345 1615 349 1619 ne
rect 349 1615 429 1619
tri 429 1615 433 1619 nw
tri 349 1610 354 1615 ne
rect 354 1610 424 1615
tri 424 1610 429 1615 nw
rect 602 1610 648 1657
tri 354 1598 366 1610 ne
rect 127 1537 136 1554
rect 170 1537 179 1554
tri 23 1456 39 1472 sw
rect 127 1468 179 1485
rect 17 1440 39 1456
rect -23 1422 39 1440
tri 39 1422 73 1456 sw
rect -23 1410 73 1422
tri 73 1410 85 1422 sw
rect 127 1410 179 1416
rect 366 1582 412 1610
tri 412 1598 424 1610 nw
rect 366 1548 372 1582
rect 406 1548 412 1582
rect 366 1510 412 1548
rect 366 1476 372 1510
rect 406 1476 412 1510
rect 602 1576 608 1610
rect 642 1576 648 1610
rect 602 1528 648 1576
rect 602 1494 608 1528
rect 642 1494 648 1528
rect 602 1482 648 1494
rect 726 1691 772 1703
rect 726 1657 732 1691
rect 766 1657 772 1691
rect 726 1610 772 1657
rect 919 1693 1509 1703
rect 919 1659 931 1693
rect 965 1659 1003 1693
rect 1037 1691 1509 1693
rect 1037 1659 1469 1691
rect 919 1657 1469 1659
rect 1503 1657 1509 1691
rect 919 1653 1509 1657
tri 919 1651 921 1653 ne
rect 921 1651 1509 1653
tri 921 1634 938 1651 ne
rect 938 1634 1025 1651
tri 1025 1634 1042 1651 nw
tri 1438 1634 1455 1651 ne
rect 1455 1634 1509 1651
tri 938 1626 946 1634 ne
rect 946 1626 1017 1634
tri 1017 1626 1025 1634 nw
tri 1455 1626 1463 1634 ne
tri 946 1619 953 1626 ne
rect 953 1619 1010 1626
tri 1010 1619 1017 1626 nw
tri 953 1615 957 1619 ne
rect 957 1615 1008 1619
tri 1008 1617 1010 1619 nw
tri 957 1610 962 1615 ne
rect 726 1576 732 1610
rect 766 1576 772 1610
rect 726 1528 772 1576
rect 726 1494 732 1528
rect 766 1494 772 1528
rect 726 1482 772 1494
rect 962 1604 1008 1615
rect 962 1570 968 1604
rect 1002 1570 1008 1604
rect 1463 1615 1509 1634
rect 1463 1581 1469 1615
rect 1503 1581 1509 1615
rect 962 1532 1008 1570
rect 962 1498 968 1532
rect 1002 1498 1008 1532
rect 1348 1564 1394 1576
rect 1463 1569 1509 1581
rect 1915 1653 1967 1665
rect 1915 1619 1924 1653
rect 1958 1619 1967 1653
rect 1348 1530 1354 1564
rect 1388 1530 1394 1564
rect 962 1486 1008 1498
rect 1265 1511 1317 1517
rect 366 1449 412 1476
tri 412 1449 438 1475 sw
tri 1239 1449 1265 1475 se
rect 1265 1449 1317 1459
rect 366 1441 438 1449
tri 438 1441 446 1449 sw
tri 1231 1441 1239 1449 se
rect 1239 1447 1317 1449
rect 1239 1441 1265 1447
rect 366 1438 1265 1441
rect -23 1404 85 1410
tri 85 1404 91 1410 sw
rect 366 1404 372 1438
rect 406 1404 1265 1438
rect -23 1402 91 1404
tri 91 1402 93 1404 sw
rect -23 1368 -17 1402
rect 17 1389 93 1402
tri 93 1389 106 1402 sw
rect 366 1395 1265 1404
rect 366 1389 1317 1395
rect 1348 1483 1394 1530
rect 1721 1566 1767 1578
rect 1721 1532 1727 1566
rect 1761 1532 1767 1566
rect 1348 1449 1354 1483
rect 1388 1449 1394 1483
rect 1348 1402 1394 1449
rect 17 1368 106 1389
tri 106 1368 127 1389 sw
rect 1348 1368 1354 1402
rect 1388 1368 1394 1402
rect 1634 1499 1686 1505
rect 1634 1433 1686 1447
rect 1721 1490 1767 1532
rect 1915 1577 1967 1619
rect 1915 1543 1924 1577
rect 1958 1543 1967 1577
rect 1915 1531 1967 1543
rect 1721 1456 1727 1490
rect 1761 1456 1767 1490
rect 1721 1444 1767 1456
rect 1634 1375 1686 1381
rect -23 1355 127 1368
tri 127 1355 140 1368 sw
tri -43 1330 -23 1350 se
rect -23 1330 140 1355
tri -49 1324 -43 1330 se
rect -43 1324 -17 1330
rect -49 1296 -17 1324
rect 17 1321 140 1330
tri 140 1321 174 1355 sw
tri 1314 1321 1348 1355 se
rect 1348 1321 1394 1368
tri 1394 1321 1428 1355 sw
rect 17 1315 1354 1321
rect 17 1296 997 1315
rect -49 1263 997 1296
rect 1049 1287 1354 1315
rect 1388 1309 2077 1321
rect 1388 1287 1749 1309
rect 1049 1263 1749 1287
rect -49 1251 1749 1263
rect -49 1234 997 1251
rect -49 1200 217 1234
rect 251 1200 603 1234
rect 637 1200 775 1234
rect 809 1200 947 1234
rect 981 1200 997 1234
rect -49 1199 997 1200
rect 1049 1234 1749 1251
rect 1049 1200 1119 1234
rect 1153 1200 1291 1234
rect 1325 1203 1749 1234
rect 1855 1203 2077 1309
rect 1325 1200 2077 1203
rect 1049 1199 2077 1200
rect -49 1187 2077 1199
rect -49 1162 997 1187
rect -49 1128 217 1162
rect 251 1128 603 1162
rect 637 1128 775 1162
rect 809 1128 947 1162
rect 981 1135 997 1162
rect 1049 1162 2077 1187
rect 1049 1135 1119 1162
rect 981 1128 1119 1135
rect 1153 1128 1291 1162
rect 1325 1128 2077 1162
rect -49 1122 2077 1128
rect 71 1039 77 1091
rect 129 1039 141 1091
rect 193 1085 199 1091
tri 199 1085 205 1091 sw
rect 193 1079 581 1085
rect 193 1045 463 1079
rect 497 1045 535 1079
rect 569 1045 581 1079
rect 193 1039 581 1045
rect 725 1079 777 1085
tri 721 1039 725 1043 se
tri 719 1037 721 1039 se
rect 721 1037 725 1039
tri 692 1010 719 1037 se
rect 719 1027 725 1037
rect 719 1015 777 1027
rect 719 1010 725 1015
tri 691 1009 692 1010 se
rect 692 1009 725 1010
rect 29 999 725 1009
rect 29 965 41 999
rect 75 965 113 999
rect 147 965 725 999
rect 29 963 725 965
rect 29 957 777 963
rect 805 1077 1870 1083
rect 857 1031 1818 1077
rect 857 1025 869 1031
rect 805 1013 869 1025
rect 857 1010 869 1013
tri 869 1010 890 1031 nw
tri 1790 1010 1811 1031 ne
rect 1811 1025 1818 1031
rect 1811 1011 1870 1025
rect 1811 1010 1818 1011
rect 857 1009 868 1010
tri 868 1009 869 1010 nw
tri 1811 1009 1812 1010 ne
rect 1812 1009 1818 1010
rect 857 999 858 1009
tri 858 999 868 1009 nw
tri 1812 1003 1818 1009 ne
tri 857 998 858 999 nw
rect 805 955 857 961
rect 1021 988 1459 1000
rect 1021 954 1033 988
rect 1067 954 1108 988
rect 1142 954 1183 988
rect 1217 954 1258 988
rect 1292 954 1459 988
rect 1021 948 1459 954
rect 1511 948 1523 1000
rect 1575 991 1666 1000
rect 1582 957 1620 991
rect 1654 957 1666 991
rect 1575 948 1666 957
rect 1818 953 1870 959
rect 1975 1082 2021 1094
rect 1975 1048 1981 1082
rect 2015 1048 2021 1082
rect 1975 1010 2021 1048
rect 1975 976 1981 1010
rect 2015 976 2021 1010
tri 1973 953 1975 955 se
rect 1975 953 2021 976
tri 1968 948 1973 953 se
rect 1973 948 2021 953
tri 1940 920 1968 948 se
rect 1968 920 2021 948
rect 67 919 2021 920
rect 67 912 1598 919
rect 67 911 519 912
rect 67 877 83 911
rect 117 877 155 911
rect 189 878 519 911
rect 553 878 591 912
rect 625 878 1598 912
rect 189 877 1598 878
rect 67 867 1598 877
rect 1650 867 1662 919
rect 1714 867 2021 919
rect 171 819 2016 825
rect 171 813 1456 819
rect 171 779 247 813
rect 281 779 319 813
rect 353 779 1045 813
rect 1079 779 1117 813
rect 1151 785 1456 813
rect 1490 785 1528 819
rect 1562 817 2016 819
rect 1562 785 1898 817
rect 1151 783 1898 785
rect 1932 783 1970 817
rect 2004 783 2016 817
rect 1151 779 2016 783
rect 171 773 2016 779
tri 1077 745 1105 773 ne
rect 1105 745 1157 773
rect 805 739 935 745
tri 1105 739 1111 745 ne
rect 857 705 889 739
rect 923 705 935 739
rect 857 693 935 705
rect 857 692 890 693
tri 890 692 891 693 nw
rect 857 687 884 692
rect 805 686 884 687
tri 884 686 890 692 nw
rect 34 680 481 686
rect 34 646 363 680
rect 397 646 435 680
rect 469 646 481 680
rect 34 640 481 646
rect 609 679 777 685
rect 609 666 725 679
rect 609 632 703 666
rect 609 627 725 632
rect 609 615 777 627
rect 805 681 879 686
tri 879 681 884 686 nw
rect 1111 681 1157 745
tri 1157 739 1191 773 nw
rect 1375 732 1421 744
rect 805 675 857 681
tri 857 659 879 681 nw
rect 805 617 857 623
rect 997 648 1049 656
rect 609 594 725 615
rect 609 560 703 594
rect 737 560 777 563
rect 609 554 777 560
rect 997 584 1049 596
rect 1111 647 1117 681
rect 1151 647 1157 681
rect 1111 609 1157 647
rect 1111 575 1117 609
rect 1151 575 1157 609
rect 1111 563 1157 575
rect 1265 698 1339 704
rect 1317 692 1339 698
rect 1333 658 1339 692
rect 1317 646 1339 658
rect 1265 634 1339 646
rect 1317 620 1339 634
rect 1333 586 1339 620
rect 1375 698 1381 732
rect 1415 698 1421 732
rect 1375 656 1421 698
rect 1375 622 1381 656
rect 1415 622 1421 656
rect 1375 610 1421 622
rect 1508 637 1560 643
rect 1317 582 1339 586
rect 1265 574 1339 582
rect 1508 570 1560 585
rect 997 526 1049 532
rect 1508 512 1560 518
rect 0 354 1594 484
rect 0 314 1594 326
rect 0 280 85 314
rect 119 280 527 314
rect 561 280 819 314
rect 853 280 1594 314
rect 0 242 1594 280
rect 0 208 85 242
rect 119 208 527 242
rect 561 208 819 242
rect 853 208 1594 242
rect 0 170 1594 208
rect 0 136 85 170
rect 119 136 527 170
rect 561 136 819 170
rect 853 136 1594 170
rect 0 124 1594 136
rect 823 43 829 95
rect 881 43 893 95
rect 945 43 1509 95
rect 1044 -571 1050 -519
rect 1102 -571 1114 -519
rect 1166 -528 1284 -519
rect 1181 -562 1238 -528
rect 1272 -562 1284 -528
rect 1166 -571 1284 -562
tri 1773 -597 1785 -585 se
rect 1785 -597 1791 -585
rect 1305 -603 1435 -597
rect 1305 -637 1317 -603
rect 1351 -637 1389 -603
rect 1423 -609 1435 -603
tri 1435 -609 1447 -597 sw
tri 1761 -609 1773 -597 se
rect 1773 -609 1791 -597
rect 1423 -637 1791 -609
rect 1843 -637 1855 -585
rect 1907 -637 1913 -585
rect 1305 -643 1435 -637
tri 1435 -643 1441 -637 nw
tri 1803 -643 1809 -637 ne
rect 1809 -643 1863 -637
tri 1809 -665 1831 -643 ne
rect 1831 -665 1863 -643
rect 1467 -717 1473 -665
rect 1525 -671 1537 -665
rect 1589 -669 1617 -665
tri 1617 -669 1621 -665 sw
tri 1831 -669 1835 -665 ne
rect 1589 -671 1621 -669
rect 1533 -705 1537 -671
rect 1605 -683 1621 -671
tri 1621 -683 1635 -669 sw
rect 1605 -705 1807 -683
rect 1525 -717 1537 -705
rect 1589 -711 1807 -705
rect 1589 -717 1595 -711
tri 1595 -717 1601 -711 nw
tri 1742 -717 1748 -711 ne
rect 1748 -717 1807 -711
tri 1748 -726 1757 -717 ne
rect 1757 -726 1807 -717
rect 1044 -732 1284 -726
rect 1044 -766 1056 -732
rect 1090 -766 1147 -732
rect 1181 -766 1238 -732
rect 1272 -766 1284 -732
tri 1757 -748 1779 -726 ne
rect 1044 -772 1284 -766
rect 1487 -793 1605 -787
rect 1487 -827 1499 -793
rect 1533 -827 1571 -793
rect 1487 -839 1605 -827
rect 1657 -839 1669 -787
rect 1721 -839 1727 -787
tri 1635 -849 1645 -839 ne
rect 1645 -849 1727 -839
tri 1645 -850 1646 -849 ne
rect 1646 -850 1727 -849
rect 1321 -856 1451 -850
rect 1321 -890 1333 -856
rect 1367 -890 1405 -856
rect 1439 -890 1451 -856
tri 1646 -874 1670 -850 ne
rect 1670 -874 1727 -850
tri 1670 -878 1674 -874 ne
rect 1321 -893 1451 -890
tri 1451 -893 1463 -881 sw
rect 1321 -896 1463 -893
tri 1391 -940 1435 -896 ne
rect 1435 -1076 1463 -896
tri 1631 -978 1674 -935 se
rect 1674 -978 1727 -874
tri 1616 -993 1631 -978 se
rect 1631 -993 1727 -978
tri 1615 -994 1616 -993 se
rect 1616 -994 1727 -993
rect 1572 -1000 1727 -994
rect 1572 -1034 1584 -1000
rect 1618 -1034 1656 -1000
rect 1690 -1034 1727 -1000
rect 1572 -1040 1727 -1034
rect 1779 -978 1807 -726
rect 1835 -839 1863 -665
tri 1863 -671 1897 -637 nw
tri 1863 -839 1871 -831 sw
rect 1835 -846 1871 -839
tri 1835 -849 1838 -846 ne
rect 1838 -849 1871 -846
tri 1871 -849 1881 -839 sw
tri 1838 -874 1863 -849 ne
rect 1863 -874 1881 -849
tri 1863 -881 1870 -874 ne
rect 1870 -881 1881 -874
tri 1881 -881 1913 -849 sw
tri 1870 -892 1881 -881 ne
rect 1881 -892 1913 -881
tri 1913 -892 1924 -881 sw
tri 1881 -935 1924 -892 ne
tri 1924 -935 1967 -892 sw
tri 1924 -962 1951 -935 ne
rect 1951 -962 1967 -935
tri 1807 -978 1823 -962 sw
tri 1951 -978 1967 -962 ne
tri 1967 -978 2010 -935 sw
rect 1779 -993 1823 -978
tri 1823 -993 1838 -978 sw
tri 1967 -993 1982 -978 ne
rect 1779 -994 1838 -993
tri 1838 -994 1839 -993 sw
rect 1779 -1000 1939 -994
rect 1779 -1034 1821 -1000
rect 1855 -1034 1893 -1000
rect 1927 -1034 1939 -1000
rect 1779 -1040 1939 -1034
tri 1962 -1060 1982 -1040 se
rect 1982 -1060 2010 -978
tri 1463 -1076 1479 -1060 sw
tri 1952 -1070 1962 -1060 se
rect 1962 -1070 2010 -1060
tri 1566 -1076 1572 -1070 se
rect 1572 -1076 1702 -1070
tri 1946 -1076 1952 -1070 se
rect 1952 -1076 2010 -1070
rect 1435 -1088 1479 -1076
tri 1479 -1088 1491 -1076 sw
tri 1554 -1088 1566 -1076 se
rect 1566 -1088 1584 -1076
rect 1435 -1110 1584 -1088
rect 1618 -1110 1656 -1076
rect 1690 -1110 1702 -1076
rect 1435 -1116 1702 -1110
rect 1867 -1082 2010 -1076
rect 1867 -1116 1879 -1082
rect 1913 -1116 1951 -1082
rect 1985 -1116 2010 -1082
rect 1867 -1122 2010 -1116
rect 1767 -1156 1813 -1144
rect 1767 -1190 1773 -1156
rect 1807 -1190 1813 -1156
rect 1767 -1228 1813 -1190
rect 1767 -1262 1773 -1228
rect 1807 -1262 1813 -1228
rect 1767 -1274 1813 -1262
<< via1 >>
rect 127 1668 179 1674
rect 127 1634 136 1668
rect 136 1634 170 1668
rect 170 1634 179 1668
rect 127 1622 179 1634
rect 127 1562 179 1606
rect 127 1554 136 1562
rect 136 1554 170 1562
rect 170 1554 179 1562
rect 127 1528 136 1537
rect 136 1528 170 1537
rect 170 1528 179 1537
rect 127 1485 179 1528
rect 127 1456 179 1468
rect 127 1422 136 1456
rect 136 1422 170 1456
rect 170 1422 179 1456
rect 127 1416 179 1422
rect 1265 1459 1317 1511
rect 1265 1395 1317 1447
rect 1634 1493 1686 1499
rect 1634 1459 1645 1493
rect 1645 1459 1679 1493
rect 1679 1459 1686 1493
rect 1634 1447 1686 1459
rect 1634 1421 1686 1433
rect 1634 1387 1645 1421
rect 1645 1387 1679 1421
rect 1679 1387 1686 1421
rect 1634 1381 1686 1387
rect 997 1263 1049 1315
rect 997 1199 1049 1251
rect 997 1135 1049 1187
rect 77 1039 129 1091
rect 141 1039 193 1091
rect 725 1027 777 1079
rect 725 963 777 1015
rect 805 1025 857 1077
rect 1818 1071 1870 1077
rect 1818 1037 1830 1071
rect 1830 1037 1864 1071
rect 1864 1037 1870 1071
rect 805 961 857 1013
rect 1818 1025 1870 1037
rect 1459 948 1511 1000
rect 1523 991 1575 1000
rect 1523 957 1548 991
rect 1548 957 1575 991
rect 1523 948 1575 957
rect 1818 999 1870 1011
rect 1818 965 1830 999
rect 1830 965 1864 999
rect 1864 965 1870 999
rect 1818 959 1870 965
rect 1598 867 1650 919
rect 1662 867 1714 919
rect 805 705 817 739
rect 817 705 851 739
rect 851 705 857 739
rect 805 687 857 705
rect 725 666 777 679
rect 725 632 737 666
rect 737 632 777 666
rect 725 627 777 632
rect 805 623 857 675
rect 997 644 1049 648
rect 725 594 777 615
rect 725 563 737 594
rect 737 563 777 594
rect 997 610 1006 644
rect 1006 610 1040 644
rect 1040 610 1049 644
rect 997 596 1049 610
rect 997 572 1049 584
rect 997 538 1006 572
rect 1006 538 1040 572
rect 1040 538 1049 572
rect 1265 692 1317 698
rect 1265 658 1299 692
rect 1299 658 1317 692
rect 1265 646 1317 658
rect 1265 620 1317 634
rect 1265 586 1299 620
rect 1299 586 1317 620
rect 1265 582 1317 586
rect 1508 585 1560 637
rect 997 532 1049 538
rect 1508 518 1560 570
rect 829 43 881 95
rect 893 43 945 95
rect 1050 -528 1102 -519
rect 1050 -562 1056 -528
rect 1056 -562 1090 -528
rect 1090 -562 1102 -528
rect 1050 -571 1102 -562
rect 1114 -528 1166 -519
rect 1114 -562 1147 -528
rect 1147 -562 1166 -528
rect 1114 -571 1166 -562
rect 1791 -637 1843 -585
rect 1855 -637 1907 -585
rect 1473 -671 1525 -665
rect 1537 -671 1589 -665
rect 1473 -705 1499 -671
rect 1499 -705 1525 -671
rect 1537 -705 1571 -671
rect 1571 -705 1589 -671
rect 1473 -717 1525 -705
rect 1537 -717 1589 -705
rect 1605 -839 1657 -787
rect 1669 -839 1721 -787
<< metal2 >>
rect 127 1674 179 1680
rect 127 1606 179 1622
rect 127 1537 179 1554
rect 127 1468 179 1485
tri 115 1135 127 1147 se
rect 127 1135 179 1416
rect 1265 1511 1317 1517
rect 1265 1447 1317 1459
tri 112 1132 115 1135 se
rect 115 1132 179 1135
tri 91 1111 112 1132 se
rect 112 1111 179 1132
rect 997 1315 1049 1321
rect 997 1251 1049 1263
rect 997 1187 1049 1199
tri 71 1091 91 1111 se
rect 91 1091 179 1111
tri 179 1091 199 1111 sw
rect 71 1039 77 1091
rect 129 1039 141 1091
rect 193 1039 199 1091
rect 725 1079 777 1085
rect 725 1015 777 1027
rect 725 679 777 963
rect 725 615 777 627
rect 805 1077 857 1083
rect 805 1013 857 1025
rect 805 739 857 961
rect 805 675 857 687
rect 805 617 857 623
rect 997 648 1049 1135
rect 997 584 1049 596
rect 725 557 777 563
tri 972 557 997 582 se
tri 947 532 972 557 se
rect 972 532 997 557
rect 1265 698 1317 1395
rect 1634 1499 1686 1505
rect 1634 1433 1686 1447
rect 1453 948 1459 1000
rect 1511 948 1523 1000
rect 1575 948 1581 1000
tri 1453 919 1482 948 ne
rect 1482 919 1560 948
tri 1560 927 1581 948 nw
tri 1610 927 1634 951 se
rect 1634 927 1686 1381
rect 1818 1077 1870 1083
rect 1818 1011 1870 1025
tri 1602 919 1610 927 se
rect 1610 919 1686 927
tri 1686 919 1720 953 sw
tri 1482 893 1508 919 ne
rect 1265 634 1317 646
rect 1265 576 1317 582
rect 1508 637 1560 919
rect 1592 867 1598 919
rect 1650 867 1662 919
rect 1714 867 1720 919
tri 941 526 947 532 se
rect 947 526 1049 532
rect 1508 570 1560 585
tri 933 518 941 526 se
rect 941 518 1007 526
tri 1007 518 1015 526 nw
tri 927 512 933 518 se
rect 933 512 1001 518
tri 1001 512 1007 518 nw
tri 923 508 927 512 se
rect 927 508 997 512
tri 997 508 1001 512 nw
tri 861 446 923 508 se
rect 923 446 935 508
tri 935 446 997 508 nw
tri 823 131 861 169 se
rect 861 131 913 446
tri 913 424 935 446 nw
tri 913 131 951 169 sw
rect 823 95 951 131
rect 823 43 829 95
rect 881 43 893 95
rect 945 43 951 95
rect 1044 -571 1050 -519
rect 1102 -571 1114 -519
rect 1166 -571 1172 -519
tri 1502 -630 1508 -624 se
rect 1508 -630 1560 518
tri 1785 -585 1818 -552 se
rect 1818 -585 1870 959
tri 1870 -585 1913 -542 sw
tri 1495 -637 1502 -630 se
rect 1502 -637 1560 -630
tri 1560 -637 1567 -630 sw
rect 1785 -637 1791 -585
rect 1843 -637 1855 -585
rect 1907 -637 1913 -585
tri 1467 -665 1495 -637 se
rect 1495 -665 1567 -637
tri 1567 -665 1595 -637 sw
rect 1467 -717 1473 -665
rect 1525 -717 1537 -665
rect 1589 -717 1595 -665
rect 1599 -839 1605 -787
rect 1657 -839 1669 -787
rect 1721 -839 1727 -787
use sky130_fd_pr__nfet_01v8__example_55959141808379  sky130_fd_pr__nfet_01v8__example_55959141808379_0
timestamp 1649977179
transform -1 0 206 0 -1 1190
box -28 0 148 97
use sky130_fd_pr__nfet_01v8__example_55959141808380  sky130_fd_pr__nfet_01v8__example_55959141808380_0
timestamp 1649977179
transform 1 0 262 0 -1 1190
box -28 0 148 97
use sky130_fd_pr__nfet_01v8__example_55959141808382  sky130_fd_pr__nfet_01v8__example_55959141808382_0
timestamp 1649977179
transform -1 0 1810 0 1 1289
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808383  sky130_fd_pr__nfet_01v8__example_55959141808383_0
timestamp 1649977179
transform 1 0 1866 0 1 1289
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808423  sky130_fd_pr__nfet_01v8__example_55959141808423_0
timestamp 1649977179
transform -1 0 1868 0 1 -1276
box -28 0 184 97
use sky130_fd_pr__nfet_01v8__example_55959141808424  sky130_fd_pr__nfet_01v8__example_55959141808424_0
timestamp 1649977179
transform -1 0 1970 0 -1 1095
box -28 0 484 63
use sky130_fd_pr__nfet_01v8__example_55959141808426  sky130_fd_pr__nfet_01v8__example_55959141808426_0
timestamp 1649977179
transform 1 0 181 0 1 1685
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808426  sky130_fd_pr__nfet_01v8__example_55959141808426_1
timestamp 1649977179
transform 1 0 181 0 1 1391
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808426  sky130_fd_pr__nfet_01v8__example_55959141808426_2
timestamp 1649977179
transform 1 0 777 0 1 1391
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808426  sky130_fd_pr__nfet_01v8__example_55959141808426_3
timestamp 1649977179
transform 1 0 777 0 -1 1889
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808427  sky130_fd_pr__nfet_01v8__example_55959141808427_0
timestamp 1649977179
transform -1 0 1280 0 -1 1237
box -28 0 316 97
use sky130_fd_pr__nfet_01v8__example_55959141808427  sky130_fd_pr__nfet_01v8__example_55959141808427_1
timestamp 1649977179
transform -1 0 936 0 -1 1237
box -28 0 316 97
use sky130_fd_pr__nfet_01v8__example_55959141808428  sky130_fd_pr__nfet_01v8__example_55959141808428_0
timestamp 1649977179
transform -1 0 1634 0 1 1289
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808429  sky130_fd_pr__nfet_01v8__example_55959141808429_0
timestamp 1649977179
transform -1 0 1288 0 -1 681
box -28 0 148 267
use sky130_fd_pr__pfet_01v8__example_55959141808431  sky130_fd_pr__pfet_01v8__example_55959141808431_0
timestamp 1649977179
transform -1 0 516 0 -1 676
box -28 0 148 267
use sky130_fd_pr__pfet_01v8__example_55959141808432  sky130_fd_pr__pfet_01v8__example_55959141808432_0
timestamp 1649977179
transform 1 0 572 0 -1 676
box -28 0 148 267
use sky130_fd_pr__pfet_01v8__example_55959141808433  sky130_fd_pr__pfet_01v8__example_55959141808433_0
timestamp 1649977179
transform 1 0 130 0 -1 357
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808435  sky130_fd_pr__pfet_01v8__example_55959141808435_0
timestamp 1649977179
transform 1 0 130 0 -1 676
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808617  sky130_fd_pr__pfet_01v8__example_55959141808617_0
timestamp 1649977179
transform 0 -1 1350 -1 0 -777
box -28 0 78 97
use sky130_fd_pr__pfet_01v8__example_55959141808617  sky130_fd_pr__pfet_01v8__example_55959141808617_1
timestamp 1649977179
transform 0 -1 1350 1 0 -721
box -28 0 78 97
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1649977179
transform -1 0 1037 0 -1 1693
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1649977179
transform -1 0 448 0 -1 1674
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1649977179
transform 0 -1 1002 1 0 1498
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1649977179
transform 0 -1 1333 -1 0 692
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1649977179
transform 1 0 83 0 1 877
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1649977179
transform -1 0 147 0 -1 999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1649977179
transform 1 0 363 0 1 646
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1649977179
transform 1 0 247 0 1 779
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1649977179
transform 0 -1 1864 -1 0 1071
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1649977179
transform 1 0 817 0 1 705
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1649977179
transform 0 -1 2015 -1 0 1082
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1649977179
transform 0 -1 1151 1 0 575
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1649977179
transform 1 0 1898 0 -1 817
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1649977179
transform 1 0 1045 0 1 779
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1649977179
transform 0 -1 1040 -1 0 644
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1649977179
transform 1 0 519 0 1 878
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1649977179
transform 0 -1 1855 1 0 1203
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1649977179
transform -1 0 637 0 1 1128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1649977179
transform -1 0 809 0 1 1128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_2
timestamp 1649977179
transform -1 0 981 0 1 1128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_3
timestamp 1649977179
transform -1 0 1153 0 1 1128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_4
timestamp 1649977179
transform -1 0 251 0 1 1128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_5
timestamp 1649977179
transform 1 0 703 0 -1 666
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_6
timestamp 1649977179
transform -1 0 1325 0 1 1128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1649977179
transform 0 -1 406 1 0 1404
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1649977179
transform 0 -1 853 1 0 136
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1649977179
transform 0 -1 119 1 0 136
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1649977179
transform 0 -1 561 1 0 136
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_0
timestamp 1649977179
transform 0 -1 17 1 0 1296
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808440  sky130_fd_pr__via_l1m1__example_55959141808440_0
timestamp 1649977179
transform 0 -1 1181 -1 0 1990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1649977179
transform 0 -1 857 -1 0 1083
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1649977179
transform 0 -1 1317 -1 0 704
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1649977179
transform 0 -1 1317 -1 0 1517
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1649977179
transform 0 -1 777 1 0 957
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1649977179
transform 0 -1 777 1 0 557
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1649977179
transform 0 -1 857 -1 0 745
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1649977179
transform 1 0 823 0 1 43
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1649977179
transform 0 1 997 -1 0 654
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_0
timestamp 1649977179
transform 0 1 997 -1 0 1321
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1649977179
transform 0 -1 1970 -1 0 1185
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1649977179
transform 0 -1 1336 -1 0 779
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1649977179
transform 0 -1 1687 -1 0 1195
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1649977179
transform 0 -1 1640 -1 0 1987
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1649977179
transform 0 -1 1817 -1 0 1981
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1649977179
transform 0 -1 949 -1 0 923
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_1
timestamp 1649977179
transform 0 -1 1293 -1 0 1004
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808394  sky130_fd_pr__via_pol1__example_55959141808394_0
timestamp 1649977179
transform 0 -1 1145 1 0 1940
box 0 0 1 1
<< labels >>
flabel metal2 s 1675 -839 1727 -787 3 FreeSans 520 90 0 0 DM[1]
port 1 nsew
flabel metal2 s 1701 -813 1701 -813 3 FreeSans 520 90 0 0 DM[1]
port 1 nsew
flabel metal1 s 0 124 34 326 3 FreeSans 400 0 0 0 VCC_IO
port 2 nsew
flabel metal1 s 0 354 34 484 3 FreeSans 400 0 0 0 VPB
port 3 nsew
flabel metal1 s 35 960 69 1005 3 FreeSans 400 0 0 0 OUT_H_N
port 4 nsew
flabel metal1 s 352 640 386 686 3 FreeSans 400 0 0 0 OUT_H
port 5 nsew
flabel metal1 s 1726 1462 1760 1496 0 FreeSans 400 180 0 0 RST_H
port 6 nsew
flabel metal1 s 1926 1593 1960 1627 0 FreeSans 400 180 0 0 SET_H
port 7 nsew
flabel metal1 s 0 1826 34 2016 3 FreeSans 400 0 0 0 VPWR
port 8 nsew
flabel metal1 s 1384 636 1418 669 0 FreeSans 200 180 0 0 HLD_H_N
port 9 nsew
flabel comment s 1553 982 1553 982 0 FreeSans 200 180 0 0 IN_I_N
flabel comment s 398 1292 398 1292 0 FreeSans 200 180 0 0 VGND
flabel comment s 1661 1384 1661 1384 0 FreeSans 200 180 0 0 FBK_N
flabel comment s 1840 1382 1840 1382 0 FreeSans 200 180 0 0 VGND
flabel comment s 2016 2012 2016 2012 0 FreeSans 200 0 0 0 RST_H
flabel comment s 1807 2012 1807 2012 0 FreeSans 200 0 0 0 SET_H
flabel comment s 626 991 626 991 0 FreeSans 200 0 0 0 OUT_H
flabel comment s 1357 800 1357 800 0 FreeSans 200 0 0 0 FBK_N
flabel comment s 1741 1078 1741 1078 0 FreeSans 200 0 0 0 VGND
flabel comment s 824 992 824 992 0 FreeSans 200 180 0 0 IN_I
flabel comment s 1472 1078 1472 1078 0 FreeSans 200 180 0 0 IN_I_N
flabel comment s 1525 600 1525 600 0 FreeSans 440 0 0 0 1
<< properties >>
string GDS_END 7787470
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7754000
<< end >>
