magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< locali >>
rect 59399 66138 59433 66154
rect 59399 66088 59433 66104
rect 59870 65435 59904 65469
rect 59399 64724 59433 64740
rect 59399 64674 59433 64690
rect 59399 63310 59433 63326
rect 59399 63260 59433 63276
rect 11510 60571 11689 60605
rect 54197 60591 54213 60625
rect 54247 60605 54373 60625
rect 54247 60591 54518 60605
rect 54339 60571 54518 60591
rect 11655 60405 11689 60571
rect 11655 60371 11781 60405
rect 11815 60371 11831 60405
rect 11655 60275 11781 60309
rect 11815 60275 11831 60309
rect 11655 60109 11689 60275
rect 11510 60075 11689 60109
rect 54339 60089 54518 60109
rect 54197 60055 54213 60089
rect 54247 60075 54518 60089
rect 54247 60055 54373 60075
rect 11510 59781 11689 59815
rect 54197 59801 54213 59835
rect 54247 59815 54373 59835
rect 54247 59801 54518 59815
rect 54339 59781 54518 59801
rect 11655 59615 11689 59781
rect 11655 59581 11781 59615
rect 11815 59581 11831 59615
rect 11655 59485 11781 59519
rect 11815 59485 11831 59519
rect 11655 59319 11689 59485
rect 11510 59285 11689 59319
rect 54339 59299 54518 59319
rect 54197 59265 54213 59299
rect 54247 59285 54518 59299
rect 54247 59265 54373 59285
rect 11510 58991 11689 59025
rect 54197 59011 54213 59045
rect 54247 59025 54373 59045
rect 54247 59011 54518 59025
rect 54339 58991 54518 59011
rect 11655 58825 11689 58991
rect 11655 58791 11781 58825
rect 11815 58791 11831 58825
rect 11655 58695 11781 58729
rect 11815 58695 11831 58729
rect 11655 58529 11689 58695
rect 11510 58495 11689 58529
rect 54339 58509 54518 58529
rect 54197 58475 54213 58509
rect 54247 58495 54518 58509
rect 54247 58475 54373 58495
rect 11510 58201 11689 58235
rect 54197 58221 54213 58255
rect 54247 58235 54373 58255
rect 54247 58221 54518 58235
rect 54339 58201 54518 58221
rect 11655 58035 11689 58201
rect 11655 58001 11781 58035
rect 11815 58001 11831 58035
rect 11655 57905 11781 57939
rect 11815 57905 11831 57939
rect 11655 57739 11689 57905
rect 11510 57705 11689 57739
rect 54339 57719 54518 57739
rect 54197 57685 54213 57719
rect 54247 57705 54518 57719
rect 54247 57685 54373 57705
rect 11510 57411 11689 57445
rect 54197 57431 54213 57465
rect 54247 57445 54373 57465
rect 54247 57431 54518 57445
rect 54339 57411 54518 57431
rect 11655 57245 11689 57411
rect 11655 57211 11781 57245
rect 11815 57211 11831 57245
rect 11655 57115 11781 57149
rect 11815 57115 11831 57149
rect 11655 56949 11689 57115
rect 11510 56915 11689 56949
rect 54339 56929 54518 56949
rect 54197 56895 54213 56929
rect 54247 56915 54518 56929
rect 54247 56895 54373 56915
rect 11510 56621 11689 56655
rect 54197 56641 54213 56675
rect 54247 56655 54373 56675
rect 54247 56641 54518 56655
rect 54339 56621 54518 56641
rect 11655 56455 11689 56621
rect 11655 56421 11781 56455
rect 11815 56421 11831 56455
rect 11655 56325 11781 56359
rect 11815 56325 11831 56359
rect 11655 56159 11689 56325
rect 11510 56125 11689 56159
rect 54339 56139 54518 56159
rect 54197 56105 54213 56139
rect 54247 56125 54518 56139
rect 54247 56105 54373 56125
rect 11510 55831 11689 55865
rect 54197 55851 54213 55885
rect 54247 55865 54373 55885
rect 54247 55851 54518 55865
rect 54339 55831 54518 55851
rect 11655 55665 11689 55831
rect 11655 55631 11781 55665
rect 11815 55631 11831 55665
rect 11655 55535 11781 55569
rect 11815 55535 11831 55569
rect 11655 55369 11689 55535
rect 11510 55335 11689 55369
rect 54339 55349 54518 55369
rect 54197 55315 54213 55349
rect 54247 55335 54518 55349
rect 54247 55315 54373 55335
rect 11510 55041 11689 55075
rect 54197 55061 54213 55095
rect 54247 55075 54373 55095
rect 54247 55061 54518 55075
rect 54339 55041 54518 55061
rect 11655 54875 11689 55041
rect 11655 54841 11781 54875
rect 11815 54841 11831 54875
rect 11655 54745 11781 54779
rect 11815 54745 11831 54779
rect 11655 54579 11689 54745
rect 11510 54545 11689 54579
rect 54339 54559 54518 54579
rect 54197 54525 54213 54559
rect 54247 54545 54518 54559
rect 54247 54525 54373 54545
rect 11510 54251 11689 54285
rect 54197 54271 54213 54305
rect 54247 54285 54373 54305
rect 54247 54271 54518 54285
rect 54339 54251 54518 54271
rect 11655 54085 11689 54251
rect 11655 54051 11781 54085
rect 11815 54051 11831 54085
rect 11655 53955 11781 53989
rect 11815 53955 11831 53989
rect 11655 53789 11689 53955
rect 11510 53755 11689 53789
rect 54339 53769 54518 53789
rect 54197 53735 54213 53769
rect 54247 53755 54518 53769
rect 54247 53735 54373 53755
rect 11510 53461 11689 53495
rect 54197 53481 54213 53515
rect 54247 53495 54373 53515
rect 54247 53481 54518 53495
rect 54339 53461 54518 53481
rect 11655 53295 11689 53461
rect 11655 53261 11781 53295
rect 11815 53261 11831 53295
rect 11655 53165 11781 53199
rect 11815 53165 11831 53199
rect 11655 52999 11689 53165
rect 11510 52965 11689 52999
rect 54339 52979 54518 52999
rect 54197 52945 54213 52979
rect 54247 52965 54518 52979
rect 54247 52945 54373 52965
rect 11510 52671 11689 52705
rect 54197 52691 54213 52725
rect 54247 52705 54373 52725
rect 54247 52691 54518 52705
rect 54339 52671 54518 52691
rect 11655 52505 11689 52671
rect 11655 52471 11781 52505
rect 11815 52471 11831 52505
rect 11655 52375 11781 52409
rect 11815 52375 11831 52409
rect 11655 52209 11689 52375
rect 11510 52175 11689 52209
rect 54339 52189 54518 52209
rect 54197 52155 54213 52189
rect 54247 52175 54518 52189
rect 54247 52155 54373 52175
rect 11510 51881 11689 51915
rect 54197 51901 54213 51935
rect 54247 51915 54373 51935
rect 54247 51901 54518 51915
rect 54339 51881 54518 51901
rect 11655 51715 11689 51881
rect 11655 51681 11781 51715
rect 11815 51681 11831 51715
rect 11655 51585 11781 51619
rect 11815 51585 11831 51619
rect 11655 51419 11689 51585
rect 11510 51385 11689 51419
rect 54339 51399 54518 51419
rect 54197 51365 54213 51399
rect 54247 51385 54518 51399
rect 54247 51365 54373 51385
rect 11510 51091 11689 51125
rect 54197 51111 54213 51145
rect 54247 51125 54373 51145
rect 54247 51111 54518 51125
rect 54339 51091 54518 51111
rect 11655 50925 11689 51091
rect 11655 50891 11781 50925
rect 11815 50891 11831 50925
rect 11655 50795 11781 50829
rect 11815 50795 11831 50829
rect 11655 50629 11689 50795
rect 11510 50595 11689 50629
rect 54339 50609 54518 50629
rect 54197 50575 54213 50609
rect 54247 50595 54518 50609
rect 54247 50575 54373 50595
rect 11510 50301 11689 50335
rect 54197 50321 54213 50355
rect 54247 50335 54373 50355
rect 54247 50321 54518 50335
rect 54339 50301 54518 50321
rect 11655 50135 11689 50301
rect 11655 50101 11781 50135
rect 11815 50101 11831 50135
rect 11655 50005 11781 50039
rect 11815 50005 11831 50039
rect 11655 49839 11689 50005
rect 11510 49805 11689 49839
rect 54339 49819 54518 49839
rect 54197 49785 54213 49819
rect 54247 49805 54518 49819
rect 54247 49785 54373 49805
rect 11510 49511 11689 49545
rect 54197 49531 54213 49565
rect 54247 49545 54373 49565
rect 54247 49531 54518 49545
rect 54339 49511 54518 49531
rect 11655 49345 11689 49511
rect 11655 49311 11781 49345
rect 11815 49311 11831 49345
rect 11655 49215 11781 49249
rect 11815 49215 11831 49249
rect 11655 49049 11689 49215
rect 11510 49015 11689 49049
rect 54339 49029 54518 49049
rect 54197 48995 54213 49029
rect 54247 49015 54518 49029
rect 54247 48995 54373 49015
rect 11510 48721 11689 48755
rect 54197 48741 54213 48775
rect 54247 48755 54373 48775
rect 54247 48741 54518 48755
rect 54339 48721 54518 48741
rect 11655 48555 11689 48721
rect 11655 48521 11781 48555
rect 11815 48521 11831 48555
rect 11655 48425 11781 48459
rect 11815 48425 11831 48459
rect 11655 48259 11689 48425
rect 11510 48225 11689 48259
rect 54339 48239 54518 48259
rect 54197 48205 54213 48239
rect 54247 48225 54518 48239
rect 54247 48205 54373 48225
rect 11510 47931 11689 47965
rect 54197 47951 54213 47985
rect 54247 47965 54373 47985
rect 54247 47951 54518 47965
rect 54339 47931 54518 47951
rect 11655 47765 11689 47931
rect 11655 47731 11781 47765
rect 11815 47731 11831 47765
rect 11655 47635 11781 47669
rect 11815 47635 11831 47669
rect 11655 47469 11689 47635
rect 11510 47435 11689 47469
rect 54339 47449 54518 47469
rect 54197 47415 54213 47449
rect 54247 47435 54518 47449
rect 54247 47415 54373 47435
rect 11510 47141 11689 47175
rect 54197 47161 54213 47195
rect 54247 47175 54373 47195
rect 54247 47161 54518 47175
rect 54339 47141 54518 47161
rect 11655 46975 11689 47141
rect 11655 46941 11781 46975
rect 11815 46941 11831 46975
rect 11655 46845 11781 46879
rect 11815 46845 11831 46879
rect 11655 46679 11689 46845
rect 11510 46645 11689 46679
rect 54339 46659 54518 46679
rect 54197 46625 54213 46659
rect 54247 46645 54518 46659
rect 54247 46625 54373 46645
rect 11510 46351 11689 46385
rect 54197 46371 54213 46405
rect 54247 46385 54373 46405
rect 54247 46371 54518 46385
rect 54339 46351 54518 46371
rect 11655 46185 11689 46351
rect 11655 46151 11781 46185
rect 11815 46151 11831 46185
rect 11655 46055 11781 46089
rect 11815 46055 11831 46089
rect 11655 45889 11689 46055
rect 11510 45855 11689 45889
rect 54339 45869 54518 45889
rect 54197 45835 54213 45869
rect 54247 45855 54518 45869
rect 54247 45835 54373 45855
rect 11510 45561 11689 45595
rect 54197 45581 54213 45615
rect 54247 45595 54373 45615
rect 54247 45581 54518 45595
rect 54339 45561 54518 45581
rect 11655 45395 11689 45561
rect 11655 45361 11781 45395
rect 11815 45361 11831 45395
rect 11655 45265 11781 45299
rect 11815 45265 11831 45299
rect 11655 45099 11689 45265
rect 11510 45065 11689 45099
rect 54339 45079 54518 45099
rect 54197 45045 54213 45079
rect 54247 45065 54518 45079
rect 54247 45045 54373 45065
rect 11510 44771 11689 44805
rect 54197 44791 54213 44825
rect 54247 44805 54373 44825
rect 54247 44791 54518 44805
rect 54339 44771 54518 44791
rect 11655 44605 11689 44771
rect 11655 44571 11781 44605
rect 11815 44571 11831 44605
rect 11655 44475 11781 44509
rect 11815 44475 11831 44509
rect 11655 44309 11689 44475
rect 11510 44275 11689 44309
rect 54339 44289 54518 44309
rect 54197 44255 54213 44289
rect 54247 44275 54518 44289
rect 54247 44255 54373 44275
rect 11510 43981 11689 44015
rect 54197 44001 54213 44035
rect 54247 44015 54373 44035
rect 54247 44001 54518 44015
rect 54339 43981 54518 44001
rect 11655 43815 11689 43981
rect 11655 43781 11781 43815
rect 11815 43781 11831 43815
rect 11655 43685 11781 43719
rect 11815 43685 11831 43719
rect 11655 43519 11689 43685
rect 11510 43485 11689 43519
rect 54339 43499 54518 43519
rect 54197 43465 54213 43499
rect 54247 43485 54518 43499
rect 54247 43465 54373 43485
rect 11510 43191 11689 43225
rect 54197 43211 54213 43245
rect 54247 43225 54373 43245
rect 54247 43211 54518 43225
rect 54339 43191 54518 43211
rect 11655 43025 11689 43191
rect 11655 42991 11781 43025
rect 11815 42991 11831 43025
rect 11655 42895 11781 42929
rect 11815 42895 11831 42929
rect 11655 42729 11689 42895
rect 11510 42695 11689 42729
rect 54339 42709 54518 42729
rect 54197 42675 54213 42709
rect 54247 42695 54518 42709
rect 54247 42675 54373 42695
rect 11510 42401 11689 42435
rect 54197 42421 54213 42455
rect 54247 42435 54373 42455
rect 54247 42421 54518 42435
rect 54339 42401 54518 42421
rect 11655 42235 11689 42401
rect 11655 42201 11781 42235
rect 11815 42201 11831 42235
rect 11655 42105 11781 42139
rect 11815 42105 11831 42139
rect 11655 41939 11689 42105
rect 11510 41905 11689 41939
rect 54339 41919 54518 41939
rect 54197 41885 54213 41919
rect 54247 41905 54518 41919
rect 54247 41885 54373 41905
rect 11510 41611 11689 41645
rect 54197 41631 54213 41665
rect 54247 41645 54373 41665
rect 54247 41631 54518 41645
rect 54339 41611 54518 41631
rect 11655 41445 11689 41611
rect 11655 41411 11781 41445
rect 11815 41411 11831 41445
rect 11655 41315 11781 41349
rect 11815 41315 11831 41349
rect 11655 41149 11689 41315
rect 11510 41115 11689 41149
rect 54339 41129 54518 41149
rect 54197 41095 54213 41129
rect 54247 41115 54518 41129
rect 54247 41095 54373 41115
rect 11510 40821 11689 40855
rect 54197 40841 54213 40875
rect 54247 40855 54373 40875
rect 54247 40841 54518 40855
rect 54339 40821 54518 40841
rect 11655 40655 11689 40821
rect 11655 40621 11781 40655
rect 11815 40621 11831 40655
rect 11655 40525 11781 40559
rect 11815 40525 11831 40559
rect 11655 40359 11689 40525
rect 11510 40325 11689 40359
rect 54339 40339 54518 40359
rect 54197 40305 54213 40339
rect 54247 40325 54518 40339
rect 54247 40305 54373 40325
rect 11510 40031 11689 40065
rect 54197 40051 54213 40085
rect 54247 40065 54373 40085
rect 54247 40051 54518 40065
rect 54339 40031 54518 40051
rect 11655 39865 11689 40031
rect 11655 39831 11781 39865
rect 11815 39831 11831 39865
rect 11655 39735 11781 39769
rect 11815 39735 11831 39769
rect 11655 39569 11689 39735
rect 11510 39535 11689 39569
rect 54339 39549 54518 39569
rect 54197 39515 54213 39549
rect 54247 39535 54518 39549
rect 54247 39515 54373 39535
rect 11510 39241 11689 39275
rect 54197 39261 54213 39295
rect 54247 39275 54373 39295
rect 54247 39261 54518 39275
rect 54339 39241 54518 39261
rect 11655 39075 11689 39241
rect 11655 39041 11781 39075
rect 11815 39041 11831 39075
rect 11655 38945 11781 38979
rect 11815 38945 11831 38979
rect 11655 38779 11689 38945
rect 11510 38745 11689 38779
rect 54339 38759 54518 38779
rect 54197 38725 54213 38759
rect 54247 38745 54518 38759
rect 54247 38725 54373 38745
rect 11510 38451 11689 38485
rect 54197 38471 54213 38505
rect 54247 38485 54373 38505
rect 54247 38471 54518 38485
rect 54339 38451 54518 38471
rect 11655 38285 11689 38451
rect 11655 38251 11781 38285
rect 11815 38251 11831 38285
rect 11655 38155 11781 38189
rect 11815 38155 11831 38189
rect 11655 37989 11689 38155
rect 11510 37955 11689 37989
rect 54339 37969 54518 37989
rect 54197 37935 54213 37969
rect 54247 37955 54518 37969
rect 54247 37935 54373 37955
rect 11510 37661 11689 37695
rect 54197 37681 54213 37715
rect 54247 37695 54373 37715
rect 54247 37681 54518 37695
rect 54339 37661 54518 37681
rect 11655 37495 11689 37661
rect 11655 37461 11781 37495
rect 11815 37461 11831 37495
rect 11655 37365 11781 37399
rect 11815 37365 11831 37399
rect 11655 37199 11689 37365
rect 11510 37165 11689 37199
rect 54339 37179 54518 37199
rect 54197 37145 54213 37179
rect 54247 37165 54518 37179
rect 54247 37145 54373 37165
rect 11510 36871 11689 36905
rect 54197 36891 54213 36925
rect 54247 36905 54373 36925
rect 54247 36891 54518 36905
rect 54339 36871 54518 36891
rect 11655 36705 11689 36871
rect 11655 36671 11781 36705
rect 11815 36671 11831 36705
rect 11655 36575 11781 36609
rect 11815 36575 11831 36609
rect 11655 36409 11689 36575
rect 11510 36375 11689 36409
rect 54339 36389 54518 36409
rect 54197 36355 54213 36389
rect 54247 36375 54518 36389
rect 54247 36355 54373 36375
rect 11510 36081 11689 36115
rect 54197 36101 54213 36135
rect 54247 36115 54373 36135
rect 54247 36101 54518 36115
rect 54339 36081 54518 36101
rect 11655 35915 11689 36081
rect 11655 35881 11781 35915
rect 11815 35881 11831 35915
rect 11655 35785 11781 35819
rect 11815 35785 11831 35819
rect 11655 35619 11689 35785
rect 11510 35585 11689 35619
rect 54339 35599 54518 35619
rect 54197 35565 54213 35599
rect 54247 35585 54518 35599
rect 54247 35565 54373 35585
rect 11510 35291 11689 35325
rect 54197 35311 54213 35345
rect 54247 35325 54373 35345
rect 54247 35311 54518 35325
rect 54339 35291 54518 35311
rect 11655 35125 11689 35291
rect 11655 35091 11781 35125
rect 11815 35091 11831 35125
rect 11655 34995 11781 35029
rect 11815 34995 11831 35029
rect 11655 34829 11689 34995
rect 11510 34795 11689 34829
rect 54339 34809 54518 34829
rect 54197 34775 54213 34809
rect 54247 34795 54518 34809
rect 54247 34775 54373 34795
rect 11510 34501 11689 34535
rect 54197 34521 54213 34555
rect 54247 34535 54373 34555
rect 54247 34521 54518 34535
rect 54339 34501 54518 34521
rect 11655 34335 11689 34501
rect 11655 34301 11781 34335
rect 11815 34301 11831 34335
rect 11655 34205 11781 34239
rect 11815 34205 11831 34239
rect 11655 34039 11689 34205
rect 11510 34005 11689 34039
rect 54339 34019 54518 34039
rect 54197 33985 54213 34019
rect 54247 34005 54518 34019
rect 54247 33985 54373 34005
rect 11510 33711 11689 33745
rect 54197 33731 54213 33765
rect 54247 33745 54373 33765
rect 54247 33731 54518 33745
rect 54339 33711 54518 33731
rect 11655 33545 11689 33711
rect 11655 33511 11781 33545
rect 11815 33511 11831 33545
rect 11655 33415 11781 33449
rect 11815 33415 11831 33449
rect 11655 33249 11689 33415
rect 11510 33215 11689 33249
rect 54339 33229 54518 33249
rect 54197 33195 54213 33229
rect 54247 33215 54518 33229
rect 54247 33195 54373 33215
rect 11510 32921 11689 32955
rect 54197 32941 54213 32975
rect 54247 32955 54373 32975
rect 54247 32941 54518 32955
rect 54339 32921 54518 32941
rect 11655 32755 11689 32921
rect 11655 32721 11781 32755
rect 11815 32721 11831 32755
rect 11655 32625 11781 32659
rect 11815 32625 11831 32659
rect 11655 32459 11689 32625
rect 11510 32425 11689 32459
rect 54339 32439 54518 32459
rect 54197 32405 54213 32439
rect 54247 32425 54518 32439
rect 54247 32405 54373 32425
rect 11510 32131 11689 32165
rect 54197 32151 54213 32185
rect 54247 32165 54373 32185
rect 54247 32151 54518 32165
rect 54339 32131 54518 32151
rect 11655 31965 11689 32131
rect 11655 31931 11781 31965
rect 11815 31931 11831 31965
rect 11655 31835 11781 31869
rect 11815 31835 11831 31869
rect 11655 31669 11689 31835
rect 11510 31635 11689 31669
rect 54339 31649 54518 31669
rect 54197 31615 54213 31649
rect 54247 31635 54518 31649
rect 54247 31615 54373 31635
rect 11510 31341 11689 31375
rect 54197 31361 54213 31395
rect 54247 31375 54373 31395
rect 54247 31361 54518 31375
rect 54339 31341 54518 31361
rect 11655 31175 11689 31341
rect 11655 31141 11781 31175
rect 11815 31141 11831 31175
rect 11655 31045 11781 31079
rect 11815 31045 11831 31079
rect 11655 30879 11689 31045
rect 11510 30845 11689 30879
rect 54339 30859 54518 30879
rect 54197 30825 54213 30859
rect 54247 30845 54518 30859
rect 54247 30825 54373 30845
rect 11510 30551 11689 30585
rect 54197 30571 54213 30605
rect 54247 30585 54373 30605
rect 54247 30571 54518 30585
rect 54339 30551 54518 30571
rect 11655 30385 11689 30551
rect 11655 30351 11781 30385
rect 11815 30351 11831 30385
rect 11655 30255 11781 30289
rect 11815 30255 11831 30289
rect 11655 30089 11689 30255
rect 11510 30055 11689 30089
rect 54339 30069 54518 30089
rect 54197 30035 54213 30069
rect 54247 30055 54518 30069
rect 54247 30035 54373 30055
rect 11510 29761 11689 29795
rect 54197 29781 54213 29815
rect 54247 29795 54373 29815
rect 54247 29781 54518 29795
rect 54339 29761 54518 29781
rect 11655 29595 11689 29761
rect 11655 29561 11781 29595
rect 11815 29561 11831 29595
rect 11655 29465 11781 29499
rect 11815 29465 11831 29499
rect 11655 29299 11689 29465
rect 11510 29265 11689 29299
rect 54339 29279 54518 29299
rect 54197 29245 54213 29279
rect 54247 29265 54518 29279
rect 54247 29245 54373 29265
rect 11510 28971 11689 29005
rect 54197 28991 54213 29025
rect 54247 29005 54373 29025
rect 54247 28991 54518 29005
rect 54339 28971 54518 28991
rect 11655 28805 11689 28971
rect 11655 28771 11781 28805
rect 11815 28771 11831 28805
rect 11655 28675 11781 28709
rect 11815 28675 11831 28709
rect 11655 28509 11689 28675
rect 11510 28475 11689 28509
rect 54339 28489 54518 28509
rect 54197 28455 54213 28489
rect 54247 28475 54518 28489
rect 54247 28455 54373 28475
rect 11510 28181 11689 28215
rect 54197 28201 54213 28235
rect 54247 28215 54373 28235
rect 54247 28201 54518 28215
rect 54339 28181 54518 28201
rect 11655 28015 11689 28181
rect 11655 27981 11781 28015
rect 11815 27981 11831 28015
rect 11655 27885 11781 27919
rect 11815 27885 11831 27919
rect 11655 27719 11689 27885
rect 11510 27685 11689 27719
rect 54339 27699 54518 27719
rect 54197 27665 54213 27699
rect 54247 27685 54518 27699
rect 54247 27665 54373 27685
rect 11510 27391 11689 27425
rect 54197 27411 54213 27445
rect 54247 27425 54373 27445
rect 54247 27411 54518 27425
rect 54339 27391 54518 27411
rect 11655 27225 11689 27391
rect 11655 27191 11781 27225
rect 11815 27191 11831 27225
rect 11655 27095 11781 27129
rect 11815 27095 11831 27129
rect 11655 26929 11689 27095
rect 11510 26895 11689 26929
rect 54339 26909 54518 26929
rect 54197 26875 54213 26909
rect 54247 26895 54518 26909
rect 54247 26875 54373 26895
rect 11510 26601 11689 26635
rect 54197 26621 54213 26655
rect 54247 26635 54373 26655
rect 54247 26621 54518 26635
rect 54339 26601 54518 26621
rect 11655 26435 11689 26601
rect 11655 26401 11781 26435
rect 11815 26401 11831 26435
rect 11655 26305 11781 26339
rect 11815 26305 11831 26339
rect 11655 26139 11689 26305
rect 11510 26105 11689 26139
rect 54339 26119 54518 26139
rect 54197 26085 54213 26119
rect 54247 26105 54518 26119
rect 54247 26085 54373 26105
rect 11510 25811 11689 25845
rect 54197 25831 54213 25865
rect 54247 25845 54373 25865
rect 54247 25831 54518 25845
rect 54339 25811 54518 25831
rect 11655 25645 11689 25811
rect 11655 25611 11781 25645
rect 11815 25611 11831 25645
rect 11655 25515 11781 25549
rect 11815 25515 11831 25549
rect 11655 25349 11689 25515
rect 11510 25315 11689 25349
rect 54339 25329 54518 25349
rect 54197 25295 54213 25329
rect 54247 25315 54518 25329
rect 54247 25295 54373 25315
rect 11510 25021 11689 25055
rect 54197 25041 54213 25075
rect 54247 25055 54373 25075
rect 54247 25041 54518 25055
rect 54339 25021 54518 25041
rect 11655 24855 11689 25021
rect 11655 24821 11781 24855
rect 11815 24821 11831 24855
rect 11655 24725 11781 24759
rect 11815 24725 11831 24759
rect 11655 24559 11689 24725
rect 11510 24525 11689 24559
rect 54339 24539 54518 24559
rect 54197 24505 54213 24539
rect 54247 24525 54518 24539
rect 54247 24505 54373 24525
rect 11510 24231 11689 24265
rect 54197 24251 54213 24285
rect 54247 24265 54373 24285
rect 54247 24251 54518 24265
rect 54339 24231 54518 24251
rect 11655 24065 11689 24231
rect 11655 24031 11781 24065
rect 11815 24031 11831 24065
rect 11655 23935 11781 23969
rect 11815 23935 11831 23969
rect 11655 23769 11689 23935
rect 11510 23735 11689 23769
rect 54339 23749 54518 23769
rect 54197 23715 54213 23749
rect 54247 23735 54518 23749
rect 54247 23715 54373 23735
rect 11510 23441 11689 23475
rect 54197 23461 54213 23495
rect 54247 23475 54373 23495
rect 54247 23461 54518 23475
rect 54339 23441 54518 23461
rect 11655 23275 11689 23441
rect 11655 23241 11781 23275
rect 11815 23241 11831 23275
rect 11655 23145 11781 23179
rect 11815 23145 11831 23179
rect 11655 22979 11689 23145
rect 11510 22945 11689 22979
rect 54339 22959 54518 22979
rect 54197 22925 54213 22959
rect 54247 22945 54518 22959
rect 54247 22925 54373 22945
rect 11510 22651 11689 22685
rect 54197 22671 54213 22705
rect 54247 22685 54373 22705
rect 54247 22671 54518 22685
rect 54339 22651 54518 22671
rect 11655 22485 11689 22651
rect 11655 22451 11781 22485
rect 11815 22451 11831 22485
rect 11655 22355 11781 22389
rect 11815 22355 11831 22389
rect 11655 22189 11689 22355
rect 11510 22155 11689 22189
rect 54339 22169 54518 22189
rect 54197 22135 54213 22169
rect 54247 22155 54518 22169
rect 54247 22135 54373 22155
rect 11510 21861 11689 21895
rect 54197 21881 54213 21915
rect 54247 21895 54373 21915
rect 54247 21881 54518 21895
rect 54339 21861 54518 21881
rect 11655 21695 11689 21861
rect 11655 21661 11781 21695
rect 11815 21661 11831 21695
rect 11655 21565 11781 21599
rect 11815 21565 11831 21599
rect 11655 21399 11689 21565
rect 11510 21365 11689 21399
rect 54339 21379 54518 21399
rect 54197 21345 54213 21379
rect 54247 21365 54518 21379
rect 54247 21345 54373 21365
rect 11510 21071 11689 21105
rect 54197 21091 54213 21125
rect 54247 21105 54373 21125
rect 54247 21091 54518 21105
rect 54339 21071 54518 21091
rect 11655 20905 11689 21071
rect 11655 20871 11781 20905
rect 11815 20871 11831 20905
rect 11655 20775 11781 20809
rect 11815 20775 11831 20809
rect 11655 20609 11689 20775
rect 11510 20575 11689 20609
rect 54339 20589 54518 20609
rect 54197 20555 54213 20589
rect 54247 20575 54518 20589
rect 54247 20555 54373 20575
rect 11510 20281 11689 20315
rect 54197 20301 54213 20335
rect 54247 20315 54373 20335
rect 54247 20301 54518 20315
rect 54339 20281 54518 20301
rect 11655 20115 11689 20281
rect 11655 20081 11781 20115
rect 11815 20081 11831 20115
rect 11655 19985 11781 20019
rect 11815 19985 11831 20019
rect 11655 19819 11689 19985
rect 11510 19785 11689 19819
rect 54339 19799 54518 19819
rect 54197 19765 54213 19799
rect 54247 19785 54518 19799
rect 54247 19765 54373 19785
rect 11510 19491 11689 19525
rect 54197 19511 54213 19545
rect 54247 19525 54373 19545
rect 54247 19511 54518 19525
rect 54339 19491 54518 19511
rect 11655 19325 11689 19491
rect 11655 19291 11781 19325
rect 11815 19291 11831 19325
rect 11655 19195 11781 19229
rect 11815 19195 11831 19229
rect 11655 19029 11689 19195
rect 11510 18995 11689 19029
rect 54339 19009 54518 19029
rect 54197 18975 54213 19009
rect 54247 18995 54518 19009
rect 54247 18975 54373 18995
rect 11510 18701 11689 18735
rect 54197 18721 54213 18755
rect 54247 18735 54373 18755
rect 54247 18721 54518 18735
rect 54339 18701 54518 18721
rect 11655 18535 11689 18701
rect 11655 18501 11781 18535
rect 11815 18501 11831 18535
rect 11655 18405 11781 18439
rect 11815 18405 11831 18439
rect 11655 18239 11689 18405
rect 11510 18205 11689 18239
rect 54339 18219 54518 18239
rect 54197 18185 54213 18219
rect 54247 18205 54518 18219
rect 54247 18185 54373 18205
rect 11510 17911 11689 17945
rect 54197 17931 54213 17965
rect 54247 17945 54373 17965
rect 54247 17931 54518 17945
rect 54339 17911 54518 17931
rect 11655 17745 11689 17911
rect 11655 17711 11781 17745
rect 11815 17711 11831 17745
rect 11655 17615 11781 17649
rect 11815 17615 11831 17649
rect 11655 17449 11689 17615
rect 11510 17415 11689 17449
rect 54339 17429 54518 17449
rect 54197 17395 54213 17429
rect 54247 17415 54518 17429
rect 54247 17395 54373 17415
rect 11510 17121 11689 17155
rect 54197 17141 54213 17175
rect 54247 17155 54373 17175
rect 54247 17141 54518 17155
rect 54339 17121 54518 17141
rect 11655 16955 11689 17121
rect 11655 16921 11781 16955
rect 11815 16921 11831 16955
rect 11655 16825 11781 16859
rect 11815 16825 11831 16859
rect 11655 16659 11689 16825
rect 11510 16625 11689 16659
rect 54339 16639 54518 16659
rect 54197 16605 54213 16639
rect 54247 16625 54518 16639
rect 54247 16605 54373 16625
rect 11510 16331 11689 16365
rect 54197 16351 54213 16385
rect 54247 16365 54373 16385
rect 54247 16351 54518 16365
rect 54339 16331 54518 16351
rect 11655 16165 11689 16331
rect 11655 16131 11781 16165
rect 11815 16131 11831 16165
rect 11655 16035 11781 16069
rect 11815 16035 11831 16069
rect 11655 15869 11689 16035
rect 11510 15835 11689 15869
rect 54339 15849 54518 15869
rect 54197 15815 54213 15849
rect 54247 15835 54518 15849
rect 54247 15815 54373 15835
rect 11510 15541 11689 15575
rect 54197 15561 54213 15595
rect 54247 15575 54373 15595
rect 54247 15561 54518 15575
rect 54339 15541 54518 15561
rect 11655 15375 11689 15541
rect 11655 15341 11781 15375
rect 11815 15341 11831 15375
rect 11655 15245 11781 15279
rect 11815 15245 11831 15279
rect 11655 15079 11689 15245
rect 11510 15045 11689 15079
rect 54339 15059 54518 15079
rect 54197 15025 54213 15059
rect 54247 15045 54518 15059
rect 54247 15025 54373 15045
rect 11510 14751 11689 14785
rect 54197 14771 54213 14805
rect 54247 14785 54373 14805
rect 54247 14771 54518 14785
rect 54339 14751 54518 14771
rect 11655 14585 11689 14751
rect 11655 14551 11781 14585
rect 11815 14551 11831 14585
rect 11655 14455 11781 14489
rect 11815 14455 11831 14489
rect 11655 14289 11689 14455
rect 11510 14255 11689 14289
rect 54339 14269 54518 14289
rect 54197 14235 54213 14269
rect 54247 14255 54518 14269
rect 54247 14235 54373 14255
rect 11510 13961 11689 13995
rect 54197 13981 54213 14015
rect 54247 13995 54373 14015
rect 54247 13981 54518 13995
rect 54339 13961 54518 13981
rect 11655 13795 11689 13961
rect 11655 13761 11781 13795
rect 11815 13761 11831 13795
rect 11655 13665 11781 13699
rect 11815 13665 11831 13699
rect 11655 13499 11689 13665
rect 11510 13465 11689 13499
rect 54339 13479 54518 13499
rect 54197 13445 54213 13479
rect 54247 13465 54518 13479
rect 54247 13445 54373 13465
rect 11510 13171 11689 13205
rect 54197 13191 54213 13225
rect 54247 13205 54373 13225
rect 54247 13191 54518 13205
rect 54339 13171 54518 13191
rect 11655 13005 11689 13171
rect 11655 12971 11781 13005
rect 11815 12971 11831 13005
rect 11655 12875 11781 12909
rect 11815 12875 11831 12909
rect 11655 12709 11689 12875
rect 11510 12675 11689 12709
rect 54339 12689 54518 12709
rect 54197 12655 54213 12689
rect 54247 12675 54518 12689
rect 54247 12655 54373 12675
rect 11510 12381 11689 12415
rect 54197 12401 54213 12435
rect 54247 12415 54373 12435
rect 54247 12401 54518 12415
rect 54339 12381 54518 12401
rect 11655 12215 11689 12381
rect 11655 12181 11781 12215
rect 11815 12181 11831 12215
rect 11655 12085 11781 12119
rect 11815 12085 11831 12119
rect 11655 11919 11689 12085
rect 11510 11885 11689 11919
rect 54339 11899 54518 11919
rect 54197 11865 54213 11899
rect 54247 11885 54518 11899
rect 54247 11865 54373 11885
rect 11510 11591 11689 11625
rect 54197 11611 54213 11645
rect 54247 11625 54373 11645
rect 54247 11611 54518 11625
rect 54339 11591 54518 11611
rect 11655 11425 11689 11591
rect 11655 11391 11781 11425
rect 11815 11391 11831 11425
rect 11655 11295 11781 11329
rect 11815 11295 11831 11329
rect 11655 11129 11689 11295
rect 11510 11095 11689 11129
rect 54339 11109 54518 11129
rect 54197 11075 54213 11109
rect 54247 11095 54518 11109
rect 54247 11075 54373 11095
rect 11510 10801 11689 10835
rect 54197 10821 54213 10855
rect 54247 10835 54373 10855
rect 54247 10821 54518 10835
rect 54339 10801 54518 10821
rect 11655 10635 11689 10801
rect 11655 10601 11781 10635
rect 11815 10601 11831 10635
rect 11655 10505 11781 10539
rect 11815 10505 11831 10539
rect 11655 10339 11689 10505
rect 11510 10305 11689 10339
rect 54339 10319 54518 10339
rect 54197 10285 54213 10319
rect 54247 10305 54518 10319
rect 54247 10285 54373 10305
rect 6471 7634 6505 7650
rect 6471 7584 6505 7600
rect 6471 6220 6505 6236
rect 6471 6170 6505 6186
rect 6000 5441 6034 5475
rect 6471 4806 6505 4822
rect 6471 4756 6505 4772
<< viali >>
rect 59399 66104 59433 66138
rect 59399 64690 59433 64724
rect 59399 63276 59433 63310
rect 54213 60591 54247 60625
rect 11781 60371 11815 60405
rect 11781 60275 11815 60309
rect 54213 60055 54247 60089
rect 54213 59801 54247 59835
rect 11781 59581 11815 59615
rect 11781 59485 11815 59519
rect 54213 59265 54247 59299
rect 54213 59011 54247 59045
rect 11781 58791 11815 58825
rect 11781 58695 11815 58729
rect 54213 58475 54247 58509
rect 54213 58221 54247 58255
rect 11781 58001 11815 58035
rect 11781 57905 11815 57939
rect 54213 57685 54247 57719
rect 54213 57431 54247 57465
rect 11781 57211 11815 57245
rect 11781 57115 11815 57149
rect 54213 56895 54247 56929
rect 54213 56641 54247 56675
rect 11781 56421 11815 56455
rect 11781 56325 11815 56359
rect 54213 56105 54247 56139
rect 54213 55851 54247 55885
rect 11781 55631 11815 55665
rect 11781 55535 11815 55569
rect 54213 55315 54247 55349
rect 54213 55061 54247 55095
rect 11781 54841 11815 54875
rect 11781 54745 11815 54779
rect 54213 54525 54247 54559
rect 54213 54271 54247 54305
rect 11781 54051 11815 54085
rect 11781 53955 11815 53989
rect 54213 53735 54247 53769
rect 54213 53481 54247 53515
rect 11781 53261 11815 53295
rect 11781 53165 11815 53199
rect 54213 52945 54247 52979
rect 54213 52691 54247 52725
rect 11781 52471 11815 52505
rect 11781 52375 11815 52409
rect 54213 52155 54247 52189
rect 54213 51901 54247 51935
rect 11781 51681 11815 51715
rect 11781 51585 11815 51619
rect 54213 51365 54247 51399
rect 54213 51111 54247 51145
rect 11781 50891 11815 50925
rect 11781 50795 11815 50829
rect 54213 50575 54247 50609
rect 54213 50321 54247 50355
rect 11781 50101 11815 50135
rect 11781 50005 11815 50039
rect 54213 49785 54247 49819
rect 54213 49531 54247 49565
rect 11781 49311 11815 49345
rect 11781 49215 11815 49249
rect 54213 48995 54247 49029
rect 54213 48741 54247 48775
rect 11781 48521 11815 48555
rect 11781 48425 11815 48459
rect 54213 48205 54247 48239
rect 54213 47951 54247 47985
rect 11781 47731 11815 47765
rect 11781 47635 11815 47669
rect 54213 47415 54247 47449
rect 54213 47161 54247 47195
rect 11781 46941 11815 46975
rect 11781 46845 11815 46879
rect 54213 46625 54247 46659
rect 54213 46371 54247 46405
rect 11781 46151 11815 46185
rect 11781 46055 11815 46089
rect 54213 45835 54247 45869
rect 54213 45581 54247 45615
rect 11781 45361 11815 45395
rect 11781 45265 11815 45299
rect 54213 45045 54247 45079
rect 54213 44791 54247 44825
rect 11781 44571 11815 44605
rect 11781 44475 11815 44509
rect 54213 44255 54247 44289
rect 54213 44001 54247 44035
rect 11781 43781 11815 43815
rect 11781 43685 11815 43719
rect 54213 43465 54247 43499
rect 54213 43211 54247 43245
rect 11781 42991 11815 43025
rect 11781 42895 11815 42929
rect 54213 42675 54247 42709
rect 54213 42421 54247 42455
rect 11781 42201 11815 42235
rect 11781 42105 11815 42139
rect 54213 41885 54247 41919
rect 54213 41631 54247 41665
rect 11781 41411 11815 41445
rect 11781 41315 11815 41349
rect 54213 41095 54247 41129
rect 54213 40841 54247 40875
rect 11781 40621 11815 40655
rect 11781 40525 11815 40559
rect 54213 40305 54247 40339
rect 54213 40051 54247 40085
rect 11781 39831 11815 39865
rect 11781 39735 11815 39769
rect 54213 39515 54247 39549
rect 54213 39261 54247 39295
rect 11781 39041 11815 39075
rect 11781 38945 11815 38979
rect 54213 38725 54247 38759
rect 54213 38471 54247 38505
rect 11781 38251 11815 38285
rect 11781 38155 11815 38189
rect 54213 37935 54247 37969
rect 54213 37681 54247 37715
rect 11781 37461 11815 37495
rect 11781 37365 11815 37399
rect 54213 37145 54247 37179
rect 54213 36891 54247 36925
rect 11781 36671 11815 36705
rect 11781 36575 11815 36609
rect 54213 36355 54247 36389
rect 54213 36101 54247 36135
rect 11781 35881 11815 35915
rect 11781 35785 11815 35819
rect 54213 35565 54247 35599
rect 54213 35311 54247 35345
rect 11781 35091 11815 35125
rect 11781 34995 11815 35029
rect 54213 34775 54247 34809
rect 54213 34521 54247 34555
rect 11781 34301 11815 34335
rect 11781 34205 11815 34239
rect 54213 33985 54247 34019
rect 54213 33731 54247 33765
rect 11781 33511 11815 33545
rect 11781 33415 11815 33449
rect 54213 33195 54247 33229
rect 54213 32941 54247 32975
rect 11781 32721 11815 32755
rect 11781 32625 11815 32659
rect 54213 32405 54247 32439
rect 54213 32151 54247 32185
rect 11781 31931 11815 31965
rect 11781 31835 11815 31869
rect 54213 31615 54247 31649
rect 54213 31361 54247 31395
rect 11781 31141 11815 31175
rect 11781 31045 11815 31079
rect 54213 30825 54247 30859
rect 54213 30571 54247 30605
rect 11781 30351 11815 30385
rect 11781 30255 11815 30289
rect 54213 30035 54247 30069
rect 54213 29781 54247 29815
rect 11781 29561 11815 29595
rect 11781 29465 11815 29499
rect 54213 29245 54247 29279
rect 54213 28991 54247 29025
rect 11781 28771 11815 28805
rect 11781 28675 11815 28709
rect 54213 28455 54247 28489
rect 54213 28201 54247 28235
rect 11781 27981 11815 28015
rect 11781 27885 11815 27919
rect 54213 27665 54247 27699
rect 54213 27411 54247 27445
rect 11781 27191 11815 27225
rect 11781 27095 11815 27129
rect 54213 26875 54247 26909
rect 54213 26621 54247 26655
rect 11781 26401 11815 26435
rect 11781 26305 11815 26339
rect 54213 26085 54247 26119
rect 54213 25831 54247 25865
rect 11781 25611 11815 25645
rect 11781 25515 11815 25549
rect 54213 25295 54247 25329
rect 54213 25041 54247 25075
rect 11781 24821 11815 24855
rect 11781 24725 11815 24759
rect 54213 24505 54247 24539
rect 54213 24251 54247 24285
rect 11781 24031 11815 24065
rect 11781 23935 11815 23969
rect 54213 23715 54247 23749
rect 54213 23461 54247 23495
rect 11781 23241 11815 23275
rect 11781 23145 11815 23179
rect 54213 22925 54247 22959
rect 54213 22671 54247 22705
rect 11781 22451 11815 22485
rect 11781 22355 11815 22389
rect 54213 22135 54247 22169
rect 54213 21881 54247 21915
rect 11781 21661 11815 21695
rect 11781 21565 11815 21599
rect 54213 21345 54247 21379
rect 54213 21091 54247 21125
rect 11781 20871 11815 20905
rect 11781 20775 11815 20809
rect 54213 20555 54247 20589
rect 54213 20301 54247 20335
rect 11781 20081 11815 20115
rect 11781 19985 11815 20019
rect 54213 19765 54247 19799
rect 54213 19511 54247 19545
rect 11781 19291 11815 19325
rect 11781 19195 11815 19229
rect 54213 18975 54247 19009
rect 54213 18721 54247 18755
rect 11781 18501 11815 18535
rect 11781 18405 11815 18439
rect 54213 18185 54247 18219
rect 54213 17931 54247 17965
rect 11781 17711 11815 17745
rect 11781 17615 11815 17649
rect 54213 17395 54247 17429
rect 54213 17141 54247 17175
rect 11781 16921 11815 16955
rect 11781 16825 11815 16859
rect 54213 16605 54247 16639
rect 54213 16351 54247 16385
rect 11781 16131 11815 16165
rect 11781 16035 11815 16069
rect 54213 15815 54247 15849
rect 54213 15561 54247 15595
rect 11781 15341 11815 15375
rect 11781 15245 11815 15279
rect 54213 15025 54247 15059
rect 54213 14771 54247 14805
rect 11781 14551 11815 14585
rect 11781 14455 11815 14489
rect 54213 14235 54247 14269
rect 54213 13981 54247 14015
rect 11781 13761 11815 13795
rect 11781 13665 11815 13699
rect 54213 13445 54247 13479
rect 54213 13191 54247 13225
rect 11781 12971 11815 13005
rect 11781 12875 11815 12909
rect 54213 12655 54247 12689
rect 54213 12401 54247 12435
rect 11781 12181 11815 12215
rect 11781 12085 11815 12119
rect 54213 11865 54247 11899
rect 54213 11611 54247 11645
rect 11781 11391 11815 11425
rect 11781 11295 11815 11329
rect 54213 11075 54247 11109
rect 54213 10821 54247 10855
rect 11781 10601 11815 10635
rect 11781 10505 11815 10539
rect 54213 10285 54247 10319
rect 6471 7600 6505 7634
rect 6471 6186 6505 6220
rect 6471 4772 6505 4806
<< metal1 >>
rect 13150 67021 13196 67275
rect 14398 67021 14444 67275
rect 15646 67021 15692 67275
rect 16894 67021 16940 67275
rect 18142 67021 18188 67275
rect 19390 67021 19436 67275
rect 20638 67021 20684 67275
rect 21886 67021 21932 67275
rect 23134 67021 23180 67275
rect 24382 67021 24428 67275
rect 25630 67021 25676 67275
rect 26878 67021 26924 67275
rect 28126 67021 28172 67275
rect 29374 67021 29420 67275
rect 30622 67021 30668 67275
rect 31870 67021 31916 67275
rect 33118 67021 33164 67275
rect 34366 67021 34412 67275
rect 35614 67021 35660 67275
rect 36862 67021 36908 67275
rect 38110 67021 38156 67275
rect 39358 67021 39404 67275
rect 40606 67021 40652 67275
rect 41854 67021 41900 67275
rect 43102 67021 43148 67275
rect 44350 67021 44396 67275
rect 45598 67021 45644 67275
rect 46846 67021 46892 67275
rect 48094 67021 48140 67275
rect 49342 67021 49388 67275
rect 50590 67021 50636 67275
rect 51838 67021 51884 67275
rect 59384 66095 59390 66147
rect 59442 66095 59448 66147
rect 59384 64681 59390 64733
rect 59442 64681 59448 64733
rect 59384 63267 59390 63319
rect 59442 63267 59448 63319
rect 53030 62629 53036 62681
rect 53088 62629 53094 62681
rect 53048 62531 53076 62629
rect 13112 61665 13140 61777
rect 13576 61665 13604 61777
rect 13112 61637 13372 61665
rect 13344 61525 13372 61637
rect 13416 61637 13604 61665
rect 13736 61665 13764 61777
rect 14200 61665 14228 61777
rect 13736 61637 13924 61665
rect 13416 61525 13444 61637
rect 13896 61525 13924 61637
rect 13968 61637 14228 61665
rect 14360 61665 14388 61777
rect 14824 61665 14852 61777
rect 14360 61637 14620 61665
rect 13968 61525 13996 61637
rect 14592 61525 14620 61637
rect 14664 61637 14852 61665
rect 14984 61665 15012 61777
rect 15448 61665 15476 61777
rect 14984 61637 15172 61665
rect 14664 61525 14692 61637
rect 15144 61525 15172 61637
rect 15216 61637 15476 61665
rect 15608 61665 15636 61777
rect 16072 61665 16100 61777
rect 15608 61637 15868 61665
rect 15216 61525 15244 61637
rect 15840 61525 15868 61637
rect 15912 61637 16100 61665
rect 16232 61665 16260 61777
rect 16696 61665 16724 61777
rect 16232 61637 16420 61665
rect 15912 61525 15940 61637
rect 16392 61525 16420 61637
rect 16464 61637 16724 61665
rect 16856 61665 16884 61777
rect 17320 61665 17348 61777
rect 16856 61637 17116 61665
rect 16464 61525 16492 61637
rect 17088 61525 17116 61637
rect 17160 61637 17348 61665
rect 17480 61665 17508 61777
rect 17944 61665 17972 61777
rect 17480 61637 17668 61665
rect 17160 61525 17188 61637
rect 17640 61525 17668 61637
rect 17712 61637 17972 61665
rect 18104 61665 18132 61777
rect 18568 61665 18596 61777
rect 18104 61637 18364 61665
rect 17712 61525 17740 61637
rect 18336 61525 18364 61637
rect 18408 61637 18596 61665
rect 18728 61665 18756 61777
rect 19192 61665 19220 61777
rect 18728 61637 18916 61665
rect 18408 61525 18436 61637
rect 18888 61525 18916 61637
rect 18960 61637 19220 61665
rect 19352 61665 19380 61777
rect 19816 61665 19844 61777
rect 19352 61637 19612 61665
rect 18960 61525 18988 61637
rect 19584 61525 19612 61637
rect 19656 61637 19844 61665
rect 19976 61665 20004 61777
rect 20440 61665 20468 61777
rect 19976 61637 20164 61665
rect 19656 61525 19684 61637
rect 20136 61525 20164 61637
rect 20208 61637 20468 61665
rect 20600 61665 20628 61777
rect 21064 61665 21092 61777
rect 20600 61637 20860 61665
rect 20208 61525 20236 61637
rect 20832 61525 20860 61637
rect 20904 61637 21092 61665
rect 21224 61665 21252 61777
rect 21688 61665 21716 61777
rect 21224 61637 21412 61665
rect 20904 61525 20932 61637
rect 21384 61525 21412 61637
rect 21456 61637 21716 61665
rect 21848 61665 21876 61777
rect 22312 61665 22340 61777
rect 21848 61637 22108 61665
rect 21456 61525 21484 61637
rect 22080 61525 22108 61637
rect 22152 61637 22340 61665
rect 22472 61665 22500 61777
rect 22936 61665 22964 61777
rect 22472 61637 22660 61665
rect 22152 61525 22180 61637
rect 22632 61525 22660 61637
rect 22704 61637 22964 61665
rect 23096 61665 23124 61777
rect 23560 61665 23588 61777
rect 23096 61637 23356 61665
rect 22704 61525 22732 61637
rect 23328 61525 23356 61637
rect 23400 61637 23588 61665
rect 23720 61665 23748 61777
rect 24184 61665 24212 61777
rect 23720 61637 23908 61665
rect 23400 61525 23428 61637
rect 23880 61525 23908 61637
rect 23952 61637 24212 61665
rect 24344 61665 24372 61777
rect 24808 61665 24836 61777
rect 24344 61637 24604 61665
rect 23952 61525 23980 61637
rect 24576 61525 24604 61637
rect 24648 61637 24836 61665
rect 24968 61665 24996 61777
rect 25432 61665 25460 61777
rect 24968 61637 25156 61665
rect 24648 61525 24676 61637
rect 25128 61525 25156 61637
rect 25200 61637 25460 61665
rect 25592 61665 25620 61777
rect 26056 61665 26084 61777
rect 25592 61637 25852 61665
rect 25200 61525 25228 61637
rect 25824 61525 25852 61637
rect 25896 61637 26084 61665
rect 26216 61665 26244 61777
rect 26680 61665 26708 61777
rect 26216 61637 26404 61665
rect 25896 61525 25924 61637
rect 26376 61525 26404 61637
rect 26448 61637 26708 61665
rect 26840 61665 26868 61777
rect 27304 61665 27332 61777
rect 26840 61637 27100 61665
rect 26448 61525 26476 61637
rect 27072 61525 27100 61637
rect 27144 61637 27332 61665
rect 27464 61665 27492 61777
rect 27928 61665 27956 61777
rect 27464 61637 27652 61665
rect 27144 61525 27172 61637
rect 27624 61525 27652 61637
rect 27696 61637 27956 61665
rect 28088 61665 28116 61777
rect 28552 61665 28580 61777
rect 28088 61637 28348 61665
rect 27696 61525 27724 61637
rect 28320 61525 28348 61637
rect 28392 61637 28580 61665
rect 28712 61665 28740 61777
rect 29176 61665 29204 61777
rect 28712 61637 28900 61665
rect 28392 61525 28420 61637
rect 28872 61525 28900 61637
rect 28944 61637 29204 61665
rect 29336 61665 29364 61777
rect 29800 61665 29828 61777
rect 29336 61637 29596 61665
rect 28944 61525 28972 61637
rect 29568 61525 29596 61637
rect 29640 61637 29828 61665
rect 29960 61665 29988 61777
rect 30424 61665 30452 61777
rect 29960 61637 30148 61665
rect 29640 61525 29668 61637
rect 30120 61525 30148 61637
rect 30192 61637 30452 61665
rect 30584 61665 30612 61777
rect 31048 61665 31076 61777
rect 30584 61637 30844 61665
rect 30192 61525 30220 61637
rect 30816 61525 30844 61637
rect 30888 61637 31076 61665
rect 31208 61665 31236 61777
rect 31672 61665 31700 61777
rect 31208 61637 31396 61665
rect 30888 61525 30916 61637
rect 31368 61525 31396 61637
rect 31440 61637 31700 61665
rect 31832 61665 31860 61777
rect 32296 61665 32324 61777
rect 31832 61637 32092 61665
rect 31440 61525 31468 61637
rect 32064 61525 32092 61637
rect 32136 61637 32324 61665
rect 32456 61665 32484 61777
rect 32920 61665 32948 61777
rect 32456 61637 32644 61665
rect 32136 61525 32164 61637
rect 32616 61525 32644 61637
rect 32688 61637 32948 61665
rect 33080 61665 33108 61777
rect 33544 61665 33572 61777
rect 33080 61637 33340 61665
rect 32688 61525 32716 61637
rect 33312 61525 33340 61637
rect 33384 61637 33572 61665
rect 33704 61665 33732 61777
rect 34168 61665 34196 61777
rect 33704 61637 33892 61665
rect 33384 61525 33412 61637
rect 33864 61525 33892 61637
rect 33936 61637 34196 61665
rect 34328 61665 34356 61777
rect 34792 61665 34820 61777
rect 34328 61637 34588 61665
rect 33936 61525 33964 61637
rect 34560 61525 34588 61637
rect 34632 61637 34820 61665
rect 34952 61665 34980 61777
rect 35416 61665 35444 61777
rect 34952 61637 35140 61665
rect 34632 61525 34660 61637
rect 35112 61525 35140 61637
rect 35184 61637 35444 61665
rect 35576 61665 35604 61777
rect 36040 61665 36068 61777
rect 35576 61637 35836 61665
rect 35184 61525 35212 61637
rect 35808 61525 35836 61637
rect 35880 61637 36068 61665
rect 36200 61665 36228 61777
rect 36664 61665 36692 61777
rect 36200 61637 36388 61665
rect 35880 61525 35908 61637
rect 36360 61525 36388 61637
rect 36432 61637 36692 61665
rect 36824 61665 36852 61777
rect 37288 61665 37316 61777
rect 36824 61637 37084 61665
rect 36432 61525 36460 61637
rect 37056 61525 37084 61637
rect 37128 61637 37316 61665
rect 37448 61665 37476 61777
rect 37912 61665 37940 61777
rect 37448 61637 37636 61665
rect 37128 61525 37156 61637
rect 37608 61525 37636 61637
rect 37680 61637 37940 61665
rect 38072 61665 38100 61777
rect 38536 61665 38564 61777
rect 38072 61637 38332 61665
rect 37680 61525 37708 61637
rect 38304 61525 38332 61637
rect 38376 61637 38564 61665
rect 38696 61665 38724 61777
rect 39160 61665 39188 61777
rect 38696 61637 38884 61665
rect 38376 61525 38404 61637
rect 38856 61525 38884 61637
rect 38928 61637 39188 61665
rect 39320 61665 39348 61777
rect 39784 61665 39812 61777
rect 39320 61637 39580 61665
rect 38928 61525 38956 61637
rect 39552 61525 39580 61637
rect 39624 61637 39812 61665
rect 39944 61665 39972 61777
rect 40408 61665 40436 61777
rect 39944 61637 40132 61665
rect 39624 61525 39652 61637
rect 40104 61525 40132 61637
rect 40176 61637 40436 61665
rect 40568 61665 40596 61777
rect 41032 61665 41060 61777
rect 40568 61637 40828 61665
rect 40176 61525 40204 61637
rect 40800 61525 40828 61637
rect 40872 61637 41060 61665
rect 41192 61665 41220 61777
rect 41656 61665 41684 61777
rect 41192 61637 41380 61665
rect 40872 61525 40900 61637
rect 41352 61525 41380 61637
rect 41424 61637 41684 61665
rect 41816 61665 41844 61777
rect 42280 61665 42308 61777
rect 41816 61637 42076 61665
rect 41424 61525 41452 61637
rect 42048 61525 42076 61637
rect 42120 61637 42308 61665
rect 42440 61665 42468 61777
rect 42904 61665 42932 61777
rect 42440 61637 42628 61665
rect 42120 61525 42148 61637
rect 42600 61525 42628 61637
rect 42672 61637 42932 61665
rect 43064 61665 43092 61777
rect 43528 61665 43556 61777
rect 43064 61637 43324 61665
rect 42672 61525 42700 61637
rect 43296 61525 43324 61637
rect 43368 61637 43556 61665
rect 43688 61665 43716 61777
rect 44152 61665 44180 61777
rect 43688 61637 43876 61665
rect 43368 61525 43396 61637
rect 43848 61525 43876 61637
rect 43920 61637 44180 61665
rect 44312 61665 44340 61777
rect 44776 61665 44804 61777
rect 44312 61637 44572 61665
rect 43920 61525 43948 61637
rect 44544 61525 44572 61637
rect 44616 61637 44804 61665
rect 44936 61665 44964 61777
rect 45400 61665 45428 61777
rect 44936 61637 45124 61665
rect 44616 61525 44644 61637
rect 45096 61525 45124 61637
rect 45168 61637 45428 61665
rect 45560 61665 45588 61777
rect 46024 61665 46052 61777
rect 45560 61637 45820 61665
rect 45168 61525 45196 61637
rect 45792 61525 45820 61637
rect 45864 61637 46052 61665
rect 46184 61665 46212 61777
rect 46648 61665 46676 61777
rect 46184 61637 46372 61665
rect 45864 61525 45892 61637
rect 46344 61525 46372 61637
rect 46416 61637 46676 61665
rect 46808 61665 46836 61777
rect 47272 61665 47300 61777
rect 46808 61637 47068 61665
rect 46416 61525 46444 61637
rect 47040 61525 47068 61637
rect 47112 61637 47300 61665
rect 47432 61665 47460 61777
rect 47896 61665 47924 61777
rect 47432 61637 47620 61665
rect 47112 61525 47140 61637
rect 47592 61525 47620 61637
rect 47664 61637 47924 61665
rect 48056 61665 48084 61777
rect 48520 61665 48548 61777
rect 48056 61637 48316 61665
rect 47664 61525 47692 61637
rect 48288 61525 48316 61637
rect 48360 61637 48548 61665
rect 48680 61665 48708 61777
rect 49144 61665 49172 61777
rect 48680 61637 48868 61665
rect 48360 61525 48388 61637
rect 48840 61525 48868 61637
rect 48912 61637 49172 61665
rect 49304 61665 49332 61777
rect 49768 61665 49796 61777
rect 49304 61637 49564 61665
rect 48912 61525 48940 61637
rect 49536 61525 49564 61637
rect 49608 61637 49796 61665
rect 49928 61665 49956 61777
rect 50392 61665 50420 61777
rect 49928 61637 50116 61665
rect 49608 61525 49636 61637
rect 50088 61525 50116 61637
rect 50160 61637 50420 61665
rect 50552 61665 50580 61777
rect 51016 61665 51044 61777
rect 50552 61637 50812 61665
rect 50160 61525 50188 61637
rect 50784 61525 50812 61637
rect 50856 61637 51044 61665
rect 51176 61665 51204 61777
rect 51640 61665 51668 61777
rect 51176 61637 51364 61665
rect 50856 61525 50884 61637
rect 51336 61525 51364 61637
rect 51408 61637 51668 61665
rect 51800 61665 51828 61777
rect 52264 61665 52292 61777
rect 51800 61637 52060 61665
rect 51408 61525 51436 61637
rect 52032 61525 52060 61637
rect 52104 61637 52292 61665
rect 52424 61665 52452 61777
rect 52888 61665 52916 61777
rect 52424 61637 52612 61665
rect 52104 61525 52132 61637
rect 52584 61525 52612 61637
rect 52656 61637 52916 61665
rect 53048 61665 53076 61777
rect 53512 61665 53540 61777
rect 53048 61637 53308 61665
rect 52656 61525 52684 61637
rect 53280 61525 53308 61637
rect 53352 61637 53540 61665
rect 53352 61525 53380 61637
rect 54336 61213 54342 61265
rect 54394 61253 54400 61265
rect 58400 61253 58406 61265
rect 54394 61225 58406 61253
rect 54394 61213 54400 61225
rect 58400 61213 58406 61225
rect 58458 61213 58464 61265
rect 54198 60582 54204 60634
rect 54256 60582 54262 60634
rect 11766 60362 11772 60414
rect 11824 60362 11830 60414
rect 11766 60266 11772 60318
rect 11824 60266 11830 60318
rect 54198 60046 54204 60098
rect 54256 60046 54262 60098
rect 54198 59792 54204 59844
rect 54256 59792 54262 59844
rect 11766 59572 11772 59624
rect 11824 59572 11830 59624
rect 11766 59476 11772 59528
rect 11824 59476 11830 59528
rect 54198 59256 54204 59308
rect 54256 59256 54262 59308
rect 54198 59002 54204 59054
rect 54256 59002 54262 59054
rect 11766 58782 11772 58834
rect 11824 58782 11830 58834
rect 11766 58686 11772 58738
rect 11824 58686 11830 58738
rect 54198 58466 54204 58518
rect 54256 58466 54262 58518
rect 54198 58212 54204 58264
rect 54256 58212 54262 58264
rect 11766 57992 11772 58044
rect 11824 57992 11830 58044
rect 11766 57896 11772 57948
rect 11824 57896 11830 57948
rect 54198 57676 54204 57728
rect 54256 57676 54262 57728
rect 54198 57422 54204 57474
rect 54256 57422 54262 57474
rect 11766 57202 11772 57254
rect 11824 57202 11830 57254
rect 11766 57106 11772 57158
rect 11824 57106 11830 57158
rect 54198 56886 54204 56938
rect 54256 56886 54262 56938
rect 54198 56632 54204 56684
rect 54256 56632 54262 56684
rect 11766 56412 11772 56464
rect 11824 56412 11830 56464
rect 11766 56316 11772 56368
rect 11824 56316 11830 56368
rect 54198 56096 54204 56148
rect 54256 56096 54262 56148
rect 54198 55842 54204 55894
rect 54256 55842 54262 55894
rect 11766 55622 11772 55674
rect 11824 55622 11830 55674
rect 11766 55526 11772 55578
rect 11824 55526 11830 55578
rect 54198 55306 54204 55358
rect 54256 55306 54262 55358
rect 54198 55052 54204 55104
rect 54256 55052 54262 55104
rect 11766 54832 11772 54884
rect 11824 54832 11830 54884
rect 11766 54736 11772 54788
rect 11824 54736 11830 54788
rect 54198 54516 54204 54568
rect 54256 54516 54262 54568
rect 54198 54262 54204 54314
rect 54256 54262 54262 54314
rect 11766 54042 11772 54094
rect 11824 54042 11830 54094
rect 11766 53946 11772 53998
rect 11824 53946 11830 53998
rect 54198 53726 54204 53778
rect 54256 53726 54262 53778
rect 54198 53472 54204 53524
rect 54256 53472 54262 53524
rect 11766 53252 11772 53304
rect 11824 53252 11830 53304
rect 11766 53156 11772 53208
rect 11824 53156 11830 53208
rect 54198 52936 54204 52988
rect 54256 52936 54262 52988
rect 54198 52682 54204 52734
rect 54256 52682 54262 52734
rect 11766 52462 11772 52514
rect 11824 52462 11830 52514
rect 11766 52366 11772 52418
rect 11824 52366 11830 52418
rect 54198 52146 54204 52198
rect 54256 52146 54262 52198
rect 54198 51892 54204 51944
rect 54256 51892 54262 51944
rect 11766 51672 11772 51724
rect 11824 51672 11830 51724
rect 11766 51576 11772 51628
rect 11824 51576 11830 51628
rect 54198 51356 54204 51408
rect 54256 51356 54262 51408
rect 54198 51102 54204 51154
rect 54256 51102 54262 51154
rect 11766 50882 11772 50934
rect 11824 50882 11830 50934
rect 11766 50786 11772 50838
rect 11824 50786 11830 50838
rect 54198 50566 54204 50618
rect 54256 50566 54262 50618
rect 54198 50312 54204 50364
rect 54256 50312 54262 50364
rect 11766 50092 11772 50144
rect 11824 50092 11830 50144
rect 11766 49996 11772 50048
rect 11824 49996 11830 50048
rect 54198 49776 54204 49828
rect 54256 49776 54262 49828
rect 54198 49522 54204 49574
rect 54256 49522 54262 49574
rect 11766 49302 11772 49354
rect 11824 49302 11830 49354
rect 11766 49206 11772 49258
rect 11824 49206 11830 49258
rect 54198 48986 54204 49038
rect 54256 48986 54262 49038
rect 54198 48732 54204 48784
rect 54256 48732 54262 48784
rect 11766 48512 11772 48564
rect 11824 48512 11830 48564
rect 11766 48416 11772 48468
rect 11824 48416 11830 48468
rect 54198 48196 54204 48248
rect 54256 48196 54262 48248
rect 54198 47942 54204 47994
rect 54256 47942 54262 47994
rect 11766 47722 11772 47774
rect 11824 47722 11830 47774
rect 11766 47626 11772 47678
rect 11824 47626 11830 47678
rect 54198 47406 54204 47458
rect 54256 47406 54262 47458
rect 54198 47152 54204 47204
rect 54256 47152 54262 47204
rect 11766 46932 11772 46984
rect 11824 46932 11830 46984
rect 11766 46836 11772 46888
rect 11824 46836 11830 46888
rect 54198 46616 54204 46668
rect 54256 46616 54262 46668
rect 54198 46362 54204 46414
rect 54256 46362 54262 46414
rect 11766 46142 11772 46194
rect 11824 46142 11830 46194
rect 11766 46046 11772 46098
rect 11824 46046 11830 46098
rect 54198 45826 54204 45878
rect 54256 45826 54262 45878
rect 54198 45572 54204 45624
rect 54256 45572 54262 45624
rect 11766 45352 11772 45404
rect 11824 45352 11830 45404
rect 11766 45256 11772 45308
rect 11824 45256 11830 45308
rect 54198 45036 54204 45088
rect 54256 45036 54262 45088
rect 54198 44782 54204 44834
rect 54256 44782 54262 44834
rect 11766 44562 11772 44614
rect 11824 44562 11830 44614
rect 11766 44466 11772 44518
rect 11824 44466 11830 44518
rect 54198 44246 54204 44298
rect 54256 44246 54262 44298
rect 54198 43992 54204 44044
rect 54256 43992 54262 44044
rect 11766 43772 11772 43824
rect 11824 43772 11830 43824
rect 11766 43676 11772 43728
rect 11824 43676 11830 43728
rect 54198 43456 54204 43508
rect 54256 43456 54262 43508
rect 54198 43202 54204 43254
rect 54256 43202 54262 43254
rect 11766 42982 11772 43034
rect 11824 42982 11830 43034
rect 11766 42886 11772 42938
rect 11824 42886 11830 42938
rect 54198 42666 54204 42718
rect 54256 42666 54262 42718
rect 54198 42412 54204 42464
rect 54256 42412 54262 42464
rect 11766 42192 11772 42244
rect 11824 42192 11830 42244
rect 11766 42096 11772 42148
rect 11824 42096 11830 42148
rect 54198 41876 54204 41928
rect 54256 41876 54262 41928
rect 54198 41622 54204 41674
rect 54256 41622 54262 41674
rect 11766 41402 11772 41454
rect 11824 41402 11830 41454
rect 11766 41306 11772 41358
rect 11824 41306 11830 41358
rect 54198 41086 54204 41138
rect 54256 41086 54262 41138
rect 54198 40832 54204 40884
rect 54256 40832 54262 40884
rect 11766 40612 11772 40664
rect 11824 40612 11830 40664
rect 11766 40516 11772 40568
rect 11824 40516 11830 40568
rect 54198 40296 54204 40348
rect 54256 40296 54262 40348
rect 54198 40042 54204 40094
rect 54256 40042 54262 40094
rect 11766 39822 11772 39874
rect 11824 39822 11830 39874
rect 11766 39726 11772 39778
rect 11824 39726 11830 39778
rect 54198 39506 54204 39558
rect 54256 39506 54262 39558
rect 54198 39252 54204 39304
rect 54256 39252 54262 39304
rect 11766 39032 11772 39084
rect 11824 39032 11830 39084
rect 11766 38936 11772 38988
rect 11824 38936 11830 38988
rect 54198 38716 54204 38768
rect 54256 38716 54262 38768
rect 54198 38462 54204 38514
rect 54256 38462 54262 38514
rect 11766 38242 11772 38294
rect 11824 38242 11830 38294
rect 11766 38146 11772 38198
rect 11824 38146 11830 38198
rect 54198 37926 54204 37978
rect 54256 37926 54262 37978
rect 54198 37672 54204 37724
rect 54256 37672 54262 37724
rect 11766 37452 11772 37504
rect 11824 37452 11830 37504
rect 11766 37356 11772 37408
rect 11824 37356 11830 37408
rect 54198 37136 54204 37188
rect 54256 37136 54262 37188
rect 54198 36882 54204 36934
rect 54256 36882 54262 36934
rect 11766 36662 11772 36714
rect 11824 36662 11830 36714
rect 11766 36566 11772 36618
rect 11824 36566 11830 36618
rect 54198 36346 54204 36398
rect 54256 36346 54262 36398
rect 54198 36092 54204 36144
rect 54256 36092 54262 36144
rect 11766 35872 11772 35924
rect 11824 35872 11830 35924
rect 11766 35776 11772 35828
rect 11824 35776 11830 35828
rect 54198 35556 54204 35608
rect 54256 35556 54262 35608
rect 54198 35302 54204 35354
rect 54256 35302 54262 35354
rect 11766 35082 11772 35134
rect 11824 35082 11830 35134
rect 11766 34986 11772 35038
rect 11824 34986 11830 35038
rect 54198 34766 54204 34818
rect 54256 34766 54262 34818
rect 54198 34512 54204 34564
rect 54256 34512 54262 34564
rect 11766 34292 11772 34344
rect 11824 34292 11830 34344
rect 11766 34196 11772 34248
rect 11824 34196 11830 34248
rect 54198 33976 54204 34028
rect 54256 33976 54262 34028
rect 54198 33722 54204 33774
rect 54256 33722 54262 33774
rect 11766 33502 11772 33554
rect 11824 33502 11830 33554
rect 11766 33406 11772 33458
rect 11824 33406 11830 33458
rect 54198 33186 54204 33238
rect 54256 33186 54262 33238
rect 54198 32932 54204 32984
rect 54256 32932 54262 32984
rect 11766 32712 11772 32764
rect 11824 32712 11830 32764
rect 11766 32616 11772 32668
rect 11824 32616 11830 32668
rect 54198 32396 54204 32448
rect 54256 32396 54262 32448
rect 54198 32142 54204 32194
rect 54256 32142 54262 32194
rect 11766 31922 11772 31974
rect 11824 31922 11830 31974
rect 11766 31826 11772 31878
rect 11824 31826 11830 31878
rect 54198 31606 54204 31658
rect 54256 31606 54262 31658
rect 54198 31352 54204 31404
rect 54256 31352 54262 31404
rect 11766 31132 11772 31184
rect 11824 31132 11830 31184
rect 11766 31036 11772 31088
rect 11824 31036 11830 31088
rect 54198 30816 54204 30868
rect 54256 30816 54262 30868
rect 54198 30562 54204 30614
rect 54256 30562 54262 30614
rect 11766 30342 11772 30394
rect 11824 30342 11830 30394
rect 11766 30246 11772 30298
rect 11824 30246 11830 30298
rect 54198 30026 54204 30078
rect 54256 30026 54262 30078
rect 54198 29772 54204 29824
rect 54256 29772 54262 29824
rect 11766 29552 11772 29604
rect 11824 29552 11830 29604
rect 11766 29456 11772 29508
rect 11824 29456 11830 29508
rect 54198 29236 54204 29288
rect 54256 29236 54262 29288
rect 54198 28982 54204 29034
rect 54256 28982 54262 29034
rect 11766 28762 11772 28814
rect 11824 28762 11830 28814
rect 11766 28666 11772 28718
rect 11824 28666 11830 28718
rect 54198 28446 54204 28498
rect 54256 28446 54262 28498
rect 54198 28192 54204 28244
rect 54256 28192 54262 28244
rect 11766 27972 11772 28024
rect 11824 27972 11830 28024
rect 11766 27876 11772 27928
rect 11824 27876 11830 27928
rect 54198 27656 54204 27708
rect 54256 27656 54262 27708
rect 54198 27402 54204 27454
rect 54256 27402 54262 27454
rect 11766 27182 11772 27234
rect 11824 27182 11830 27234
rect 11766 27086 11772 27138
rect 11824 27086 11830 27138
rect 54198 26866 54204 26918
rect 54256 26866 54262 26918
rect 54198 26612 54204 26664
rect 54256 26612 54262 26664
rect 11766 26392 11772 26444
rect 11824 26392 11830 26444
rect 11766 26296 11772 26348
rect 11824 26296 11830 26348
rect 54198 26076 54204 26128
rect 54256 26076 54262 26128
rect 54198 25822 54204 25874
rect 54256 25822 54262 25874
rect 11766 25602 11772 25654
rect 11824 25602 11830 25654
rect 11766 25506 11772 25558
rect 11824 25506 11830 25558
rect 54198 25286 54204 25338
rect 54256 25286 54262 25338
rect 54198 25032 54204 25084
rect 54256 25032 54262 25084
rect 11766 24812 11772 24864
rect 11824 24812 11830 24864
rect 11766 24716 11772 24768
rect 11824 24716 11830 24768
rect 54198 24496 54204 24548
rect 54256 24496 54262 24548
rect 54198 24242 54204 24294
rect 54256 24242 54262 24294
rect 11766 24022 11772 24074
rect 11824 24022 11830 24074
rect 11766 23926 11772 23978
rect 11824 23926 11830 23978
rect 54198 23706 54204 23758
rect 54256 23706 54262 23758
rect 54198 23452 54204 23504
rect 54256 23452 54262 23504
rect 11766 23232 11772 23284
rect 11824 23232 11830 23284
rect 11766 23136 11772 23188
rect 11824 23136 11830 23188
rect 54198 22916 54204 22968
rect 54256 22916 54262 22968
rect 54198 22662 54204 22714
rect 54256 22662 54262 22714
rect 11766 22442 11772 22494
rect 11824 22442 11830 22494
rect 11766 22346 11772 22398
rect 11824 22346 11830 22398
rect 54198 22126 54204 22178
rect 54256 22126 54262 22178
rect 54198 21872 54204 21924
rect 54256 21872 54262 21924
rect 11766 21652 11772 21704
rect 11824 21652 11830 21704
rect 11766 21556 11772 21608
rect 11824 21556 11830 21608
rect 54198 21336 54204 21388
rect 54256 21336 54262 21388
rect 54198 21082 54204 21134
rect 54256 21082 54262 21134
rect 11766 20862 11772 20914
rect 11824 20862 11830 20914
rect 11766 20766 11772 20818
rect 11824 20766 11830 20818
rect 54198 20546 54204 20598
rect 54256 20546 54262 20598
rect 54198 20292 54204 20344
rect 54256 20292 54262 20344
rect 11766 20072 11772 20124
rect 11824 20072 11830 20124
rect 11766 19976 11772 20028
rect 11824 19976 11830 20028
rect 54198 19756 54204 19808
rect 54256 19756 54262 19808
rect 54198 19502 54204 19554
rect 54256 19502 54262 19554
rect 11766 19282 11772 19334
rect 11824 19282 11830 19334
rect 11766 19186 11772 19238
rect 11824 19186 11830 19238
rect 54198 18966 54204 19018
rect 54256 18966 54262 19018
rect 54198 18712 54204 18764
rect 54256 18712 54262 18764
rect 11766 18492 11772 18544
rect 11824 18492 11830 18544
rect 11766 18396 11772 18448
rect 11824 18396 11830 18448
rect 54198 18176 54204 18228
rect 54256 18176 54262 18228
rect 18 10204 46 18104
rect 98 10204 126 18104
rect 178 10204 206 18104
rect 258 10204 286 18104
rect 338 10204 366 18104
rect 418 10204 446 18104
rect 498 10204 526 18104
rect 54198 17922 54204 17974
rect 54256 17922 54262 17974
rect 11766 17702 11772 17754
rect 11824 17702 11830 17754
rect 11766 17606 11772 17658
rect 11824 17606 11830 17658
rect 54198 17386 54204 17438
rect 54256 17386 54262 17438
rect 54198 17132 54204 17184
rect 54256 17132 54262 17184
rect 11766 16912 11772 16964
rect 11824 16912 11830 16964
rect 11766 16816 11772 16868
rect 11824 16816 11830 16868
rect 54198 16596 54204 16648
rect 54256 16596 54262 16648
rect 54198 16342 54204 16394
rect 54256 16342 54262 16394
rect 11766 16122 11772 16174
rect 11824 16122 11830 16174
rect 11766 16026 11772 16078
rect 11824 16026 11830 16078
rect 54198 15806 54204 15858
rect 54256 15806 54262 15858
rect 54198 15552 54204 15604
rect 54256 15552 54262 15604
rect 11766 15332 11772 15384
rect 11824 15332 11830 15384
rect 11766 15236 11772 15288
rect 11824 15236 11830 15288
rect 54198 15016 54204 15068
rect 54256 15016 54262 15068
rect 54198 14762 54204 14814
rect 54256 14762 54262 14814
rect 11766 14542 11772 14594
rect 11824 14542 11830 14594
rect 11766 14446 11772 14498
rect 11824 14446 11830 14498
rect 54198 14226 54204 14278
rect 54256 14226 54262 14278
rect 54198 13972 54204 14024
rect 54256 13972 54262 14024
rect 11766 13752 11772 13804
rect 11824 13752 11830 13804
rect 11766 13656 11772 13708
rect 11824 13656 11830 13708
rect 54198 13436 54204 13488
rect 54256 13436 54262 13488
rect 54198 13182 54204 13234
rect 54256 13182 54262 13234
rect 11766 12962 11772 13014
rect 11824 12962 11830 13014
rect 11766 12866 11772 12918
rect 11824 12866 11830 12918
rect 54198 12646 54204 12698
rect 54256 12646 54262 12698
rect 54198 12392 54204 12444
rect 54256 12392 54262 12444
rect 11766 12172 11772 12224
rect 11824 12172 11830 12224
rect 11766 12076 11772 12128
rect 11824 12076 11830 12128
rect 54198 11856 54204 11908
rect 54256 11856 54262 11908
rect 54198 11602 54204 11654
rect 54256 11602 54262 11654
rect 11766 11382 11772 11434
rect 11824 11382 11830 11434
rect 11766 11286 11772 11338
rect 11824 11286 11830 11338
rect 54198 11066 54204 11118
rect 54256 11066 54262 11118
rect 54198 10812 54204 10864
rect 54256 10812 54262 10864
rect 11766 10592 11772 10644
rect 11824 10592 11830 10644
rect 11766 10496 11772 10548
rect 11824 10496 11830 10548
rect 54198 10276 54204 10328
rect 54256 10276 54262 10328
rect 65502 10204 65530 18104
rect 65582 10204 65610 18104
rect 65662 10204 65690 18104
rect 65742 10204 65770 18104
rect 65822 10204 65850 18104
rect 65902 10204 65930 18104
rect 65982 10204 66010 18104
rect 7564 9645 7570 9697
rect 7622 9685 7628 9697
rect 11532 9685 11538 9697
rect 7622 9657 11538 9685
rect 7622 9645 7628 9657
rect 11532 9645 11538 9657
rect 11590 9645 11596 9697
rect 12864 9273 12892 9385
rect 12488 9245 12892 9273
rect 12936 9273 12964 9385
rect 13128 9273 13156 9385
rect 12936 9245 12980 9273
rect 12488 9133 12516 9245
rect 12952 9133 12980 9245
rect 13112 9245 13156 9273
rect 13200 9273 13228 9385
rect 14112 9273 14140 9385
rect 13200 9245 13604 9273
rect 13112 9133 13140 9245
rect 13576 9133 13604 9245
rect 13736 9245 14140 9273
rect 14184 9273 14212 9385
rect 14376 9273 14404 9385
rect 14184 9245 14228 9273
rect 13736 9133 13764 9245
rect 14200 9133 14228 9245
rect 14360 9245 14404 9273
rect 14448 9273 14476 9385
rect 15360 9273 15388 9385
rect 14448 9245 14852 9273
rect 14360 9133 14388 9245
rect 14824 9133 14852 9245
rect 14984 9245 15388 9273
rect 15432 9273 15460 9385
rect 15624 9273 15652 9385
rect 15432 9245 15476 9273
rect 14984 9133 15012 9245
rect 15448 9133 15476 9245
rect 15608 9245 15652 9273
rect 15696 9273 15724 9385
rect 16608 9273 16636 9385
rect 15696 9245 16100 9273
rect 15608 9133 15636 9245
rect 16072 9133 16100 9245
rect 16232 9245 16636 9273
rect 16680 9273 16708 9385
rect 16872 9273 16900 9385
rect 16680 9245 16724 9273
rect 16232 9133 16260 9245
rect 16696 9133 16724 9245
rect 16856 9245 16900 9273
rect 16944 9273 16972 9385
rect 17856 9273 17884 9385
rect 16944 9245 17348 9273
rect 16856 9133 16884 9245
rect 17320 9133 17348 9245
rect 17480 9245 17884 9273
rect 17928 9273 17956 9385
rect 18120 9273 18148 9385
rect 17928 9245 17972 9273
rect 17480 9133 17508 9245
rect 17944 9133 17972 9245
rect 18104 9245 18148 9273
rect 18192 9273 18220 9385
rect 19104 9273 19132 9385
rect 18192 9245 18596 9273
rect 18104 9133 18132 9245
rect 18568 9133 18596 9245
rect 18728 9245 19132 9273
rect 19176 9273 19204 9385
rect 19368 9273 19396 9385
rect 19176 9245 19220 9273
rect 18728 9133 18756 9245
rect 19192 9133 19220 9245
rect 19352 9245 19396 9273
rect 19440 9273 19468 9385
rect 20352 9273 20380 9385
rect 19440 9245 19844 9273
rect 19352 9133 19380 9245
rect 19816 9133 19844 9245
rect 19976 9245 20380 9273
rect 20424 9273 20452 9385
rect 20616 9273 20644 9385
rect 20424 9245 20468 9273
rect 19976 9133 20004 9245
rect 20440 9133 20468 9245
rect 20600 9245 20644 9273
rect 20688 9273 20716 9385
rect 21600 9273 21628 9385
rect 20688 9245 21092 9273
rect 20600 9133 20628 9245
rect 21064 9133 21092 9245
rect 21224 9245 21628 9273
rect 21672 9273 21700 9385
rect 21864 9273 21892 9385
rect 21672 9245 21716 9273
rect 21224 9133 21252 9245
rect 21688 9133 21716 9245
rect 21848 9245 21892 9273
rect 21936 9273 21964 9385
rect 22848 9273 22876 9385
rect 21936 9245 22340 9273
rect 21848 9133 21876 9245
rect 22312 9133 22340 9245
rect 22472 9245 22876 9273
rect 22920 9273 22948 9385
rect 23112 9273 23140 9385
rect 22920 9245 22964 9273
rect 22472 9133 22500 9245
rect 22936 9133 22964 9245
rect 23096 9245 23140 9273
rect 23184 9273 23212 9385
rect 24096 9273 24124 9385
rect 23184 9245 23588 9273
rect 23096 9133 23124 9245
rect 23560 9133 23588 9245
rect 23720 9245 24124 9273
rect 24168 9273 24196 9385
rect 24360 9273 24388 9385
rect 24168 9245 24212 9273
rect 23720 9133 23748 9245
rect 24184 9133 24212 9245
rect 24344 9245 24388 9273
rect 24432 9273 24460 9385
rect 25344 9273 25372 9385
rect 24432 9245 24836 9273
rect 24344 9133 24372 9245
rect 24808 9133 24836 9245
rect 24968 9245 25372 9273
rect 25416 9273 25444 9385
rect 25608 9273 25636 9385
rect 25416 9245 25460 9273
rect 24968 9133 24996 9245
rect 25432 9133 25460 9245
rect 25592 9245 25636 9273
rect 25680 9273 25708 9385
rect 26592 9273 26620 9385
rect 25680 9245 26084 9273
rect 25592 9133 25620 9245
rect 26056 9133 26084 9245
rect 26216 9245 26620 9273
rect 26664 9273 26692 9385
rect 26856 9273 26884 9385
rect 26664 9245 26708 9273
rect 26216 9133 26244 9245
rect 26680 9133 26708 9245
rect 26840 9245 26884 9273
rect 26928 9273 26956 9385
rect 27840 9273 27868 9385
rect 26928 9245 27332 9273
rect 26840 9133 26868 9245
rect 27304 9133 27332 9245
rect 27464 9245 27868 9273
rect 27912 9273 27940 9385
rect 28104 9273 28132 9385
rect 27912 9245 27956 9273
rect 27464 9133 27492 9245
rect 27928 9133 27956 9245
rect 28088 9245 28132 9273
rect 28176 9273 28204 9385
rect 29088 9273 29116 9385
rect 28176 9245 28580 9273
rect 28088 9133 28116 9245
rect 28552 9133 28580 9245
rect 28712 9245 29116 9273
rect 29160 9273 29188 9385
rect 29352 9273 29380 9385
rect 29160 9245 29204 9273
rect 28712 9133 28740 9245
rect 29176 9133 29204 9245
rect 29336 9245 29380 9273
rect 29424 9273 29452 9385
rect 30336 9273 30364 9385
rect 29424 9245 29828 9273
rect 29336 9133 29364 9245
rect 29800 9133 29828 9245
rect 29960 9245 30364 9273
rect 30408 9273 30436 9385
rect 30600 9273 30628 9385
rect 30408 9245 30452 9273
rect 29960 9133 29988 9245
rect 30424 9133 30452 9245
rect 30584 9245 30628 9273
rect 30672 9273 30700 9385
rect 31584 9273 31612 9385
rect 30672 9245 31076 9273
rect 30584 9133 30612 9245
rect 31048 9133 31076 9245
rect 31208 9245 31612 9273
rect 31656 9273 31684 9385
rect 31848 9273 31876 9385
rect 31656 9245 31700 9273
rect 31208 9133 31236 9245
rect 31672 9133 31700 9245
rect 31832 9245 31876 9273
rect 31920 9273 31948 9385
rect 32832 9273 32860 9385
rect 31920 9245 32324 9273
rect 31832 9133 31860 9245
rect 32296 9133 32324 9245
rect 32456 9245 32860 9273
rect 32904 9273 32932 9385
rect 33096 9273 33124 9385
rect 32904 9245 32948 9273
rect 32456 9133 32484 9245
rect 32920 9133 32948 9245
rect 33080 9245 33124 9273
rect 33168 9273 33196 9385
rect 34080 9273 34108 9385
rect 33168 9245 33572 9273
rect 33080 9133 33108 9245
rect 33544 9133 33572 9245
rect 33704 9245 34108 9273
rect 34152 9273 34180 9385
rect 34344 9273 34372 9385
rect 34152 9245 34196 9273
rect 33704 9133 33732 9245
rect 34168 9133 34196 9245
rect 34328 9245 34372 9273
rect 34416 9273 34444 9385
rect 35328 9273 35356 9385
rect 34416 9245 34820 9273
rect 34328 9133 34356 9245
rect 34792 9133 34820 9245
rect 34952 9245 35356 9273
rect 35400 9273 35428 9385
rect 35592 9273 35620 9385
rect 35400 9245 35444 9273
rect 34952 9133 34980 9245
rect 35416 9133 35444 9245
rect 35576 9245 35620 9273
rect 35664 9273 35692 9385
rect 36576 9273 36604 9385
rect 35664 9245 36068 9273
rect 35576 9133 35604 9245
rect 36040 9133 36068 9245
rect 36200 9245 36604 9273
rect 36648 9273 36676 9385
rect 36840 9273 36868 9385
rect 36648 9245 36692 9273
rect 36200 9133 36228 9245
rect 36664 9133 36692 9245
rect 36824 9245 36868 9273
rect 36912 9273 36940 9385
rect 37824 9273 37852 9385
rect 36912 9245 37316 9273
rect 36824 9133 36852 9245
rect 37288 9133 37316 9245
rect 37448 9245 37852 9273
rect 37896 9273 37924 9385
rect 38088 9273 38116 9385
rect 37896 9245 37940 9273
rect 37448 9133 37476 9245
rect 37912 9133 37940 9245
rect 38072 9245 38116 9273
rect 38160 9273 38188 9385
rect 39072 9273 39100 9385
rect 38160 9245 38564 9273
rect 38072 9133 38100 9245
rect 38536 9133 38564 9245
rect 38696 9245 39100 9273
rect 39144 9273 39172 9385
rect 39336 9273 39364 9385
rect 39144 9245 39188 9273
rect 38696 9133 38724 9245
rect 39160 9133 39188 9245
rect 39320 9245 39364 9273
rect 39408 9273 39436 9385
rect 40320 9273 40348 9385
rect 39408 9245 39812 9273
rect 39320 9133 39348 9245
rect 39784 9133 39812 9245
rect 39944 9245 40348 9273
rect 40392 9273 40420 9385
rect 40584 9273 40612 9385
rect 40392 9245 40436 9273
rect 39944 9133 39972 9245
rect 40408 9133 40436 9245
rect 40568 9245 40612 9273
rect 40656 9273 40684 9385
rect 41568 9273 41596 9385
rect 40656 9245 41060 9273
rect 40568 9133 40596 9245
rect 41032 9133 41060 9245
rect 41192 9245 41596 9273
rect 41640 9273 41668 9385
rect 41832 9273 41860 9385
rect 41640 9245 41684 9273
rect 41192 9133 41220 9245
rect 41656 9133 41684 9245
rect 41816 9245 41860 9273
rect 41904 9273 41932 9385
rect 42816 9273 42844 9385
rect 41904 9245 42308 9273
rect 41816 9133 41844 9245
rect 42280 9133 42308 9245
rect 42440 9245 42844 9273
rect 42888 9273 42916 9385
rect 43080 9273 43108 9385
rect 42888 9245 42932 9273
rect 42440 9133 42468 9245
rect 42904 9133 42932 9245
rect 43064 9245 43108 9273
rect 43152 9273 43180 9385
rect 44064 9273 44092 9385
rect 43152 9245 43556 9273
rect 43064 9133 43092 9245
rect 43528 9133 43556 9245
rect 43688 9245 44092 9273
rect 44136 9273 44164 9385
rect 44328 9273 44356 9385
rect 44136 9245 44180 9273
rect 43688 9133 43716 9245
rect 44152 9133 44180 9245
rect 44312 9245 44356 9273
rect 44400 9273 44428 9385
rect 45312 9273 45340 9385
rect 44400 9245 44804 9273
rect 44312 9133 44340 9245
rect 44776 9133 44804 9245
rect 44936 9245 45340 9273
rect 45384 9273 45412 9385
rect 45576 9273 45604 9385
rect 45384 9245 45428 9273
rect 44936 9133 44964 9245
rect 45400 9133 45428 9245
rect 45560 9245 45604 9273
rect 45648 9273 45676 9385
rect 46560 9273 46588 9385
rect 45648 9245 46052 9273
rect 45560 9133 45588 9245
rect 46024 9133 46052 9245
rect 46184 9245 46588 9273
rect 46632 9273 46660 9385
rect 46824 9273 46852 9385
rect 46632 9245 46676 9273
rect 46184 9133 46212 9245
rect 46648 9133 46676 9245
rect 46808 9245 46852 9273
rect 46896 9273 46924 9385
rect 47808 9273 47836 9385
rect 46896 9245 47300 9273
rect 46808 9133 46836 9245
rect 47272 9133 47300 9245
rect 47432 9245 47836 9273
rect 47880 9273 47908 9385
rect 48072 9273 48100 9385
rect 47880 9245 47924 9273
rect 47432 9133 47460 9245
rect 47896 9133 47924 9245
rect 48056 9245 48100 9273
rect 48144 9273 48172 9385
rect 49056 9273 49084 9385
rect 48144 9245 48548 9273
rect 48056 9133 48084 9245
rect 48520 9133 48548 9245
rect 48680 9245 49084 9273
rect 49128 9273 49156 9385
rect 49320 9273 49348 9385
rect 49128 9245 49172 9273
rect 48680 9133 48708 9245
rect 49144 9133 49172 9245
rect 49304 9245 49348 9273
rect 49392 9273 49420 9385
rect 50304 9273 50332 9385
rect 49392 9245 49796 9273
rect 49304 9133 49332 9245
rect 49768 9133 49796 9245
rect 49928 9245 50332 9273
rect 50376 9273 50404 9385
rect 50568 9273 50596 9385
rect 50376 9245 50420 9273
rect 49928 9133 49956 9245
rect 50392 9133 50420 9245
rect 50552 9245 50596 9273
rect 50640 9273 50668 9385
rect 51552 9273 51580 9385
rect 50640 9245 51044 9273
rect 50552 9133 50580 9245
rect 51016 9133 51044 9245
rect 51176 9245 51580 9273
rect 51624 9273 51652 9385
rect 51816 9273 51844 9385
rect 51624 9245 51668 9273
rect 51176 9133 51204 9245
rect 51640 9133 51668 9245
rect 51800 9245 51844 9273
rect 51888 9273 51916 9385
rect 52800 9273 52828 9385
rect 51888 9245 52292 9273
rect 51800 9133 51828 9245
rect 52264 9133 52292 9245
rect 52424 9245 52828 9273
rect 52872 9273 52900 9385
rect 52872 9245 52916 9273
rect 52424 9133 52452 9245
rect 52888 9133 52916 9245
rect 12952 8281 12980 8379
rect 12934 8229 12940 8281
rect 12992 8229 12998 8281
rect 6456 7591 6462 7643
rect 6514 7591 6520 7643
rect 6456 6177 6462 6229
rect 6514 6177 6520 6229
rect 6456 4763 6462 4815
rect 6514 4763 6520 4815
rect 13150 3635 13196 3889
rect 14398 3635 14444 3889
rect 15646 3635 15692 3889
rect 16894 3635 16940 3889
rect 18142 3635 18188 3889
rect 19390 3635 19436 3889
rect 20638 3635 20684 3889
rect 21886 3635 21932 3889
rect 23134 3635 23180 3889
rect 24382 3635 24428 3889
rect 25630 3635 25676 3889
rect 26878 3635 26924 3889
rect 28126 3635 28172 3889
rect 29374 3635 29420 3889
rect 30622 3635 30668 3889
rect 31870 3635 31916 3889
rect 33118 3635 33164 3889
rect 34366 3635 34412 3889
rect 35614 3635 35660 3889
rect 36862 3635 36908 3889
rect 38110 3635 38156 3889
rect 39358 3635 39404 3889
rect 40606 3635 40652 3889
rect 41854 3635 41900 3889
rect 43102 3635 43148 3889
rect 44350 3635 44396 3889
rect 45598 3635 45644 3889
rect 46846 3635 46892 3889
rect 48094 3635 48140 3889
rect 49342 3635 49388 3889
rect 50590 3635 50636 3889
rect 51838 3635 51884 3889
rect 13301 1376 13361 1432
rect 14549 1376 14609 1432
rect 15797 1376 15857 1432
rect 17045 1376 17105 1432
rect 18293 1376 18353 1432
rect 19541 1376 19601 1432
rect 20789 1376 20849 1432
rect 22037 1376 22097 1432
rect 23285 1376 23345 1432
rect 24533 1376 24593 1432
rect 25781 1376 25841 1432
rect 27029 1376 27089 1432
rect 28277 1376 28337 1432
rect 29525 1376 29585 1432
rect 30773 1376 30833 1432
rect 32021 1376 32081 1432
rect 33269 1376 33329 1432
rect 34517 1376 34577 1432
rect 35765 1376 35825 1432
rect 37013 1376 37073 1432
rect 38261 1376 38321 1432
rect 39509 1376 39569 1432
rect 40757 1376 40817 1432
rect 42005 1376 42065 1432
rect 43253 1376 43313 1432
rect 44501 1376 44561 1432
rect 45749 1376 45809 1432
rect 46997 1376 47057 1432
rect 48245 1376 48305 1432
rect 49493 1376 49553 1432
rect 50741 1376 50801 1432
rect 51989 1376 52049 1432
<< via1 >>
rect 59390 66138 59442 66147
rect 59390 66104 59399 66138
rect 59399 66104 59433 66138
rect 59433 66104 59442 66138
rect 59390 66095 59442 66104
rect 59390 64724 59442 64733
rect 59390 64690 59399 64724
rect 59399 64690 59433 64724
rect 59433 64690 59442 64724
rect 59390 64681 59442 64690
rect 59390 63310 59442 63319
rect 59390 63276 59399 63310
rect 59399 63276 59433 63310
rect 59433 63276 59442 63310
rect 59390 63267 59442 63276
rect 53036 62629 53088 62681
rect 54342 61213 54394 61265
rect 58406 61213 58458 61265
rect 54204 60625 54256 60634
rect 54204 60591 54213 60625
rect 54213 60591 54247 60625
rect 54247 60591 54256 60625
rect 54204 60582 54256 60591
rect 11772 60405 11824 60414
rect 11772 60371 11781 60405
rect 11781 60371 11815 60405
rect 11815 60371 11824 60405
rect 11772 60362 11824 60371
rect 11772 60309 11824 60318
rect 11772 60275 11781 60309
rect 11781 60275 11815 60309
rect 11815 60275 11824 60309
rect 11772 60266 11824 60275
rect 54204 60089 54256 60098
rect 54204 60055 54213 60089
rect 54213 60055 54247 60089
rect 54247 60055 54256 60089
rect 54204 60046 54256 60055
rect 54204 59835 54256 59844
rect 54204 59801 54213 59835
rect 54213 59801 54247 59835
rect 54247 59801 54256 59835
rect 54204 59792 54256 59801
rect 11772 59615 11824 59624
rect 11772 59581 11781 59615
rect 11781 59581 11815 59615
rect 11815 59581 11824 59615
rect 11772 59572 11824 59581
rect 11772 59519 11824 59528
rect 11772 59485 11781 59519
rect 11781 59485 11815 59519
rect 11815 59485 11824 59519
rect 11772 59476 11824 59485
rect 54204 59299 54256 59308
rect 54204 59265 54213 59299
rect 54213 59265 54247 59299
rect 54247 59265 54256 59299
rect 54204 59256 54256 59265
rect 54204 59045 54256 59054
rect 54204 59011 54213 59045
rect 54213 59011 54247 59045
rect 54247 59011 54256 59045
rect 54204 59002 54256 59011
rect 11772 58825 11824 58834
rect 11772 58791 11781 58825
rect 11781 58791 11815 58825
rect 11815 58791 11824 58825
rect 11772 58782 11824 58791
rect 11772 58729 11824 58738
rect 11772 58695 11781 58729
rect 11781 58695 11815 58729
rect 11815 58695 11824 58729
rect 11772 58686 11824 58695
rect 54204 58509 54256 58518
rect 54204 58475 54213 58509
rect 54213 58475 54247 58509
rect 54247 58475 54256 58509
rect 54204 58466 54256 58475
rect 54204 58255 54256 58264
rect 54204 58221 54213 58255
rect 54213 58221 54247 58255
rect 54247 58221 54256 58255
rect 54204 58212 54256 58221
rect 11772 58035 11824 58044
rect 11772 58001 11781 58035
rect 11781 58001 11815 58035
rect 11815 58001 11824 58035
rect 11772 57992 11824 58001
rect 11772 57939 11824 57948
rect 11772 57905 11781 57939
rect 11781 57905 11815 57939
rect 11815 57905 11824 57939
rect 11772 57896 11824 57905
rect 54204 57719 54256 57728
rect 54204 57685 54213 57719
rect 54213 57685 54247 57719
rect 54247 57685 54256 57719
rect 54204 57676 54256 57685
rect 54204 57465 54256 57474
rect 54204 57431 54213 57465
rect 54213 57431 54247 57465
rect 54247 57431 54256 57465
rect 54204 57422 54256 57431
rect 11772 57245 11824 57254
rect 11772 57211 11781 57245
rect 11781 57211 11815 57245
rect 11815 57211 11824 57245
rect 11772 57202 11824 57211
rect 11772 57149 11824 57158
rect 11772 57115 11781 57149
rect 11781 57115 11815 57149
rect 11815 57115 11824 57149
rect 11772 57106 11824 57115
rect 54204 56929 54256 56938
rect 54204 56895 54213 56929
rect 54213 56895 54247 56929
rect 54247 56895 54256 56929
rect 54204 56886 54256 56895
rect 54204 56675 54256 56684
rect 54204 56641 54213 56675
rect 54213 56641 54247 56675
rect 54247 56641 54256 56675
rect 54204 56632 54256 56641
rect 11772 56455 11824 56464
rect 11772 56421 11781 56455
rect 11781 56421 11815 56455
rect 11815 56421 11824 56455
rect 11772 56412 11824 56421
rect 11772 56359 11824 56368
rect 11772 56325 11781 56359
rect 11781 56325 11815 56359
rect 11815 56325 11824 56359
rect 11772 56316 11824 56325
rect 54204 56139 54256 56148
rect 54204 56105 54213 56139
rect 54213 56105 54247 56139
rect 54247 56105 54256 56139
rect 54204 56096 54256 56105
rect 54204 55885 54256 55894
rect 54204 55851 54213 55885
rect 54213 55851 54247 55885
rect 54247 55851 54256 55885
rect 54204 55842 54256 55851
rect 11772 55665 11824 55674
rect 11772 55631 11781 55665
rect 11781 55631 11815 55665
rect 11815 55631 11824 55665
rect 11772 55622 11824 55631
rect 11772 55569 11824 55578
rect 11772 55535 11781 55569
rect 11781 55535 11815 55569
rect 11815 55535 11824 55569
rect 11772 55526 11824 55535
rect 54204 55349 54256 55358
rect 54204 55315 54213 55349
rect 54213 55315 54247 55349
rect 54247 55315 54256 55349
rect 54204 55306 54256 55315
rect 54204 55095 54256 55104
rect 54204 55061 54213 55095
rect 54213 55061 54247 55095
rect 54247 55061 54256 55095
rect 54204 55052 54256 55061
rect 11772 54875 11824 54884
rect 11772 54841 11781 54875
rect 11781 54841 11815 54875
rect 11815 54841 11824 54875
rect 11772 54832 11824 54841
rect 11772 54779 11824 54788
rect 11772 54745 11781 54779
rect 11781 54745 11815 54779
rect 11815 54745 11824 54779
rect 11772 54736 11824 54745
rect 54204 54559 54256 54568
rect 54204 54525 54213 54559
rect 54213 54525 54247 54559
rect 54247 54525 54256 54559
rect 54204 54516 54256 54525
rect 54204 54305 54256 54314
rect 54204 54271 54213 54305
rect 54213 54271 54247 54305
rect 54247 54271 54256 54305
rect 54204 54262 54256 54271
rect 11772 54085 11824 54094
rect 11772 54051 11781 54085
rect 11781 54051 11815 54085
rect 11815 54051 11824 54085
rect 11772 54042 11824 54051
rect 11772 53989 11824 53998
rect 11772 53955 11781 53989
rect 11781 53955 11815 53989
rect 11815 53955 11824 53989
rect 11772 53946 11824 53955
rect 54204 53769 54256 53778
rect 54204 53735 54213 53769
rect 54213 53735 54247 53769
rect 54247 53735 54256 53769
rect 54204 53726 54256 53735
rect 54204 53515 54256 53524
rect 54204 53481 54213 53515
rect 54213 53481 54247 53515
rect 54247 53481 54256 53515
rect 54204 53472 54256 53481
rect 11772 53295 11824 53304
rect 11772 53261 11781 53295
rect 11781 53261 11815 53295
rect 11815 53261 11824 53295
rect 11772 53252 11824 53261
rect 11772 53199 11824 53208
rect 11772 53165 11781 53199
rect 11781 53165 11815 53199
rect 11815 53165 11824 53199
rect 11772 53156 11824 53165
rect 54204 52979 54256 52988
rect 54204 52945 54213 52979
rect 54213 52945 54247 52979
rect 54247 52945 54256 52979
rect 54204 52936 54256 52945
rect 54204 52725 54256 52734
rect 54204 52691 54213 52725
rect 54213 52691 54247 52725
rect 54247 52691 54256 52725
rect 54204 52682 54256 52691
rect 11772 52505 11824 52514
rect 11772 52471 11781 52505
rect 11781 52471 11815 52505
rect 11815 52471 11824 52505
rect 11772 52462 11824 52471
rect 11772 52409 11824 52418
rect 11772 52375 11781 52409
rect 11781 52375 11815 52409
rect 11815 52375 11824 52409
rect 11772 52366 11824 52375
rect 54204 52189 54256 52198
rect 54204 52155 54213 52189
rect 54213 52155 54247 52189
rect 54247 52155 54256 52189
rect 54204 52146 54256 52155
rect 54204 51935 54256 51944
rect 54204 51901 54213 51935
rect 54213 51901 54247 51935
rect 54247 51901 54256 51935
rect 54204 51892 54256 51901
rect 11772 51715 11824 51724
rect 11772 51681 11781 51715
rect 11781 51681 11815 51715
rect 11815 51681 11824 51715
rect 11772 51672 11824 51681
rect 11772 51619 11824 51628
rect 11772 51585 11781 51619
rect 11781 51585 11815 51619
rect 11815 51585 11824 51619
rect 11772 51576 11824 51585
rect 54204 51399 54256 51408
rect 54204 51365 54213 51399
rect 54213 51365 54247 51399
rect 54247 51365 54256 51399
rect 54204 51356 54256 51365
rect 54204 51145 54256 51154
rect 54204 51111 54213 51145
rect 54213 51111 54247 51145
rect 54247 51111 54256 51145
rect 54204 51102 54256 51111
rect 11772 50925 11824 50934
rect 11772 50891 11781 50925
rect 11781 50891 11815 50925
rect 11815 50891 11824 50925
rect 11772 50882 11824 50891
rect 11772 50829 11824 50838
rect 11772 50795 11781 50829
rect 11781 50795 11815 50829
rect 11815 50795 11824 50829
rect 11772 50786 11824 50795
rect 54204 50609 54256 50618
rect 54204 50575 54213 50609
rect 54213 50575 54247 50609
rect 54247 50575 54256 50609
rect 54204 50566 54256 50575
rect 54204 50355 54256 50364
rect 54204 50321 54213 50355
rect 54213 50321 54247 50355
rect 54247 50321 54256 50355
rect 54204 50312 54256 50321
rect 11772 50135 11824 50144
rect 11772 50101 11781 50135
rect 11781 50101 11815 50135
rect 11815 50101 11824 50135
rect 11772 50092 11824 50101
rect 11772 50039 11824 50048
rect 11772 50005 11781 50039
rect 11781 50005 11815 50039
rect 11815 50005 11824 50039
rect 11772 49996 11824 50005
rect 54204 49819 54256 49828
rect 54204 49785 54213 49819
rect 54213 49785 54247 49819
rect 54247 49785 54256 49819
rect 54204 49776 54256 49785
rect 54204 49565 54256 49574
rect 54204 49531 54213 49565
rect 54213 49531 54247 49565
rect 54247 49531 54256 49565
rect 54204 49522 54256 49531
rect 11772 49345 11824 49354
rect 11772 49311 11781 49345
rect 11781 49311 11815 49345
rect 11815 49311 11824 49345
rect 11772 49302 11824 49311
rect 11772 49249 11824 49258
rect 11772 49215 11781 49249
rect 11781 49215 11815 49249
rect 11815 49215 11824 49249
rect 11772 49206 11824 49215
rect 54204 49029 54256 49038
rect 54204 48995 54213 49029
rect 54213 48995 54247 49029
rect 54247 48995 54256 49029
rect 54204 48986 54256 48995
rect 54204 48775 54256 48784
rect 54204 48741 54213 48775
rect 54213 48741 54247 48775
rect 54247 48741 54256 48775
rect 54204 48732 54256 48741
rect 11772 48555 11824 48564
rect 11772 48521 11781 48555
rect 11781 48521 11815 48555
rect 11815 48521 11824 48555
rect 11772 48512 11824 48521
rect 11772 48459 11824 48468
rect 11772 48425 11781 48459
rect 11781 48425 11815 48459
rect 11815 48425 11824 48459
rect 11772 48416 11824 48425
rect 54204 48239 54256 48248
rect 54204 48205 54213 48239
rect 54213 48205 54247 48239
rect 54247 48205 54256 48239
rect 54204 48196 54256 48205
rect 54204 47985 54256 47994
rect 54204 47951 54213 47985
rect 54213 47951 54247 47985
rect 54247 47951 54256 47985
rect 54204 47942 54256 47951
rect 11772 47765 11824 47774
rect 11772 47731 11781 47765
rect 11781 47731 11815 47765
rect 11815 47731 11824 47765
rect 11772 47722 11824 47731
rect 11772 47669 11824 47678
rect 11772 47635 11781 47669
rect 11781 47635 11815 47669
rect 11815 47635 11824 47669
rect 11772 47626 11824 47635
rect 54204 47449 54256 47458
rect 54204 47415 54213 47449
rect 54213 47415 54247 47449
rect 54247 47415 54256 47449
rect 54204 47406 54256 47415
rect 54204 47195 54256 47204
rect 54204 47161 54213 47195
rect 54213 47161 54247 47195
rect 54247 47161 54256 47195
rect 54204 47152 54256 47161
rect 11772 46975 11824 46984
rect 11772 46941 11781 46975
rect 11781 46941 11815 46975
rect 11815 46941 11824 46975
rect 11772 46932 11824 46941
rect 11772 46879 11824 46888
rect 11772 46845 11781 46879
rect 11781 46845 11815 46879
rect 11815 46845 11824 46879
rect 11772 46836 11824 46845
rect 54204 46659 54256 46668
rect 54204 46625 54213 46659
rect 54213 46625 54247 46659
rect 54247 46625 54256 46659
rect 54204 46616 54256 46625
rect 54204 46405 54256 46414
rect 54204 46371 54213 46405
rect 54213 46371 54247 46405
rect 54247 46371 54256 46405
rect 54204 46362 54256 46371
rect 11772 46185 11824 46194
rect 11772 46151 11781 46185
rect 11781 46151 11815 46185
rect 11815 46151 11824 46185
rect 11772 46142 11824 46151
rect 11772 46089 11824 46098
rect 11772 46055 11781 46089
rect 11781 46055 11815 46089
rect 11815 46055 11824 46089
rect 11772 46046 11824 46055
rect 54204 45869 54256 45878
rect 54204 45835 54213 45869
rect 54213 45835 54247 45869
rect 54247 45835 54256 45869
rect 54204 45826 54256 45835
rect 54204 45615 54256 45624
rect 54204 45581 54213 45615
rect 54213 45581 54247 45615
rect 54247 45581 54256 45615
rect 54204 45572 54256 45581
rect 11772 45395 11824 45404
rect 11772 45361 11781 45395
rect 11781 45361 11815 45395
rect 11815 45361 11824 45395
rect 11772 45352 11824 45361
rect 11772 45299 11824 45308
rect 11772 45265 11781 45299
rect 11781 45265 11815 45299
rect 11815 45265 11824 45299
rect 11772 45256 11824 45265
rect 54204 45079 54256 45088
rect 54204 45045 54213 45079
rect 54213 45045 54247 45079
rect 54247 45045 54256 45079
rect 54204 45036 54256 45045
rect 54204 44825 54256 44834
rect 54204 44791 54213 44825
rect 54213 44791 54247 44825
rect 54247 44791 54256 44825
rect 54204 44782 54256 44791
rect 11772 44605 11824 44614
rect 11772 44571 11781 44605
rect 11781 44571 11815 44605
rect 11815 44571 11824 44605
rect 11772 44562 11824 44571
rect 11772 44509 11824 44518
rect 11772 44475 11781 44509
rect 11781 44475 11815 44509
rect 11815 44475 11824 44509
rect 11772 44466 11824 44475
rect 54204 44289 54256 44298
rect 54204 44255 54213 44289
rect 54213 44255 54247 44289
rect 54247 44255 54256 44289
rect 54204 44246 54256 44255
rect 54204 44035 54256 44044
rect 54204 44001 54213 44035
rect 54213 44001 54247 44035
rect 54247 44001 54256 44035
rect 54204 43992 54256 44001
rect 11772 43815 11824 43824
rect 11772 43781 11781 43815
rect 11781 43781 11815 43815
rect 11815 43781 11824 43815
rect 11772 43772 11824 43781
rect 11772 43719 11824 43728
rect 11772 43685 11781 43719
rect 11781 43685 11815 43719
rect 11815 43685 11824 43719
rect 11772 43676 11824 43685
rect 54204 43499 54256 43508
rect 54204 43465 54213 43499
rect 54213 43465 54247 43499
rect 54247 43465 54256 43499
rect 54204 43456 54256 43465
rect 54204 43245 54256 43254
rect 54204 43211 54213 43245
rect 54213 43211 54247 43245
rect 54247 43211 54256 43245
rect 54204 43202 54256 43211
rect 11772 43025 11824 43034
rect 11772 42991 11781 43025
rect 11781 42991 11815 43025
rect 11815 42991 11824 43025
rect 11772 42982 11824 42991
rect 11772 42929 11824 42938
rect 11772 42895 11781 42929
rect 11781 42895 11815 42929
rect 11815 42895 11824 42929
rect 11772 42886 11824 42895
rect 54204 42709 54256 42718
rect 54204 42675 54213 42709
rect 54213 42675 54247 42709
rect 54247 42675 54256 42709
rect 54204 42666 54256 42675
rect 54204 42455 54256 42464
rect 54204 42421 54213 42455
rect 54213 42421 54247 42455
rect 54247 42421 54256 42455
rect 54204 42412 54256 42421
rect 11772 42235 11824 42244
rect 11772 42201 11781 42235
rect 11781 42201 11815 42235
rect 11815 42201 11824 42235
rect 11772 42192 11824 42201
rect 11772 42139 11824 42148
rect 11772 42105 11781 42139
rect 11781 42105 11815 42139
rect 11815 42105 11824 42139
rect 11772 42096 11824 42105
rect 54204 41919 54256 41928
rect 54204 41885 54213 41919
rect 54213 41885 54247 41919
rect 54247 41885 54256 41919
rect 54204 41876 54256 41885
rect 54204 41665 54256 41674
rect 54204 41631 54213 41665
rect 54213 41631 54247 41665
rect 54247 41631 54256 41665
rect 54204 41622 54256 41631
rect 11772 41445 11824 41454
rect 11772 41411 11781 41445
rect 11781 41411 11815 41445
rect 11815 41411 11824 41445
rect 11772 41402 11824 41411
rect 11772 41349 11824 41358
rect 11772 41315 11781 41349
rect 11781 41315 11815 41349
rect 11815 41315 11824 41349
rect 11772 41306 11824 41315
rect 54204 41129 54256 41138
rect 54204 41095 54213 41129
rect 54213 41095 54247 41129
rect 54247 41095 54256 41129
rect 54204 41086 54256 41095
rect 54204 40875 54256 40884
rect 54204 40841 54213 40875
rect 54213 40841 54247 40875
rect 54247 40841 54256 40875
rect 54204 40832 54256 40841
rect 11772 40655 11824 40664
rect 11772 40621 11781 40655
rect 11781 40621 11815 40655
rect 11815 40621 11824 40655
rect 11772 40612 11824 40621
rect 11772 40559 11824 40568
rect 11772 40525 11781 40559
rect 11781 40525 11815 40559
rect 11815 40525 11824 40559
rect 11772 40516 11824 40525
rect 54204 40339 54256 40348
rect 54204 40305 54213 40339
rect 54213 40305 54247 40339
rect 54247 40305 54256 40339
rect 54204 40296 54256 40305
rect 54204 40085 54256 40094
rect 54204 40051 54213 40085
rect 54213 40051 54247 40085
rect 54247 40051 54256 40085
rect 54204 40042 54256 40051
rect 11772 39865 11824 39874
rect 11772 39831 11781 39865
rect 11781 39831 11815 39865
rect 11815 39831 11824 39865
rect 11772 39822 11824 39831
rect 11772 39769 11824 39778
rect 11772 39735 11781 39769
rect 11781 39735 11815 39769
rect 11815 39735 11824 39769
rect 11772 39726 11824 39735
rect 54204 39549 54256 39558
rect 54204 39515 54213 39549
rect 54213 39515 54247 39549
rect 54247 39515 54256 39549
rect 54204 39506 54256 39515
rect 54204 39295 54256 39304
rect 54204 39261 54213 39295
rect 54213 39261 54247 39295
rect 54247 39261 54256 39295
rect 54204 39252 54256 39261
rect 11772 39075 11824 39084
rect 11772 39041 11781 39075
rect 11781 39041 11815 39075
rect 11815 39041 11824 39075
rect 11772 39032 11824 39041
rect 11772 38979 11824 38988
rect 11772 38945 11781 38979
rect 11781 38945 11815 38979
rect 11815 38945 11824 38979
rect 11772 38936 11824 38945
rect 54204 38759 54256 38768
rect 54204 38725 54213 38759
rect 54213 38725 54247 38759
rect 54247 38725 54256 38759
rect 54204 38716 54256 38725
rect 54204 38505 54256 38514
rect 54204 38471 54213 38505
rect 54213 38471 54247 38505
rect 54247 38471 54256 38505
rect 54204 38462 54256 38471
rect 11772 38285 11824 38294
rect 11772 38251 11781 38285
rect 11781 38251 11815 38285
rect 11815 38251 11824 38285
rect 11772 38242 11824 38251
rect 11772 38189 11824 38198
rect 11772 38155 11781 38189
rect 11781 38155 11815 38189
rect 11815 38155 11824 38189
rect 11772 38146 11824 38155
rect 54204 37969 54256 37978
rect 54204 37935 54213 37969
rect 54213 37935 54247 37969
rect 54247 37935 54256 37969
rect 54204 37926 54256 37935
rect 54204 37715 54256 37724
rect 54204 37681 54213 37715
rect 54213 37681 54247 37715
rect 54247 37681 54256 37715
rect 54204 37672 54256 37681
rect 11772 37495 11824 37504
rect 11772 37461 11781 37495
rect 11781 37461 11815 37495
rect 11815 37461 11824 37495
rect 11772 37452 11824 37461
rect 11772 37399 11824 37408
rect 11772 37365 11781 37399
rect 11781 37365 11815 37399
rect 11815 37365 11824 37399
rect 11772 37356 11824 37365
rect 54204 37179 54256 37188
rect 54204 37145 54213 37179
rect 54213 37145 54247 37179
rect 54247 37145 54256 37179
rect 54204 37136 54256 37145
rect 54204 36925 54256 36934
rect 54204 36891 54213 36925
rect 54213 36891 54247 36925
rect 54247 36891 54256 36925
rect 54204 36882 54256 36891
rect 11772 36705 11824 36714
rect 11772 36671 11781 36705
rect 11781 36671 11815 36705
rect 11815 36671 11824 36705
rect 11772 36662 11824 36671
rect 11772 36609 11824 36618
rect 11772 36575 11781 36609
rect 11781 36575 11815 36609
rect 11815 36575 11824 36609
rect 11772 36566 11824 36575
rect 54204 36389 54256 36398
rect 54204 36355 54213 36389
rect 54213 36355 54247 36389
rect 54247 36355 54256 36389
rect 54204 36346 54256 36355
rect 54204 36135 54256 36144
rect 54204 36101 54213 36135
rect 54213 36101 54247 36135
rect 54247 36101 54256 36135
rect 54204 36092 54256 36101
rect 11772 35915 11824 35924
rect 11772 35881 11781 35915
rect 11781 35881 11815 35915
rect 11815 35881 11824 35915
rect 11772 35872 11824 35881
rect 11772 35819 11824 35828
rect 11772 35785 11781 35819
rect 11781 35785 11815 35819
rect 11815 35785 11824 35819
rect 11772 35776 11824 35785
rect 54204 35599 54256 35608
rect 54204 35565 54213 35599
rect 54213 35565 54247 35599
rect 54247 35565 54256 35599
rect 54204 35556 54256 35565
rect 54204 35345 54256 35354
rect 54204 35311 54213 35345
rect 54213 35311 54247 35345
rect 54247 35311 54256 35345
rect 54204 35302 54256 35311
rect 11772 35125 11824 35134
rect 11772 35091 11781 35125
rect 11781 35091 11815 35125
rect 11815 35091 11824 35125
rect 11772 35082 11824 35091
rect 11772 35029 11824 35038
rect 11772 34995 11781 35029
rect 11781 34995 11815 35029
rect 11815 34995 11824 35029
rect 11772 34986 11824 34995
rect 54204 34809 54256 34818
rect 54204 34775 54213 34809
rect 54213 34775 54247 34809
rect 54247 34775 54256 34809
rect 54204 34766 54256 34775
rect 54204 34555 54256 34564
rect 54204 34521 54213 34555
rect 54213 34521 54247 34555
rect 54247 34521 54256 34555
rect 54204 34512 54256 34521
rect 11772 34335 11824 34344
rect 11772 34301 11781 34335
rect 11781 34301 11815 34335
rect 11815 34301 11824 34335
rect 11772 34292 11824 34301
rect 11772 34239 11824 34248
rect 11772 34205 11781 34239
rect 11781 34205 11815 34239
rect 11815 34205 11824 34239
rect 11772 34196 11824 34205
rect 54204 34019 54256 34028
rect 54204 33985 54213 34019
rect 54213 33985 54247 34019
rect 54247 33985 54256 34019
rect 54204 33976 54256 33985
rect 54204 33765 54256 33774
rect 54204 33731 54213 33765
rect 54213 33731 54247 33765
rect 54247 33731 54256 33765
rect 54204 33722 54256 33731
rect 11772 33545 11824 33554
rect 11772 33511 11781 33545
rect 11781 33511 11815 33545
rect 11815 33511 11824 33545
rect 11772 33502 11824 33511
rect 11772 33449 11824 33458
rect 11772 33415 11781 33449
rect 11781 33415 11815 33449
rect 11815 33415 11824 33449
rect 11772 33406 11824 33415
rect 54204 33229 54256 33238
rect 54204 33195 54213 33229
rect 54213 33195 54247 33229
rect 54247 33195 54256 33229
rect 54204 33186 54256 33195
rect 54204 32975 54256 32984
rect 54204 32941 54213 32975
rect 54213 32941 54247 32975
rect 54247 32941 54256 32975
rect 54204 32932 54256 32941
rect 11772 32755 11824 32764
rect 11772 32721 11781 32755
rect 11781 32721 11815 32755
rect 11815 32721 11824 32755
rect 11772 32712 11824 32721
rect 11772 32659 11824 32668
rect 11772 32625 11781 32659
rect 11781 32625 11815 32659
rect 11815 32625 11824 32659
rect 11772 32616 11824 32625
rect 54204 32439 54256 32448
rect 54204 32405 54213 32439
rect 54213 32405 54247 32439
rect 54247 32405 54256 32439
rect 54204 32396 54256 32405
rect 54204 32185 54256 32194
rect 54204 32151 54213 32185
rect 54213 32151 54247 32185
rect 54247 32151 54256 32185
rect 54204 32142 54256 32151
rect 11772 31965 11824 31974
rect 11772 31931 11781 31965
rect 11781 31931 11815 31965
rect 11815 31931 11824 31965
rect 11772 31922 11824 31931
rect 11772 31869 11824 31878
rect 11772 31835 11781 31869
rect 11781 31835 11815 31869
rect 11815 31835 11824 31869
rect 11772 31826 11824 31835
rect 54204 31649 54256 31658
rect 54204 31615 54213 31649
rect 54213 31615 54247 31649
rect 54247 31615 54256 31649
rect 54204 31606 54256 31615
rect 54204 31395 54256 31404
rect 54204 31361 54213 31395
rect 54213 31361 54247 31395
rect 54247 31361 54256 31395
rect 54204 31352 54256 31361
rect 11772 31175 11824 31184
rect 11772 31141 11781 31175
rect 11781 31141 11815 31175
rect 11815 31141 11824 31175
rect 11772 31132 11824 31141
rect 11772 31079 11824 31088
rect 11772 31045 11781 31079
rect 11781 31045 11815 31079
rect 11815 31045 11824 31079
rect 11772 31036 11824 31045
rect 54204 30859 54256 30868
rect 54204 30825 54213 30859
rect 54213 30825 54247 30859
rect 54247 30825 54256 30859
rect 54204 30816 54256 30825
rect 54204 30605 54256 30614
rect 54204 30571 54213 30605
rect 54213 30571 54247 30605
rect 54247 30571 54256 30605
rect 54204 30562 54256 30571
rect 11772 30385 11824 30394
rect 11772 30351 11781 30385
rect 11781 30351 11815 30385
rect 11815 30351 11824 30385
rect 11772 30342 11824 30351
rect 11772 30289 11824 30298
rect 11772 30255 11781 30289
rect 11781 30255 11815 30289
rect 11815 30255 11824 30289
rect 11772 30246 11824 30255
rect 54204 30069 54256 30078
rect 54204 30035 54213 30069
rect 54213 30035 54247 30069
rect 54247 30035 54256 30069
rect 54204 30026 54256 30035
rect 54204 29815 54256 29824
rect 54204 29781 54213 29815
rect 54213 29781 54247 29815
rect 54247 29781 54256 29815
rect 54204 29772 54256 29781
rect 11772 29595 11824 29604
rect 11772 29561 11781 29595
rect 11781 29561 11815 29595
rect 11815 29561 11824 29595
rect 11772 29552 11824 29561
rect 11772 29499 11824 29508
rect 11772 29465 11781 29499
rect 11781 29465 11815 29499
rect 11815 29465 11824 29499
rect 11772 29456 11824 29465
rect 54204 29279 54256 29288
rect 54204 29245 54213 29279
rect 54213 29245 54247 29279
rect 54247 29245 54256 29279
rect 54204 29236 54256 29245
rect 54204 29025 54256 29034
rect 54204 28991 54213 29025
rect 54213 28991 54247 29025
rect 54247 28991 54256 29025
rect 54204 28982 54256 28991
rect 11772 28805 11824 28814
rect 11772 28771 11781 28805
rect 11781 28771 11815 28805
rect 11815 28771 11824 28805
rect 11772 28762 11824 28771
rect 11772 28709 11824 28718
rect 11772 28675 11781 28709
rect 11781 28675 11815 28709
rect 11815 28675 11824 28709
rect 11772 28666 11824 28675
rect 54204 28489 54256 28498
rect 54204 28455 54213 28489
rect 54213 28455 54247 28489
rect 54247 28455 54256 28489
rect 54204 28446 54256 28455
rect 54204 28235 54256 28244
rect 54204 28201 54213 28235
rect 54213 28201 54247 28235
rect 54247 28201 54256 28235
rect 54204 28192 54256 28201
rect 11772 28015 11824 28024
rect 11772 27981 11781 28015
rect 11781 27981 11815 28015
rect 11815 27981 11824 28015
rect 11772 27972 11824 27981
rect 11772 27919 11824 27928
rect 11772 27885 11781 27919
rect 11781 27885 11815 27919
rect 11815 27885 11824 27919
rect 11772 27876 11824 27885
rect 54204 27699 54256 27708
rect 54204 27665 54213 27699
rect 54213 27665 54247 27699
rect 54247 27665 54256 27699
rect 54204 27656 54256 27665
rect 54204 27445 54256 27454
rect 54204 27411 54213 27445
rect 54213 27411 54247 27445
rect 54247 27411 54256 27445
rect 54204 27402 54256 27411
rect 11772 27225 11824 27234
rect 11772 27191 11781 27225
rect 11781 27191 11815 27225
rect 11815 27191 11824 27225
rect 11772 27182 11824 27191
rect 11772 27129 11824 27138
rect 11772 27095 11781 27129
rect 11781 27095 11815 27129
rect 11815 27095 11824 27129
rect 11772 27086 11824 27095
rect 54204 26909 54256 26918
rect 54204 26875 54213 26909
rect 54213 26875 54247 26909
rect 54247 26875 54256 26909
rect 54204 26866 54256 26875
rect 54204 26655 54256 26664
rect 54204 26621 54213 26655
rect 54213 26621 54247 26655
rect 54247 26621 54256 26655
rect 54204 26612 54256 26621
rect 11772 26435 11824 26444
rect 11772 26401 11781 26435
rect 11781 26401 11815 26435
rect 11815 26401 11824 26435
rect 11772 26392 11824 26401
rect 11772 26339 11824 26348
rect 11772 26305 11781 26339
rect 11781 26305 11815 26339
rect 11815 26305 11824 26339
rect 11772 26296 11824 26305
rect 54204 26119 54256 26128
rect 54204 26085 54213 26119
rect 54213 26085 54247 26119
rect 54247 26085 54256 26119
rect 54204 26076 54256 26085
rect 54204 25865 54256 25874
rect 54204 25831 54213 25865
rect 54213 25831 54247 25865
rect 54247 25831 54256 25865
rect 54204 25822 54256 25831
rect 11772 25645 11824 25654
rect 11772 25611 11781 25645
rect 11781 25611 11815 25645
rect 11815 25611 11824 25645
rect 11772 25602 11824 25611
rect 11772 25549 11824 25558
rect 11772 25515 11781 25549
rect 11781 25515 11815 25549
rect 11815 25515 11824 25549
rect 11772 25506 11824 25515
rect 54204 25329 54256 25338
rect 54204 25295 54213 25329
rect 54213 25295 54247 25329
rect 54247 25295 54256 25329
rect 54204 25286 54256 25295
rect 54204 25075 54256 25084
rect 54204 25041 54213 25075
rect 54213 25041 54247 25075
rect 54247 25041 54256 25075
rect 54204 25032 54256 25041
rect 11772 24855 11824 24864
rect 11772 24821 11781 24855
rect 11781 24821 11815 24855
rect 11815 24821 11824 24855
rect 11772 24812 11824 24821
rect 11772 24759 11824 24768
rect 11772 24725 11781 24759
rect 11781 24725 11815 24759
rect 11815 24725 11824 24759
rect 11772 24716 11824 24725
rect 54204 24539 54256 24548
rect 54204 24505 54213 24539
rect 54213 24505 54247 24539
rect 54247 24505 54256 24539
rect 54204 24496 54256 24505
rect 54204 24285 54256 24294
rect 54204 24251 54213 24285
rect 54213 24251 54247 24285
rect 54247 24251 54256 24285
rect 54204 24242 54256 24251
rect 11772 24065 11824 24074
rect 11772 24031 11781 24065
rect 11781 24031 11815 24065
rect 11815 24031 11824 24065
rect 11772 24022 11824 24031
rect 11772 23969 11824 23978
rect 11772 23935 11781 23969
rect 11781 23935 11815 23969
rect 11815 23935 11824 23969
rect 11772 23926 11824 23935
rect 54204 23749 54256 23758
rect 54204 23715 54213 23749
rect 54213 23715 54247 23749
rect 54247 23715 54256 23749
rect 54204 23706 54256 23715
rect 54204 23495 54256 23504
rect 54204 23461 54213 23495
rect 54213 23461 54247 23495
rect 54247 23461 54256 23495
rect 54204 23452 54256 23461
rect 11772 23275 11824 23284
rect 11772 23241 11781 23275
rect 11781 23241 11815 23275
rect 11815 23241 11824 23275
rect 11772 23232 11824 23241
rect 11772 23179 11824 23188
rect 11772 23145 11781 23179
rect 11781 23145 11815 23179
rect 11815 23145 11824 23179
rect 11772 23136 11824 23145
rect 54204 22959 54256 22968
rect 54204 22925 54213 22959
rect 54213 22925 54247 22959
rect 54247 22925 54256 22959
rect 54204 22916 54256 22925
rect 54204 22705 54256 22714
rect 54204 22671 54213 22705
rect 54213 22671 54247 22705
rect 54247 22671 54256 22705
rect 54204 22662 54256 22671
rect 11772 22485 11824 22494
rect 11772 22451 11781 22485
rect 11781 22451 11815 22485
rect 11815 22451 11824 22485
rect 11772 22442 11824 22451
rect 11772 22389 11824 22398
rect 11772 22355 11781 22389
rect 11781 22355 11815 22389
rect 11815 22355 11824 22389
rect 11772 22346 11824 22355
rect 54204 22169 54256 22178
rect 54204 22135 54213 22169
rect 54213 22135 54247 22169
rect 54247 22135 54256 22169
rect 54204 22126 54256 22135
rect 54204 21915 54256 21924
rect 54204 21881 54213 21915
rect 54213 21881 54247 21915
rect 54247 21881 54256 21915
rect 54204 21872 54256 21881
rect 11772 21695 11824 21704
rect 11772 21661 11781 21695
rect 11781 21661 11815 21695
rect 11815 21661 11824 21695
rect 11772 21652 11824 21661
rect 11772 21599 11824 21608
rect 11772 21565 11781 21599
rect 11781 21565 11815 21599
rect 11815 21565 11824 21599
rect 11772 21556 11824 21565
rect 54204 21379 54256 21388
rect 54204 21345 54213 21379
rect 54213 21345 54247 21379
rect 54247 21345 54256 21379
rect 54204 21336 54256 21345
rect 54204 21125 54256 21134
rect 54204 21091 54213 21125
rect 54213 21091 54247 21125
rect 54247 21091 54256 21125
rect 54204 21082 54256 21091
rect 11772 20905 11824 20914
rect 11772 20871 11781 20905
rect 11781 20871 11815 20905
rect 11815 20871 11824 20905
rect 11772 20862 11824 20871
rect 11772 20809 11824 20818
rect 11772 20775 11781 20809
rect 11781 20775 11815 20809
rect 11815 20775 11824 20809
rect 11772 20766 11824 20775
rect 54204 20589 54256 20598
rect 54204 20555 54213 20589
rect 54213 20555 54247 20589
rect 54247 20555 54256 20589
rect 54204 20546 54256 20555
rect 54204 20335 54256 20344
rect 54204 20301 54213 20335
rect 54213 20301 54247 20335
rect 54247 20301 54256 20335
rect 54204 20292 54256 20301
rect 11772 20115 11824 20124
rect 11772 20081 11781 20115
rect 11781 20081 11815 20115
rect 11815 20081 11824 20115
rect 11772 20072 11824 20081
rect 11772 20019 11824 20028
rect 11772 19985 11781 20019
rect 11781 19985 11815 20019
rect 11815 19985 11824 20019
rect 11772 19976 11824 19985
rect 54204 19799 54256 19808
rect 54204 19765 54213 19799
rect 54213 19765 54247 19799
rect 54247 19765 54256 19799
rect 54204 19756 54256 19765
rect 54204 19545 54256 19554
rect 54204 19511 54213 19545
rect 54213 19511 54247 19545
rect 54247 19511 54256 19545
rect 54204 19502 54256 19511
rect 11772 19325 11824 19334
rect 11772 19291 11781 19325
rect 11781 19291 11815 19325
rect 11815 19291 11824 19325
rect 11772 19282 11824 19291
rect 11772 19229 11824 19238
rect 11772 19195 11781 19229
rect 11781 19195 11815 19229
rect 11815 19195 11824 19229
rect 11772 19186 11824 19195
rect 54204 19009 54256 19018
rect 54204 18975 54213 19009
rect 54213 18975 54247 19009
rect 54247 18975 54256 19009
rect 54204 18966 54256 18975
rect 54204 18755 54256 18764
rect 54204 18721 54213 18755
rect 54213 18721 54247 18755
rect 54247 18721 54256 18755
rect 54204 18712 54256 18721
rect 11772 18535 11824 18544
rect 11772 18501 11781 18535
rect 11781 18501 11815 18535
rect 11815 18501 11824 18535
rect 11772 18492 11824 18501
rect 11772 18439 11824 18448
rect 11772 18405 11781 18439
rect 11781 18405 11815 18439
rect 11815 18405 11824 18439
rect 11772 18396 11824 18405
rect 54204 18219 54256 18228
rect 54204 18185 54213 18219
rect 54213 18185 54247 18219
rect 54247 18185 54256 18219
rect 54204 18176 54256 18185
rect 54204 17965 54256 17974
rect 54204 17931 54213 17965
rect 54213 17931 54247 17965
rect 54247 17931 54256 17965
rect 54204 17922 54256 17931
rect 11772 17745 11824 17754
rect 11772 17711 11781 17745
rect 11781 17711 11815 17745
rect 11815 17711 11824 17745
rect 11772 17702 11824 17711
rect 11772 17649 11824 17658
rect 11772 17615 11781 17649
rect 11781 17615 11815 17649
rect 11815 17615 11824 17649
rect 11772 17606 11824 17615
rect 54204 17429 54256 17438
rect 54204 17395 54213 17429
rect 54213 17395 54247 17429
rect 54247 17395 54256 17429
rect 54204 17386 54256 17395
rect 54204 17175 54256 17184
rect 54204 17141 54213 17175
rect 54213 17141 54247 17175
rect 54247 17141 54256 17175
rect 54204 17132 54256 17141
rect 11772 16955 11824 16964
rect 11772 16921 11781 16955
rect 11781 16921 11815 16955
rect 11815 16921 11824 16955
rect 11772 16912 11824 16921
rect 11772 16859 11824 16868
rect 11772 16825 11781 16859
rect 11781 16825 11815 16859
rect 11815 16825 11824 16859
rect 11772 16816 11824 16825
rect 54204 16639 54256 16648
rect 54204 16605 54213 16639
rect 54213 16605 54247 16639
rect 54247 16605 54256 16639
rect 54204 16596 54256 16605
rect 54204 16385 54256 16394
rect 54204 16351 54213 16385
rect 54213 16351 54247 16385
rect 54247 16351 54256 16385
rect 54204 16342 54256 16351
rect 11772 16165 11824 16174
rect 11772 16131 11781 16165
rect 11781 16131 11815 16165
rect 11815 16131 11824 16165
rect 11772 16122 11824 16131
rect 11772 16069 11824 16078
rect 11772 16035 11781 16069
rect 11781 16035 11815 16069
rect 11815 16035 11824 16069
rect 11772 16026 11824 16035
rect 54204 15849 54256 15858
rect 54204 15815 54213 15849
rect 54213 15815 54247 15849
rect 54247 15815 54256 15849
rect 54204 15806 54256 15815
rect 54204 15595 54256 15604
rect 54204 15561 54213 15595
rect 54213 15561 54247 15595
rect 54247 15561 54256 15595
rect 54204 15552 54256 15561
rect 11772 15375 11824 15384
rect 11772 15341 11781 15375
rect 11781 15341 11815 15375
rect 11815 15341 11824 15375
rect 11772 15332 11824 15341
rect 11772 15279 11824 15288
rect 11772 15245 11781 15279
rect 11781 15245 11815 15279
rect 11815 15245 11824 15279
rect 11772 15236 11824 15245
rect 54204 15059 54256 15068
rect 54204 15025 54213 15059
rect 54213 15025 54247 15059
rect 54247 15025 54256 15059
rect 54204 15016 54256 15025
rect 54204 14805 54256 14814
rect 54204 14771 54213 14805
rect 54213 14771 54247 14805
rect 54247 14771 54256 14805
rect 54204 14762 54256 14771
rect 11772 14585 11824 14594
rect 11772 14551 11781 14585
rect 11781 14551 11815 14585
rect 11815 14551 11824 14585
rect 11772 14542 11824 14551
rect 11772 14489 11824 14498
rect 11772 14455 11781 14489
rect 11781 14455 11815 14489
rect 11815 14455 11824 14489
rect 11772 14446 11824 14455
rect 54204 14269 54256 14278
rect 54204 14235 54213 14269
rect 54213 14235 54247 14269
rect 54247 14235 54256 14269
rect 54204 14226 54256 14235
rect 54204 14015 54256 14024
rect 54204 13981 54213 14015
rect 54213 13981 54247 14015
rect 54247 13981 54256 14015
rect 54204 13972 54256 13981
rect 11772 13795 11824 13804
rect 11772 13761 11781 13795
rect 11781 13761 11815 13795
rect 11815 13761 11824 13795
rect 11772 13752 11824 13761
rect 11772 13699 11824 13708
rect 11772 13665 11781 13699
rect 11781 13665 11815 13699
rect 11815 13665 11824 13699
rect 11772 13656 11824 13665
rect 54204 13479 54256 13488
rect 54204 13445 54213 13479
rect 54213 13445 54247 13479
rect 54247 13445 54256 13479
rect 54204 13436 54256 13445
rect 54204 13225 54256 13234
rect 54204 13191 54213 13225
rect 54213 13191 54247 13225
rect 54247 13191 54256 13225
rect 54204 13182 54256 13191
rect 11772 13005 11824 13014
rect 11772 12971 11781 13005
rect 11781 12971 11815 13005
rect 11815 12971 11824 13005
rect 11772 12962 11824 12971
rect 11772 12909 11824 12918
rect 11772 12875 11781 12909
rect 11781 12875 11815 12909
rect 11815 12875 11824 12909
rect 11772 12866 11824 12875
rect 54204 12689 54256 12698
rect 54204 12655 54213 12689
rect 54213 12655 54247 12689
rect 54247 12655 54256 12689
rect 54204 12646 54256 12655
rect 54204 12435 54256 12444
rect 54204 12401 54213 12435
rect 54213 12401 54247 12435
rect 54247 12401 54256 12435
rect 54204 12392 54256 12401
rect 11772 12215 11824 12224
rect 11772 12181 11781 12215
rect 11781 12181 11815 12215
rect 11815 12181 11824 12215
rect 11772 12172 11824 12181
rect 11772 12119 11824 12128
rect 11772 12085 11781 12119
rect 11781 12085 11815 12119
rect 11815 12085 11824 12119
rect 11772 12076 11824 12085
rect 54204 11899 54256 11908
rect 54204 11865 54213 11899
rect 54213 11865 54247 11899
rect 54247 11865 54256 11899
rect 54204 11856 54256 11865
rect 54204 11645 54256 11654
rect 54204 11611 54213 11645
rect 54213 11611 54247 11645
rect 54247 11611 54256 11645
rect 54204 11602 54256 11611
rect 11772 11425 11824 11434
rect 11772 11391 11781 11425
rect 11781 11391 11815 11425
rect 11815 11391 11824 11425
rect 11772 11382 11824 11391
rect 11772 11329 11824 11338
rect 11772 11295 11781 11329
rect 11781 11295 11815 11329
rect 11815 11295 11824 11329
rect 11772 11286 11824 11295
rect 54204 11109 54256 11118
rect 54204 11075 54213 11109
rect 54213 11075 54247 11109
rect 54247 11075 54256 11109
rect 54204 11066 54256 11075
rect 54204 10855 54256 10864
rect 54204 10821 54213 10855
rect 54213 10821 54247 10855
rect 54247 10821 54256 10855
rect 54204 10812 54256 10821
rect 11772 10635 11824 10644
rect 11772 10601 11781 10635
rect 11781 10601 11815 10635
rect 11815 10601 11824 10635
rect 11772 10592 11824 10601
rect 11772 10539 11824 10548
rect 11772 10505 11781 10539
rect 11781 10505 11815 10539
rect 11815 10505 11824 10539
rect 11772 10496 11824 10505
rect 54204 10319 54256 10328
rect 54204 10285 54213 10319
rect 54213 10285 54247 10319
rect 54247 10285 54256 10319
rect 54204 10276 54256 10285
rect 7570 9645 7622 9697
rect 11538 9645 11590 9697
rect 12940 8229 12992 8281
rect 6462 7634 6514 7643
rect 6462 7600 6471 7634
rect 6471 7600 6505 7634
rect 6505 7600 6514 7634
rect 6462 7591 6514 7600
rect 6462 6220 6514 6229
rect 6462 6186 6471 6220
rect 6471 6186 6505 6220
rect 6505 6186 6514 6220
rect 6462 6177 6514 6186
rect 6462 4806 6514 4815
rect 6462 4772 6471 4806
rect 6471 4772 6505 4806
rect 6505 4772 6514 4806
rect 6462 4763 6514 4772
<< metal2 >>
rect 53034 62683 53090 62692
rect 53034 62618 53090 62627
rect 54354 61271 54382 67359
rect 54478 62543 54506 67359
rect 54602 65118 54630 67359
rect 59388 66149 59444 66158
rect 59388 66084 59444 66093
rect 54588 65109 54644 65118
rect 54588 65044 54644 65053
rect 54464 62534 54520 62543
rect 54464 62469 54520 62478
rect 54342 61265 54394 61271
rect 54342 61207 54394 61213
rect 54354 60876 54382 61207
rect 54478 60895 54506 62469
rect 54602 60895 54630 65044
rect 59388 64735 59444 64744
rect 59388 64670 59444 64679
rect 59388 63321 59444 63330
rect 59388 63256 59444 63265
rect 58406 61265 58458 61271
rect 58406 61207 58458 61213
rect 33014 60848 54382 60876
rect 58418 60735 58446 61207
rect 54198 60582 54204 60634
rect 54256 60582 54262 60634
rect 11766 60362 11772 60414
rect 11824 60362 11830 60414
rect 11766 60266 11772 60318
rect 11824 60266 11830 60318
rect 54198 60046 54204 60098
rect 54256 60046 54262 60098
rect 54198 59792 54204 59844
rect 54256 59792 54262 59844
rect 11766 59572 11772 59624
rect 11824 59572 11830 59624
rect 11766 59476 11772 59528
rect 11824 59476 11830 59528
rect 54198 59256 54204 59308
rect 54256 59256 54262 59308
rect 54198 59002 54204 59054
rect 54256 59002 54262 59054
rect 11766 58782 11772 58834
rect 11824 58782 11830 58834
rect 11766 58686 11772 58738
rect 11824 58686 11830 58738
rect 54198 58466 54204 58518
rect 54256 58466 54262 58518
rect 54198 58212 54204 58264
rect 54256 58212 54262 58264
rect 11766 57992 11772 58044
rect 11824 57992 11830 58044
rect 11766 57896 11772 57948
rect 11824 57896 11830 57948
rect 54198 57676 54204 57728
rect 54256 57676 54262 57728
rect 54198 57422 54204 57474
rect 54256 57422 54262 57474
rect 11766 57202 11772 57254
rect 11824 57202 11830 57254
rect 11766 57106 11772 57158
rect 11824 57106 11830 57158
rect 54198 56886 54204 56938
rect 54256 56886 54262 56938
rect 54198 56632 54204 56684
rect 54256 56632 54262 56684
rect 11766 56412 11772 56464
rect 11824 56412 11830 56464
rect 11766 56316 11772 56368
rect 11824 56316 11830 56368
rect 54198 56096 54204 56148
rect 54256 56096 54262 56148
rect 54198 55842 54204 55894
rect 54256 55842 54262 55894
rect 11766 55622 11772 55674
rect 11824 55622 11830 55674
rect 11766 55526 11772 55578
rect 11824 55526 11830 55578
rect 54198 55306 54204 55358
rect 54256 55306 54262 55358
rect 54198 55052 54204 55104
rect 54256 55052 54262 55104
rect 11766 54832 11772 54884
rect 11824 54832 11830 54884
rect 11766 54736 11772 54788
rect 11824 54736 11830 54788
rect 54198 54516 54204 54568
rect 54256 54516 54262 54568
rect 54198 54262 54204 54314
rect 54256 54262 54262 54314
rect 11766 54042 11772 54094
rect 11824 54042 11830 54094
rect 11766 53946 11772 53998
rect 11824 53946 11830 53998
rect 54198 53726 54204 53778
rect 54256 53726 54262 53778
rect 54198 53472 54204 53524
rect 54256 53472 54262 53524
rect 11766 53252 11772 53304
rect 11824 53252 11830 53304
rect 11766 53156 11772 53208
rect 11824 53156 11830 53208
rect 54198 52936 54204 52988
rect 54256 52936 54262 52988
rect 54198 52682 54204 52734
rect 54256 52682 54262 52734
rect 11766 52462 11772 52514
rect 11824 52462 11830 52514
rect 11766 52366 11772 52418
rect 11824 52366 11830 52418
rect 54198 52146 54204 52198
rect 54256 52146 54262 52198
rect 54198 51892 54204 51944
rect 54256 51892 54262 51944
rect 11766 51672 11772 51724
rect 11824 51672 11830 51724
rect 11766 51576 11772 51628
rect 11824 51576 11830 51628
rect 54198 51356 54204 51408
rect 54256 51356 54262 51408
rect 54198 51102 54204 51154
rect 54256 51102 54262 51154
rect 11766 50882 11772 50934
rect 11824 50882 11830 50934
rect 11766 50786 11772 50838
rect 11824 50786 11830 50838
rect 54198 50566 54204 50618
rect 54256 50566 54262 50618
rect 54198 50312 54204 50364
rect 54256 50312 54262 50364
rect 11766 50092 11772 50144
rect 11824 50092 11830 50144
rect 11766 49996 11772 50048
rect 11824 49996 11830 50048
rect 54198 49776 54204 49828
rect 54256 49776 54262 49828
rect 54198 49522 54204 49574
rect 54256 49522 54262 49574
rect 11766 49302 11772 49354
rect 11824 49302 11830 49354
rect 11766 49206 11772 49258
rect 11824 49206 11830 49258
rect 54198 48986 54204 49038
rect 54256 48986 54262 49038
rect 54198 48732 54204 48784
rect 54256 48732 54262 48784
rect 11766 48512 11772 48564
rect 11824 48512 11830 48564
rect 11766 48416 11772 48468
rect 11824 48416 11830 48468
rect 54198 48196 54204 48248
rect 54256 48196 54262 48248
rect 54198 47942 54204 47994
rect 54256 47942 54262 47994
rect 11766 47722 11772 47774
rect 11824 47722 11830 47774
rect 11766 47626 11772 47678
rect 11824 47626 11830 47678
rect 54198 47406 54204 47458
rect 54256 47406 54262 47458
rect 54198 47152 54204 47204
rect 54256 47152 54262 47204
rect 11766 46932 11772 46984
rect 11824 46932 11830 46984
rect 11766 46836 11772 46888
rect 11824 46836 11830 46888
rect 54198 46616 54204 46668
rect 54256 46616 54262 46668
rect 54198 46362 54204 46414
rect 54256 46362 54262 46414
rect 11766 46142 11772 46194
rect 11824 46142 11830 46194
rect 11766 46046 11772 46098
rect 11824 46046 11830 46098
rect 54198 45826 54204 45878
rect 54256 45826 54262 45878
rect 54198 45572 54204 45624
rect 54256 45572 54262 45624
rect 11766 45352 11772 45404
rect 11824 45352 11830 45404
rect 11766 45256 11772 45308
rect 11824 45256 11830 45308
rect 54198 45036 54204 45088
rect 54256 45036 54262 45088
rect 54198 44782 54204 44834
rect 54256 44782 54262 44834
rect 11766 44562 11772 44614
rect 11824 44562 11830 44614
rect 11766 44466 11772 44518
rect 11824 44466 11830 44518
rect 54198 44246 54204 44298
rect 54256 44246 54262 44298
rect 54198 43992 54204 44044
rect 54256 43992 54262 44044
rect 11766 43772 11772 43824
rect 11824 43772 11830 43824
rect 11766 43676 11772 43728
rect 11824 43676 11830 43728
rect 54198 43456 54204 43508
rect 54256 43456 54262 43508
rect 54198 43202 54204 43254
rect 54256 43202 54262 43254
rect 11766 42982 11772 43034
rect 11824 42982 11830 43034
rect 11766 42886 11772 42938
rect 11824 42886 11830 42938
rect 54198 42666 54204 42718
rect 54256 42666 54262 42718
rect 54198 42412 54204 42464
rect 54256 42412 54262 42464
rect 11766 42192 11772 42244
rect 11824 42192 11830 42244
rect 11766 42096 11772 42148
rect 11824 42096 11830 42148
rect 54198 41876 54204 41928
rect 54256 41876 54262 41928
rect 54198 41622 54204 41674
rect 54256 41622 54262 41674
rect 11766 41402 11772 41454
rect 11824 41402 11830 41454
rect 11766 41306 11772 41358
rect 11824 41306 11830 41358
rect 54198 41086 54204 41138
rect 54256 41086 54262 41138
rect 54198 40832 54204 40884
rect 54256 40832 54262 40884
rect 11766 40612 11772 40664
rect 11824 40612 11830 40664
rect 11766 40516 11772 40568
rect 11824 40516 11830 40568
rect 54198 40296 54204 40348
rect 54256 40296 54262 40348
rect 54198 40042 54204 40094
rect 54256 40042 54262 40094
rect 11766 39822 11772 39874
rect 11824 39822 11830 39874
rect 11766 39726 11772 39778
rect 11824 39726 11830 39778
rect 54198 39506 54204 39558
rect 54256 39506 54262 39558
rect 54198 39252 54204 39304
rect 54256 39252 54262 39304
rect 11766 39032 11772 39084
rect 11824 39032 11830 39084
rect 11766 38936 11772 38988
rect 11824 38936 11830 38988
rect 54198 38716 54204 38768
rect 54256 38716 54262 38768
rect 54198 38462 54204 38514
rect 54256 38462 54262 38514
rect 11766 38242 11772 38294
rect 11824 38242 11830 38294
rect 11766 38146 11772 38198
rect 11824 38146 11830 38198
rect 54198 37926 54204 37978
rect 54256 37926 54262 37978
rect 54198 37672 54204 37724
rect 54256 37672 54262 37724
rect 11766 37452 11772 37504
rect 11824 37452 11830 37504
rect 11766 37356 11772 37408
rect 11824 37356 11830 37408
rect 54198 37136 54204 37188
rect 54256 37136 54262 37188
rect 54198 36882 54204 36934
rect 54256 36882 54262 36934
rect 11766 36662 11772 36714
rect 11824 36662 11830 36714
rect 11766 36566 11772 36618
rect 11824 36566 11830 36618
rect 54198 36346 54204 36398
rect 54256 36346 54262 36398
rect 54198 36092 54204 36144
rect 54256 36092 54262 36144
rect 11766 35872 11772 35924
rect 11824 35872 11830 35924
rect 11766 35776 11772 35828
rect 11824 35776 11830 35828
rect 54198 35556 54204 35608
rect 54256 35556 54262 35608
rect 54198 35302 54204 35354
rect 54256 35302 54262 35354
rect 11766 35082 11772 35134
rect 11824 35082 11830 35134
rect 11766 34986 11772 35038
rect 11824 34986 11830 35038
rect 54198 34766 54204 34818
rect 54256 34766 54262 34818
rect 54198 34512 54204 34564
rect 54256 34512 54262 34564
rect 11766 34292 11772 34344
rect 11824 34292 11830 34344
rect 11766 34196 11772 34248
rect 11824 34196 11830 34248
rect 54198 33976 54204 34028
rect 54256 33976 54262 34028
rect 54198 33722 54204 33774
rect 54256 33722 54262 33774
rect 11766 33502 11772 33554
rect 11824 33502 11830 33554
rect 11766 33406 11772 33458
rect 11824 33406 11830 33458
rect 54198 33186 54204 33238
rect 54256 33186 54262 33238
rect 54198 32932 54204 32984
rect 54256 32932 54262 32984
rect 11766 32712 11772 32764
rect 11824 32712 11830 32764
rect 11766 32616 11772 32668
rect 11824 32616 11830 32668
rect 54198 32396 54204 32448
rect 54256 32396 54262 32448
rect 54198 32142 54204 32194
rect 54256 32142 54262 32194
rect 11766 31922 11772 31974
rect 11824 31922 11830 31974
rect 11766 31826 11772 31878
rect 11824 31826 11830 31878
rect 54198 31606 54204 31658
rect 54256 31606 54262 31658
rect 54198 31352 54204 31404
rect 54256 31352 54262 31404
rect 11766 31132 11772 31184
rect 11824 31132 11830 31184
rect 11766 31036 11772 31088
rect 11824 31036 11830 31088
rect 54198 30816 54204 30868
rect 54256 30816 54262 30868
rect 54198 30562 54204 30614
rect 54256 30562 54262 30614
rect 11766 30342 11772 30394
rect 11824 30342 11830 30394
rect 11766 30246 11772 30298
rect 11824 30246 11830 30298
rect 54198 30026 54204 30078
rect 54256 30026 54262 30078
rect 54198 29772 54204 29824
rect 54256 29772 54262 29824
rect 11766 29552 11772 29604
rect 11824 29552 11830 29604
rect 11766 29456 11772 29508
rect 11824 29456 11830 29508
rect 54198 29236 54204 29288
rect 54256 29236 54262 29288
rect 54198 28982 54204 29034
rect 54256 28982 54262 29034
rect 11766 28762 11772 28814
rect 11824 28762 11830 28814
rect 11766 28666 11772 28718
rect 11824 28666 11830 28718
rect 54198 28446 54204 28498
rect 54256 28446 54262 28498
rect 54198 28192 54204 28244
rect 54256 28192 54262 28244
rect 11766 27972 11772 28024
rect 11824 27972 11830 28024
rect 11766 27876 11772 27928
rect 11824 27876 11830 27928
rect 54198 27656 54204 27708
rect 54256 27656 54262 27708
rect 54198 27402 54204 27454
rect 54256 27402 54262 27454
rect 11766 27182 11772 27234
rect 11824 27182 11830 27234
rect 11766 27086 11772 27138
rect 11824 27086 11830 27138
rect 54198 26866 54204 26918
rect 54256 26866 54262 26918
rect 54198 26612 54204 26664
rect 54256 26612 54262 26664
rect 11766 26392 11772 26444
rect 11824 26392 11830 26444
rect 11766 26296 11772 26348
rect 11824 26296 11830 26348
rect 54198 26076 54204 26128
rect 54256 26076 54262 26128
rect 54198 25822 54204 25874
rect 54256 25822 54262 25874
rect 11766 25602 11772 25654
rect 11824 25602 11830 25654
rect 11766 25506 11772 25558
rect 11824 25506 11830 25558
rect 54198 25286 54204 25338
rect 54256 25286 54262 25338
rect 54198 25032 54204 25084
rect 54256 25032 54262 25084
rect 11766 24812 11772 24864
rect 11824 24812 11830 24864
rect 11766 24716 11772 24768
rect 11824 24716 11830 24768
rect 54198 24496 54204 24548
rect 54256 24496 54262 24548
rect 54198 24242 54204 24294
rect 54256 24242 54262 24294
rect 11766 24022 11772 24074
rect 11824 24022 11830 24074
rect 11766 23926 11772 23978
rect 11824 23926 11830 23978
rect 54198 23706 54204 23758
rect 54256 23706 54262 23758
rect 54198 23452 54204 23504
rect 54256 23452 54262 23504
rect 11766 23232 11772 23284
rect 11824 23232 11830 23284
rect 11766 23136 11772 23188
rect 11824 23136 11830 23188
rect 54198 22916 54204 22968
rect 54256 22916 54262 22968
rect 54198 22662 54204 22714
rect 54256 22662 54262 22714
rect 11766 22442 11772 22494
rect 11824 22442 11830 22494
rect 11766 22346 11772 22398
rect 11824 22346 11830 22398
rect 54198 22126 54204 22178
rect 54256 22126 54262 22178
rect 54198 21872 54204 21924
rect 54256 21872 54262 21924
rect 11766 21652 11772 21704
rect 11824 21652 11830 21704
rect 11766 21556 11772 21608
rect 11824 21556 11830 21608
rect 54198 21336 54204 21388
rect 54256 21336 54262 21388
rect 54198 21082 54204 21134
rect 54256 21082 54262 21134
rect 11766 20862 11772 20914
rect 11824 20862 11830 20914
rect 11766 20766 11772 20818
rect 11824 20766 11830 20818
rect 54198 20546 54204 20598
rect 54256 20546 54262 20598
rect 54198 20292 54204 20344
rect 54256 20292 54262 20344
rect 11766 20072 11772 20124
rect 11824 20072 11830 20124
rect 11766 19976 11772 20028
rect 11824 19976 11830 20028
rect 54198 19756 54204 19808
rect 54256 19756 54262 19808
rect 54198 19502 54204 19554
rect 54256 19502 54262 19554
rect 11766 19282 11772 19334
rect 11824 19282 11830 19334
rect 11766 19186 11772 19238
rect 11824 19186 11830 19238
rect 54198 18966 54204 19018
rect 54256 18966 54262 19018
rect 54198 18712 54204 18764
rect 54256 18712 54262 18764
rect 11766 18492 11772 18544
rect 11824 18492 11830 18544
rect 11766 18396 11772 18448
rect 11824 18396 11830 18448
rect 54198 18176 54204 18228
rect 54256 18176 54262 18228
rect 54198 17922 54204 17974
rect 54256 17922 54262 17974
rect 11766 17702 11772 17754
rect 11824 17702 11830 17754
rect 11766 17606 11772 17658
rect 11824 17606 11830 17658
rect 54198 17386 54204 17438
rect 54256 17386 54262 17438
rect 54198 17132 54204 17184
rect 54256 17132 54262 17184
rect 11766 16912 11772 16964
rect 11824 16912 11830 16964
rect 11766 16816 11772 16868
rect 11824 16816 11830 16868
rect 54198 16596 54204 16648
rect 54256 16596 54262 16648
rect 54198 16342 54204 16394
rect 54256 16342 54262 16394
rect 11766 16122 11772 16174
rect 11824 16122 11830 16174
rect 11766 16026 11772 16078
rect 11824 16026 11830 16078
rect 54198 15806 54204 15858
rect 54256 15806 54262 15858
rect 54198 15552 54204 15604
rect 54256 15552 54262 15604
rect 11766 15332 11772 15384
rect 11824 15332 11830 15384
rect 11766 15236 11772 15288
rect 11824 15236 11830 15288
rect 54198 15016 54204 15068
rect 54256 15016 54262 15068
rect 54198 14762 54204 14814
rect 54256 14762 54262 14814
rect 11766 14542 11772 14594
rect 11824 14542 11830 14594
rect 11766 14446 11772 14498
rect 11824 14446 11830 14498
rect 54198 14226 54204 14278
rect 54256 14226 54262 14278
rect 54198 13972 54204 14024
rect 54256 13972 54262 14024
rect 11766 13752 11772 13804
rect 11824 13752 11830 13804
rect 11766 13656 11772 13708
rect 11824 13656 11830 13708
rect 54198 13436 54204 13488
rect 54256 13436 54262 13488
rect 54198 13182 54204 13234
rect 54256 13182 54262 13234
rect 11766 12962 11772 13014
rect 11824 12962 11830 13014
rect 11766 12866 11772 12918
rect 11824 12866 11830 12918
rect 54198 12646 54204 12698
rect 54256 12646 54262 12698
rect 54198 12392 54204 12444
rect 54256 12392 54262 12444
rect 11766 12172 11772 12224
rect 11824 12172 11830 12224
rect 11766 12076 11772 12128
rect 11824 12076 11830 12128
rect 54198 11856 54204 11908
rect 54256 11856 54262 11908
rect 54198 11602 54204 11654
rect 54256 11602 54262 11654
rect 11766 11382 11772 11434
rect 11824 11382 11830 11434
rect 11766 11286 11772 11338
rect 11824 11286 11830 11338
rect 54198 11066 54204 11118
rect 54256 11066 54262 11118
rect 54198 10812 54204 10864
rect 54256 10812 54262 10864
rect 11766 10592 11772 10644
rect 11824 10592 11830 10644
rect 11766 10496 11772 10548
rect 11824 10496 11830 10548
rect 54198 10276 54204 10328
rect 54256 10276 54262 10328
rect 7582 9703 7610 10175
rect 7570 9697 7622 9703
rect 7570 9639 7622 9645
rect 6460 7645 6516 7654
rect 6460 7580 6516 7589
rect 6460 6231 6516 6240
rect 6460 6166 6516 6175
rect 11178 5866 11206 10015
rect 11164 5857 11220 5866
rect 11164 5792 11220 5801
rect 6460 4817 6516 4826
rect 6460 4752 6516 4761
rect 11178 0 11206 5792
rect 11302 555 11330 10015
rect 11426 8441 11454 10015
rect 11550 9842 11578 10015
rect 11550 9814 33014 9842
rect 11550 9703 11578 9814
rect 11538 9697 11590 9703
rect 11538 9639 11590 9645
rect 11412 8432 11468 8441
rect 11412 8367 11468 8376
rect 11288 546 11344 555
rect 11288 481 11344 490
rect 11302 0 11330 481
rect 11426 0 11454 8367
rect 11550 0 11578 9639
rect 12938 8283 12994 8292
rect 12938 8218 12994 8227
rect 13032 256 13060 284
rect 23016 256 23044 284
rect 33000 256 33028 284
rect 42984 256 43012 284
<< via2 >>
rect 53034 62681 53090 62683
rect 53034 62629 53036 62681
rect 53036 62629 53088 62681
rect 53088 62629 53090 62681
rect 53034 62627 53090 62629
rect 59388 66147 59444 66149
rect 59388 66095 59390 66147
rect 59390 66095 59442 66147
rect 59442 66095 59444 66147
rect 59388 66093 59444 66095
rect 54588 65053 54644 65109
rect 54464 62478 54520 62534
rect 59388 64733 59444 64735
rect 59388 64681 59390 64733
rect 59390 64681 59442 64733
rect 59442 64681 59444 64733
rect 59388 64679 59444 64681
rect 59388 63319 59444 63321
rect 59388 63267 59390 63319
rect 59390 63267 59442 63319
rect 59442 63267 59444 63319
rect 59388 63265 59444 63267
rect 6460 7643 6516 7645
rect 6460 7591 6462 7643
rect 6462 7591 6514 7643
rect 6514 7591 6516 7643
rect 6460 7589 6516 7591
rect 6460 6229 6516 6231
rect 6460 6177 6462 6229
rect 6462 6177 6514 6229
rect 6514 6177 6516 6229
rect 6460 6175 6516 6177
rect 11164 5801 11220 5857
rect 6460 4815 6516 4817
rect 6460 4763 6462 4815
rect 6462 4763 6514 4815
rect 6514 4763 6516 4815
rect 6460 4761 6516 4763
rect 11412 8376 11468 8432
rect 11288 490 11344 546
rect 12938 8281 12994 8283
rect 12938 8229 12940 8281
rect 12940 8229 12992 8281
rect 12992 8229 12994 8281
rect 12938 8227 12994 8229
<< metal3 >>
rect 13378 67118 13476 67216
rect 14626 67118 14724 67216
rect 15874 67118 15972 67216
rect 17122 67118 17220 67216
rect 18370 67118 18468 67216
rect 19618 67118 19716 67216
rect 20866 67118 20964 67216
rect 22114 67118 22212 67216
rect 23362 67118 23460 67216
rect 24610 67118 24708 67216
rect 25858 67118 25956 67216
rect 27106 67118 27204 67216
rect 28354 67118 28452 67216
rect 29602 67118 29700 67216
rect 30850 67118 30948 67216
rect 32098 67118 32196 67216
rect 33346 67118 33444 67216
rect 34594 67118 34692 67216
rect 35842 67118 35940 67216
rect 37090 67118 37188 67216
rect 38338 67118 38436 67216
rect 39586 67118 39684 67216
rect 40834 67118 40932 67216
rect 42082 67118 42180 67216
rect 43330 67118 43428 67216
rect 44578 67118 44676 67216
rect 45826 67118 45924 67216
rect 47074 67118 47172 67216
rect 48322 67118 48420 67216
rect 49570 67118 49668 67216
rect 50818 67118 50916 67216
rect 52066 67118 52164 67216
rect 13378 66796 13476 66894
rect 14626 66796 14724 66894
rect 15874 66796 15972 66894
rect 17122 66796 17220 66894
rect 18370 66796 18468 66894
rect 19618 66796 19716 66894
rect 20866 66796 20964 66894
rect 22114 66796 22212 66894
rect 23362 66796 23460 66894
rect 24610 66796 24708 66894
rect 25858 66796 25956 66894
rect 27106 66796 27204 66894
rect 28354 66796 28452 66894
rect 29602 66796 29700 66894
rect 30850 66796 30948 66894
rect 32098 66796 32196 66894
rect 33346 66796 33444 66894
rect 34594 66796 34692 66894
rect 35842 66796 35940 66894
rect 37090 66796 37188 66894
rect 38338 66796 38436 66894
rect 39586 66796 39684 66894
rect 40834 66796 40932 66894
rect 42082 66796 42180 66894
rect 43330 66796 43428 66894
rect 44578 66796 44676 66894
rect 45826 66796 45924 66894
rect 47074 66796 47172 66894
rect 48322 66796 48420 66894
rect 49570 66796 49668 66894
rect 50818 66796 50916 66894
rect 52066 66796 52164 66894
rect 59367 66149 59465 66170
rect 59367 66093 59388 66149
rect 59444 66093 59465 66149
rect 59367 66072 59465 66093
rect 13366 65958 13464 66056
rect 14614 65958 14712 66056
rect 15862 65958 15960 66056
rect 17110 65958 17208 66056
rect 18358 65958 18456 66056
rect 19606 65958 19704 66056
rect 20854 65958 20952 66056
rect 22102 65958 22200 66056
rect 23350 65958 23448 66056
rect 24598 65958 24696 66056
rect 25846 65958 25944 66056
rect 27094 65958 27192 66056
rect 28342 65958 28440 66056
rect 29590 65958 29688 66056
rect 30838 65958 30936 66056
rect 32086 65958 32184 66056
rect 33334 65958 33432 66056
rect 34582 65958 34680 66056
rect 35830 65958 35928 66056
rect 37078 65958 37176 66056
rect 38326 65958 38424 66056
rect 39574 65958 39672 66056
rect 40822 65958 40920 66056
rect 42070 65958 42168 66056
rect 43318 65958 43416 66056
rect 44566 65958 44664 66056
rect 45814 65958 45912 66056
rect 47062 65958 47160 66056
rect 48310 65958 48408 66056
rect 49558 65958 49656 66056
rect 50806 65958 50904 66056
rect 52054 65958 52152 66056
rect 13448 65184 13546 65282
rect 14696 65184 14794 65282
rect 15944 65184 16042 65282
rect 17192 65184 17290 65282
rect 18440 65184 18538 65282
rect 19688 65184 19786 65282
rect 20936 65184 21034 65282
rect 22184 65184 22282 65282
rect 23432 65184 23530 65282
rect 24680 65184 24778 65282
rect 25928 65184 26026 65282
rect 27176 65184 27274 65282
rect 28424 65184 28522 65282
rect 29672 65184 29770 65282
rect 30920 65184 31018 65282
rect 32168 65184 32266 65282
rect 33416 65184 33514 65282
rect 34664 65184 34762 65282
rect 35912 65184 36010 65282
rect 37160 65184 37258 65282
rect 38408 65184 38506 65282
rect 39656 65184 39754 65282
rect 40904 65184 41002 65282
rect 42152 65184 42250 65282
rect 43400 65184 43498 65282
rect 44648 65184 44746 65282
rect 45896 65184 45994 65282
rect 47144 65184 47242 65282
rect 48392 65184 48490 65282
rect 49640 65184 49738 65282
rect 50888 65184 50986 65282
rect 52136 65184 52234 65282
rect 54583 65111 54649 65114
rect 33014 65109 54649 65111
rect 33014 65053 54588 65109
rect 54644 65053 54649 65109
rect 33014 65051 54649 65053
rect 54583 65048 54649 65051
rect 59367 64735 59465 64756
rect 59367 64679 59388 64735
rect 59444 64679 59465 64735
rect 59367 64658 59465 64679
rect 13621 63411 13719 63509
rect 14869 63411 14967 63509
rect 16117 63411 16215 63509
rect 17365 63411 17463 63509
rect 18613 63411 18711 63509
rect 19861 63411 19959 63509
rect 21109 63411 21207 63509
rect 22357 63411 22455 63509
rect 23605 63411 23703 63509
rect 24853 63411 24951 63509
rect 26101 63411 26199 63509
rect 27349 63411 27447 63509
rect 28597 63411 28695 63509
rect 29845 63411 29943 63509
rect 31093 63411 31191 63509
rect 32341 63411 32439 63509
rect 33589 63411 33687 63509
rect 34837 63411 34935 63509
rect 36085 63411 36183 63509
rect 37333 63411 37431 63509
rect 38581 63411 38679 63509
rect 39829 63411 39927 63509
rect 41077 63411 41175 63509
rect 42325 63411 42423 63509
rect 43573 63411 43671 63509
rect 44821 63411 44919 63509
rect 46069 63411 46167 63509
rect 47317 63411 47415 63509
rect 48565 63411 48663 63509
rect 49813 63411 49911 63509
rect 51061 63411 51159 63509
rect 52309 63411 52407 63509
rect 59367 63321 59465 63342
rect 59367 63265 59388 63321
rect 59444 63265 59465 63321
rect 59367 63244 59465 63265
rect 53029 62685 53095 62688
rect 53029 62683 66112 62685
rect 53029 62627 53034 62683
rect 53090 62627 66112 62683
rect 53029 62625 66112 62627
rect 53029 62622 53095 62625
rect 54459 62536 54525 62539
rect 33326 62534 54525 62536
rect 33326 62478 54464 62534
rect 54520 62478 54525 62534
rect 33326 62476 54525 62478
rect 54459 62473 54525 62476
rect 13190 61838 13288 61936
rect 14052 61838 14150 61936
rect 14438 61838 14536 61936
rect 15300 61838 15398 61936
rect 15686 61838 15784 61936
rect 16548 61838 16646 61936
rect 16934 61838 17032 61936
rect 17796 61838 17894 61936
rect 18182 61838 18280 61936
rect 19044 61838 19142 61936
rect 19430 61838 19528 61936
rect 20292 61838 20390 61936
rect 20678 61838 20776 61936
rect 21540 61838 21638 61936
rect 21926 61838 22024 61936
rect 22788 61838 22886 61936
rect 23174 61838 23272 61936
rect 24036 61838 24134 61936
rect 24422 61838 24520 61936
rect 25284 61838 25382 61936
rect 25670 61838 25768 61936
rect 26532 61838 26630 61936
rect 26918 61838 27016 61936
rect 27780 61838 27878 61936
rect 28166 61838 28264 61936
rect 29028 61838 29126 61936
rect 29414 61838 29512 61936
rect 30276 61838 30374 61936
rect 30662 61838 30760 61936
rect 31524 61838 31622 61936
rect 31910 61838 32008 61936
rect 32772 61838 32870 61936
rect 33158 61838 33256 61936
rect 34020 61838 34118 61936
rect 34406 61838 34504 61936
rect 35268 61838 35366 61936
rect 35654 61838 35752 61936
rect 36516 61838 36614 61936
rect 36902 61838 37000 61936
rect 37764 61838 37862 61936
rect 38150 61838 38248 61936
rect 39012 61838 39110 61936
rect 39398 61838 39496 61936
rect 40260 61838 40358 61936
rect 40646 61838 40744 61936
rect 41508 61838 41606 61936
rect 41894 61838 41992 61936
rect 42756 61838 42854 61936
rect 43142 61838 43240 61936
rect 44004 61838 44102 61936
rect 44390 61838 44488 61936
rect 45252 61838 45350 61936
rect 45638 61838 45736 61936
rect 46500 61838 46598 61936
rect 46886 61838 46984 61936
rect 47748 61838 47846 61936
rect 48134 61838 48232 61936
rect 48996 61838 49094 61936
rect 49382 61838 49480 61936
rect 50244 61838 50342 61936
rect 50630 61838 50728 61936
rect 51492 61838 51590 61936
rect 51878 61838 51976 61936
rect 52740 61838 52838 61936
rect 53126 61838 53224 61936
rect 12685 61247 12783 61345
rect 13328 61266 13388 61326
rect 13952 61266 14012 61326
rect 14576 61266 14636 61326
rect 15200 61266 15260 61326
rect 15824 61266 15884 61326
rect 16448 61266 16508 61326
rect 17072 61266 17132 61326
rect 17696 61266 17756 61326
rect 18320 61266 18380 61326
rect 18944 61266 19004 61326
rect 19568 61266 19628 61326
rect 20192 61266 20252 61326
rect 20816 61266 20876 61326
rect 21440 61266 21500 61326
rect 22064 61266 22124 61326
rect 22688 61266 22748 61326
rect 23312 61266 23372 61326
rect 23936 61266 23996 61326
rect 24560 61266 24620 61326
rect 25184 61266 25244 61326
rect 25808 61266 25868 61326
rect 26432 61266 26492 61326
rect 27056 61266 27116 61326
rect 27680 61266 27740 61326
rect 28304 61266 28364 61326
rect 28928 61266 28988 61326
rect 29552 61266 29612 61326
rect 30176 61266 30236 61326
rect 30800 61266 30860 61326
rect 31424 61266 31484 61326
rect 32048 61266 32108 61326
rect 32672 61266 32732 61326
rect 33296 61266 33356 61326
rect 33920 61266 33980 61326
rect 34544 61266 34604 61326
rect 35168 61266 35228 61326
rect 35792 61266 35852 61326
rect 36416 61266 36476 61326
rect 37040 61266 37100 61326
rect 37664 61266 37724 61326
rect 38288 61266 38348 61326
rect 38912 61266 38972 61326
rect 39536 61266 39596 61326
rect 40160 61266 40220 61326
rect 40784 61266 40844 61326
rect 41408 61266 41468 61326
rect 42032 61266 42092 61326
rect 42656 61266 42716 61326
rect 43280 61266 43340 61326
rect 43904 61266 43964 61326
rect 44528 61266 44588 61326
rect 45152 61266 45212 61326
rect 45776 61266 45836 61326
rect 46400 61266 46460 61326
rect 47024 61266 47084 61326
rect 47648 61266 47708 61326
rect 48272 61266 48332 61326
rect 48896 61266 48956 61326
rect 49520 61266 49580 61326
rect 50144 61266 50204 61326
rect 50768 61266 50828 61326
rect 51392 61266 51452 61326
rect 52016 61266 52076 61326
rect 52640 61266 52700 61326
rect 53245 61247 53343 61345
rect 12008 60942 12068 61002
rect 53960 60942 54020 61002
rect 12008 60705 12068 60765
rect 53960 60705 54020 60765
rect 12008 60468 12068 60528
rect 53960 60468 54020 60528
rect 5776 60343 5874 60441
rect 6201 60343 6299 60441
rect 6633 60343 6731 60441
rect 7015 60320 7113 60418
rect 7287 60320 7385 60418
rect 58643 60320 58741 60418
rect 58915 60320 59013 60418
rect 59297 60343 59395 60441
rect 59729 60343 59827 60441
rect 60154 60343 60252 60441
rect 12008 60152 12068 60212
rect 53960 60152 54020 60212
rect 5776 59969 5874 60067
rect 6201 59911 6299 60009
rect 6633 59911 6731 60009
rect 7015 59925 7113 60023
rect 7287 59925 7385 60023
rect 12008 59915 12068 59975
rect 53960 59915 54020 59975
rect 58643 59925 58741 60023
rect 58915 59925 59013 60023
rect 59297 59911 59395 60009
rect 59729 59911 59827 60009
rect 60154 59969 60252 60067
rect 12008 59678 12068 59738
rect 53960 59678 54020 59738
rect 5776 59553 5874 59651
rect 6201 59553 6299 59651
rect 6633 59553 6731 59651
rect 7015 59530 7113 59628
rect 7287 59530 7382 59628
rect 58643 59530 58741 59628
rect 58915 59530 59013 59628
rect 59297 59553 59395 59651
rect 59729 59553 59827 59651
rect 60154 59553 60252 59651
rect 12008 59362 12068 59422
rect 53960 59362 54020 59422
rect 5776 59179 5874 59277
rect 6201 59121 6299 59219
rect 6633 59121 6731 59219
rect 7015 59135 7113 59233
rect 7287 59135 7385 59233
rect 12008 59125 12068 59185
rect 53960 59125 54020 59185
rect 58643 59135 58741 59233
rect 58915 59135 59013 59233
rect 59297 59121 59395 59219
rect 59729 59121 59827 59219
rect 60154 59179 60252 59277
rect 12008 58888 12068 58948
rect 53960 58888 54020 58948
rect 5776 58763 5874 58861
rect 6201 58763 6299 58861
rect 6633 58763 6731 58861
rect 7015 58740 7113 58838
rect 7287 58740 7385 58838
rect 58643 58740 58741 58838
rect 58915 58740 59013 58838
rect 59297 58763 59395 58861
rect 59729 58763 59827 58861
rect 60154 58763 60252 58861
rect 12008 58572 12068 58632
rect 53960 58572 54020 58632
rect 5776 58389 5874 58487
rect 6201 58331 6299 58429
rect 6633 58331 6731 58429
rect 7015 58345 7113 58443
rect 7287 58345 7385 58443
rect 12008 58335 12068 58395
rect 53960 58335 54020 58395
rect 58643 58345 58741 58443
rect 58915 58345 59013 58443
rect 59297 58331 59395 58429
rect 59729 58331 59827 58429
rect 60154 58389 60252 58487
rect 12008 58098 12068 58158
rect 53960 58098 54020 58158
rect 5776 57973 5874 58071
rect 6201 57973 6299 58071
rect 6633 57973 6731 58071
rect 7015 57950 7113 58048
rect 7287 57950 7385 58048
rect 58643 57950 58741 58048
rect 58915 57950 59013 58048
rect 59297 57973 59395 58071
rect 59729 57973 59827 58071
rect 60154 57973 60252 58071
rect 12008 57782 12068 57842
rect 53960 57782 54020 57842
rect 5776 57599 5874 57697
rect 6201 57541 6299 57639
rect 6633 57541 6731 57639
rect 7015 57555 7113 57653
rect 7287 57555 7385 57653
rect 12008 57545 12068 57605
rect 53960 57545 54020 57605
rect 58643 57555 58741 57653
rect 58915 57555 59013 57653
rect 59297 57541 59395 57639
rect 59729 57541 59827 57639
rect 60154 57599 60252 57697
rect 12008 57308 12068 57368
rect 53960 57308 54020 57368
rect 5776 57183 5874 57281
rect 6201 57183 6299 57281
rect 6633 57183 6731 57281
rect 7015 57160 7113 57258
rect 7287 57160 7385 57258
rect 58643 57160 58741 57258
rect 58915 57160 59013 57258
rect 59297 57183 59395 57281
rect 59729 57183 59827 57281
rect 60154 57183 60252 57281
rect 12008 56992 12068 57052
rect 53960 56992 54020 57052
rect 5776 56809 5874 56907
rect 6201 56751 6299 56849
rect 6633 56751 6731 56849
rect 7015 56765 7113 56863
rect 7287 56765 7385 56863
rect 12008 56755 12068 56815
rect 53960 56755 54020 56815
rect 58643 56765 58741 56863
rect 58915 56765 59013 56863
rect 59297 56751 59395 56849
rect 59729 56751 59827 56849
rect 60154 56809 60252 56907
rect 12008 56518 12068 56578
rect 53960 56518 54020 56578
rect 5776 56393 5874 56491
rect 6201 56393 6299 56491
rect 6633 56393 6731 56491
rect 7015 56370 7113 56468
rect 7287 56370 7385 56468
rect 58643 56370 58741 56468
rect 58915 56370 59013 56468
rect 59297 56393 59395 56491
rect 59729 56393 59827 56491
rect 60154 56393 60252 56491
rect 12008 56202 12068 56262
rect 53960 56202 54020 56262
rect 5776 56019 5874 56117
rect 6201 55961 6299 56059
rect 6633 55961 6731 56059
rect 7015 55975 7113 56073
rect 7287 55975 7385 56073
rect 12008 55965 12068 56025
rect 53960 55965 54020 56025
rect 58643 55975 58741 56073
rect 58915 55975 59013 56073
rect 59297 55961 59395 56059
rect 59729 55961 59827 56059
rect 60154 56019 60252 56117
rect 12008 55728 12068 55788
rect 53960 55728 54020 55788
rect 5776 55603 5874 55701
rect 6201 55603 6299 55701
rect 6633 55603 6731 55701
rect 7015 55580 7113 55678
rect 7287 55580 7385 55678
rect 58643 55580 58741 55678
rect 58915 55580 59013 55678
rect 59297 55603 59395 55701
rect 59729 55603 59827 55701
rect 60154 55603 60252 55701
rect 12008 55412 12068 55472
rect 53960 55412 54020 55472
rect 5776 55229 5874 55327
rect 6201 55171 6299 55269
rect 6633 55171 6731 55269
rect 7015 55185 7113 55283
rect 7287 55185 7385 55283
rect 12008 55175 12068 55235
rect 53960 55175 54020 55235
rect 58643 55185 58741 55283
rect 58915 55185 59013 55283
rect 59297 55171 59395 55269
rect 59729 55171 59827 55269
rect 60154 55229 60252 55327
rect 12008 54938 12068 54998
rect 53960 54938 54020 54998
rect 5776 54813 5874 54911
rect 6201 54813 6299 54911
rect 6633 54813 6731 54911
rect 7015 54790 7113 54888
rect 7287 54790 7385 54888
rect 58643 54790 58741 54888
rect 58915 54790 59013 54888
rect 59297 54813 59395 54911
rect 59729 54813 59827 54911
rect 60154 54813 60252 54911
rect 12008 54622 12068 54682
rect 53960 54622 54020 54682
rect 5776 54439 5874 54537
rect 6201 54381 6299 54479
rect 6633 54381 6731 54479
rect 7015 54395 7113 54493
rect 7287 54395 7385 54493
rect 12008 54385 12068 54445
rect 53960 54385 54020 54445
rect 58643 54395 58741 54493
rect 58915 54395 59013 54493
rect 59297 54381 59395 54479
rect 59729 54381 59827 54479
rect 60154 54439 60252 54537
rect 12008 54148 12068 54208
rect 53960 54148 54020 54208
rect 5776 54023 5874 54121
rect 6201 54023 6299 54121
rect 6633 54023 6731 54121
rect 7015 54000 7113 54098
rect 7287 54000 7385 54098
rect 58643 54000 58741 54098
rect 58915 54000 59013 54098
rect 59297 54023 59395 54121
rect 59729 54023 59827 54121
rect 60154 54023 60252 54121
rect 12008 53832 12068 53892
rect 53960 53832 54020 53892
rect 5776 53649 5874 53747
rect 6201 53591 6299 53689
rect 6633 53591 6731 53689
rect 7015 53605 7113 53703
rect 7287 53605 7385 53703
rect 12008 53595 12068 53655
rect 53960 53595 54020 53655
rect 58643 53605 58741 53703
rect 58915 53605 59013 53703
rect 59297 53591 59395 53689
rect 59729 53591 59827 53689
rect 60154 53649 60252 53747
rect 12008 53358 12068 53418
rect 53960 53358 54020 53418
rect 5776 53233 5874 53331
rect 6201 53233 6299 53331
rect 6633 53233 6731 53331
rect 7015 53210 7113 53308
rect 7287 53210 7385 53308
rect 58643 53210 58741 53308
rect 58915 53210 59013 53308
rect 59297 53233 59395 53331
rect 59729 53233 59827 53331
rect 60154 53233 60252 53331
rect 12008 53042 12068 53102
rect 53960 53042 54020 53102
rect 5776 52859 5874 52957
rect 6201 52801 6299 52899
rect 6633 52801 6731 52899
rect 7015 52815 7113 52913
rect 7287 52815 7385 52913
rect 12008 52805 12068 52865
rect 53960 52805 54020 52865
rect 58643 52815 58741 52913
rect 58915 52815 59013 52913
rect 59297 52801 59395 52899
rect 59729 52801 59827 52899
rect 60154 52859 60252 52957
rect 12008 52568 12068 52628
rect 53960 52568 54020 52628
rect 5776 52443 5874 52541
rect 6201 52443 6299 52541
rect 6633 52443 6731 52541
rect 7015 52420 7113 52518
rect 7287 52420 7385 52518
rect 58643 52420 58741 52518
rect 58915 52420 59013 52518
rect 59297 52443 59395 52541
rect 59729 52443 59827 52541
rect 60154 52443 60252 52541
rect 12008 52252 12068 52312
rect 53960 52252 54020 52312
rect 5776 52069 5874 52167
rect 6201 52011 6299 52109
rect 6633 52011 6731 52109
rect 7015 52025 7113 52123
rect 7287 52025 7385 52123
rect 12008 52015 12068 52075
rect 53960 52015 54020 52075
rect 58643 52025 58741 52123
rect 58915 52025 59013 52123
rect 59297 52011 59395 52109
rect 59729 52011 59827 52109
rect 60154 52069 60252 52167
rect 12008 51778 12068 51838
rect 53960 51778 54020 51838
rect 5776 51653 5874 51751
rect 6201 51653 6299 51751
rect 6633 51653 6731 51751
rect 7015 51630 7113 51728
rect 7287 51630 7385 51728
rect 58643 51630 58741 51728
rect 58915 51630 59013 51728
rect 59297 51653 59395 51751
rect 59729 51653 59827 51751
rect 60154 51653 60252 51751
rect 12008 51462 12068 51522
rect 53960 51462 54020 51522
rect 5776 51279 5874 51377
rect 6201 51221 6299 51319
rect 6633 51221 6731 51319
rect 7015 51235 7113 51333
rect 7287 51235 7385 51333
rect 12008 51225 12068 51285
rect 53960 51225 54020 51285
rect 58643 51235 58741 51333
rect 58915 51235 59013 51333
rect 59297 51221 59395 51319
rect 59729 51221 59827 51319
rect 60154 51279 60252 51377
rect 12008 50988 12068 51048
rect 53960 50988 54020 51048
rect 5776 50863 5874 50961
rect 6201 50863 6299 50961
rect 6633 50863 6731 50961
rect 7015 50840 7113 50938
rect 7287 50840 7385 50938
rect 58643 50840 58741 50938
rect 58915 50840 59013 50938
rect 59297 50863 59395 50961
rect 59729 50863 59827 50961
rect 60154 50863 60252 50961
rect 12008 50672 12068 50732
rect 53960 50672 54020 50732
rect 5776 50489 5874 50587
rect 6201 50431 6299 50529
rect 6633 50431 6731 50529
rect 7015 50445 7113 50543
rect 7287 50445 7385 50543
rect 12008 50435 12068 50495
rect 53960 50435 54020 50495
rect 58643 50445 58741 50543
rect 58915 50445 59013 50543
rect 59297 50431 59395 50529
rect 59729 50431 59827 50529
rect 60154 50489 60252 50587
rect 12008 50198 12068 50258
rect 53960 50198 54020 50258
rect 5776 50073 5874 50171
rect 6201 50073 6299 50171
rect 6633 50073 6731 50171
rect 7015 50050 7113 50148
rect 7287 50050 7385 50148
rect 58643 50050 58741 50148
rect 58915 50050 59013 50148
rect 59297 50073 59395 50171
rect 59729 50073 59827 50171
rect 60154 50073 60252 50171
rect 12008 49882 12068 49942
rect 53960 49882 54020 49942
rect 5776 49699 5874 49797
rect 6201 49641 6299 49739
rect 6633 49641 6731 49739
rect 7015 49655 7113 49753
rect 7287 49655 7385 49753
rect 12008 49645 12068 49705
rect 53960 49645 54020 49705
rect 58643 49655 58741 49753
rect 58915 49655 59013 49753
rect 59297 49641 59395 49739
rect 59729 49641 59827 49739
rect 60154 49699 60252 49797
rect 12008 49408 12068 49468
rect 53960 49408 54020 49468
rect 5776 49283 5874 49381
rect 6201 49283 6299 49381
rect 6633 49283 6731 49381
rect 7015 49260 7113 49358
rect 7287 49260 7385 49358
rect 58643 49260 58741 49358
rect 58915 49260 59013 49358
rect 59297 49283 59395 49381
rect 59729 49283 59827 49381
rect 60154 49283 60252 49381
rect 12008 49092 12068 49152
rect 53960 49092 54020 49152
rect 5776 48909 5874 49007
rect 6201 48851 6299 48949
rect 6633 48851 6731 48949
rect 7015 48865 7113 48963
rect 7287 48865 7385 48963
rect 12008 48855 12068 48915
rect 53960 48855 54020 48915
rect 58643 48865 58741 48963
rect 58915 48865 59013 48963
rect 59297 48851 59395 48949
rect 59729 48851 59827 48949
rect 60154 48909 60252 49007
rect 12008 48618 12068 48678
rect 53960 48618 54020 48678
rect 5776 48493 5874 48591
rect 6201 48493 6299 48591
rect 6633 48493 6731 48591
rect 7015 48470 7113 48568
rect 7287 48470 7385 48568
rect 58643 48470 58741 48568
rect 58915 48470 59013 48568
rect 59297 48493 59395 48591
rect 59729 48493 59827 48591
rect 60154 48493 60252 48591
rect 12008 48302 12068 48362
rect 53960 48302 54020 48362
rect 5776 48119 5874 48217
rect 6201 48061 6299 48159
rect 6633 48061 6731 48159
rect 7015 48075 7113 48173
rect 7287 48075 7385 48173
rect 12008 48065 12068 48125
rect 53960 48065 54020 48125
rect 58643 48075 58741 48173
rect 58915 48075 59013 48173
rect 59297 48061 59395 48159
rect 59729 48061 59827 48159
rect 60154 48119 60252 48217
rect 12008 47828 12068 47888
rect 53960 47828 54020 47888
rect 5776 47703 5874 47801
rect 6201 47703 6299 47801
rect 6633 47703 6731 47801
rect 7015 47680 7113 47778
rect 7287 47680 7385 47778
rect 58643 47680 58741 47778
rect 58915 47680 59013 47778
rect 59297 47703 59395 47801
rect 59729 47703 59827 47801
rect 60154 47703 60252 47801
rect 12008 47512 12068 47572
rect 53960 47512 54020 47572
rect 5776 47329 5874 47427
rect 6201 47271 6299 47369
rect 6633 47271 6731 47369
rect 7015 47285 7113 47383
rect 7287 47285 7385 47383
rect 12008 47275 12068 47335
rect 53960 47275 54020 47335
rect 58643 47285 58741 47383
rect 58915 47285 59013 47383
rect 59297 47271 59395 47369
rect 59729 47271 59827 47369
rect 60154 47329 60252 47427
rect 12008 47038 12068 47098
rect 53960 47038 54020 47098
rect 5776 46913 5874 47011
rect 6201 46913 6299 47011
rect 6633 46913 6731 47011
rect 7015 46890 7113 46988
rect 7287 46890 7385 46988
rect 58643 46890 58741 46988
rect 58915 46890 59013 46988
rect 59297 46913 59395 47011
rect 59729 46913 59827 47011
rect 60154 46913 60252 47011
rect 12008 46722 12068 46782
rect 53960 46722 54020 46782
rect 5776 46539 5874 46637
rect 6201 46481 6299 46579
rect 6633 46481 6731 46579
rect 7015 46495 7113 46593
rect 7287 46495 7385 46593
rect 12008 46485 12068 46545
rect 53960 46485 54020 46545
rect 58643 46495 58741 46593
rect 58915 46495 59013 46593
rect 59297 46481 59395 46579
rect 59729 46481 59827 46579
rect 60154 46539 60252 46637
rect 12008 46248 12068 46308
rect 53960 46248 54020 46308
rect 5776 46123 5874 46221
rect 6201 46123 6299 46221
rect 6633 46123 6731 46221
rect 7015 46100 7113 46198
rect 7287 46100 7385 46198
rect 58643 46100 58741 46198
rect 58915 46100 59013 46198
rect 59297 46123 59395 46221
rect 59729 46123 59827 46221
rect 60154 46123 60252 46221
rect 12008 45932 12068 45992
rect 53960 45932 54020 45992
rect 5776 45749 5874 45847
rect 6201 45691 6299 45789
rect 6633 45691 6731 45789
rect 7015 45705 7113 45803
rect 7287 45705 7385 45803
rect 12008 45695 12068 45755
rect 53960 45695 54020 45755
rect 58643 45705 58741 45803
rect 58915 45705 59013 45803
rect 59297 45691 59395 45789
rect 59729 45691 59827 45789
rect 60154 45749 60252 45847
rect 12008 45458 12068 45518
rect 53960 45458 54020 45518
rect 5776 45333 5874 45431
rect 6201 45333 6299 45431
rect 6633 45333 6731 45431
rect 7015 45310 7113 45408
rect 7287 45310 7385 45408
rect 58643 45310 58741 45408
rect 58915 45310 59013 45408
rect 59297 45333 59395 45431
rect 59729 45333 59827 45431
rect 60154 45333 60252 45431
rect 12008 45142 12068 45202
rect 53960 45142 54020 45202
rect 5776 44959 5874 45057
rect 6201 44901 6299 44999
rect 6633 44901 6731 44999
rect 7015 44915 7113 45013
rect 7287 44915 7385 45013
rect 12008 44905 12068 44965
rect 53960 44905 54020 44965
rect 58643 44915 58741 45013
rect 58915 44915 59013 45013
rect 59297 44901 59395 44999
rect 59729 44901 59827 44999
rect 60154 44959 60252 45057
rect 12008 44668 12068 44728
rect 53960 44668 54020 44728
rect 5776 44543 5874 44641
rect 6201 44543 6299 44641
rect 6633 44543 6731 44641
rect 7015 44520 7113 44618
rect 7287 44520 7385 44618
rect 58643 44520 58741 44618
rect 58915 44520 59013 44618
rect 59297 44543 59395 44641
rect 59729 44543 59827 44641
rect 60154 44543 60252 44641
rect 12008 44352 12068 44412
rect 53960 44352 54020 44412
rect 5776 44169 5874 44267
rect 6201 44111 6299 44209
rect 6633 44111 6731 44209
rect 7015 44125 7113 44223
rect 7287 44125 7385 44223
rect 12008 44115 12068 44175
rect 53960 44115 54020 44175
rect 58643 44125 58741 44223
rect 58915 44125 59013 44223
rect 59297 44111 59395 44209
rect 59729 44111 59827 44209
rect 60154 44169 60252 44267
rect 12008 43878 12068 43938
rect 53960 43878 54020 43938
rect 5776 43753 5874 43851
rect 6201 43753 6299 43851
rect 6633 43753 6731 43851
rect 7015 43730 7113 43828
rect 7287 43730 7385 43828
rect 58643 43730 58741 43828
rect 58915 43730 59013 43828
rect 59297 43753 59395 43851
rect 59729 43753 59827 43851
rect 60154 43753 60252 43851
rect 12008 43562 12068 43622
rect 53960 43562 54020 43622
rect 5776 43379 5874 43477
rect 6201 43321 6299 43419
rect 6633 43321 6731 43419
rect 7015 43335 7113 43433
rect 7287 43335 7385 43433
rect 12008 43325 12068 43385
rect 53960 43325 54020 43385
rect 58643 43335 58741 43433
rect 58915 43335 59013 43433
rect 59297 43321 59395 43419
rect 59729 43321 59827 43419
rect 60154 43379 60252 43477
rect 12008 43088 12068 43148
rect 53960 43088 54020 43148
rect 5776 42963 5874 43061
rect 6201 42963 6299 43061
rect 6633 42963 6731 43061
rect 7015 42940 7113 43038
rect 7287 42940 7385 43038
rect 58643 42940 58741 43038
rect 58915 42940 59013 43038
rect 59297 42963 59395 43061
rect 59729 42963 59827 43061
rect 60154 42963 60252 43061
rect 12008 42772 12068 42832
rect 53960 42772 54020 42832
rect 5776 42589 5874 42687
rect 6201 42531 6299 42629
rect 6633 42531 6731 42629
rect 7015 42545 7113 42643
rect 7287 42545 7385 42643
rect 12008 42535 12068 42595
rect 53960 42535 54020 42595
rect 58643 42545 58741 42643
rect 58915 42545 59013 42643
rect 59297 42531 59395 42629
rect 59729 42531 59827 42629
rect 60154 42589 60252 42687
rect 12008 42298 12068 42358
rect 53960 42298 54020 42358
rect 5776 42173 5874 42271
rect 6201 42173 6299 42271
rect 6633 42173 6731 42271
rect 7015 42150 7113 42248
rect 7287 42150 7385 42248
rect 58643 42150 58741 42248
rect 58915 42150 59013 42248
rect 59297 42173 59395 42271
rect 59729 42173 59827 42271
rect 60154 42173 60252 42271
rect 12008 41982 12068 42042
rect 53960 41982 54020 42042
rect 5776 41799 5874 41897
rect 6201 41741 6299 41839
rect 6633 41741 6731 41839
rect 7015 41755 7113 41853
rect 7287 41755 7385 41853
rect 12008 41745 12068 41805
rect 53960 41745 54020 41805
rect 58643 41755 58741 41853
rect 58915 41755 59013 41853
rect 59297 41741 59395 41839
rect 59729 41741 59827 41839
rect 60154 41799 60252 41897
rect 12008 41508 12068 41568
rect 53960 41508 54020 41568
rect 5776 41383 5874 41481
rect 6201 41383 6299 41481
rect 6633 41383 6731 41481
rect 7015 41360 7113 41458
rect 7287 41360 7385 41458
rect 58643 41360 58741 41458
rect 58915 41360 59013 41458
rect 59297 41383 59395 41481
rect 59729 41383 59827 41481
rect 60154 41383 60252 41481
rect 12008 41192 12068 41252
rect 53960 41192 54020 41252
rect 5776 41009 5874 41107
rect 6201 40951 6299 41049
rect 6633 40951 6731 41049
rect 7015 40965 7113 41063
rect 7287 40965 7385 41063
rect 12008 40955 12068 41015
rect 53960 40955 54020 41015
rect 58643 40965 58741 41063
rect 58915 40965 59013 41063
rect 59297 40951 59395 41049
rect 59729 40951 59827 41049
rect 60154 41009 60252 41107
rect 12008 40718 12068 40778
rect 53960 40718 54020 40778
rect 5776 40593 5874 40691
rect 6201 40593 6299 40691
rect 6633 40593 6731 40691
rect 7015 40570 7113 40668
rect 7287 40570 7385 40668
rect 58643 40570 58741 40668
rect 58915 40570 59013 40668
rect 59297 40593 59395 40691
rect 59729 40593 59827 40691
rect 60154 40593 60252 40691
rect 12008 40402 12068 40462
rect 53960 40402 54020 40462
rect 5776 40219 5874 40317
rect 6201 40161 6299 40259
rect 6633 40161 6731 40259
rect 7015 40175 7113 40273
rect 7287 40175 7385 40273
rect 12008 40165 12068 40225
rect 53960 40165 54020 40225
rect 58643 40175 58741 40273
rect 58915 40175 59013 40273
rect 59297 40161 59395 40259
rect 59729 40161 59827 40259
rect 60154 40219 60252 40317
rect 12008 39928 12068 39988
rect 53960 39928 54020 39988
rect 5776 39803 5874 39901
rect 6201 39803 6299 39901
rect 6633 39803 6731 39901
rect 7015 39780 7113 39878
rect 7287 39780 7385 39878
rect 58643 39780 58741 39878
rect 58915 39780 59013 39878
rect 59297 39803 59395 39901
rect 59729 39803 59827 39901
rect 60154 39803 60252 39901
rect 12008 39612 12068 39672
rect 53960 39612 54020 39672
rect 5776 39429 5874 39527
rect 6201 39371 6299 39469
rect 6633 39371 6731 39469
rect 7015 39385 7113 39483
rect 7287 39385 7385 39483
rect 12008 39375 12068 39435
rect 53960 39375 54020 39435
rect 58643 39385 58741 39483
rect 58915 39385 59013 39483
rect 59297 39371 59395 39469
rect 59729 39371 59827 39469
rect 60154 39429 60252 39527
rect 12008 39138 12068 39198
rect 53960 39138 54020 39198
rect 5776 39013 5874 39111
rect 6201 39013 6299 39111
rect 6633 39013 6731 39111
rect 7015 38990 7113 39088
rect 7287 38990 7385 39088
rect 58643 38990 58741 39088
rect 58915 38990 59013 39088
rect 59297 39013 59395 39111
rect 59729 39013 59827 39111
rect 60154 39013 60252 39111
rect 12008 38822 12068 38882
rect 53960 38822 54020 38882
rect 5776 38639 5874 38737
rect 6201 38581 6299 38679
rect 6633 38581 6731 38679
rect 7015 38595 7113 38693
rect 7287 38595 7385 38693
rect 12008 38585 12068 38645
rect 53960 38585 54020 38645
rect 58643 38595 58741 38693
rect 58915 38595 59013 38693
rect 59297 38581 59395 38679
rect 59729 38581 59827 38679
rect 60154 38639 60252 38737
rect 12008 38348 12068 38408
rect 53960 38348 54020 38408
rect 5776 38223 5874 38321
rect 6201 38223 6299 38321
rect 6633 38223 6731 38321
rect 7015 38200 7113 38298
rect 7287 38200 7385 38298
rect 58643 38200 58741 38298
rect 58915 38200 59013 38298
rect 59297 38223 59395 38321
rect 59729 38223 59827 38321
rect 60154 38223 60252 38321
rect 12008 38032 12068 38092
rect 53960 38032 54020 38092
rect 5776 37849 5874 37947
rect 6201 37791 6299 37889
rect 6633 37791 6731 37889
rect 7015 37805 7113 37903
rect 7287 37805 7385 37903
rect 12008 37795 12068 37855
rect 53960 37795 54020 37855
rect 58643 37805 58741 37903
rect 58915 37805 59013 37903
rect 59297 37791 59395 37889
rect 59729 37791 59827 37889
rect 60154 37849 60252 37947
rect 12008 37558 12068 37618
rect 53960 37558 54020 37618
rect 5776 37433 5874 37531
rect 6201 37433 6299 37531
rect 6633 37433 6731 37531
rect 7015 37410 7113 37508
rect 7287 37410 7385 37508
rect 58643 37410 58741 37508
rect 58915 37410 59013 37508
rect 59297 37433 59395 37531
rect 59729 37433 59827 37531
rect 60154 37433 60252 37531
rect 12008 37242 12068 37302
rect 53960 37242 54020 37302
rect 5776 37059 5874 37157
rect 6201 37001 6299 37099
rect 6633 37001 6731 37099
rect 7015 37015 7113 37113
rect 7287 37015 7385 37113
rect 12008 37005 12068 37065
rect 53960 37005 54020 37065
rect 58643 37015 58741 37113
rect 58915 37015 59013 37113
rect 59297 37001 59395 37099
rect 59729 37001 59827 37099
rect 60154 37059 60252 37157
rect 12008 36768 12068 36828
rect 53960 36768 54020 36828
rect 5776 36643 5874 36741
rect 6201 36643 6299 36741
rect 6633 36643 6731 36741
rect 7015 36620 7113 36718
rect 7287 36620 7385 36718
rect 58643 36620 58741 36718
rect 58915 36620 59013 36718
rect 59297 36643 59395 36741
rect 59729 36643 59827 36741
rect 60154 36643 60252 36741
rect 12008 36452 12068 36512
rect 53960 36452 54020 36512
rect 5776 36269 5874 36367
rect 6201 36211 6299 36309
rect 6633 36211 6731 36309
rect 7015 36225 7113 36323
rect 7287 36225 7385 36323
rect 12008 36215 12068 36275
rect 53960 36215 54020 36275
rect 58643 36225 58741 36323
rect 58915 36225 59013 36323
rect 59297 36211 59395 36309
rect 59729 36211 59827 36309
rect 60154 36269 60252 36367
rect 12008 35978 12068 36038
rect 53960 35978 54020 36038
rect 5776 35853 5874 35951
rect 6201 35853 6299 35951
rect 6633 35853 6731 35951
rect 7015 35830 7113 35928
rect 7287 35830 7385 35928
rect 58643 35830 58741 35928
rect 58915 35830 59013 35928
rect 59297 35853 59395 35951
rect 59729 35853 59827 35951
rect 60154 35853 60252 35951
rect 12008 35662 12068 35722
rect 53960 35662 54020 35722
rect 5776 35479 5874 35577
rect 6201 35421 6299 35519
rect 6633 35421 6731 35519
rect 7015 35435 7113 35533
rect 7287 35435 7385 35533
rect 7733 35391 7831 35489
rect 8158 35390 8256 35488
rect 9201 35406 9299 35504
rect 10725 35406 10823 35504
rect 12008 35425 12068 35485
rect 53960 35425 54020 35485
rect 55205 35406 55303 35504
rect 56729 35406 56827 35504
rect 57772 35390 57870 35488
rect 58197 35391 58295 35489
rect 58643 35435 58741 35533
rect 58915 35435 59013 35533
rect 59297 35421 59395 35519
rect 59729 35421 59827 35519
rect 60154 35479 60252 35577
rect 12008 35188 12068 35248
rect 53960 35188 54020 35248
rect 5776 35063 5874 35161
rect 6201 35063 6299 35161
rect 6633 35063 6731 35161
rect 7015 35040 7113 35138
rect 7287 35040 7385 35138
rect 58643 35040 58741 35138
rect 58915 35040 59013 35138
rect 59297 35063 59395 35161
rect 59729 35063 59827 35161
rect 60154 35063 60252 35161
rect 12008 34872 12068 34932
rect 53960 34872 54020 34932
rect 5776 34689 5874 34787
rect 6201 34631 6299 34729
rect 6633 34631 6731 34729
rect 7015 34645 7113 34743
rect 7287 34645 7385 34743
rect 12008 34635 12068 34695
rect 53960 34635 54020 34695
rect 58643 34645 58741 34743
rect 58915 34645 59013 34743
rect 59297 34631 59395 34729
rect 59729 34631 59827 34729
rect 60154 34689 60252 34787
rect 12008 34398 12068 34458
rect 53960 34398 54020 34458
rect 5776 34273 5874 34371
rect 6201 34273 6299 34371
rect 6633 34273 6731 34371
rect 7015 34250 7113 34348
rect 7287 34250 7385 34348
rect 58643 34250 58741 34348
rect 58915 34250 59013 34348
rect 59297 34273 59395 34371
rect 59729 34273 59827 34371
rect 60154 34273 60252 34371
rect 12008 34082 12068 34142
rect 53960 34082 54020 34142
rect 5776 33899 5874 33997
rect 6201 33841 6299 33939
rect 6633 33841 6731 33939
rect 7015 33855 7113 33953
rect 7287 33855 7385 33953
rect 12008 33845 12068 33905
rect 53960 33845 54020 33905
rect 58643 33855 58741 33953
rect 58915 33855 59013 33953
rect 59297 33841 59395 33939
rect 59729 33841 59827 33939
rect 60154 33899 60252 33997
rect 12008 33608 12068 33668
rect 53960 33608 54020 33668
rect 5776 33483 5874 33581
rect 6201 33483 6299 33581
rect 6633 33483 6731 33581
rect 7015 33460 7113 33558
rect 7287 33460 7385 33558
rect 58643 33460 58741 33558
rect 58915 33460 59013 33558
rect 59297 33483 59395 33581
rect 59729 33483 59827 33581
rect 60154 33483 60252 33581
rect 12008 33292 12068 33352
rect 53960 33292 54020 33352
rect 5776 33109 5874 33207
rect 6201 33051 6299 33149
rect 6633 33051 6731 33149
rect 7015 33065 7113 33163
rect 7287 33065 7385 33163
rect 12008 33055 12068 33115
rect 53960 33055 54020 33115
rect 58643 33065 58741 33163
rect 58915 33065 59013 33163
rect 59297 33051 59395 33149
rect 59729 33051 59827 33149
rect 60154 33109 60252 33207
rect 12008 32818 12068 32878
rect 53960 32818 54020 32878
rect 5776 32693 5874 32791
rect 6201 32693 6299 32791
rect 6633 32693 6731 32791
rect 7015 32670 7113 32768
rect 7287 32670 7385 32768
rect 58643 32670 58741 32768
rect 58915 32670 59013 32768
rect 59297 32693 59395 32791
rect 59729 32693 59827 32791
rect 60154 32693 60252 32791
rect 12008 32502 12068 32562
rect 53960 32502 54020 32562
rect 5776 32319 5874 32417
rect 6201 32261 6299 32359
rect 6633 32261 6731 32359
rect 7015 32275 7113 32373
rect 7287 32275 7385 32373
rect 12008 32265 12068 32325
rect 53960 32265 54020 32325
rect 58643 32275 58741 32373
rect 58915 32275 59013 32373
rect 59297 32261 59395 32359
rect 59729 32261 59827 32359
rect 60154 32319 60252 32417
rect 12008 32028 12068 32088
rect 53960 32028 54020 32088
rect 5776 31903 5874 32001
rect 6201 31903 6299 32001
rect 6633 31903 6731 32001
rect 7015 31880 7113 31978
rect 7287 31880 7385 31978
rect 58643 31880 58741 31978
rect 58915 31880 59013 31978
rect 59297 31903 59395 32001
rect 59729 31903 59827 32001
rect 60154 31903 60252 32001
rect 12008 31712 12068 31772
rect 53960 31712 54020 31772
rect 5776 31529 5874 31627
rect 6201 31471 6299 31569
rect 6633 31471 6731 31569
rect 7015 31485 7113 31583
rect 7287 31485 7385 31583
rect 12008 31475 12068 31535
rect 53960 31475 54020 31535
rect 58643 31485 58741 31583
rect 58915 31485 59013 31583
rect 59297 31471 59395 31569
rect 59729 31471 59827 31569
rect 60154 31529 60252 31627
rect 12008 31238 12068 31298
rect 53960 31238 54020 31298
rect 5776 31113 5874 31211
rect 6201 31113 6299 31211
rect 6633 31113 6731 31211
rect 7015 31090 7113 31188
rect 7287 31090 7385 31188
rect 58643 31090 58741 31188
rect 58915 31090 59013 31188
rect 59297 31113 59395 31211
rect 59729 31113 59827 31211
rect 60154 31113 60252 31211
rect 12008 30922 12068 30982
rect 53960 30922 54020 30982
rect 5776 30739 5874 30837
rect 6201 30681 6299 30779
rect 6633 30681 6731 30779
rect 7015 30695 7113 30793
rect 7287 30695 7385 30793
rect 12008 30685 12068 30745
rect 53960 30685 54020 30745
rect 58643 30695 58741 30793
rect 58915 30695 59013 30793
rect 59297 30681 59395 30779
rect 59729 30681 59827 30779
rect 60154 30739 60252 30837
rect 12008 30448 12068 30508
rect 53960 30448 54020 30508
rect 5776 30323 5874 30421
rect 6201 30323 6299 30421
rect 6633 30323 6731 30421
rect 7015 30300 7113 30398
rect 7287 30300 7385 30398
rect 58643 30300 58741 30398
rect 58915 30300 59013 30398
rect 59297 30323 59395 30421
rect 59729 30323 59827 30421
rect 60154 30323 60252 30421
rect 12008 30132 12068 30192
rect 53960 30132 54020 30192
rect 5776 29949 5874 30047
rect 6201 29891 6299 29989
rect 6633 29891 6731 29989
rect 7015 29905 7113 30003
rect 7287 29905 7385 30003
rect 12008 29895 12068 29955
rect 53960 29895 54020 29955
rect 58643 29905 58741 30003
rect 58915 29905 59013 30003
rect 59297 29891 59395 29989
rect 59729 29891 59827 29989
rect 60154 29949 60252 30047
rect 12008 29658 12068 29718
rect 53960 29658 54020 29718
rect 5776 29533 5874 29631
rect 6201 29533 6299 29631
rect 6633 29533 6731 29631
rect 7015 29510 7113 29608
rect 7287 29510 7385 29608
rect 58643 29510 58741 29608
rect 58915 29510 59013 29608
rect 59297 29533 59395 29631
rect 59729 29533 59827 29631
rect 60154 29533 60252 29631
rect 12008 29342 12068 29402
rect 53960 29342 54020 29402
rect 5776 29159 5874 29257
rect 6201 29101 6299 29199
rect 6633 29101 6731 29199
rect 7015 29115 7113 29213
rect 7287 29115 7385 29213
rect 12008 29105 12068 29165
rect 53960 29105 54020 29165
rect 58643 29115 58741 29213
rect 58915 29115 59013 29213
rect 59297 29101 59395 29199
rect 59729 29101 59827 29199
rect 60154 29159 60252 29257
rect 12008 28868 12068 28928
rect 53960 28868 54020 28928
rect 5776 28743 5874 28841
rect 6201 28743 6299 28841
rect 6633 28743 6731 28841
rect 7015 28720 7113 28818
rect 7287 28720 7385 28818
rect 58643 28720 58741 28818
rect 58915 28720 59013 28818
rect 59297 28743 59395 28841
rect 59729 28743 59827 28841
rect 60154 28743 60252 28841
rect 12008 28552 12068 28612
rect 53960 28552 54020 28612
rect 5776 28369 5874 28467
rect 6201 28311 6299 28409
rect 6633 28311 6731 28409
rect 7015 28325 7113 28423
rect 7287 28325 7385 28423
rect 12008 28315 12068 28375
rect 53960 28315 54020 28375
rect 58643 28325 58741 28423
rect 58915 28325 59013 28423
rect 59297 28311 59395 28409
rect 59729 28311 59827 28409
rect 60154 28369 60252 28467
rect 12008 28078 12068 28138
rect 53960 28078 54020 28138
rect 5776 27953 5874 28051
rect 6201 27953 6299 28051
rect 6633 27953 6731 28051
rect 7015 27930 7113 28028
rect 7287 27930 7385 28028
rect 58643 27930 58741 28028
rect 58915 27930 59013 28028
rect 59297 27953 59395 28051
rect 59729 27953 59827 28051
rect 60154 27953 60252 28051
rect 12008 27762 12068 27822
rect 53960 27762 54020 27822
rect 5776 27579 5874 27677
rect 6201 27521 6299 27619
rect 6633 27521 6731 27619
rect 7015 27535 7113 27633
rect 7287 27535 7385 27633
rect 12008 27525 12068 27585
rect 53960 27525 54020 27585
rect 58643 27535 58741 27633
rect 58915 27535 59013 27633
rect 59297 27521 59395 27619
rect 59729 27521 59827 27619
rect 60154 27579 60252 27677
rect 12008 27288 12068 27348
rect 53960 27288 54020 27348
rect 5776 27163 5874 27261
rect 6201 27163 6299 27261
rect 6633 27163 6731 27261
rect 7015 27140 7113 27238
rect 7287 27140 7382 27238
rect 58643 27140 58741 27238
rect 58915 27140 59013 27238
rect 59297 27163 59395 27261
rect 59729 27163 59827 27261
rect 60154 27163 60252 27261
rect 12008 26972 12068 27032
rect 53960 26972 54020 27032
rect 5776 26789 5874 26887
rect 6201 26731 6299 26829
rect 6633 26731 6731 26829
rect 7015 26745 7113 26843
rect 7287 26745 7385 26843
rect 12008 26735 12068 26795
rect 53960 26735 54020 26795
rect 58643 26745 58741 26843
rect 58915 26745 59013 26843
rect 59297 26731 59395 26829
rect 59729 26731 59827 26829
rect 60154 26789 60252 26887
rect 12008 26498 12068 26558
rect 53960 26498 54020 26558
rect 5776 26373 5874 26471
rect 6201 26373 6299 26471
rect 6633 26373 6731 26471
rect 7015 26350 7113 26448
rect 7287 26350 7385 26448
rect 58643 26350 58741 26448
rect 58915 26350 59013 26448
rect 59297 26373 59395 26471
rect 59729 26373 59827 26471
rect 60154 26373 60252 26471
rect 12008 26182 12068 26242
rect 53960 26182 54020 26242
rect 5776 25999 5874 26097
rect 6201 25941 6299 26039
rect 6633 25941 6731 26039
rect 7015 25955 7113 26053
rect 7287 25955 7385 26053
rect 12008 25945 12068 26005
rect 53960 25945 54020 26005
rect 58643 25955 58741 26053
rect 58915 25955 59013 26053
rect 59297 25941 59395 26039
rect 59729 25941 59827 26039
rect 60154 25999 60252 26097
rect 12008 25708 12068 25768
rect 53960 25708 54020 25768
rect 5776 25583 5874 25681
rect 6201 25583 6299 25681
rect 6633 25583 6731 25681
rect 7015 25560 7113 25658
rect 7287 25560 7385 25658
rect 58643 25560 58741 25658
rect 58915 25560 59013 25658
rect 59297 25583 59395 25681
rect 59729 25583 59827 25681
rect 60154 25583 60252 25681
rect 12008 25392 12068 25452
rect 53960 25392 54020 25452
rect 5776 25209 5874 25307
rect 6201 25151 6299 25249
rect 6633 25151 6731 25249
rect 7015 25165 7113 25263
rect 7287 25165 7385 25263
rect 12008 25155 12068 25215
rect 53960 25155 54020 25215
rect 58643 25165 58741 25263
rect 58915 25165 59013 25263
rect 59297 25151 59395 25249
rect 59729 25151 59827 25249
rect 60154 25209 60252 25307
rect 12008 24918 12068 24978
rect 53960 24918 54020 24978
rect 5776 24793 5874 24891
rect 6201 24793 6299 24891
rect 6633 24793 6731 24891
rect 7015 24770 7113 24868
rect 7287 24770 7385 24868
rect 58643 24770 58741 24868
rect 58915 24770 59013 24868
rect 59297 24793 59395 24891
rect 59729 24793 59827 24891
rect 60154 24793 60252 24891
rect 12008 24602 12068 24662
rect 53960 24602 54020 24662
rect 5776 24419 5874 24517
rect 6201 24361 6299 24459
rect 6633 24361 6731 24459
rect 7015 24375 7113 24473
rect 7287 24375 7385 24473
rect 12008 24365 12068 24425
rect 53960 24365 54020 24425
rect 58643 24375 58741 24473
rect 58915 24375 59013 24473
rect 59297 24361 59395 24459
rect 59729 24361 59827 24459
rect 60154 24419 60252 24517
rect 12008 24128 12068 24188
rect 53960 24128 54020 24188
rect 5776 24003 5874 24101
rect 6201 24003 6299 24101
rect 6633 24003 6731 24101
rect 7015 23980 7113 24078
rect 7287 23980 7385 24078
rect 58643 23980 58741 24078
rect 58915 23980 59013 24078
rect 59297 24003 59395 24101
rect 59729 24003 59827 24101
rect 60154 24003 60252 24101
rect 12008 23812 12068 23872
rect 53960 23812 54020 23872
rect 5776 23629 5874 23727
rect 6201 23571 6299 23669
rect 6633 23571 6731 23669
rect 7015 23585 7113 23683
rect 7287 23585 7385 23683
rect 12008 23575 12068 23635
rect 53960 23575 54020 23635
rect 58643 23585 58741 23683
rect 58915 23585 59013 23683
rect 59297 23571 59395 23669
rect 59729 23571 59827 23669
rect 60154 23629 60252 23727
rect 12008 23338 12068 23398
rect 53960 23338 54020 23398
rect 5776 23213 5874 23311
rect 6201 23213 6299 23311
rect 6633 23213 6731 23311
rect 7015 23190 7113 23288
rect 7287 23190 7385 23288
rect 58643 23190 58741 23288
rect 58915 23190 59013 23288
rect 59297 23213 59395 23311
rect 59729 23213 59827 23311
rect 60154 23213 60252 23311
rect 12008 23022 12068 23082
rect 53960 23022 54020 23082
rect 5776 22839 5874 22937
rect 6201 22781 6299 22879
rect 6633 22781 6731 22879
rect 7015 22795 7113 22893
rect 7287 22795 7385 22893
rect 12008 22785 12068 22845
rect 53960 22785 54020 22845
rect 58643 22795 58741 22893
rect 58915 22795 59013 22893
rect 59297 22781 59395 22879
rect 59729 22781 59827 22879
rect 60154 22839 60252 22937
rect 12008 22548 12068 22608
rect 53960 22548 54020 22608
rect 5776 22423 5874 22521
rect 6201 22423 6299 22521
rect 6633 22423 6731 22521
rect 7015 22400 7113 22498
rect 7287 22400 7385 22498
rect 58643 22400 58741 22498
rect 58915 22400 59013 22498
rect 59297 22423 59395 22521
rect 59729 22423 59827 22521
rect 60154 22423 60252 22521
rect 12008 22232 12068 22292
rect 53960 22232 54020 22292
rect 5776 22049 5874 22147
rect 6201 21991 6299 22089
rect 6633 21991 6731 22089
rect 7015 22005 7113 22103
rect 7287 22005 7385 22103
rect 12008 21995 12068 22055
rect 53960 21995 54020 22055
rect 58643 22005 58741 22103
rect 58915 22005 59013 22103
rect 59297 21991 59395 22089
rect 59729 21991 59827 22089
rect 60154 22049 60252 22147
rect 12008 21758 12068 21818
rect 53960 21758 54020 21818
rect 5776 21633 5874 21731
rect 6201 21633 6299 21731
rect 6633 21633 6731 21731
rect 7015 21610 7113 21708
rect 7287 21610 7385 21708
rect 58643 21610 58741 21708
rect 58915 21610 59013 21708
rect 59297 21633 59395 21731
rect 59729 21633 59827 21731
rect 60154 21633 60252 21731
rect 12008 21442 12068 21502
rect 53960 21442 54020 21502
rect 5776 21259 5874 21357
rect 6201 21201 6299 21299
rect 6633 21201 6731 21299
rect 7015 21215 7113 21313
rect 7287 21215 7385 21313
rect 12008 21205 12068 21265
rect 53960 21205 54020 21265
rect 58643 21215 58741 21313
rect 58915 21215 59013 21313
rect 59297 21201 59395 21299
rect 59729 21201 59827 21299
rect 60154 21259 60252 21357
rect 12008 20968 12068 21028
rect 53960 20968 54020 21028
rect 5776 20843 5874 20941
rect 6201 20843 6299 20941
rect 6633 20843 6731 20941
rect 7015 20820 7113 20918
rect 7287 20820 7385 20918
rect 58643 20820 58741 20918
rect 58915 20820 59013 20918
rect 59297 20843 59395 20941
rect 59729 20843 59827 20941
rect 60154 20843 60252 20941
rect 12008 20652 12068 20712
rect 53960 20652 54020 20712
rect 5776 20469 5874 20567
rect 6201 20411 6299 20509
rect 6633 20411 6731 20509
rect 7015 20425 7113 20523
rect 7287 20425 7385 20523
rect 12008 20415 12068 20475
rect 53960 20415 54020 20475
rect 58643 20425 58741 20523
rect 58915 20425 59013 20523
rect 59297 20411 59395 20509
rect 59729 20411 59827 20509
rect 60154 20469 60252 20567
rect 12008 20178 12068 20238
rect 53960 20178 54020 20238
rect 5776 20053 5874 20151
rect 6201 20053 6299 20151
rect 6633 20053 6731 20151
rect 7015 20030 7113 20128
rect 7287 20030 7385 20128
rect 58643 20030 58741 20128
rect 58915 20030 59013 20128
rect 59297 20053 59395 20151
rect 59729 20053 59827 20151
rect 60154 20053 60252 20151
rect 12008 19862 12068 19922
rect 53960 19862 54020 19922
rect 5776 19679 5874 19777
rect 6201 19621 6299 19719
rect 6633 19621 6731 19719
rect 7015 19635 7113 19733
rect 7287 19635 7385 19733
rect 12008 19625 12068 19685
rect 53960 19625 54020 19685
rect 58643 19635 58741 19733
rect 58915 19635 59013 19733
rect 59297 19621 59395 19719
rect 59729 19621 59827 19719
rect 60154 19679 60252 19777
rect 12008 19388 12068 19448
rect 53960 19388 54020 19448
rect 5776 19263 5874 19361
rect 6201 19263 6299 19361
rect 6633 19263 6731 19361
rect 7015 19240 7113 19338
rect 7287 19240 7385 19338
rect 58643 19240 58741 19338
rect 58915 19240 59013 19338
rect 59297 19263 59395 19361
rect 59729 19263 59827 19361
rect 60154 19263 60252 19361
rect 12008 19072 12068 19132
rect 53960 19072 54020 19132
rect 5776 18889 5874 18987
rect 6201 18831 6299 18929
rect 6633 18831 6731 18929
rect 7015 18845 7113 18943
rect 7287 18845 7385 18943
rect 12008 18835 12068 18895
rect 53960 18835 54020 18895
rect 58643 18845 58741 18943
rect 58915 18845 59013 18943
rect 59297 18831 59395 18929
rect 59729 18831 59827 18929
rect 60154 18889 60252 18987
rect 12008 18598 12068 18658
rect 53960 18598 54020 18658
rect 5776 18473 5874 18571
rect 6201 18473 6299 18571
rect 6633 18473 6731 18571
rect 7015 18450 7113 18548
rect 7287 18450 7385 18548
rect 58643 18450 58741 18548
rect 58915 18450 59013 18548
rect 59297 18473 59395 18571
rect 59729 18473 59827 18571
rect 60154 18473 60252 18571
rect 12008 18282 12068 18342
rect 53960 18282 54020 18342
rect 5776 18099 5874 18197
rect 6201 18041 6299 18139
rect 6633 18041 6731 18139
rect 7015 18055 7113 18153
rect 7287 18055 7385 18153
rect 12008 18045 12068 18105
rect 53960 18045 54020 18105
rect 58643 18055 58741 18153
rect 58915 18055 59013 18153
rect 59297 18041 59395 18139
rect 59729 18041 59827 18139
rect 60154 18099 60252 18197
rect 12008 17808 12068 17868
rect 53960 17808 54020 17868
rect 2486 17683 2584 17781
rect 2911 17683 3009 17781
rect 3343 17683 3441 17781
rect 3725 17660 3823 17758
rect 3997 17660 4095 17758
rect 5776 17683 5874 17781
rect 6201 17683 6299 17781
rect 6633 17683 6731 17781
rect 7015 17660 7113 17758
rect 7287 17660 7385 17758
rect 58643 17660 58741 17758
rect 58915 17660 59013 17758
rect 59297 17683 59395 17781
rect 59729 17683 59827 17781
rect 60154 17683 60252 17781
rect 61933 17660 62031 17758
rect 62205 17660 62303 17758
rect 62587 17683 62685 17781
rect 63019 17683 63117 17781
rect 63444 17683 63542 17781
rect 12008 17492 12068 17552
rect 53960 17492 54020 17552
rect 5776 17309 5874 17407
rect 6201 17251 6299 17349
rect 6633 17251 6731 17349
rect 7015 17265 7113 17363
rect 7287 17265 7385 17363
rect 12008 17255 12068 17315
rect 53960 17255 54020 17315
rect 58643 17265 58741 17363
rect 58915 17265 59013 17363
rect 59297 17251 59395 17349
rect 59729 17251 59827 17349
rect 60154 17309 60252 17407
rect 12008 17018 12068 17078
rect 53960 17018 54020 17078
rect 2486 16893 2584 16991
rect 2911 16893 3009 16991
rect 3343 16893 3441 16991
rect 3725 16870 3823 16968
rect 3997 16870 4095 16968
rect 5776 16893 5874 16991
rect 6201 16893 6299 16991
rect 6633 16893 6731 16991
rect 7015 16870 7113 16968
rect 7287 16870 7385 16968
rect 58643 16870 58741 16968
rect 58915 16870 59013 16968
rect 59297 16893 59395 16991
rect 59729 16893 59827 16991
rect 60154 16893 60252 16991
rect 61933 16870 62031 16968
rect 62205 16870 62303 16968
rect 62587 16893 62685 16991
rect 63019 16893 63117 16991
rect 63444 16893 63542 16991
rect 12008 16702 12068 16762
rect 53960 16702 54020 16762
rect 5776 16519 5874 16617
rect 6201 16461 6299 16559
rect 6633 16461 6731 16559
rect 7015 16475 7113 16573
rect 7287 16475 7385 16573
rect 12008 16465 12068 16525
rect 53960 16465 54020 16525
rect 58643 16475 58741 16573
rect 58915 16475 59013 16573
rect 59297 16461 59395 16559
rect 59729 16461 59827 16559
rect 60154 16519 60252 16617
rect 12008 16228 12068 16288
rect 53960 16228 54020 16288
rect 2486 16103 2584 16201
rect 2911 16103 3009 16201
rect 3343 16103 3441 16201
rect 3725 16080 3823 16178
rect 3997 16080 4095 16178
rect 5776 16103 5874 16201
rect 6201 16103 6299 16201
rect 6633 16103 6731 16201
rect 7015 16080 7113 16178
rect 7287 16080 7385 16178
rect 58643 16080 58741 16178
rect 58915 16080 59013 16178
rect 59297 16103 59395 16201
rect 59729 16103 59827 16201
rect 60154 16103 60252 16201
rect 61933 16080 62031 16178
rect 62205 16080 62303 16178
rect 62587 16103 62685 16201
rect 63019 16103 63117 16201
rect 63444 16103 63542 16201
rect 12008 15912 12068 15972
rect 53960 15912 54020 15972
rect 5776 15729 5874 15827
rect 6201 15671 6299 15769
rect 6633 15671 6731 15769
rect 7015 15685 7113 15783
rect 7287 15685 7385 15783
rect 12008 15675 12068 15735
rect 53960 15675 54020 15735
rect 58643 15685 58741 15783
rect 58915 15685 59013 15783
rect 59297 15671 59395 15769
rect 59729 15671 59827 15769
rect 60154 15729 60252 15827
rect 12008 15438 12068 15498
rect 53960 15438 54020 15498
rect 1155 15290 1253 15388
rect 1427 15290 1525 15388
rect 2486 15313 2584 15411
rect 2911 15313 3009 15411
rect 3343 15313 3441 15411
rect 3725 15290 3823 15388
rect 3997 15290 4095 15388
rect 5776 15313 5874 15411
rect 6201 15313 6299 15411
rect 6633 15313 6731 15411
rect 7015 15290 7113 15388
rect 7287 15290 7385 15388
rect 58643 15290 58741 15388
rect 58915 15290 59013 15388
rect 59297 15313 59395 15411
rect 59729 15313 59827 15411
rect 60154 15313 60252 15411
rect 61933 15290 62031 15388
rect 62205 15290 62303 15388
rect 62587 15313 62685 15411
rect 63019 15313 63117 15411
rect 63444 15313 63542 15411
rect 64503 15290 64601 15388
rect 64775 15290 64873 15388
rect 12008 15122 12068 15182
rect 53960 15122 54020 15182
rect 5776 14939 5874 15037
rect 6201 14881 6299 14979
rect 6633 14881 6731 14979
rect 7015 14895 7113 14993
rect 7287 14895 7385 14993
rect 12008 14885 12068 14945
rect 53960 14885 54020 14945
rect 58643 14895 58741 14993
rect 58915 14895 59013 14993
rect 59297 14881 59395 14979
rect 59729 14881 59827 14979
rect 60154 14939 60252 15037
rect 12008 14648 12068 14708
rect 53960 14648 54020 14708
rect 5776 14523 5874 14621
rect 6201 14523 6299 14621
rect 6633 14523 6731 14621
rect 7015 14500 7113 14598
rect 7287 14500 7385 14598
rect 58643 14500 58741 14598
rect 58915 14500 59013 14598
rect 59297 14523 59395 14621
rect 59729 14523 59827 14621
rect 60154 14523 60252 14621
rect 12008 14332 12068 14392
rect 53960 14332 54020 14392
rect 5776 14149 5874 14247
rect 6201 14091 6299 14189
rect 6633 14091 6731 14189
rect 7015 14105 7113 14203
rect 7287 14105 7385 14203
rect 12008 14095 12068 14155
rect 53960 14095 54020 14155
rect 58643 14105 58741 14203
rect 58915 14105 59013 14203
rect 59297 14091 59395 14189
rect 59729 14091 59827 14189
rect 60154 14149 60252 14247
rect 12008 13858 12068 13918
rect 53960 13858 54020 13918
rect 2921 13717 3019 13815
rect 3346 13717 3444 13815
rect 3725 13710 3823 13808
rect 3997 13710 4095 13808
rect 5776 13733 5874 13831
rect 6201 13733 6299 13831
rect 6633 13733 6731 13831
rect 7015 13710 7113 13808
rect 7287 13710 7385 13808
rect 58643 13710 58741 13808
rect 58915 13710 59013 13808
rect 59297 13733 59395 13831
rect 59729 13733 59827 13831
rect 60154 13733 60252 13831
rect 61933 13710 62031 13808
rect 62205 13710 62303 13808
rect 62584 13717 62682 13815
rect 63009 13717 63107 13815
rect 12008 13542 12068 13602
rect 53960 13542 54020 13602
rect 5776 13359 5874 13457
rect 6201 13301 6299 13399
rect 6633 13301 6731 13399
rect 7015 13315 7113 13413
rect 7287 13315 7385 13413
rect 12008 13305 12068 13365
rect 53960 13305 54020 13365
rect 58643 13315 58741 13413
rect 58915 13315 59013 13413
rect 59297 13301 59395 13399
rect 59729 13301 59827 13399
rect 60154 13359 60252 13457
rect 12008 13068 12068 13128
rect 53960 13068 54020 13128
rect 1751 12920 1849 13018
rect 2023 12920 2121 13018
rect 2921 12927 3019 13025
rect 3346 12927 3444 13025
rect 3725 12920 3823 13018
rect 3997 12920 4095 13018
rect 5776 12943 5874 13041
rect 6201 12943 6299 13041
rect 6633 12943 6731 13041
rect 7015 12920 7113 13018
rect 7287 12920 7385 13018
rect 58643 12920 58741 13018
rect 58915 12920 59013 13018
rect 59297 12943 59395 13041
rect 59729 12943 59827 13041
rect 60154 12943 60252 13041
rect 61933 12920 62031 13018
rect 62205 12920 62303 13018
rect 62584 12927 62682 13025
rect 63009 12927 63107 13025
rect 63907 12920 64005 13018
rect 64179 12920 64277 13018
rect 12008 12752 12068 12812
rect 53960 12752 54020 12812
rect 5776 12569 5874 12667
rect 6201 12511 6299 12609
rect 6633 12511 6731 12609
rect 7015 12525 7113 12623
rect 7287 12525 7385 12623
rect 12008 12515 12068 12575
rect 53960 12515 54020 12575
rect 58643 12525 58741 12623
rect 58915 12525 59013 12623
rect 59297 12511 59395 12609
rect 59729 12511 59827 12609
rect 60154 12569 60252 12667
rect 12008 12278 12068 12338
rect 53960 12278 54020 12338
rect 5776 12153 5874 12251
rect 6201 12153 6299 12251
rect 6633 12153 6731 12251
rect 7015 12130 7113 12228
rect 7287 12130 7385 12228
rect 58643 12130 58741 12228
rect 58915 12130 59013 12228
rect 59297 12153 59395 12251
rect 59729 12153 59827 12251
rect 60154 12153 60252 12251
rect 12008 11962 12068 12022
rect 53960 11962 54020 12022
rect 5776 11779 5874 11877
rect 6201 11721 6299 11819
rect 6633 11721 6731 11819
rect 7015 11735 7113 11833
rect 7287 11735 7385 11833
rect 12008 11725 12068 11785
rect 53960 11725 54020 11785
rect 58643 11735 58741 11833
rect 58915 11735 59013 11833
rect 59297 11721 59395 11819
rect 59729 11721 59827 11819
rect 60154 11779 60252 11877
rect 12008 11488 12068 11548
rect 53960 11488 54020 11548
rect 2921 11347 3019 11445
rect 3346 11347 3444 11445
rect 3725 11340 3823 11438
rect 3997 11340 4095 11438
rect 5776 11363 5874 11461
rect 6201 11363 6299 11461
rect 6633 11363 6731 11461
rect 7015 11340 7113 11438
rect 7287 11340 7385 11438
rect 58643 11340 58741 11438
rect 58915 11340 59013 11438
rect 59297 11363 59395 11461
rect 59729 11363 59827 11461
rect 60154 11363 60252 11461
rect 61933 11340 62031 11438
rect 62205 11340 62303 11438
rect 62584 11347 62682 11445
rect 63009 11347 63107 11445
rect 12008 11172 12068 11232
rect 53960 11172 54020 11232
rect 5776 10989 5874 11087
rect 6201 10931 6299 11029
rect 6633 10931 6731 11029
rect 7015 10945 7113 11043
rect 7287 10945 7385 11043
rect 12008 10935 12068 10995
rect 53960 10935 54020 10995
rect 58643 10945 58741 11043
rect 58915 10945 59013 11043
rect 59297 10931 59395 11029
rect 59729 10931 59827 11029
rect 60154 10989 60252 11087
rect 12008 10698 12068 10758
rect 53960 10698 54020 10758
rect 1751 10550 1849 10648
rect 2023 10550 2121 10648
rect 2921 10557 3019 10655
rect 3346 10557 3444 10655
rect 3725 10550 3823 10648
rect 3997 10550 4095 10648
rect 5776 10573 5874 10671
rect 6201 10573 6299 10671
rect 6633 10573 6731 10671
rect 7015 10550 7113 10648
rect 7287 10550 7385 10648
rect 58643 10550 58741 10648
rect 58915 10550 59013 10648
rect 59297 10573 59395 10671
rect 59729 10573 59827 10671
rect 60154 10573 60252 10671
rect 61933 10550 62031 10648
rect 62205 10550 62303 10648
rect 62584 10557 62682 10655
rect 63009 10557 63107 10655
rect 63907 10550 64005 10648
rect 64179 10550 64277 10648
rect 12008 10382 12068 10442
rect 53960 10382 54020 10442
rect 12008 10145 12068 10205
rect 53960 10145 54020 10205
rect 12008 9908 12068 9968
rect 53960 9908 54020 9968
rect 12685 9565 12783 9663
rect 13328 9584 13388 9644
rect 13952 9584 14012 9644
rect 14576 9584 14636 9644
rect 15200 9584 15260 9644
rect 15824 9584 15884 9644
rect 16448 9584 16508 9644
rect 17072 9584 17132 9644
rect 17696 9584 17756 9644
rect 18320 9584 18380 9644
rect 18944 9584 19004 9644
rect 19568 9584 19628 9644
rect 20192 9584 20252 9644
rect 20816 9584 20876 9644
rect 21440 9584 21500 9644
rect 22064 9584 22124 9644
rect 22688 9584 22748 9644
rect 23312 9584 23372 9644
rect 23936 9584 23996 9644
rect 24560 9584 24620 9644
rect 25184 9584 25244 9644
rect 25808 9584 25868 9644
rect 26432 9584 26492 9644
rect 27056 9584 27116 9644
rect 27680 9584 27740 9644
rect 28304 9584 28364 9644
rect 28928 9584 28988 9644
rect 29552 9584 29612 9644
rect 30176 9584 30236 9644
rect 30800 9584 30860 9644
rect 31424 9584 31484 9644
rect 32048 9584 32108 9644
rect 32672 9584 32732 9644
rect 33296 9584 33356 9644
rect 33920 9584 33980 9644
rect 34544 9584 34604 9644
rect 35168 9584 35228 9644
rect 35792 9584 35852 9644
rect 36416 9584 36476 9644
rect 37040 9584 37100 9644
rect 37664 9584 37724 9644
rect 38288 9584 38348 9644
rect 38912 9584 38972 9644
rect 39536 9584 39596 9644
rect 40160 9584 40220 9644
rect 40784 9584 40844 9644
rect 41408 9584 41468 9644
rect 42032 9584 42092 9644
rect 42656 9584 42716 9644
rect 43280 9584 43340 9644
rect 43904 9584 43964 9644
rect 44528 9584 44588 9644
rect 45152 9584 45212 9644
rect 45776 9584 45836 9644
rect 46400 9584 46460 9644
rect 47024 9584 47084 9644
rect 47648 9584 47708 9644
rect 48272 9584 48332 9644
rect 48896 9584 48956 9644
rect 49520 9584 49580 9644
rect 50144 9584 50204 9644
rect 50768 9584 50828 9644
rect 51392 9584 51452 9644
rect 52016 9584 52076 9644
rect 52640 9584 52700 9644
rect 53245 9565 53343 9663
rect 12804 8974 12902 9072
rect 13190 8974 13288 9072
rect 14052 8974 14150 9072
rect 14438 8974 14536 9072
rect 15300 8974 15398 9072
rect 15686 8974 15784 9072
rect 16548 8974 16646 9072
rect 16934 8974 17032 9072
rect 17796 8974 17894 9072
rect 18182 8974 18280 9072
rect 19044 8974 19142 9072
rect 19430 8974 19528 9072
rect 20292 8974 20390 9072
rect 20678 8974 20776 9072
rect 21540 8974 21638 9072
rect 21926 8974 22024 9072
rect 22788 8974 22886 9072
rect 23174 8974 23272 9072
rect 24036 8974 24134 9072
rect 24422 8974 24520 9072
rect 25284 8974 25382 9072
rect 25670 8974 25768 9072
rect 26532 8974 26630 9072
rect 26918 8974 27016 9072
rect 27780 8974 27878 9072
rect 28166 8974 28264 9072
rect 29028 8974 29126 9072
rect 29414 8974 29512 9072
rect 30276 8974 30374 9072
rect 30662 8974 30760 9072
rect 31524 8974 31622 9072
rect 31910 8974 32008 9072
rect 32772 8974 32870 9072
rect 33158 8974 33256 9072
rect 34020 8974 34118 9072
rect 34406 8974 34504 9072
rect 35268 8974 35366 9072
rect 35654 8974 35752 9072
rect 36516 8974 36614 9072
rect 36902 8974 37000 9072
rect 37764 8974 37862 9072
rect 38150 8974 38248 9072
rect 39012 8974 39110 9072
rect 39398 8974 39496 9072
rect 40260 8974 40358 9072
rect 40646 8974 40744 9072
rect 41508 8974 41606 9072
rect 41894 8974 41992 9072
rect 42756 8974 42854 9072
rect 43142 8974 43240 9072
rect 44004 8974 44102 9072
rect 44390 8974 44488 9072
rect 45252 8974 45350 9072
rect 45638 8974 45736 9072
rect 46500 8974 46598 9072
rect 46886 8974 46984 9072
rect 47748 8974 47846 9072
rect 48134 8974 48232 9072
rect 48996 8974 49094 9072
rect 49382 8974 49480 9072
rect 50244 8974 50342 9072
rect 50630 8974 50728 9072
rect 51492 8974 51590 9072
rect 51878 8974 51976 9072
rect 52740 8974 52838 9072
rect 11407 8434 11473 8437
rect 11407 8432 32702 8434
rect 11407 8376 11412 8432
rect 11468 8376 32702 8432
rect 11407 8374 32702 8376
rect 11407 8371 11473 8374
rect 12933 8285 12999 8288
rect 0 8283 12999 8285
rect 0 8227 12938 8283
rect 12994 8227 12999 8283
rect 0 8225 12999 8227
rect 12933 8222 12999 8225
rect 6439 7645 6537 7666
rect 6439 7589 6460 7645
rect 6516 7589 6537 7645
rect 6439 7568 6537 7589
rect 13621 7401 13719 7499
rect 14869 7401 14967 7499
rect 16117 7401 16215 7499
rect 17365 7401 17463 7499
rect 18613 7401 18711 7499
rect 19861 7401 19959 7499
rect 21109 7401 21207 7499
rect 22357 7401 22455 7499
rect 23605 7401 23703 7499
rect 24853 7401 24951 7499
rect 26101 7401 26199 7499
rect 27349 7401 27447 7499
rect 28597 7401 28695 7499
rect 29845 7401 29943 7499
rect 31093 7401 31191 7499
rect 32341 7401 32439 7499
rect 33589 7401 33687 7499
rect 34837 7401 34935 7499
rect 36085 7401 36183 7499
rect 37333 7401 37431 7499
rect 38581 7401 38679 7499
rect 39829 7401 39927 7499
rect 41077 7401 41175 7499
rect 42325 7401 42423 7499
rect 43573 7401 43671 7499
rect 44821 7401 44919 7499
rect 46069 7401 46167 7499
rect 47317 7401 47415 7499
rect 48565 7401 48663 7499
rect 49813 7401 49911 7499
rect 51061 7401 51159 7499
rect 52309 7401 52407 7499
rect 6439 6231 6537 6252
rect 6439 6175 6460 6231
rect 6516 6175 6537 6231
rect 6439 6154 6537 6175
rect 11159 5859 11225 5862
rect 11159 5857 33014 5859
rect 11159 5801 11164 5857
rect 11220 5801 33014 5857
rect 11159 5799 33014 5801
rect 11159 5796 11225 5799
rect 13448 5628 13546 5726
rect 14696 5628 14794 5726
rect 15944 5628 16042 5726
rect 17192 5628 17290 5726
rect 18440 5628 18538 5726
rect 19688 5628 19786 5726
rect 20936 5628 21034 5726
rect 22184 5628 22282 5726
rect 23432 5628 23530 5726
rect 24680 5628 24778 5726
rect 25928 5628 26026 5726
rect 27176 5628 27274 5726
rect 28424 5628 28522 5726
rect 29672 5628 29770 5726
rect 30920 5628 31018 5726
rect 32168 5628 32266 5726
rect 33416 5628 33514 5726
rect 34664 5628 34762 5726
rect 35912 5628 36010 5726
rect 37160 5628 37258 5726
rect 38408 5628 38506 5726
rect 39656 5628 39754 5726
rect 40904 5628 41002 5726
rect 42152 5628 42250 5726
rect 43400 5628 43498 5726
rect 44648 5628 44746 5726
rect 45896 5628 45994 5726
rect 47144 5628 47242 5726
rect 48392 5628 48490 5726
rect 49640 5628 49738 5726
rect 50888 5628 50986 5726
rect 52136 5628 52234 5726
rect 13366 4854 13464 4952
rect 14614 4854 14712 4952
rect 15862 4854 15960 4952
rect 17110 4854 17208 4952
rect 18358 4854 18456 4952
rect 19606 4854 19704 4952
rect 20854 4854 20952 4952
rect 22102 4854 22200 4952
rect 23350 4854 23448 4952
rect 24598 4854 24696 4952
rect 25846 4854 25944 4952
rect 27094 4854 27192 4952
rect 28342 4854 28440 4952
rect 29590 4854 29688 4952
rect 30838 4854 30936 4952
rect 32086 4854 32184 4952
rect 33334 4854 33432 4952
rect 34582 4854 34680 4952
rect 35830 4854 35928 4952
rect 37078 4854 37176 4952
rect 38326 4854 38424 4952
rect 39574 4854 39672 4952
rect 40822 4854 40920 4952
rect 42070 4854 42168 4952
rect 43318 4854 43416 4952
rect 44566 4854 44664 4952
rect 45814 4854 45912 4952
rect 47062 4854 47160 4952
rect 48310 4854 48408 4952
rect 49558 4854 49656 4952
rect 50806 4854 50904 4952
rect 52054 4854 52152 4952
rect 6439 4817 6537 4838
rect 6439 4761 6460 4817
rect 6516 4761 6537 4817
rect 6439 4740 6537 4761
rect 13378 4016 13476 4114
rect 14626 4016 14724 4114
rect 15874 4016 15972 4114
rect 17122 4016 17220 4114
rect 18370 4016 18468 4114
rect 19618 4016 19716 4114
rect 20866 4016 20964 4114
rect 22114 4016 22212 4114
rect 23362 4016 23460 4114
rect 24610 4016 24708 4114
rect 25858 4016 25956 4114
rect 27106 4016 27204 4114
rect 28354 4016 28452 4114
rect 29602 4016 29700 4114
rect 30850 4016 30948 4114
rect 32098 4016 32196 4114
rect 33346 4016 33444 4114
rect 34594 4016 34692 4114
rect 35842 4016 35940 4114
rect 37090 4016 37188 4114
rect 38338 4016 38436 4114
rect 39586 4016 39684 4114
rect 40834 4016 40932 4114
rect 42082 4016 42180 4114
rect 43330 4016 43428 4114
rect 44578 4016 44676 4114
rect 45826 4016 45924 4114
rect 47074 4016 47172 4114
rect 48322 4016 48420 4114
rect 49570 4016 49668 4114
rect 50818 4016 50916 4114
rect 52066 4016 52164 4114
rect 13378 3694 13476 3792
rect 14626 3694 14724 3792
rect 15874 3694 15972 3792
rect 17122 3694 17220 3792
rect 18370 3694 18468 3792
rect 19618 3694 19716 3792
rect 20866 3694 20964 3792
rect 22114 3694 22212 3792
rect 23362 3694 23460 3792
rect 24610 3694 24708 3792
rect 25858 3694 25956 3792
rect 27106 3694 27204 3792
rect 28354 3694 28452 3792
rect 29602 3694 29700 3792
rect 30850 3694 30948 3792
rect 32098 3694 32196 3792
rect 33346 3694 33444 3792
rect 34594 3694 34692 3792
rect 35842 3694 35940 3792
rect 37090 3694 37188 3792
rect 38338 3694 38436 3792
rect 39586 3694 39684 3792
rect 40834 3694 40932 3792
rect 42082 3694 42180 3792
rect 43330 3694 43428 3792
rect 44578 3694 44676 3792
rect 45826 3694 45924 3792
rect 47074 3694 47172 3792
rect 48322 3694 48420 3792
rect 49570 3694 49668 3792
rect 50818 3694 50916 3792
rect 52066 3694 52164 3792
rect 13264 2901 13362 2999
rect 14512 2901 14610 2999
rect 15760 2901 15858 2999
rect 17008 2901 17106 2999
rect 18256 2901 18354 2999
rect 19504 2901 19602 2999
rect 20752 2901 20850 2999
rect 22000 2901 22098 2999
rect 23248 2901 23346 2999
rect 24496 2901 24594 2999
rect 25744 2901 25842 2999
rect 26992 2901 27090 2999
rect 28240 2901 28338 2999
rect 29488 2901 29586 2999
rect 30736 2901 30834 2999
rect 31984 2901 32082 2999
rect 33232 2901 33330 2999
rect 34480 2901 34578 2999
rect 35728 2901 35826 2999
rect 36976 2901 37074 2999
rect 38224 2901 38322 2999
rect 39472 2901 39570 2999
rect 40720 2901 40818 2999
rect 41968 2901 42066 2999
rect 43216 2901 43314 2999
rect 44464 2901 44562 2999
rect 45712 2901 45810 2999
rect 46960 2901 47058 2999
rect 48208 2901 48306 2999
rect 49456 2901 49554 2999
rect 50704 2901 50802 2999
rect 51952 2901 52050 2999
rect 13253 2464 13351 2562
rect 14501 2464 14599 2562
rect 15749 2464 15847 2562
rect 16997 2464 17095 2562
rect 18245 2464 18343 2562
rect 19493 2464 19591 2562
rect 20741 2464 20839 2562
rect 21989 2464 22087 2562
rect 23237 2464 23335 2562
rect 24485 2464 24583 2562
rect 25733 2464 25831 2562
rect 26981 2464 27079 2562
rect 28229 2464 28327 2562
rect 29477 2464 29575 2562
rect 30725 2464 30823 2562
rect 31973 2464 32071 2562
rect 33221 2464 33319 2562
rect 34469 2464 34567 2562
rect 35717 2464 35815 2562
rect 36965 2464 37063 2562
rect 38213 2464 38311 2562
rect 39461 2464 39559 2562
rect 40709 2464 40807 2562
rect 41957 2464 42055 2562
rect 43205 2464 43303 2562
rect 44453 2464 44551 2562
rect 45701 2464 45799 2562
rect 46949 2464 47047 2562
rect 48197 2464 48295 2562
rect 49445 2464 49543 2562
rect 50693 2464 50791 2562
rect 51941 2464 52039 2562
rect 13374 2132 13472 2230
rect 14622 2132 14720 2230
rect 15870 2132 15968 2230
rect 17118 2132 17216 2230
rect 18366 2132 18464 2230
rect 19614 2132 19712 2230
rect 20862 2132 20960 2230
rect 22110 2132 22208 2230
rect 23358 2132 23456 2230
rect 24606 2132 24704 2230
rect 25854 2132 25952 2230
rect 27102 2132 27200 2230
rect 28350 2132 28448 2230
rect 29598 2132 29696 2230
rect 30846 2132 30944 2230
rect 32094 2132 32192 2230
rect 33342 2132 33440 2230
rect 34590 2132 34688 2230
rect 35838 2132 35936 2230
rect 37086 2132 37184 2230
rect 38334 2132 38432 2230
rect 39582 2132 39680 2230
rect 40830 2132 40928 2230
rect 42078 2132 42176 2230
rect 43326 2132 43424 2230
rect 44574 2132 44672 2230
rect 45822 2132 45920 2230
rect 47070 2132 47168 2230
rect 48318 2132 48416 2230
rect 49566 2132 49664 2230
rect 50814 2132 50912 2230
rect 52062 2132 52160 2230
rect 13259 1930 13357 2028
rect 14507 1930 14605 2028
rect 15755 1930 15853 2028
rect 17003 1930 17101 2028
rect 18251 1930 18349 2028
rect 19499 1930 19597 2028
rect 20747 1930 20845 2028
rect 21995 1930 22093 2028
rect 23243 1930 23341 2028
rect 24491 1930 24589 2028
rect 25739 1930 25837 2028
rect 26987 1930 27085 2028
rect 28235 1930 28333 2028
rect 29483 1930 29581 2028
rect 30731 1930 30829 2028
rect 31979 1930 32077 2028
rect 33227 1930 33325 2028
rect 34475 1930 34573 2028
rect 35723 1930 35821 2028
rect 36971 1930 37069 2028
rect 38219 1930 38317 2028
rect 39467 1930 39565 2028
rect 40715 1930 40813 2028
rect 41963 1930 42061 2028
rect 43211 1930 43309 2028
rect 44459 1930 44557 2028
rect 45707 1930 45805 2028
rect 46955 1930 47053 2028
rect 48203 1930 48301 2028
rect 49451 1930 49549 2028
rect 50699 1930 50797 2028
rect 51947 1930 52045 2028
rect 13273 1514 13371 1612
rect 14521 1514 14619 1612
rect 15769 1514 15867 1612
rect 17017 1514 17115 1612
rect 18265 1514 18363 1612
rect 19513 1514 19611 1612
rect 20761 1514 20859 1612
rect 22009 1514 22107 1612
rect 23257 1514 23355 1612
rect 24505 1514 24603 1612
rect 25753 1514 25851 1612
rect 27001 1514 27099 1612
rect 28249 1514 28347 1612
rect 29497 1514 29595 1612
rect 30745 1514 30843 1612
rect 31993 1514 32091 1612
rect 33241 1514 33339 1612
rect 34489 1514 34587 1612
rect 35737 1514 35835 1612
rect 36985 1514 37083 1612
rect 38233 1514 38331 1612
rect 39481 1514 39579 1612
rect 40729 1514 40827 1612
rect 41977 1514 42075 1612
rect 43225 1514 43323 1612
rect 44473 1514 44571 1612
rect 45721 1514 45819 1612
rect 46969 1514 47067 1612
rect 48217 1514 48315 1612
rect 49465 1514 49563 1612
rect 50713 1514 50811 1612
rect 51961 1514 52059 1612
rect 13370 1071 13468 1169
rect 23354 1071 23452 1169
rect 33338 1071 33436 1169
rect 43322 1071 43420 1169
rect 11283 548 11349 551
rect 11283 546 33014 548
rect 11283 490 11288 546
rect 11344 490 33014 546
rect 11283 488 33014 490
rect 11283 485 11349 488
rect 13370 -49 13468 49
rect 23354 -49 23452 49
rect 33338 -49 33436 49
rect 43322 -49 43420 49
use contact_7  contact_7_0
timestamp 1649977179
transform 1 0 6459 0 1 7584
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1649977179
transform 1 0 6459 0 1 4756
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1649977179
transform 1 0 6459 0 1 6170
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1649977179
transform 1 0 59387 0 1 63260
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1649977179
transform 1 0 59387 0 1 66088
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1649977179
transform 1 0 59387 0 1 64674
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1649977179
transform 1 0 12934 0 1 8223
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1649977179
transform 1 0 6456 0 1 7585
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1649977179
transform 1 0 6456 0 1 4757
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1649977179
transform 1 0 6456 0 1 6171
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1649977179
transform 1 0 11532 0 1 9639
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1649977179
transform 1 0 7564 0 1 9639
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1649977179
transform 1 0 59384 0 1 63261
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1649977179
transform 1 0 59384 0 1 66089
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1649977179
transform 1 0 59384 0 1 64675
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1649977179
transform 1 0 54336 0 1 61207
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1649977179
transform 1 0 58400 0 1 61207
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1649977179
transform 1 0 53030 0 1 62623
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1649977179
transform 1 0 12933 0 1 8218
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1649977179
transform 1 0 6455 0 1 7580
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1649977179
transform 1 0 6455 0 1 4752
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1649977179
transform 1 0 6455 0 1 6166
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1649977179
transform 1 0 11159 0 1 5792
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1649977179
transform 1 0 11283 0 1 481
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1649977179
transform 1 0 11407 0 1 8367
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1649977179
transform 1 0 59383 0 1 63256
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1649977179
transform 1 0 59383 0 1 66084
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1649977179
transform 1 0 59383 0 1 64670
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1649977179
transform 1 0 54583 0 1 65044
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1649977179
transform 1 0 54459 0 1 62469
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1649977179
transform 1 0 53029 0 1 62618
box 0 0 1 1
use contact_28  contact_28_0
timestamp 1649977179
transform 1 0 54197 0 1 11859
box 0 0 1 1
use contact_28  contact_28_1
timestamp 1649977179
transform 1 0 54197 0 1 11605
box 0 0 1 1
use contact_28  contact_28_2
timestamp 1649977179
transform 1 0 54197 0 1 11069
box 0 0 1 1
use contact_28  contact_28_3
timestamp 1649977179
transform 1 0 54197 0 1 10815
box 0 0 1 1
use contact_28  contact_28_4
timestamp 1649977179
transform 1 0 54197 0 1 10279
box 0 0 1 1
use contact_28  contact_28_5
timestamp 1649977179
transform 1 0 54197 0 1 16599
box 0 0 1 1
use contact_28  contact_28_6
timestamp 1649977179
transform 1 0 54197 0 1 16345
box 0 0 1 1
use contact_28  contact_28_7
timestamp 1649977179
transform 1 0 54197 0 1 15809
box 0 0 1 1
use contact_28  contact_28_8
timestamp 1649977179
transform 1 0 54197 0 1 15555
box 0 0 1 1
use contact_28  contact_28_9
timestamp 1649977179
transform 1 0 54197 0 1 15019
box 0 0 1 1
use contact_28  contact_28_10
timestamp 1649977179
transform 1 0 54197 0 1 14765
box 0 0 1 1
use contact_28  contact_28_11
timestamp 1649977179
transform 1 0 54197 0 1 14229
box 0 0 1 1
use contact_28  contact_28_12
timestamp 1649977179
transform 1 0 54197 0 1 13975
box 0 0 1 1
use contact_28  contact_28_13
timestamp 1649977179
transform 1 0 54197 0 1 13439
box 0 0 1 1
use contact_28  contact_28_14
timestamp 1649977179
transform 1 0 54197 0 1 13185
box 0 0 1 1
use contact_28  contact_28_15
timestamp 1649977179
transform 1 0 54197 0 1 12649
box 0 0 1 1
use contact_28  contact_28_16
timestamp 1649977179
transform 1 0 54197 0 1 12395
box 0 0 1 1
use contact_28  contact_28_17
timestamp 1649977179
transform 1 0 54197 0 1 18715
box 0 0 1 1
use contact_28  contact_28_18
timestamp 1649977179
transform 1 0 54197 0 1 18179
box 0 0 1 1
use contact_28  contact_28_19
timestamp 1649977179
transform 1 0 54197 0 1 17925
box 0 0 1 1
use contact_28  contact_28_20
timestamp 1649977179
transform 1 0 54197 0 1 17389
box 0 0 1 1
use contact_28  contact_28_21
timestamp 1649977179
transform 1 0 54197 0 1 17135
box 0 0 1 1
use contact_28  contact_28_22
timestamp 1649977179
transform 1 0 54197 0 1 33189
box 0 0 1 1
use contact_28  contact_28_23
timestamp 1649977179
transform 1 0 54197 0 1 32935
box 0 0 1 1
use contact_28  contact_28_24
timestamp 1649977179
transform 1 0 54197 0 1 32399
box 0 0 1 1
use contact_28  contact_28_25
timestamp 1649977179
transform 1 0 54197 0 1 32145
box 0 0 1 1
use contact_28  contact_28_26
timestamp 1649977179
transform 1 0 54197 0 1 31609
box 0 0 1 1
use contact_28  contact_28_27
timestamp 1649977179
transform 1 0 54197 0 1 31355
box 0 0 1 1
use contact_28  contact_28_28
timestamp 1649977179
transform 1 0 54197 0 1 30819
box 0 0 1 1
use contact_28  contact_28_29
timestamp 1649977179
transform 1 0 54197 0 1 30565
box 0 0 1 1
use contact_28  contact_28_30
timestamp 1649977179
transform 1 0 54197 0 1 30029
box 0 0 1 1
use contact_28  contact_28_31
timestamp 1649977179
transform 1 0 54197 0 1 29775
box 0 0 1 1
use contact_28  contact_28_32
timestamp 1649977179
transform 1 0 54197 0 1 29239
box 0 0 1 1
use contact_28  contact_28_33
timestamp 1649977179
transform 1 0 54197 0 1 28985
box 0 0 1 1
use contact_28  contact_28_34
timestamp 1649977179
transform 1 0 54197 0 1 28449
box 0 0 1 1
use contact_28  contact_28_35
timestamp 1649977179
transform 1 0 54197 0 1 28195
box 0 0 1 1
use contact_28  contact_28_36
timestamp 1649977179
transform 1 0 54197 0 1 27659
box 0 0 1 1
use contact_28  contact_28_37
timestamp 1649977179
transform 1 0 54197 0 1 27405
box 0 0 1 1
use contact_28  contact_28_38
timestamp 1649977179
transform 1 0 54197 0 1 26869
box 0 0 1 1
use contact_28  contact_28_39
timestamp 1649977179
transform 1 0 54197 0 1 26615
box 0 0 1 1
use contact_28  contact_28_40
timestamp 1649977179
transform 1 0 54197 0 1 26079
box 0 0 1 1
use contact_28  contact_28_41
timestamp 1649977179
transform 1 0 54197 0 1 25825
box 0 0 1 1
use contact_28  contact_28_42
timestamp 1649977179
transform 1 0 54197 0 1 25289
box 0 0 1 1
use contact_28  contact_28_43
timestamp 1649977179
transform 1 0 54197 0 1 25035
box 0 0 1 1
use contact_28  contact_28_44
timestamp 1649977179
transform 1 0 54197 0 1 24499
box 0 0 1 1
use contact_28  contact_28_45
timestamp 1649977179
transform 1 0 54197 0 1 24245
box 0 0 1 1
use contact_28  contact_28_46
timestamp 1649977179
transform 1 0 54197 0 1 23709
box 0 0 1 1
use contact_28  contact_28_47
timestamp 1649977179
transform 1 0 54197 0 1 23455
box 0 0 1 1
use contact_28  contact_28_48
timestamp 1649977179
transform 1 0 54197 0 1 22919
box 0 0 1 1
use contact_28  contact_28_49
timestamp 1649977179
transform 1 0 54197 0 1 22665
box 0 0 1 1
use contact_28  contact_28_50
timestamp 1649977179
transform 1 0 54197 0 1 22129
box 0 0 1 1
use contact_28  contact_28_51
timestamp 1649977179
transform 1 0 54197 0 1 21875
box 0 0 1 1
use contact_28  contact_28_52
timestamp 1649977179
transform 1 0 54197 0 1 21339
box 0 0 1 1
use contact_28  contact_28_53
timestamp 1649977179
transform 1 0 54197 0 1 21085
box 0 0 1 1
use contact_28  contact_28_54
timestamp 1649977179
transform 1 0 54197 0 1 20549
box 0 0 1 1
use contact_28  contact_28_55
timestamp 1649977179
transform 1 0 54197 0 1 20295
box 0 0 1 1
use contact_28  contact_28_56
timestamp 1649977179
transform 1 0 54197 0 1 19759
box 0 0 1 1
use contact_28  contact_28_57
timestamp 1649977179
transform 1 0 54197 0 1 19505
box 0 0 1 1
use contact_28  contact_28_58
timestamp 1649977179
transform 1 0 54197 0 1 18969
box 0 0 1 1
use contact_28  contact_28_59
timestamp 1649977179
transform 1 0 11765 0 1 16125
box 0 0 1 1
use contact_28  contact_28_60
timestamp 1649977179
transform 1 0 11765 0 1 16029
box 0 0 1 1
use contact_28  contact_28_61
timestamp 1649977179
transform 1 0 11765 0 1 15335
box 0 0 1 1
use contact_28  contact_28_62
timestamp 1649977179
transform 1 0 11765 0 1 15239
box 0 0 1 1
use contact_28  contact_28_63
timestamp 1649977179
transform 1 0 11765 0 1 14545
box 0 0 1 1
use contact_28  contact_28_64
timestamp 1649977179
transform 1 0 11765 0 1 14449
box 0 0 1 1
use contact_28  contact_28_65
timestamp 1649977179
transform 1 0 11765 0 1 13755
box 0 0 1 1
use contact_28  contact_28_66
timestamp 1649977179
transform 1 0 11765 0 1 13659
box 0 0 1 1
use contact_28  contact_28_67
timestamp 1649977179
transform 1 0 11765 0 1 12965
box 0 0 1 1
use contact_28  contact_28_68
timestamp 1649977179
transform 1 0 11765 0 1 12869
box 0 0 1 1
use contact_28  contact_28_69
timestamp 1649977179
transform 1 0 11765 0 1 12175
box 0 0 1 1
use contact_28  contact_28_70
timestamp 1649977179
transform 1 0 11765 0 1 12079
box 0 0 1 1
use contact_28  contact_28_71
timestamp 1649977179
transform 1 0 11765 0 1 11385
box 0 0 1 1
use contact_28  contact_28_72
timestamp 1649977179
transform 1 0 11765 0 1 11289
box 0 0 1 1
use contact_28  contact_28_73
timestamp 1649977179
transform 1 0 11765 0 1 10595
box 0 0 1 1
use contact_28  contact_28_74
timestamp 1649977179
transform 1 0 11765 0 1 10499
box 0 0 1 1
use contact_28  contact_28_75
timestamp 1649977179
transform 1 0 11765 0 1 16915
box 0 0 1 1
use contact_28  contact_28_76
timestamp 1649977179
transform 1 0 11765 0 1 16819
box 0 0 1 1
use contact_28  contact_28_77
timestamp 1649977179
transform 1 0 11765 0 1 33505
box 0 0 1 1
use contact_28  contact_28_78
timestamp 1649977179
transform 1 0 11765 0 1 33409
box 0 0 1 1
use contact_28  contact_28_79
timestamp 1649977179
transform 1 0 11765 0 1 32715
box 0 0 1 1
use contact_28  contact_28_80
timestamp 1649977179
transform 1 0 11765 0 1 32619
box 0 0 1 1
use contact_28  contact_28_81
timestamp 1649977179
transform 1 0 11765 0 1 31925
box 0 0 1 1
use contact_28  contact_28_82
timestamp 1649977179
transform 1 0 11765 0 1 31829
box 0 0 1 1
use contact_28  contact_28_83
timestamp 1649977179
transform 1 0 11765 0 1 31135
box 0 0 1 1
use contact_28  contact_28_84
timestamp 1649977179
transform 1 0 11765 0 1 31039
box 0 0 1 1
use contact_28  contact_28_85
timestamp 1649977179
transform 1 0 11765 0 1 30345
box 0 0 1 1
use contact_28  contact_28_86
timestamp 1649977179
transform 1 0 11765 0 1 30249
box 0 0 1 1
use contact_28  contact_28_87
timestamp 1649977179
transform 1 0 11765 0 1 29555
box 0 0 1 1
use contact_28  contact_28_88
timestamp 1649977179
transform 1 0 11765 0 1 29459
box 0 0 1 1
use contact_28  contact_28_89
timestamp 1649977179
transform 1 0 11765 0 1 28765
box 0 0 1 1
use contact_28  contact_28_90
timestamp 1649977179
transform 1 0 11765 0 1 28669
box 0 0 1 1
use contact_28  contact_28_91
timestamp 1649977179
transform 1 0 11765 0 1 27975
box 0 0 1 1
use contact_28  contact_28_92
timestamp 1649977179
transform 1 0 11765 0 1 27879
box 0 0 1 1
use contact_28  contact_28_93
timestamp 1649977179
transform 1 0 11765 0 1 27185
box 0 0 1 1
use contact_28  contact_28_94
timestamp 1649977179
transform 1 0 11765 0 1 27089
box 0 0 1 1
use contact_28  contact_28_95
timestamp 1649977179
transform 1 0 11765 0 1 26395
box 0 0 1 1
use contact_28  contact_28_96
timestamp 1649977179
transform 1 0 11765 0 1 26299
box 0 0 1 1
use contact_28  contact_28_97
timestamp 1649977179
transform 1 0 11765 0 1 25605
box 0 0 1 1
use contact_28  contact_28_98
timestamp 1649977179
transform 1 0 11765 0 1 25509
box 0 0 1 1
use contact_28  contact_28_99
timestamp 1649977179
transform 1 0 11765 0 1 24815
box 0 0 1 1
use contact_28  contact_28_100
timestamp 1649977179
transform 1 0 11765 0 1 24719
box 0 0 1 1
use contact_28  contact_28_101
timestamp 1649977179
transform 1 0 11765 0 1 24025
box 0 0 1 1
use contact_28  contact_28_102
timestamp 1649977179
transform 1 0 11765 0 1 23929
box 0 0 1 1
use contact_28  contact_28_103
timestamp 1649977179
transform 1 0 11765 0 1 23235
box 0 0 1 1
use contact_28  contact_28_104
timestamp 1649977179
transform 1 0 11765 0 1 23139
box 0 0 1 1
use contact_28  contact_28_105
timestamp 1649977179
transform 1 0 11765 0 1 22445
box 0 0 1 1
use contact_28  contact_28_106
timestamp 1649977179
transform 1 0 11765 0 1 22349
box 0 0 1 1
use contact_28  contact_28_107
timestamp 1649977179
transform 1 0 11765 0 1 21655
box 0 0 1 1
use contact_28  contact_28_108
timestamp 1649977179
transform 1 0 11765 0 1 21559
box 0 0 1 1
use contact_28  contact_28_109
timestamp 1649977179
transform 1 0 11765 0 1 20865
box 0 0 1 1
use contact_28  contact_28_110
timestamp 1649977179
transform 1 0 11765 0 1 20769
box 0 0 1 1
use contact_28  contact_28_111
timestamp 1649977179
transform 1 0 11765 0 1 20075
box 0 0 1 1
use contact_28  contact_28_112
timestamp 1649977179
transform 1 0 11765 0 1 19979
box 0 0 1 1
use contact_28  contact_28_113
timestamp 1649977179
transform 1 0 11765 0 1 19285
box 0 0 1 1
use contact_28  contact_28_114
timestamp 1649977179
transform 1 0 11765 0 1 19189
box 0 0 1 1
use contact_28  contact_28_115
timestamp 1649977179
transform 1 0 11765 0 1 18495
box 0 0 1 1
use contact_28  contact_28_116
timestamp 1649977179
transform 1 0 11765 0 1 18399
box 0 0 1 1
use contact_28  contact_28_117
timestamp 1649977179
transform 1 0 11765 0 1 17705
box 0 0 1 1
use contact_28  contact_28_118
timestamp 1649977179
transform 1 0 11765 0 1 17609
box 0 0 1 1
use contact_28  contact_28_119
timestamp 1649977179
transform 1 0 11765 0 1 37359
box 0 0 1 1
use contact_28  contact_28_120
timestamp 1649977179
transform 1 0 11765 0 1 36665
box 0 0 1 1
use contact_28  contact_28_121
timestamp 1649977179
transform 1 0 11765 0 1 36569
box 0 0 1 1
use contact_28  contact_28_122
timestamp 1649977179
transform 1 0 11765 0 1 35875
box 0 0 1 1
use contact_28  contact_28_123
timestamp 1649977179
transform 1 0 11765 0 1 35779
box 0 0 1 1
use contact_28  contact_28_124
timestamp 1649977179
transform 1 0 11765 0 1 35085
box 0 0 1 1
use contact_28  contact_28_125
timestamp 1649977179
transform 1 0 11765 0 1 34989
box 0 0 1 1
use contact_28  contact_28_126
timestamp 1649977179
transform 1 0 11765 0 1 34295
box 0 0 1 1
use contact_28  contact_28_127
timestamp 1649977179
transform 1 0 11765 0 1 34199
box 0 0 1 1
use contact_28  contact_28_128
timestamp 1649977179
transform 1 0 11765 0 1 47629
box 0 0 1 1
use contact_28  contact_28_129
timestamp 1649977179
transform 1 0 11765 0 1 46935
box 0 0 1 1
use contact_28  contact_28_130
timestamp 1649977179
transform 1 0 11765 0 1 46839
box 0 0 1 1
use contact_28  contact_28_131
timestamp 1649977179
transform 1 0 11765 0 1 46145
box 0 0 1 1
use contact_28  contact_28_132
timestamp 1649977179
transform 1 0 11765 0 1 46049
box 0 0 1 1
use contact_28  contact_28_133
timestamp 1649977179
transform 1 0 11765 0 1 45355
box 0 0 1 1
use contact_28  contact_28_134
timestamp 1649977179
transform 1 0 11765 0 1 45259
box 0 0 1 1
use contact_28  contact_28_135
timestamp 1649977179
transform 1 0 11765 0 1 44565
box 0 0 1 1
use contact_28  contact_28_136
timestamp 1649977179
transform 1 0 11765 0 1 44469
box 0 0 1 1
use contact_28  contact_28_137
timestamp 1649977179
transform 1 0 11765 0 1 43775
box 0 0 1 1
use contact_28  contact_28_138
timestamp 1649977179
transform 1 0 11765 0 1 43679
box 0 0 1 1
use contact_28  contact_28_139
timestamp 1649977179
transform 1 0 11765 0 1 42985
box 0 0 1 1
use contact_28  contact_28_140
timestamp 1649977179
transform 1 0 11765 0 1 42889
box 0 0 1 1
use contact_28  contact_28_141
timestamp 1649977179
transform 1 0 11765 0 1 42195
box 0 0 1 1
use contact_28  contact_28_142
timestamp 1649977179
transform 1 0 11765 0 1 42099
box 0 0 1 1
use contact_28  contact_28_143
timestamp 1649977179
transform 1 0 11765 0 1 41405
box 0 0 1 1
use contact_28  contact_28_144
timestamp 1649977179
transform 1 0 11765 0 1 41309
box 0 0 1 1
use contact_28  contact_28_145
timestamp 1649977179
transform 1 0 11765 0 1 40615
box 0 0 1 1
use contact_28  contact_28_146
timestamp 1649977179
transform 1 0 11765 0 1 40519
box 0 0 1 1
use contact_28  contact_28_147
timestamp 1649977179
transform 1 0 11765 0 1 39825
box 0 0 1 1
use contact_28  contact_28_148
timestamp 1649977179
transform 1 0 11765 0 1 39729
box 0 0 1 1
use contact_28  contact_28_149
timestamp 1649977179
transform 1 0 11765 0 1 39035
box 0 0 1 1
use contact_28  contact_28_150
timestamp 1649977179
transform 1 0 11765 0 1 38939
box 0 0 1 1
use contact_28  contact_28_151
timestamp 1649977179
transform 1 0 11765 0 1 38245
box 0 0 1 1
use contact_28  contact_28_152
timestamp 1649977179
transform 1 0 11765 0 1 38149
box 0 0 1 1
use contact_28  contact_28_153
timestamp 1649977179
transform 1 0 11765 0 1 37455
box 0 0 1 1
use contact_28  contact_28_154
timestamp 1649977179
transform 1 0 11765 0 1 50095
box 0 0 1 1
use contact_28  contact_28_155
timestamp 1649977179
transform 1 0 11765 0 1 49999
box 0 0 1 1
use contact_28  contact_28_156
timestamp 1649977179
transform 1 0 11765 0 1 49305
box 0 0 1 1
use contact_28  contact_28_157
timestamp 1649977179
transform 1 0 11765 0 1 49209
box 0 0 1 1
use contact_28  contact_28_158
timestamp 1649977179
transform 1 0 11765 0 1 48515
box 0 0 1 1
use contact_28  contact_28_159
timestamp 1649977179
transform 1 0 11765 0 1 48419
box 0 0 1 1
use contact_28  contact_28_160
timestamp 1649977179
transform 1 0 11765 0 1 47725
box 0 0 1 1
use contact_28  contact_28_161
timestamp 1649977179
transform 1 0 11765 0 1 60365
box 0 0 1 1
use contact_28  contact_28_162
timestamp 1649977179
transform 1 0 11765 0 1 60269
box 0 0 1 1
use contact_28  contact_28_163
timestamp 1649977179
transform 1 0 11765 0 1 59575
box 0 0 1 1
use contact_28  contact_28_164
timestamp 1649977179
transform 1 0 11765 0 1 59479
box 0 0 1 1
use contact_28  contact_28_165
timestamp 1649977179
transform 1 0 11765 0 1 58785
box 0 0 1 1
use contact_28  contact_28_166
timestamp 1649977179
transform 1 0 11765 0 1 58689
box 0 0 1 1
use contact_28  contact_28_167
timestamp 1649977179
transform 1 0 11765 0 1 57995
box 0 0 1 1
use contact_28  contact_28_168
timestamp 1649977179
transform 1 0 11765 0 1 57899
box 0 0 1 1
use contact_28  contact_28_169
timestamp 1649977179
transform 1 0 11765 0 1 57205
box 0 0 1 1
use contact_28  contact_28_170
timestamp 1649977179
transform 1 0 11765 0 1 57109
box 0 0 1 1
use contact_28  contact_28_171
timestamp 1649977179
transform 1 0 11765 0 1 56415
box 0 0 1 1
use contact_28  contact_28_172
timestamp 1649977179
transform 1 0 11765 0 1 56319
box 0 0 1 1
use contact_28  contact_28_173
timestamp 1649977179
transform 1 0 11765 0 1 55625
box 0 0 1 1
use contact_28  contact_28_174
timestamp 1649977179
transform 1 0 11765 0 1 55529
box 0 0 1 1
use contact_28  contact_28_175
timestamp 1649977179
transform 1 0 11765 0 1 54835
box 0 0 1 1
use contact_28  contact_28_176
timestamp 1649977179
transform 1 0 11765 0 1 54739
box 0 0 1 1
use contact_28  contact_28_177
timestamp 1649977179
transform 1 0 11765 0 1 54045
box 0 0 1 1
use contact_28  contact_28_178
timestamp 1649977179
transform 1 0 11765 0 1 53949
box 0 0 1 1
use contact_28  contact_28_179
timestamp 1649977179
transform 1 0 11765 0 1 53255
box 0 0 1 1
use contact_28  contact_28_180
timestamp 1649977179
transform 1 0 11765 0 1 53159
box 0 0 1 1
use contact_28  contact_28_181
timestamp 1649977179
transform 1 0 11765 0 1 52465
box 0 0 1 1
use contact_28  contact_28_182
timestamp 1649977179
transform 1 0 11765 0 1 52369
box 0 0 1 1
use contact_28  contact_28_183
timestamp 1649977179
transform 1 0 11765 0 1 51675
box 0 0 1 1
use contact_28  contact_28_184
timestamp 1649977179
transform 1 0 11765 0 1 51579
box 0 0 1 1
use contact_28  contact_28_185
timestamp 1649977179
transform 1 0 11765 0 1 50885
box 0 0 1 1
use contact_28  contact_28_186
timestamp 1649977179
transform 1 0 11765 0 1 50789
box 0 0 1 1
use contact_28  contact_28_187
timestamp 1649977179
transform 1 0 54197 0 1 46365
box 0 0 1 1
use contact_28  contact_28_188
timestamp 1649977179
transform 1 0 54197 0 1 45829
box 0 0 1 1
use contact_28  contact_28_189
timestamp 1649977179
transform 1 0 54197 0 1 45575
box 0 0 1 1
use contact_28  contact_28_190
timestamp 1649977179
transform 1 0 54197 0 1 45039
box 0 0 1 1
use contact_28  contact_28_191
timestamp 1649977179
transform 1 0 54197 0 1 44785
box 0 0 1 1
use contact_28  contact_28_192
timestamp 1649977179
transform 1 0 54197 0 1 44249
box 0 0 1 1
use contact_28  contact_28_193
timestamp 1649977179
transform 1 0 54197 0 1 43995
box 0 0 1 1
use contact_28  contact_28_194
timestamp 1649977179
transform 1 0 54197 0 1 43459
box 0 0 1 1
use contact_28  contact_28_195
timestamp 1649977179
transform 1 0 54197 0 1 43205
box 0 0 1 1
use contact_28  contact_28_196
timestamp 1649977179
transform 1 0 54197 0 1 42669
box 0 0 1 1
use contact_28  contact_28_197
timestamp 1649977179
transform 1 0 54197 0 1 42415
box 0 0 1 1
use contact_28  contact_28_198
timestamp 1649977179
transform 1 0 54197 0 1 41879
box 0 0 1 1
use contact_28  contact_28_199
timestamp 1649977179
transform 1 0 54197 0 1 41625
box 0 0 1 1
use contact_28  contact_28_200
timestamp 1649977179
transform 1 0 54197 0 1 41089
box 0 0 1 1
use contact_28  contact_28_201
timestamp 1649977179
transform 1 0 54197 0 1 40835
box 0 0 1 1
use contact_28  contact_28_202
timestamp 1649977179
transform 1 0 54197 0 1 40299
box 0 0 1 1
use contact_28  contact_28_203
timestamp 1649977179
transform 1 0 54197 0 1 40045
box 0 0 1 1
use contact_28  contact_28_204
timestamp 1649977179
transform 1 0 54197 0 1 39509
box 0 0 1 1
use contact_28  contact_28_205
timestamp 1649977179
transform 1 0 54197 0 1 39255
box 0 0 1 1
use contact_28  contact_28_206
timestamp 1649977179
transform 1 0 54197 0 1 38719
box 0 0 1 1
use contact_28  contact_28_207
timestamp 1649977179
transform 1 0 54197 0 1 38465
box 0 0 1 1
use contact_28  contact_28_208
timestamp 1649977179
transform 1 0 54197 0 1 37929
box 0 0 1 1
use contact_28  contact_28_209
timestamp 1649977179
transform 1 0 54197 0 1 37675
box 0 0 1 1
use contact_28  contact_28_210
timestamp 1649977179
transform 1 0 54197 0 1 37139
box 0 0 1 1
use contact_28  contact_28_211
timestamp 1649977179
transform 1 0 54197 0 1 36885
box 0 0 1 1
use contact_28  contact_28_212
timestamp 1649977179
transform 1 0 54197 0 1 36349
box 0 0 1 1
use contact_28  contact_28_213
timestamp 1649977179
transform 1 0 54197 0 1 36095
box 0 0 1 1
use contact_28  contact_28_214
timestamp 1649977179
transform 1 0 54197 0 1 35559
box 0 0 1 1
use contact_28  contact_28_215
timestamp 1649977179
transform 1 0 54197 0 1 35305
box 0 0 1 1
use contact_28  contact_28_216
timestamp 1649977179
transform 1 0 54197 0 1 34769
box 0 0 1 1
use contact_28  contact_28_217
timestamp 1649977179
transform 1 0 54197 0 1 34515
box 0 0 1 1
use contact_28  contact_28_218
timestamp 1649977179
transform 1 0 54197 0 1 33979
box 0 0 1 1
use contact_28  contact_28_219
timestamp 1649977179
transform 1 0 54197 0 1 33725
box 0 0 1 1
use contact_28  contact_28_220
timestamp 1649977179
transform 1 0 54197 0 1 50315
box 0 0 1 1
use contact_28  contact_28_221
timestamp 1649977179
transform 1 0 54197 0 1 49779
box 0 0 1 1
use contact_28  contact_28_222
timestamp 1649977179
transform 1 0 54197 0 1 49525
box 0 0 1 1
use contact_28  contact_28_223
timestamp 1649977179
transform 1 0 54197 0 1 48989
box 0 0 1 1
use contact_28  contact_28_224
timestamp 1649977179
transform 1 0 54197 0 1 48735
box 0 0 1 1
use contact_28  contact_28_225
timestamp 1649977179
transform 1 0 54197 0 1 48199
box 0 0 1 1
use contact_28  contact_28_226
timestamp 1649977179
transform 1 0 54197 0 1 47945
box 0 0 1 1
use contact_28  contact_28_227
timestamp 1649977179
transform 1 0 54197 0 1 47409
box 0 0 1 1
use contact_28  contact_28_228
timestamp 1649977179
transform 1 0 54197 0 1 47155
box 0 0 1 1
use contact_28  contact_28_229
timestamp 1649977179
transform 1 0 54197 0 1 46619
box 0 0 1 1
use contact_28  contact_28_230
timestamp 1649977179
transform 1 0 54197 0 1 60585
box 0 0 1 1
use contact_28  contact_28_231
timestamp 1649977179
transform 1 0 54197 0 1 60049
box 0 0 1 1
use contact_28  contact_28_232
timestamp 1649977179
transform 1 0 54197 0 1 59795
box 0 0 1 1
use contact_28  contact_28_233
timestamp 1649977179
transform 1 0 54197 0 1 59259
box 0 0 1 1
use contact_28  contact_28_234
timestamp 1649977179
transform 1 0 54197 0 1 59005
box 0 0 1 1
use contact_28  contact_28_235
timestamp 1649977179
transform 1 0 54197 0 1 58469
box 0 0 1 1
use contact_28  contact_28_236
timestamp 1649977179
transform 1 0 54197 0 1 58215
box 0 0 1 1
use contact_28  contact_28_237
timestamp 1649977179
transform 1 0 54197 0 1 57679
box 0 0 1 1
use contact_28  contact_28_238
timestamp 1649977179
transform 1 0 54197 0 1 57425
box 0 0 1 1
use contact_28  contact_28_239
timestamp 1649977179
transform 1 0 54197 0 1 56889
box 0 0 1 1
use contact_28  contact_28_240
timestamp 1649977179
transform 1 0 54197 0 1 56635
box 0 0 1 1
use contact_28  contact_28_241
timestamp 1649977179
transform 1 0 54197 0 1 56099
box 0 0 1 1
use contact_28  contact_28_242
timestamp 1649977179
transform 1 0 54197 0 1 55845
box 0 0 1 1
use contact_28  contact_28_243
timestamp 1649977179
transform 1 0 54197 0 1 55309
box 0 0 1 1
use contact_28  contact_28_244
timestamp 1649977179
transform 1 0 54197 0 1 55055
box 0 0 1 1
use contact_28  contact_28_245
timestamp 1649977179
transform 1 0 54197 0 1 54519
box 0 0 1 1
use contact_28  contact_28_246
timestamp 1649977179
transform 1 0 54197 0 1 54265
box 0 0 1 1
use contact_28  contact_28_247
timestamp 1649977179
transform 1 0 54197 0 1 53729
box 0 0 1 1
use contact_28  contact_28_248
timestamp 1649977179
transform 1 0 54197 0 1 53475
box 0 0 1 1
use contact_28  contact_28_249
timestamp 1649977179
transform 1 0 54197 0 1 52939
box 0 0 1 1
use contact_28  contact_28_250
timestamp 1649977179
transform 1 0 54197 0 1 52685
box 0 0 1 1
use contact_28  contact_28_251
timestamp 1649977179
transform 1 0 54197 0 1 52149
box 0 0 1 1
use contact_28  contact_28_252
timestamp 1649977179
transform 1 0 54197 0 1 51895
box 0 0 1 1
use contact_28  contact_28_253
timestamp 1649977179
transform 1 0 54197 0 1 51359
box 0 0 1 1
use contact_28  contact_28_254
timestamp 1649977179
transform 1 0 54197 0 1 51105
box 0 0 1 1
use contact_28  contact_28_255
timestamp 1649977179
transform 1 0 54197 0 1 50569
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1649977179
transform 1 0 54198 0 1 11602
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1649977179
transform 1 0 54198 0 1 11066
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1649977179
transform 1 0 54198 0 1 10812
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1649977179
transform 1 0 54198 0 1 10276
box 0 0 1 1
use contact_29  contact_29_4
timestamp 1649977179
transform 1 0 54198 0 1 16596
box 0 0 1 1
use contact_29  contact_29_5
timestamp 1649977179
transform 1 0 54198 0 1 16342
box 0 0 1 1
use contact_29  contact_29_6
timestamp 1649977179
transform 1 0 54198 0 1 15806
box 0 0 1 1
use contact_29  contact_29_7
timestamp 1649977179
transform 1 0 54198 0 1 15552
box 0 0 1 1
use contact_29  contact_29_8
timestamp 1649977179
transform 1 0 54198 0 1 15016
box 0 0 1 1
use contact_29  contact_29_9
timestamp 1649977179
transform 1 0 54198 0 1 14762
box 0 0 1 1
use contact_29  contact_29_10
timestamp 1649977179
transform 1 0 54198 0 1 14226
box 0 0 1 1
use contact_29  contact_29_11
timestamp 1649977179
transform 1 0 54198 0 1 13972
box 0 0 1 1
use contact_29  contact_29_12
timestamp 1649977179
transform 1 0 54198 0 1 13436
box 0 0 1 1
use contact_29  contact_29_13
timestamp 1649977179
transform 1 0 54198 0 1 13182
box 0 0 1 1
use contact_29  contact_29_14
timestamp 1649977179
transform 1 0 54198 0 1 12646
box 0 0 1 1
use contact_29  contact_29_15
timestamp 1649977179
transform 1 0 54198 0 1 12392
box 0 0 1 1
use contact_29  contact_29_16
timestamp 1649977179
transform 1 0 54198 0 1 11856
box 0 0 1 1
use contact_29  contact_29_17
timestamp 1649977179
transform 1 0 54198 0 1 18176
box 0 0 1 1
use contact_29  contact_29_18
timestamp 1649977179
transform 1 0 54198 0 1 17922
box 0 0 1 1
use contact_29  contact_29_19
timestamp 1649977179
transform 1 0 54198 0 1 17386
box 0 0 1 1
use contact_29  contact_29_20
timestamp 1649977179
transform 1 0 54198 0 1 17132
box 0 0 1 1
use contact_29  contact_29_21
timestamp 1649977179
transform 1 0 54198 0 1 33186
box 0 0 1 1
use contact_29  contact_29_22
timestamp 1649977179
transform 1 0 54198 0 1 32932
box 0 0 1 1
use contact_29  contact_29_23
timestamp 1649977179
transform 1 0 54198 0 1 32396
box 0 0 1 1
use contact_29  contact_29_24
timestamp 1649977179
transform 1 0 54198 0 1 32142
box 0 0 1 1
use contact_29  contact_29_25
timestamp 1649977179
transform 1 0 54198 0 1 31606
box 0 0 1 1
use contact_29  contact_29_26
timestamp 1649977179
transform 1 0 54198 0 1 31352
box 0 0 1 1
use contact_29  contact_29_27
timestamp 1649977179
transform 1 0 54198 0 1 30816
box 0 0 1 1
use contact_29  contact_29_28
timestamp 1649977179
transform 1 0 54198 0 1 30562
box 0 0 1 1
use contact_29  contact_29_29
timestamp 1649977179
transform 1 0 54198 0 1 30026
box 0 0 1 1
use contact_29  contact_29_30
timestamp 1649977179
transform 1 0 54198 0 1 29772
box 0 0 1 1
use contact_29  contact_29_31
timestamp 1649977179
transform 1 0 54198 0 1 29236
box 0 0 1 1
use contact_29  contact_29_32
timestamp 1649977179
transform 1 0 54198 0 1 28982
box 0 0 1 1
use contact_29  contact_29_33
timestamp 1649977179
transform 1 0 54198 0 1 28446
box 0 0 1 1
use contact_29  contact_29_34
timestamp 1649977179
transform 1 0 54198 0 1 28192
box 0 0 1 1
use contact_29  contact_29_35
timestamp 1649977179
transform 1 0 54198 0 1 27656
box 0 0 1 1
use contact_29  contact_29_36
timestamp 1649977179
transform 1 0 54198 0 1 27402
box 0 0 1 1
use contact_29  contact_29_37
timestamp 1649977179
transform 1 0 54198 0 1 26866
box 0 0 1 1
use contact_29  contact_29_38
timestamp 1649977179
transform 1 0 54198 0 1 26612
box 0 0 1 1
use contact_29  contact_29_39
timestamp 1649977179
transform 1 0 54198 0 1 26076
box 0 0 1 1
use contact_29  contact_29_40
timestamp 1649977179
transform 1 0 54198 0 1 25822
box 0 0 1 1
use contact_29  contact_29_41
timestamp 1649977179
transform 1 0 54198 0 1 25286
box 0 0 1 1
use contact_29  contact_29_42
timestamp 1649977179
transform 1 0 54198 0 1 25032
box 0 0 1 1
use contact_29  contact_29_43
timestamp 1649977179
transform 1 0 54198 0 1 24496
box 0 0 1 1
use contact_29  contact_29_44
timestamp 1649977179
transform 1 0 54198 0 1 24242
box 0 0 1 1
use contact_29  contact_29_45
timestamp 1649977179
transform 1 0 54198 0 1 23706
box 0 0 1 1
use contact_29  contact_29_46
timestamp 1649977179
transform 1 0 54198 0 1 23452
box 0 0 1 1
use contact_29  contact_29_47
timestamp 1649977179
transform 1 0 54198 0 1 22916
box 0 0 1 1
use contact_29  contact_29_48
timestamp 1649977179
transform 1 0 54198 0 1 22662
box 0 0 1 1
use contact_29  contact_29_49
timestamp 1649977179
transform 1 0 54198 0 1 22126
box 0 0 1 1
use contact_29  contact_29_50
timestamp 1649977179
transform 1 0 54198 0 1 21872
box 0 0 1 1
use contact_29  contact_29_51
timestamp 1649977179
transform 1 0 54198 0 1 21336
box 0 0 1 1
use contact_29  contact_29_52
timestamp 1649977179
transform 1 0 54198 0 1 21082
box 0 0 1 1
use contact_29  contact_29_53
timestamp 1649977179
transform 1 0 54198 0 1 20546
box 0 0 1 1
use contact_29  contact_29_54
timestamp 1649977179
transform 1 0 54198 0 1 20292
box 0 0 1 1
use contact_29  contact_29_55
timestamp 1649977179
transform 1 0 54198 0 1 19756
box 0 0 1 1
use contact_29  contact_29_56
timestamp 1649977179
transform 1 0 54198 0 1 19502
box 0 0 1 1
use contact_29  contact_29_57
timestamp 1649977179
transform 1 0 54198 0 1 18966
box 0 0 1 1
use contact_29  contact_29_58
timestamp 1649977179
transform 1 0 54198 0 1 18712
box 0 0 1 1
use contact_29  contact_29_59
timestamp 1649977179
transform 1 0 11766 0 1 16122
box 0 0 1 1
use contact_29  contact_29_60
timestamp 1649977179
transform 1 0 11766 0 1 16026
box 0 0 1 1
use contact_29  contact_29_61
timestamp 1649977179
transform 1 0 11766 0 1 15332
box 0 0 1 1
use contact_29  contact_29_62
timestamp 1649977179
transform 1 0 11766 0 1 15236
box 0 0 1 1
use contact_29  contact_29_63
timestamp 1649977179
transform 1 0 11766 0 1 14542
box 0 0 1 1
use contact_29  contact_29_64
timestamp 1649977179
transform 1 0 11766 0 1 14446
box 0 0 1 1
use contact_29  contact_29_65
timestamp 1649977179
transform 1 0 11766 0 1 13752
box 0 0 1 1
use contact_29  contact_29_66
timestamp 1649977179
transform 1 0 11766 0 1 13656
box 0 0 1 1
use contact_29  contact_29_67
timestamp 1649977179
transform 1 0 11766 0 1 12962
box 0 0 1 1
use contact_29  contact_29_68
timestamp 1649977179
transform 1 0 11766 0 1 12866
box 0 0 1 1
use contact_29  contact_29_69
timestamp 1649977179
transform 1 0 11766 0 1 12172
box 0 0 1 1
use contact_29  contact_29_70
timestamp 1649977179
transform 1 0 11766 0 1 12076
box 0 0 1 1
use contact_29  contact_29_71
timestamp 1649977179
transform 1 0 11766 0 1 11382
box 0 0 1 1
use contact_29  contact_29_72
timestamp 1649977179
transform 1 0 11766 0 1 11286
box 0 0 1 1
use contact_29  contact_29_73
timestamp 1649977179
transform 1 0 11766 0 1 10592
box 0 0 1 1
use contact_29  contact_29_74
timestamp 1649977179
transform 1 0 11766 0 1 10496
box 0 0 1 1
use contact_29  contact_29_75
timestamp 1649977179
transform 1 0 11766 0 1 16816
box 0 0 1 1
use contact_29  contact_29_76
timestamp 1649977179
transform 1 0 11766 0 1 33502
box 0 0 1 1
use contact_29  contact_29_77
timestamp 1649977179
transform 1 0 11766 0 1 33406
box 0 0 1 1
use contact_29  contact_29_78
timestamp 1649977179
transform 1 0 11766 0 1 32712
box 0 0 1 1
use contact_29  contact_29_79
timestamp 1649977179
transform 1 0 11766 0 1 32616
box 0 0 1 1
use contact_29  contact_29_80
timestamp 1649977179
transform 1 0 11766 0 1 31922
box 0 0 1 1
use contact_29  contact_29_81
timestamp 1649977179
transform 1 0 11766 0 1 31826
box 0 0 1 1
use contact_29  contact_29_82
timestamp 1649977179
transform 1 0 11766 0 1 31132
box 0 0 1 1
use contact_29  contact_29_83
timestamp 1649977179
transform 1 0 11766 0 1 31036
box 0 0 1 1
use contact_29  contact_29_84
timestamp 1649977179
transform 1 0 11766 0 1 30342
box 0 0 1 1
use contact_29  contact_29_85
timestamp 1649977179
transform 1 0 11766 0 1 30246
box 0 0 1 1
use contact_29  contact_29_86
timestamp 1649977179
transform 1 0 11766 0 1 29552
box 0 0 1 1
use contact_29  contact_29_87
timestamp 1649977179
transform 1 0 11766 0 1 29456
box 0 0 1 1
use contact_29  contact_29_88
timestamp 1649977179
transform 1 0 11766 0 1 28762
box 0 0 1 1
use contact_29  contact_29_89
timestamp 1649977179
transform 1 0 11766 0 1 28666
box 0 0 1 1
use contact_29  contact_29_90
timestamp 1649977179
transform 1 0 11766 0 1 27972
box 0 0 1 1
use contact_29  contact_29_91
timestamp 1649977179
transform 1 0 11766 0 1 27876
box 0 0 1 1
use contact_29  contact_29_92
timestamp 1649977179
transform 1 0 11766 0 1 27182
box 0 0 1 1
use contact_29  contact_29_93
timestamp 1649977179
transform 1 0 11766 0 1 27086
box 0 0 1 1
use contact_29  contact_29_94
timestamp 1649977179
transform 1 0 11766 0 1 26392
box 0 0 1 1
use contact_29  contact_29_95
timestamp 1649977179
transform 1 0 11766 0 1 26296
box 0 0 1 1
use contact_29  contact_29_96
timestamp 1649977179
transform 1 0 11766 0 1 25602
box 0 0 1 1
use contact_29  contact_29_97
timestamp 1649977179
transform 1 0 11766 0 1 25506
box 0 0 1 1
use contact_29  contact_29_98
timestamp 1649977179
transform 1 0 11766 0 1 24812
box 0 0 1 1
use contact_29  contact_29_99
timestamp 1649977179
transform 1 0 11766 0 1 24716
box 0 0 1 1
use contact_29  contact_29_100
timestamp 1649977179
transform 1 0 11766 0 1 24022
box 0 0 1 1
use contact_29  contact_29_101
timestamp 1649977179
transform 1 0 11766 0 1 23926
box 0 0 1 1
use contact_29  contact_29_102
timestamp 1649977179
transform 1 0 11766 0 1 23232
box 0 0 1 1
use contact_29  contact_29_103
timestamp 1649977179
transform 1 0 11766 0 1 23136
box 0 0 1 1
use contact_29  contact_29_104
timestamp 1649977179
transform 1 0 11766 0 1 22442
box 0 0 1 1
use contact_29  contact_29_105
timestamp 1649977179
transform 1 0 11766 0 1 22346
box 0 0 1 1
use contact_29  contact_29_106
timestamp 1649977179
transform 1 0 11766 0 1 21652
box 0 0 1 1
use contact_29  contact_29_107
timestamp 1649977179
transform 1 0 11766 0 1 21556
box 0 0 1 1
use contact_29  contact_29_108
timestamp 1649977179
transform 1 0 11766 0 1 20862
box 0 0 1 1
use contact_29  contact_29_109
timestamp 1649977179
transform 1 0 11766 0 1 20766
box 0 0 1 1
use contact_29  contact_29_110
timestamp 1649977179
transform 1 0 11766 0 1 20072
box 0 0 1 1
use contact_29  contact_29_111
timestamp 1649977179
transform 1 0 11766 0 1 19976
box 0 0 1 1
use contact_29  contact_29_112
timestamp 1649977179
transform 1 0 11766 0 1 19282
box 0 0 1 1
use contact_29  contact_29_113
timestamp 1649977179
transform 1 0 11766 0 1 19186
box 0 0 1 1
use contact_29  contact_29_114
timestamp 1649977179
transform 1 0 11766 0 1 18492
box 0 0 1 1
use contact_29  contact_29_115
timestamp 1649977179
transform 1 0 11766 0 1 18396
box 0 0 1 1
use contact_29  contact_29_116
timestamp 1649977179
transform 1 0 11766 0 1 17702
box 0 0 1 1
use contact_29  contact_29_117
timestamp 1649977179
transform 1 0 11766 0 1 17606
box 0 0 1 1
use contact_29  contact_29_118
timestamp 1649977179
transform 1 0 11766 0 1 16912
box 0 0 1 1
use contact_29  contact_29_119
timestamp 1649977179
transform 1 0 11766 0 1 37356
box 0 0 1 1
use contact_29  contact_29_120
timestamp 1649977179
transform 1 0 11766 0 1 36662
box 0 0 1 1
use contact_29  contact_29_121
timestamp 1649977179
transform 1 0 11766 0 1 36566
box 0 0 1 1
use contact_29  contact_29_122
timestamp 1649977179
transform 1 0 11766 0 1 35872
box 0 0 1 1
use contact_29  contact_29_123
timestamp 1649977179
transform 1 0 11766 0 1 35776
box 0 0 1 1
use contact_29  contact_29_124
timestamp 1649977179
transform 1 0 11766 0 1 35082
box 0 0 1 1
use contact_29  contact_29_125
timestamp 1649977179
transform 1 0 11766 0 1 34986
box 0 0 1 1
use contact_29  contact_29_126
timestamp 1649977179
transform 1 0 11766 0 1 34292
box 0 0 1 1
use contact_29  contact_29_127
timestamp 1649977179
transform 1 0 11766 0 1 34196
box 0 0 1 1
use contact_29  contact_29_128
timestamp 1649977179
transform 1 0 11766 0 1 47626
box 0 0 1 1
use contact_29  contact_29_129
timestamp 1649977179
transform 1 0 11766 0 1 46932
box 0 0 1 1
use contact_29  contact_29_130
timestamp 1649977179
transform 1 0 11766 0 1 46836
box 0 0 1 1
use contact_29  contact_29_131
timestamp 1649977179
transform 1 0 11766 0 1 46142
box 0 0 1 1
use contact_29  contact_29_132
timestamp 1649977179
transform 1 0 11766 0 1 46046
box 0 0 1 1
use contact_29  contact_29_133
timestamp 1649977179
transform 1 0 11766 0 1 45352
box 0 0 1 1
use contact_29  contact_29_134
timestamp 1649977179
transform 1 0 11766 0 1 45256
box 0 0 1 1
use contact_29  contact_29_135
timestamp 1649977179
transform 1 0 11766 0 1 44562
box 0 0 1 1
use contact_29  contact_29_136
timestamp 1649977179
transform 1 0 11766 0 1 44466
box 0 0 1 1
use contact_29  contact_29_137
timestamp 1649977179
transform 1 0 11766 0 1 43772
box 0 0 1 1
use contact_29  contact_29_138
timestamp 1649977179
transform 1 0 11766 0 1 43676
box 0 0 1 1
use contact_29  contact_29_139
timestamp 1649977179
transform 1 0 11766 0 1 42982
box 0 0 1 1
use contact_29  contact_29_140
timestamp 1649977179
transform 1 0 11766 0 1 42886
box 0 0 1 1
use contact_29  contact_29_141
timestamp 1649977179
transform 1 0 11766 0 1 42192
box 0 0 1 1
use contact_29  contact_29_142
timestamp 1649977179
transform 1 0 11766 0 1 42096
box 0 0 1 1
use contact_29  contact_29_143
timestamp 1649977179
transform 1 0 11766 0 1 41402
box 0 0 1 1
use contact_29  contact_29_144
timestamp 1649977179
transform 1 0 11766 0 1 41306
box 0 0 1 1
use contact_29  contact_29_145
timestamp 1649977179
transform 1 0 11766 0 1 40612
box 0 0 1 1
use contact_29  contact_29_146
timestamp 1649977179
transform 1 0 11766 0 1 40516
box 0 0 1 1
use contact_29  contact_29_147
timestamp 1649977179
transform 1 0 11766 0 1 39822
box 0 0 1 1
use contact_29  contact_29_148
timestamp 1649977179
transform 1 0 11766 0 1 39726
box 0 0 1 1
use contact_29  contact_29_149
timestamp 1649977179
transform 1 0 11766 0 1 39032
box 0 0 1 1
use contact_29  contact_29_150
timestamp 1649977179
transform 1 0 11766 0 1 38936
box 0 0 1 1
use contact_29  contact_29_151
timestamp 1649977179
transform 1 0 11766 0 1 38242
box 0 0 1 1
use contact_29  contact_29_152
timestamp 1649977179
transform 1 0 11766 0 1 38146
box 0 0 1 1
use contact_29  contact_29_153
timestamp 1649977179
transform 1 0 11766 0 1 37452
box 0 0 1 1
use contact_29  contact_29_154
timestamp 1649977179
transform 1 0 11766 0 1 50092
box 0 0 1 1
use contact_29  contact_29_155
timestamp 1649977179
transform 1 0 11766 0 1 49996
box 0 0 1 1
use contact_29  contact_29_156
timestamp 1649977179
transform 1 0 11766 0 1 49302
box 0 0 1 1
use contact_29  contact_29_157
timestamp 1649977179
transform 1 0 11766 0 1 49206
box 0 0 1 1
use contact_29  contact_29_158
timestamp 1649977179
transform 1 0 11766 0 1 48512
box 0 0 1 1
use contact_29  contact_29_159
timestamp 1649977179
transform 1 0 11766 0 1 48416
box 0 0 1 1
use contact_29  contact_29_160
timestamp 1649977179
transform 1 0 11766 0 1 47722
box 0 0 1 1
use contact_29  contact_29_161
timestamp 1649977179
transform 1 0 11766 0 1 60362
box 0 0 1 1
use contact_29  contact_29_162
timestamp 1649977179
transform 1 0 11766 0 1 60266
box 0 0 1 1
use contact_29  contact_29_163
timestamp 1649977179
transform 1 0 11766 0 1 59572
box 0 0 1 1
use contact_29  contact_29_164
timestamp 1649977179
transform 1 0 11766 0 1 59476
box 0 0 1 1
use contact_29  contact_29_165
timestamp 1649977179
transform 1 0 11766 0 1 58782
box 0 0 1 1
use contact_29  contact_29_166
timestamp 1649977179
transform 1 0 11766 0 1 58686
box 0 0 1 1
use contact_29  contact_29_167
timestamp 1649977179
transform 1 0 11766 0 1 57992
box 0 0 1 1
use contact_29  contact_29_168
timestamp 1649977179
transform 1 0 11766 0 1 57896
box 0 0 1 1
use contact_29  contact_29_169
timestamp 1649977179
transform 1 0 11766 0 1 57202
box 0 0 1 1
use contact_29  contact_29_170
timestamp 1649977179
transform 1 0 11766 0 1 57106
box 0 0 1 1
use contact_29  contact_29_171
timestamp 1649977179
transform 1 0 11766 0 1 56412
box 0 0 1 1
use contact_29  contact_29_172
timestamp 1649977179
transform 1 0 11766 0 1 56316
box 0 0 1 1
use contact_29  contact_29_173
timestamp 1649977179
transform 1 0 11766 0 1 55622
box 0 0 1 1
use contact_29  contact_29_174
timestamp 1649977179
transform 1 0 11766 0 1 55526
box 0 0 1 1
use contact_29  contact_29_175
timestamp 1649977179
transform 1 0 11766 0 1 54832
box 0 0 1 1
use contact_29  contact_29_176
timestamp 1649977179
transform 1 0 11766 0 1 54736
box 0 0 1 1
use contact_29  contact_29_177
timestamp 1649977179
transform 1 0 11766 0 1 54042
box 0 0 1 1
use contact_29  contact_29_178
timestamp 1649977179
transform 1 0 11766 0 1 53946
box 0 0 1 1
use contact_29  contact_29_179
timestamp 1649977179
transform 1 0 11766 0 1 53252
box 0 0 1 1
use contact_29  contact_29_180
timestamp 1649977179
transform 1 0 11766 0 1 53156
box 0 0 1 1
use contact_29  contact_29_181
timestamp 1649977179
transform 1 0 11766 0 1 52462
box 0 0 1 1
use contact_29  contact_29_182
timestamp 1649977179
transform 1 0 11766 0 1 52366
box 0 0 1 1
use contact_29  contact_29_183
timestamp 1649977179
transform 1 0 11766 0 1 51672
box 0 0 1 1
use contact_29  contact_29_184
timestamp 1649977179
transform 1 0 11766 0 1 51576
box 0 0 1 1
use contact_29  contact_29_185
timestamp 1649977179
transform 1 0 11766 0 1 50882
box 0 0 1 1
use contact_29  contact_29_186
timestamp 1649977179
transform 1 0 11766 0 1 50786
box 0 0 1 1
use contact_29  contact_29_187
timestamp 1649977179
transform 1 0 54198 0 1 46362
box 0 0 1 1
use contact_29  contact_29_188
timestamp 1649977179
transform 1 0 54198 0 1 45826
box 0 0 1 1
use contact_29  contact_29_189
timestamp 1649977179
transform 1 0 54198 0 1 45572
box 0 0 1 1
use contact_29  contact_29_190
timestamp 1649977179
transform 1 0 54198 0 1 45036
box 0 0 1 1
use contact_29  contact_29_191
timestamp 1649977179
transform 1 0 54198 0 1 44782
box 0 0 1 1
use contact_29  contact_29_192
timestamp 1649977179
transform 1 0 54198 0 1 44246
box 0 0 1 1
use contact_29  contact_29_193
timestamp 1649977179
transform 1 0 54198 0 1 43992
box 0 0 1 1
use contact_29  contact_29_194
timestamp 1649977179
transform 1 0 54198 0 1 43456
box 0 0 1 1
use contact_29  contact_29_195
timestamp 1649977179
transform 1 0 54198 0 1 43202
box 0 0 1 1
use contact_29  contact_29_196
timestamp 1649977179
transform 1 0 54198 0 1 42666
box 0 0 1 1
use contact_29  contact_29_197
timestamp 1649977179
transform 1 0 54198 0 1 42412
box 0 0 1 1
use contact_29  contact_29_198
timestamp 1649977179
transform 1 0 54198 0 1 41876
box 0 0 1 1
use contact_29  contact_29_199
timestamp 1649977179
transform 1 0 54198 0 1 41622
box 0 0 1 1
use contact_29  contact_29_200
timestamp 1649977179
transform 1 0 54198 0 1 41086
box 0 0 1 1
use contact_29  contact_29_201
timestamp 1649977179
transform 1 0 54198 0 1 40832
box 0 0 1 1
use contact_29  contact_29_202
timestamp 1649977179
transform 1 0 54198 0 1 40296
box 0 0 1 1
use contact_29  contact_29_203
timestamp 1649977179
transform 1 0 54198 0 1 40042
box 0 0 1 1
use contact_29  contact_29_204
timestamp 1649977179
transform 1 0 54198 0 1 39506
box 0 0 1 1
use contact_29  contact_29_205
timestamp 1649977179
transform 1 0 54198 0 1 39252
box 0 0 1 1
use contact_29  contact_29_206
timestamp 1649977179
transform 1 0 54198 0 1 38716
box 0 0 1 1
use contact_29  contact_29_207
timestamp 1649977179
transform 1 0 54198 0 1 38462
box 0 0 1 1
use contact_29  contact_29_208
timestamp 1649977179
transform 1 0 54198 0 1 37926
box 0 0 1 1
use contact_29  contact_29_209
timestamp 1649977179
transform 1 0 54198 0 1 37672
box 0 0 1 1
use contact_29  contact_29_210
timestamp 1649977179
transform 1 0 54198 0 1 37136
box 0 0 1 1
use contact_29  contact_29_211
timestamp 1649977179
transform 1 0 54198 0 1 36882
box 0 0 1 1
use contact_29  contact_29_212
timestamp 1649977179
transform 1 0 54198 0 1 36346
box 0 0 1 1
use contact_29  contact_29_213
timestamp 1649977179
transform 1 0 54198 0 1 36092
box 0 0 1 1
use contact_29  contact_29_214
timestamp 1649977179
transform 1 0 54198 0 1 35556
box 0 0 1 1
use contact_29  contact_29_215
timestamp 1649977179
transform 1 0 54198 0 1 35302
box 0 0 1 1
use contact_29  contact_29_216
timestamp 1649977179
transform 1 0 54198 0 1 34766
box 0 0 1 1
use contact_29  contact_29_217
timestamp 1649977179
transform 1 0 54198 0 1 34512
box 0 0 1 1
use contact_29  contact_29_218
timestamp 1649977179
transform 1 0 54198 0 1 33976
box 0 0 1 1
use contact_29  contact_29_219
timestamp 1649977179
transform 1 0 54198 0 1 33722
box 0 0 1 1
use contact_29  contact_29_220
timestamp 1649977179
transform 1 0 54198 0 1 50312
box 0 0 1 1
use contact_29  contact_29_221
timestamp 1649977179
transform 1 0 54198 0 1 49776
box 0 0 1 1
use contact_29  contact_29_222
timestamp 1649977179
transform 1 0 54198 0 1 49522
box 0 0 1 1
use contact_29  contact_29_223
timestamp 1649977179
transform 1 0 54198 0 1 48986
box 0 0 1 1
use contact_29  contact_29_224
timestamp 1649977179
transform 1 0 54198 0 1 48732
box 0 0 1 1
use contact_29  contact_29_225
timestamp 1649977179
transform 1 0 54198 0 1 48196
box 0 0 1 1
use contact_29  contact_29_226
timestamp 1649977179
transform 1 0 54198 0 1 47942
box 0 0 1 1
use contact_29  contact_29_227
timestamp 1649977179
transform 1 0 54198 0 1 47406
box 0 0 1 1
use contact_29  contact_29_228
timestamp 1649977179
transform 1 0 54198 0 1 47152
box 0 0 1 1
use contact_29  contact_29_229
timestamp 1649977179
transform 1 0 54198 0 1 46616
box 0 0 1 1
use contact_29  contact_29_230
timestamp 1649977179
transform 1 0 54198 0 1 60582
box 0 0 1 1
use contact_29  contact_29_231
timestamp 1649977179
transform 1 0 54198 0 1 60046
box 0 0 1 1
use contact_29  contact_29_232
timestamp 1649977179
transform 1 0 54198 0 1 59792
box 0 0 1 1
use contact_29  contact_29_233
timestamp 1649977179
transform 1 0 54198 0 1 59256
box 0 0 1 1
use contact_29  contact_29_234
timestamp 1649977179
transform 1 0 54198 0 1 59002
box 0 0 1 1
use contact_29  contact_29_235
timestamp 1649977179
transform 1 0 54198 0 1 58466
box 0 0 1 1
use contact_29  contact_29_236
timestamp 1649977179
transform 1 0 54198 0 1 58212
box 0 0 1 1
use contact_29  contact_29_237
timestamp 1649977179
transform 1 0 54198 0 1 57676
box 0 0 1 1
use contact_29  contact_29_238
timestamp 1649977179
transform 1 0 54198 0 1 57422
box 0 0 1 1
use contact_29  contact_29_239
timestamp 1649977179
transform 1 0 54198 0 1 56886
box 0 0 1 1
use contact_29  contact_29_240
timestamp 1649977179
transform 1 0 54198 0 1 56632
box 0 0 1 1
use contact_29  contact_29_241
timestamp 1649977179
transform 1 0 54198 0 1 56096
box 0 0 1 1
use contact_29  contact_29_242
timestamp 1649977179
transform 1 0 54198 0 1 55842
box 0 0 1 1
use contact_29  contact_29_243
timestamp 1649977179
transform 1 0 54198 0 1 55306
box 0 0 1 1
use contact_29  contact_29_244
timestamp 1649977179
transform 1 0 54198 0 1 55052
box 0 0 1 1
use contact_29  contact_29_245
timestamp 1649977179
transform 1 0 54198 0 1 54516
box 0 0 1 1
use contact_29  contact_29_246
timestamp 1649977179
transform 1 0 54198 0 1 54262
box 0 0 1 1
use contact_29  contact_29_247
timestamp 1649977179
transform 1 0 54198 0 1 53726
box 0 0 1 1
use contact_29  contact_29_248
timestamp 1649977179
transform 1 0 54198 0 1 53472
box 0 0 1 1
use contact_29  contact_29_249
timestamp 1649977179
transform 1 0 54198 0 1 52936
box 0 0 1 1
use contact_29  contact_29_250
timestamp 1649977179
transform 1 0 54198 0 1 52682
box 0 0 1 1
use contact_29  contact_29_251
timestamp 1649977179
transform 1 0 54198 0 1 52146
box 0 0 1 1
use contact_29  contact_29_252
timestamp 1649977179
transform 1 0 54198 0 1 51892
box 0 0 1 1
use contact_29  contact_29_253
timestamp 1649977179
transform 1 0 54198 0 1 51356
box 0 0 1 1
use contact_29  contact_29_254
timestamp 1649977179
transform 1 0 54198 0 1 51102
box 0 0 1 1
use contact_29  contact_29_255
timestamp 1649977179
transform 1 0 54198 0 1 50566
box 0 0 1 1
use cr_0  cr_0_0
timestamp 1649977179
transform 1 0 11798 0 1 9385
box -4946 -3924 1278 -2440
use cr_1  cr_1_0
timestamp 1649977179
transform 1 0 11798 0 1 9385
box 41154 54580 47254 56064
use pinvbuf  pinvbuf_0
timestamp 1649977179
transform 1 0 5936 0 1 4789
box -36 -17 1140 2845
use pinvbuf  pinvbuf_1
timestamp 1649977179
transform -1 0 59968 0 -1 66121
box -36 -17 1140 2845
use port_address  port_address_0
timestamp 1649977179
transform -1 0 66028 0 1 10175
box 0 -56 11528 50649
use port_address  port_address_1
timestamp 1649977179
transform 1 0 0 0 1 10175
box 0 -56 11528 50649
use port_data_0  port_data_0_0
timestamp 1649977179
transform 1 0 13046 0 1 61525
box -160 238 40560 5750
use port_data  port_data_0
timestamp 1649977179
transform 1 0 12422 0 -1 9385
box 0 238 40560 9434
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1649977179
transform 1 0 11798 0 1 9385
box -42 0 42474 52140
<< labels >>
rlabel locali s 59887 65452 59887 65452 4 addr1_0
port 105 nsew
rlabel locali s 6017 5458 6017 5458 4 addr0_0
port 97 nsew
rlabel metal1 s 49365 67148 49365 67148 4 dout1_29
port 62 nsew
rlabel metal1 s 33141 67148 33141 67148 4 dout1_16
port 49 nsew
rlabel metal1 s 36885 67148 36885 67148 4 dout1_19
port 52 nsew
rlabel metal1 s 40629 67148 40629 67148 4 dout1_22
port 55 nsew
rlabel metal1 s 38133 67148 38133 67148 4 dout1_20
port 53 nsew
rlabel metal1 s 50613 67148 50613 67148 4 dout1_30
port 63 nsew
rlabel metal1 s 46869 67148 46869 67148 4 dout1_27
port 60 nsew
rlabel metal1 s 34389 67148 34389 67148 4 dout1_17
port 50 nsew
rlabel metal1 s 39381 67148 39381 67148 4 dout1_21
port 54 nsew
rlabel metal1 s 35637 67148 35637 67148 4 dout1_18
port 51 nsew
rlabel metal1 s 41877 67148 41877 67148 4 dout1_23
port 56 nsew
rlabel metal1 s 44373 67148 44373 67148 4 dout1_25
port 58 nsew
rlabel metal1 s 48117 67148 48117 67148 4 dout1_28
port 61 nsew
rlabel metal1 s 45621 67148 45621 67148 4 dout1_26
port 59 nsew
rlabel metal1 s 43125 67148 43125 67148 4 dout1_24
port 57 nsew
rlabel metal1 s 51861 67148 51861 67148 4 dout1_31
port 64 nsew
rlabel metal1 s 18165 67148 18165 67148 4 dout1_4
port 37 nsew
rlabel metal1 s 29397 67148 29397 67148 4 dout1_13
port 46 nsew
rlabel metal1 s 20661 67148 20661 67148 4 dout1_6
port 39 nsew
rlabel metal1 s 16917 67148 16917 67148 4 dout1_3
port 36 nsew
rlabel metal1 s 15669 67148 15669 67148 4 dout1_2
port 35 nsew
rlabel metal1 s 30645 67148 30645 67148 4 dout1_14
port 47 nsew
rlabel metal1 s 13173 67148 13173 67148 4 dout1_0
port 33 nsew
rlabel metal1 s 24405 67148 24405 67148 4 dout1_9
port 42 nsew
rlabel metal1 s 25653 67148 25653 67148 4 dout1_10
port 43 nsew
rlabel metal1 s 28149 67148 28149 67148 4 dout1_12
port 45 nsew
rlabel metal1 s 23157 67148 23157 67148 4 dout1_8
port 41 nsew
rlabel metal1 s 21909 67148 21909 67148 4 dout1_7
port 40 nsew
rlabel metal1 s 14421 67148 14421 67148 4 dout1_1
port 34 nsew
rlabel metal1 s 26901 67148 26901 67148 4 dout1_11
port 44 nsew
rlabel metal1 s 31893 67148 31893 67148 4 dout1_15
port 48 nsew
rlabel metal1 s 19413 67148 19413 67148 4 dout1_5
port 38 nsew
rlabel metal1 s 25653 3762 25653 3762 4 dout0_10
port 11 nsew
rlabel metal1 s 23315 1404 23315 1404 4 din0_8
port 73 nsew
rlabel metal1 s 192 14154 192 14154 4 addr0_3
port 100 nsew
rlabel metal1 s 31893 3762 31893 3762 4 dout0_15
port 16 nsew
rlabel metal1 s 29555 1404 29555 1404 4 din0_13
port 78 nsew
rlabel metal1 s 19413 3762 19413 3762 4 dout0_5
port 6 nsew
rlabel metal1 s 30803 1404 30803 1404 4 din0_14
port 79 nsew
rlabel metal1 s 14421 3762 14421 3762 4 dout0_1
port 2 nsew
rlabel metal1 s 13173 3762 13173 3762 4 dout0_0
port 1 nsew
rlabel metal1 s 20661 3762 20661 3762 4 dout0_6
port 7 nsew
rlabel metal1 s 15669 3762 15669 3762 4 dout0_2
port 3 nsew
rlabel metal1 s 30645 3762 30645 3762 4 dout0_14
port 15 nsew
rlabel metal1 s 15827 1404 15827 1404 4 din0_2
port 67 nsew
rlabel metal1 s 20819 1404 20819 1404 4 din0_6
port 71 nsew
rlabel metal1 s 432 14154 432 14154 4 addr0_6
port 103 nsew
rlabel metal1 s 14579 1404 14579 1404 4 din0_1
port 66 nsew
rlabel metal1 s 352 14154 352 14154 4 addr0_5
port 102 nsew
rlabel metal1 s 17075 1404 17075 1404 4 din0_3
port 68 nsew
rlabel metal1 s 18323 1404 18323 1404 4 din0_4
port 69 nsew
rlabel metal1 s 29397 3762 29397 3762 4 dout0_13
port 14 nsew
rlabel metal1 s 32 14154 32 14154 4 addr0_1
port 98 nsew
rlabel metal1 s 13331 1404 13331 1404 4 din0_0
port 65 nsew
rlabel metal1 s 24563 1404 24563 1404 4 din0_9
port 74 nsew
rlabel metal1 s 18165 3762 18165 3762 4 dout0_4
port 5 nsew
rlabel metal1 s 28307 1404 28307 1404 4 din0_12
port 77 nsew
rlabel metal1 s 112 14154 112 14154 4 addr0_2
port 99 nsew
rlabel metal1 s 512 14154 512 14154 4 addr0_7
port 104 nsew
rlabel metal1 s 22067 1404 22067 1404 4 din0_7
port 72 nsew
rlabel metal1 s 25811 1404 25811 1404 4 din0_10
port 75 nsew
rlabel metal1 s 26901 3762 26901 3762 4 dout0_11
port 12 nsew
rlabel metal1 s 19571 1404 19571 1404 4 din0_5
port 70 nsew
rlabel metal1 s 272 14154 272 14154 4 addr0_4
port 101 nsew
rlabel metal1 s 28149 3762 28149 3762 4 dout0_12
port 13 nsew
rlabel metal1 s 27059 1404 27059 1404 4 din0_11
port 76 nsew
rlabel metal1 s 16917 3762 16917 3762 4 dout0_3
port 4 nsew
rlabel metal1 s 24405 3762 24405 3762 4 dout0_9
port 10 nsew
rlabel metal1 s 32051 1404 32051 1404 4 din0_15
port 80 nsew
rlabel metal1 s 21909 3762 21909 3762 4 dout0_7
port 8 nsew
rlabel metal1 s 23157 3762 23157 3762 4 dout0_8
port 9 nsew
rlabel metal1 s 48117 3762 48117 3762 4 dout0_28
port 29 nsew
rlabel metal1 s 45621 3762 45621 3762 4 dout0_26
port 27 nsew
rlabel metal1 s 65916 14154 65916 14154 4 addr1_2
port 107 nsew
rlabel metal1 s 65676 14154 65676 14154 4 addr1_5
port 110 nsew
rlabel metal1 s 38291 1404 38291 1404 4 din0_20
port 85 nsew
rlabel metal1 s 65836 14154 65836 14154 4 addr1_3
port 108 nsew
rlabel metal1 s 65596 14154 65596 14154 4 addr1_6
port 111 nsew
rlabel metal1 s 49365 3762 49365 3762 4 dout0_29
port 30 nsew
rlabel metal1 s 46869 3762 46869 3762 4 dout0_27
port 28 nsew
rlabel metal1 s 37043 1404 37043 1404 4 din0_19
port 84 nsew
rlabel metal1 s 39539 1404 39539 1404 4 din0_21
port 86 nsew
rlabel metal1 s 48275 1404 48275 1404 4 din0_28
port 93 nsew
rlabel metal1 s 34547 1404 34547 1404 4 din0_17
port 82 nsew
rlabel metal1 s 34389 3762 34389 3762 4 dout0_17
port 18 nsew
rlabel metal1 s 40629 3762 40629 3762 4 dout0_22
port 23 nsew
rlabel metal1 s 65516 14154 65516 14154 4 addr1_7
port 112 nsew
rlabel metal1 s 42035 1404 42035 1404 4 din0_23
port 88 nsew
rlabel metal1 s 49523 1404 49523 1404 4 din0_29
port 94 nsew
rlabel metal1 s 35795 1404 35795 1404 4 din0_18
port 83 nsew
rlabel metal1 s 33141 3762 33141 3762 4 dout0_16
port 17 nsew
rlabel metal1 s 38133 3762 38133 3762 4 dout0_20
port 21 nsew
rlabel metal1 s 50771 1404 50771 1404 4 din0_30
port 95 nsew
rlabel metal1 s 36885 3762 36885 3762 4 dout0_19
port 20 nsew
rlabel metal1 s 43125 3762 43125 3762 4 dout0_24
port 25 nsew
rlabel metal1 s 39381 3762 39381 3762 4 dout0_21
port 22 nsew
rlabel metal1 s 50613 3762 50613 3762 4 dout0_30
port 31 nsew
rlabel metal1 s 45779 1404 45779 1404 4 din0_26
port 91 nsew
rlabel metal1 s 40787 1404 40787 1404 4 din0_22
port 87 nsew
rlabel metal1 s 43283 1404 43283 1404 4 din0_24
port 89 nsew
rlabel metal1 s 44531 1404 44531 1404 4 din0_25
port 90 nsew
rlabel metal1 s 35637 3762 35637 3762 4 dout0_18
port 19 nsew
rlabel metal1 s 52019 1404 52019 1404 4 din0_31
port 96 nsew
rlabel metal1 s 44373 3762 44373 3762 4 dout0_25
port 26 nsew
rlabel metal1 s 33299 1404 33299 1404 4 din0_16
port 81 nsew
rlabel metal1 s 47027 1404 47027 1404 4 din0_27
port 92 nsew
rlabel metal1 s 65756 14154 65756 14154 4 addr1_4
port 109 nsew
rlabel metal1 s 51861 3762 51861 3762 4 dout0_31
port 32 nsew
rlabel metal1 s 41877 3762 41877 3762 4 dout0_23
port 24 nsew
rlabel metal1 s 65996 14154 65996 14154 4 addr1_1
port 106 nsew
rlabel metal2 s 13046 270 13046 270 4 bank_wmask0_0
port 118 nsew
rlabel metal2 s 42998 270 42998 270 4 bank_wmask0_3
port 121 nsew
rlabel metal2 s 54616 64127 54616 64127 4 s_en1
port 114 nsew
rlabel metal2 s 11316 5007 11316 5007 4 w_en0
port 117 nsew
rlabel metal2 s 11440 5007 11440 5007 4 p_en_bar0
port 115 nsew
rlabel metal2 s 54368 64127 54368 64127 4 wl_en1
port 123 nsew
rlabel metal2 s 23030 270 23030 270 4 bank_wmask0_1
port 119 nsew
rlabel metal2 s 11564 5007 11564 5007 4 wl_en0
port 122 nsew
rlabel metal2 s 11192 5007 11192 5007 4 s_en0
port 113 nsew
rlabel metal2 s 33014 270 33014 270 4 bank_wmask0_2
port 120 nsew
rlabel metal2 s 54492 64127 54492 64127 4 p_en_bar1
port 116 nsew
rlabel metal3 s 59778 59170 59778 59170 4 vdd
port 124 nsew
rlabel metal3 s 59778 59602 59778 59602 4 vdd
port 124 nsew
rlabel metal3 s 58692 59579 58692 59579 4 vdd
port 124 nsew
rlabel metal3 s 59346 59602 59346 59602 4 vdd
port 124 nsew
rlabel metal3 s 59346 59960 59346 59960 4 vdd
port 124 nsew
rlabel metal3 s 59416 64707 59416 64707 4 vdd
port 124 nsew
rlabel metal3 s 58692 58789 58692 58789 4 vdd
port 124 nsew
rlabel metal3 s 59346 59170 59346 59170 4 vdd
port 124 nsew
rlabel metal3 s 59778 58812 59778 58812 4 vdd
port 124 nsew
rlabel metal3 s 58692 60369 58692 60369 4 vdd
port 124 nsew
rlabel metal3 s 58692 59184 58692 59184 4 vdd
port 124 nsew
rlabel metal3 s 58692 59974 58692 59974 4 vdd
port 124 nsew
rlabel metal3 s 59346 58812 59346 58812 4 vdd
port 124 nsew
rlabel metal3 s 59346 60392 59346 60392 4 vdd
port 124 nsew
rlabel metal3 s 59778 60392 59778 60392 4 vdd
port 124 nsew
rlabel metal3 s 59778 59960 59778 59960 4 vdd
port 124 nsew
rlabel metal3 s 59587 62655 59587 62655 4 rbl_bl1
port 125 nsew
rlabel metal3 s 60203 59602 60203 59602 4 gnd
port 125 nsew
rlabel metal3 s 60203 60392 60203 60392 4 gnd
port 125 nsew
rlabel metal3 s 59416 66121 59416 66121 4 gnd
port 125 nsew
rlabel metal3 s 58964 59974 58964 59974 4 gnd
port 125 nsew
rlabel metal3 s 60203 60018 60203 60018 4 gnd
port 125 nsew
rlabel metal3 s 58964 58789 58964 58789 4 gnd
port 125 nsew
rlabel metal3 s 58964 59184 58964 59184 4 gnd
port 125 nsew
rlabel metal3 s 58964 59579 58964 59579 4 gnd
port 125 nsew
rlabel metal3 s 60203 58812 60203 58812 4 gnd
port 125 nsew
rlabel metal3 s 59416 63293 59416 63293 4 gnd
port 125 nsew
rlabel metal3 s 58964 60369 58964 60369 4 gnd
port 125 nsew
rlabel metal3 s 60203 59228 60203 59228 4 gnd
port 125 nsew
rlabel metal3 s 49045 61887 49045 61887 4 vdd
port 124 nsew
rlabel metal3 s 51422 61296 51422 61296 4 vdd
port 124 nsew
rlabel metal3 s 50855 66007 50855 66007 4 vdd
port 124 nsew
rlabel metal3 s 49431 61887 49431 61887 4 vdd
port 124 nsew
rlabel metal3 s 49619 66845 49619 66845 4 vdd
port 124 nsew
rlabel metal3 s 52789 61887 52789 61887 4 vdd
port 124 nsew
rlabel metal3 s 49550 61296 49550 61296 4 vdd
port 124 nsew
rlabel metal3 s 51541 61887 51541 61887 4 vdd
port 124 nsew
rlabel metal3 s 52670 61296 52670 61296 4 vdd
port 124 nsew
rlabel metal3 s 48926 61296 48926 61296 4 vdd
port 124 nsew
rlabel metal3 s 52046 61296 52046 61296 4 vdd
port 124 nsew
rlabel metal3 s 50867 66845 50867 66845 4 vdd
port 124 nsew
rlabel metal3 s 51927 61887 51927 61887 4 vdd
port 124 nsew
rlabel metal3 s 50937 65233 50937 65233 4 gnd
port 125 nsew
rlabel metal3 s 50174 61296 50174 61296 4 vdd
port 124 nsew
rlabel metal3 s 52103 66007 52103 66007 4 vdd
port 124 nsew
rlabel metal3 s 50679 61887 50679 61887 4 vdd
port 124 nsew
rlabel metal3 s 49862 63460 49862 63460 4 gnd
port 125 nsew
rlabel metal3 s 49607 66007 49607 66007 4 vdd
port 124 nsew
rlabel metal3 s 52115 66845 52115 66845 4 vdd
port 124 nsew
rlabel metal3 s 49689 65233 49689 65233 4 gnd
port 125 nsew
rlabel metal3 s 53990 60972 53990 60972 4 gnd
port 125 nsew
rlabel metal3 s 52115 67167 52115 67167 4 gnd
port 125 nsew
rlabel metal3 s 50867 67167 50867 67167 4 gnd
port 125 nsew
rlabel metal3 s 53990 59155 53990 59155 4 gnd
port 125 nsew
rlabel metal3 s 51110 63460 51110 63460 4 gnd
port 125 nsew
rlabel metal3 s 53990 60735 53990 60735 4 gnd
port 125 nsew
rlabel metal3 s 53175 61887 53175 61887 4 vdd
port 124 nsew
rlabel metal3 s 52185 65233 52185 65233 4 gnd
port 125 nsew
rlabel metal3 s 53990 60182 53990 60182 4 gnd
port 125 nsew
rlabel metal3 s 53990 59392 53990 59392 4 gnd
port 125 nsew
rlabel metal3 s 50293 61887 50293 61887 4 vdd
port 124 nsew
rlabel metal3 s 50798 61296 50798 61296 4 vdd
port 124 nsew
rlabel metal3 s 53294 61296 53294 61296 4 vdd
port 124 nsew
rlabel metal3 s 49619 67167 49619 67167 4 gnd
port 125 nsew
rlabel metal3 s 53990 60498 53990 60498 4 gnd
port 125 nsew
rlabel metal3 s 53990 58918 53990 58918 4 gnd
port 125 nsew
rlabel metal3 s 53990 59945 53990 59945 4 gnd
port 125 nsew
rlabel metal3 s 52358 63460 52358 63460 4 gnd
port 125 nsew
rlabel metal3 s 53990 59708 53990 59708 4 gnd
port 125 nsew
rlabel metal3 s 53990 53862 53990 53862 4 gnd
port 125 nsew
rlabel metal3 s 53990 55995 53990 55995 4 gnd
port 125 nsew
rlabel metal3 s 53990 57338 53990 57338 4 gnd
port 125 nsew
rlabel metal3 s 53990 57812 53990 57812 4 gnd
port 125 nsew
rlabel metal3 s 53990 58128 53990 58128 4 gnd
port 125 nsew
rlabel metal3 s 53990 51255 53990 51255 4 gnd
port 125 nsew
rlabel metal3 s 53990 52835 53990 52835 4 gnd
port 125 nsew
rlabel metal3 s 53990 52282 53990 52282 4 gnd
port 125 nsew
rlabel metal3 s 53990 53625 53990 53625 4 gnd
port 125 nsew
rlabel metal3 s 53990 54178 53990 54178 4 gnd
port 125 nsew
rlabel metal3 s 53990 52045 53990 52045 4 gnd
port 125 nsew
rlabel metal3 s 53990 58365 53990 58365 4 gnd
port 125 nsew
rlabel metal3 s 53990 54415 53990 54415 4 gnd
port 125 nsew
rlabel metal3 s 53990 58602 53990 58602 4 gnd
port 125 nsew
rlabel metal3 s 53990 51808 53990 51808 4 gnd
port 125 nsew
rlabel metal3 s 53990 54652 53990 54652 4 gnd
port 125 nsew
rlabel metal3 s 53990 50702 53990 50702 4 gnd
port 125 nsew
rlabel metal3 s 53990 50465 53990 50465 4 gnd
port 125 nsew
rlabel metal3 s 53990 51492 53990 51492 4 gnd
port 125 nsew
rlabel metal3 s 53990 56548 53990 56548 4 gnd
port 125 nsew
rlabel metal3 s 53990 55758 53990 55758 4 gnd
port 125 nsew
rlabel metal3 s 53990 57575 53990 57575 4 gnd
port 125 nsew
rlabel metal3 s 53990 53388 53990 53388 4 gnd
port 125 nsew
rlabel metal3 s 53990 56232 53990 56232 4 gnd
port 125 nsew
rlabel metal3 s 53990 52598 53990 52598 4 gnd
port 125 nsew
rlabel metal3 s 53990 54968 53990 54968 4 gnd
port 125 nsew
rlabel metal3 s 53990 53072 53990 53072 4 gnd
port 125 nsew
rlabel metal3 s 53990 51018 53990 51018 4 gnd
port 125 nsew
rlabel metal3 s 53990 55442 53990 55442 4 gnd
port 125 nsew
rlabel metal3 s 53990 56785 53990 56785 4 gnd
port 125 nsew
rlabel metal3 s 53990 57022 53990 57022 4 gnd
port 125 nsew
rlabel metal3 s 53990 55205 53990 55205 4 gnd
port 125 nsew
rlabel metal3 s 60203 57648 60203 57648 4 gnd
port 125 nsew
rlabel metal3 s 59346 55652 59346 55652 4 vdd
port 124 nsew
rlabel metal3 s 60203 58438 60203 58438 4 gnd
port 125 nsew
rlabel metal3 s 58964 57209 58964 57209 4 gnd
port 125 nsew
rlabel metal3 s 59346 57590 59346 57590 4 vdd
port 124 nsew
rlabel metal3 s 59778 56800 59778 56800 4 vdd
port 124 nsew
rlabel metal3 s 58964 55234 58964 55234 4 gnd
port 125 nsew
rlabel metal3 s 59778 58022 59778 58022 4 vdd
port 124 nsew
rlabel metal3 s 58692 57604 58692 57604 4 vdd
port 124 nsew
rlabel metal3 s 60203 56442 60203 56442 4 gnd
port 125 nsew
rlabel metal3 s 58692 56024 58692 56024 4 vdd
port 124 nsew
rlabel metal3 s 58964 57604 58964 57604 4 gnd
port 125 nsew
rlabel metal3 s 59346 57232 59346 57232 4 vdd
port 124 nsew
rlabel metal3 s 58964 55629 58964 55629 4 gnd
port 125 nsew
rlabel metal3 s 59778 56442 59778 56442 4 vdd
port 124 nsew
rlabel metal3 s 59778 55220 59778 55220 4 vdd
port 124 nsew
rlabel metal3 s 59346 56442 59346 56442 4 vdd
port 124 nsew
rlabel metal3 s 58964 56024 58964 56024 4 gnd
port 125 nsew
rlabel metal3 s 58964 56419 58964 56419 4 gnd
port 125 nsew
rlabel metal3 s 59778 57232 59778 57232 4 vdd
port 124 nsew
rlabel metal3 s 58692 56814 58692 56814 4 vdd
port 124 nsew
rlabel metal3 s 58692 55629 58692 55629 4 vdd
port 124 nsew
rlabel metal3 s 60203 56068 60203 56068 4 gnd
port 125 nsew
rlabel metal3 s 58692 57209 58692 57209 4 vdd
port 124 nsew
rlabel metal3 s 59346 58022 59346 58022 4 vdd
port 124 nsew
rlabel metal3 s 58964 56814 58964 56814 4 gnd
port 125 nsew
rlabel metal3 s 58692 54839 58692 54839 4 vdd
port 124 nsew
rlabel metal3 s 58692 58394 58692 58394 4 vdd
port 124 nsew
rlabel metal3 s 60203 55278 60203 55278 4 gnd
port 125 nsew
rlabel metal3 s 59346 58380 59346 58380 4 vdd
port 124 nsew
rlabel metal3 s 59778 55652 59778 55652 4 vdd
port 124 nsew
rlabel metal3 s 58692 56419 58692 56419 4 vdd
port 124 nsew
rlabel metal3 s 60203 58022 60203 58022 4 gnd
port 125 nsew
rlabel metal3 s 60203 54862 60203 54862 4 gnd
port 125 nsew
rlabel metal3 s 58964 57999 58964 57999 4 gnd
port 125 nsew
rlabel metal3 s 59346 54862 59346 54862 4 vdd
port 124 nsew
rlabel metal3 s 59346 56800 59346 56800 4 vdd
port 124 nsew
rlabel metal3 s 59778 57590 59778 57590 4 vdd
port 124 nsew
rlabel metal3 s 58964 54839 58964 54839 4 gnd
port 125 nsew
rlabel metal3 s 59346 56010 59346 56010 4 vdd
port 124 nsew
rlabel metal3 s 59778 56010 59778 56010 4 vdd
port 124 nsew
rlabel metal3 s 59778 54862 59778 54862 4 vdd
port 124 nsew
rlabel metal3 s 59346 55220 59346 55220 4 vdd
port 124 nsew
rlabel metal3 s 60203 57232 60203 57232 4 gnd
port 125 nsew
rlabel metal3 s 58964 58394 58964 58394 4 gnd
port 125 nsew
rlabel metal3 s 58692 57999 58692 57999 4 vdd
port 124 nsew
rlabel metal3 s 58692 55234 58692 55234 4 vdd
port 124 nsew
rlabel metal3 s 59778 58380 59778 58380 4 vdd
port 124 nsew
rlabel metal3 s 60203 55652 60203 55652 4 gnd
port 125 nsew
rlabel metal3 s 60203 56858 60203 56858 4 gnd
port 125 nsew
rlabel metal3 s 60203 53282 60203 53282 4 gnd
port 125 nsew
rlabel metal3 s 60203 50538 60203 50538 4 gnd
port 125 nsew
rlabel metal3 s 58692 51284 58692 51284 4 vdd
port 124 nsew
rlabel metal3 s 59778 52850 59778 52850 4 vdd
port 124 nsew
rlabel metal3 s 59778 54430 59778 54430 4 vdd
port 124 nsew
rlabel metal3 s 59346 53282 59346 53282 4 vdd
port 124 nsew
rlabel metal3 s 58692 51679 58692 51679 4 vdd
port 124 nsew
rlabel metal3 s 58692 53654 58692 53654 4 vdd
port 124 nsew
rlabel metal3 s 59346 52060 59346 52060 4 vdd
port 124 nsew
rlabel metal3 s 59778 51702 59778 51702 4 vdd
port 124 nsew
rlabel metal3 s 59778 50912 59778 50912 4 vdd
port 124 nsew
rlabel metal3 s 58964 52469 58964 52469 4 gnd
port 125 nsew
rlabel metal3 s 58964 53259 58964 53259 4 gnd
port 125 nsew
rlabel metal3 s 60203 51328 60203 51328 4 gnd
port 125 nsew
rlabel metal3 s 60203 53698 60203 53698 4 gnd
port 125 nsew
rlabel metal3 s 60203 54072 60203 54072 4 gnd
port 125 nsew
rlabel metal3 s 58692 53259 58692 53259 4 vdd
port 124 nsew
rlabel metal3 s 59346 50480 59346 50480 4 vdd
port 124 nsew
rlabel metal3 s 58964 50494 58964 50494 4 gnd
port 125 nsew
rlabel metal3 s 58964 50889 58964 50889 4 gnd
port 125 nsew
rlabel metal3 s 59778 51270 59778 51270 4 vdd
port 124 nsew
rlabel metal3 s 59778 54072 59778 54072 4 vdd
port 124 nsew
rlabel metal3 s 59778 53282 59778 53282 4 vdd
port 124 nsew
rlabel metal3 s 58692 50494 58692 50494 4 vdd
port 124 nsew
rlabel metal3 s 60203 54488 60203 54488 4 gnd
port 125 nsew
rlabel metal3 s 59778 53640 59778 53640 4 vdd
port 124 nsew
rlabel metal3 s 59778 50480 59778 50480 4 vdd
port 124 nsew
rlabel metal3 s 59346 52492 59346 52492 4 vdd
port 124 nsew
rlabel metal3 s 59346 54430 59346 54430 4 vdd
port 124 nsew
rlabel metal3 s 59346 54072 59346 54072 4 vdd
port 124 nsew
rlabel metal3 s 60203 52492 60203 52492 4 gnd
port 125 nsew
rlabel metal3 s 59346 50912 59346 50912 4 vdd
port 124 nsew
rlabel metal3 s 58964 53654 58964 53654 4 gnd
port 125 nsew
rlabel metal3 s 58964 52864 58964 52864 4 gnd
port 125 nsew
rlabel metal3 s 58964 54049 58964 54049 4 gnd
port 125 nsew
rlabel metal3 s 59778 52492 59778 52492 4 vdd
port 124 nsew
rlabel metal3 s 60203 52908 60203 52908 4 gnd
port 125 nsew
rlabel metal3 s 58692 54444 58692 54444 4 vdd
port 124 nsew
rlabel metal3 s 58964 54444 58964 54444 4 gnd
port 125 nsew
rlabel metal3 s 59346 53640 59346 53640 4 vdd
port 124 nsew
rlabel metal3 s 60203 50912 60203 50912 4 gnd
port 125 nsew
rlabel metal3 s 59346 51270 59346 51270 4 vdd
port 124 nsew
rlabel metal3 s 59778 52060 59778 52060 4 vdd
port 124 nsew
rlabel metal3 s 59346 51702 59346 51702 4 vdd
port 124 nsew
rlabel metal3 s 58692 52074 58692 52074 4 vdd
port 124 nsew
rlabel metal3 s 58692 52469 58692 52469 4 vdd
port 124 nsew
rlabel metal3 s 58964 51679 58964 51679 4 gnd
port 125 nsew
rlabel metal3 s 59346 52850 59346 52850 4 vdd
port 124 nsew
rlabel metal3 s 58964 52074 58964 52074 4 gnd
port 125 nsew
rlabel metal3 s 60203 52118 60203 52118 4 gnd
port 125 nsew
rlabel metal3 s 60203 51702 60203 51702 4 gnd
port 125 nsew
rlabel metal3 s 58692 52864 58692 52864 4 vdd
port 124 nsew
rlabel metal3 s 58964 51284 58964 51284 4 gnd
port 125 nsew
rlabel metal3 s 58692 50889 58692 50889 4 vdd
port 124 nsew
rlabel metal3 s 58692 54049 58692 54049 4 vdd
port 124 nsew
rlabel metal3 s 45687 61887 45687 61887 4 vdd
port 124 nsew
rlabel metal3 s 48614 63460 48614 63460 4 gnd
port 125 nsew
rlabel metal3 s 44627 67167 44627 67167 4 gnd
port 125 nsew
rlabel metal3 s 42805 61887 42805 61887 4 vdd
port 124 nsew
rlabel metal3 s 42062 61296 42062 61296 4 vdd
port 124 nsew
rlabel metal3 s 44627 66845 44627 66845 4 vdd
port 124 nsew
rlabel metal3 s 42131 66845 42131 66845 4 vdd
port 124 nsew
rlabel metal3 s 44697 65233 44697 65233 4 gnd
port 125 nsew
rlabel metal3 s 45301 61887 45301 61887 4 vdd
port 124 nsew
rlabel metal3 s 48371 66845 48371 66845 4 vdd
port 124 nsew
rlabel metal3 s 44615 66007 44615 66007 4 vdd
port 124 nsew
rlabel metal3 s 42686 61296 42686 61296 4 vdd
port 124 nsew
rlabel metal3 s 45182 61296 45182 61296 4 vdd
port 124 nsew
rlabel metal3 s 46118 63460 46118 63460 4 gnd
port 125 nsew
rlabel metal3 s 43622 63460 43622 63460 4 gnd
port 125 nsew
rlabel metal3 s 48371 67167 48371 67167 4 gnd
port 125 nsew
rlabel metal3 s 45806 61296 45806 61296 4 vdd
port 124 nsew
rlabel metal3 s 45945 65233 45945 65233 4 gnd
port 125 nsew
rlabel metal3 s 44558 61296 44558 61296 4 vdd
port 124 nsew
rlabel metal3 s 46549 61887 46549 61887 4 vdd
port 124 nsew
rlabel metal3 s 43191 61887 43191 61887 4 vdd
port 124 nsew
rlabel metal3 s 48359 66007 48359 66007 4 vdd
port 124 nsew
rlabel metal3 s 44439 61887 44439 61887 4 vdd
port 124 nsew
rlabel metal3 s 41126 63460 41126 63460 4 gnd
port 125 nsew
rlabel metal3 s 43449 65233 43449 65233 4 gnd
port 125 nsew
rlabel metal3 s 43367 66007 43367 66007 4 vdd
port 124 nsew
rlabel metal3 s 48302 61296 48302 61296 4 vdd
port 124 nsew
rlabel metal3 s 41943 61887 41943 61887 4 vdd
port 124 nsew
rlabel metal3 s 42201 65233 42201 65233 4 gnd
port 125 nsew
rlabel metal3 s 47797 61887 47797 61887 4 vdd
port 124 nsew
rlabel metal3 s 47193 65233 47193 65233 4 gnd
port 125 nsew
rlabel metal3 s 46430 61296 46430 61296 4 vdd
port 124 nsew
rlabel metal3 s 42119 66007 42119 66007 4 vdd
port 124 nsew
rlabel metal3 s 44053 61887 44053 61887 4 vdd
port 124 nsew
rlabel metal3 s 45875 67167 45875 67167 4 gnd
port 125 nsew
rlabel metal3 s 43310 61296 43310 61296 4 vdd
port 124 nsew
rlabel metal3 s 45875 66845 45875 66845 4 vdd
port 124 nsew
rlabel metal3 s 47111 66007 47111 66007 4 vdd
port 124 nsew
rlabel metal3 s 44870 63460 44870 63460 4 gnd
port 125 nsew
rlabel metal3 s 41557 61887 41557 61887 4 vdd
port 124 nsew
rlabel metal3 s 47366 63460 47366 63460 4 gnd
port 125 nsew
rlabel metal3 s 41438 61296 41438 61296 4 vdd
port 124 nsew
rlabel metal3 s 47123 67167 47123 67167 4 gnd
port 125 nsew
rlabel metal3 s 48441 65233 48441 65233 4 gnd
port 125 nsew
rlabel metal3 s 47054 61296 47054 61296 4 vdd
port 124 nsew
rlabel metal3 s 42131 67167 42131 67167 4 gnd
port 125 nsew
rlabel metal3 s 43379 67167 43379 67167 4 gnd
port 125 nsew
rlabel metal3 s 47123 66845 47123 66845 4 vdd
port 124 nsew
rlabel metal3 s 43379 66845 43379 66845 4 vdd
port 124 nsew
rlabel metal3 s 42374 63460 42374 63460 4 gnd
port 125 nsew
rlabel metal3 s 46935 61887 46935 61887 4 vdd
port 124 nsew
rlabel metal3 s 43934 61296 43934 61296 4 vdd
port 124 nsew
rlabel metal3 s 48183 61887 48183 61887 4 vdd
port 124 nsew
rlabel metal3 s 45863 66007 45863 66007 4 vdd
port 124 nsew
rlabel metal3 s 47678 61296 47678 61296 4 vdd
port 124 nsew
rlabel metal3 s 40871 66007 40871 66007 4 vdd
port 124 nsew
rlabel metal3 s 33395 66845 33395 66845 4 vdd
port 124 nsew
rlabel metal3 s 37139 67167 37139 67167 4 gnd
port 125 nsew
rlabel metal3 s 34643 67167 34643 67167 4 gnd
port 125 nsew
rlabel metal3 s 37070 61296 37070 61296 4 vdd
port 124 nsew
rlabel metal3 s 35961 65233 35961 65233 4 gnd
port 125 nsew
rlabel metal3 s 38942 61296 38942 61296 4 vdd
port 124 nsew
rlabel metal3 s 33326 61296 33326 61296 4 vdd
port 124 nsew
rlabel metal3 s 35879 66007 35879 66007 4 vdd
port 124 nsew
rlabel metal3 s 39447 61887 39447 61887 4 vdd
port 124 nsew
rlabel metal3 s 34574 61296 34574 61296 4 vdd
port 124 nsew
rlabel metal3 s 34631 66007 34631 66007 4 vdd
port 124 nsew
rlabel metal3 s 40190 61296 40190 61296 4 vdd
port 124 nsew
rlabel metal3 s 36446 61296 36446 61296 4 vdd
port 124 nsew
rlabel metal3 s 39623 66007 39623 66007 4 vdd
port 124 nsew
rlabel metal3 s 34455 61887 34455 61887 4 vdd
port 124 nsew
rlabel metal3 s 33465 65233 33465 65233 4 gnd
port 125 nsew
rlabel metal3 s 38375 66007 38375 66007 4 vdd
port 124 nsew
rlabel metal3 s 36951 61887 36951 61887 4 vdd
port 124 nsew
rlabel metal3 s 37139 66845 37139 66845 4 vdd
port 124 nsew
rlabel metal3 s 35891 67167 35891 67167 4 gnd
port 125 nsew
rlabel metal3 s 39705 65233 39705 65233 4 gnd
port 125 nsew
rlabel metal3 s 34713 65233 34713 65233 4 gnd
port 125 nsew
rlabel metal3 s 38318 61296 38318 61296 4 vdd
port 124 nsew
rlabel metal3 s 40883 66845 40883 66845 4 vdd
port 124 nsew
rlabel metal3 s 35822 61296 35822 61296 4 vdd
port 124 nsew
rlabel metal3 s 33395 67167 33395 67167 4 gnd
port 125 nsew
rlabel metal3 s 36565 61887 36565 61887 4 vdd
port 124 nsew
rlabel metal3 s 35891 66845 35891 66845 4 vdd
port 124 nsew
rlabel metal3 s 34886 63460 34886 63460 4 gnd
port 125 nsew
rlabel metal3 s 37382 63460 37382 63460 4 gnd
port 125 nsew
rlabel metal3 s 40309 61887 40309 61887 4 vdd
port 124 nsew
rlabel metal3 s 37127 66007 37127 66007 4 vdd
port 124 nsew
rlabel metal3 s 33383 66007 33383 66007 4 vdd
port 124 nsew
rlabel metal3 s 37694 61296 37694 61296 4 vdd
port 124 nsew
rlabel metal3 s 40953 65233 40953 65233 4 gnd
port 125 nsew
rlabel metal3 s 38387 66845 38387 66845 4 vdd
port 124 nsew
rlabel metal3 s 35198 61296 35198 61296 4 vdd
port 124 nsew
rlabel metal3 s 33950 61296 33950 61296 4 vdd
port 124 nsew
rlabel metal3 s 40883 67167 40883 67167 4 gnd
port 125 nsew
rlabel metal3 s 36134 63460 36134 63460 4 gnd
port 125 nsew
rlabel metal3 s 39566 61296 39566 61296 4 vdd
port 124 nsew
rlabel metal3 s 39635 66845 39635 66845 4 vdd
port 124 nsew
rlabel metal3 s 38387 67167 38387 67167 4 gnd
port 125 nsew
rlabel metal3 s 40814 61296 40814 61296 4 vdd
port 124 nsew
rlabel metal3 s 37209 65233 37209 65233 4 gnd
port 125 nsew
rlabel metal3 s 35317 61887 35317 61887 4 vdd
port 124 nsew
rlabel metal3 s 34643 66845 34643 66845 4 vdd
port 124 nsew
rlabel metal3 s 38630 63460 38630 63460 4 gnd
port 125 nsew
rlabel metal3 s 40695 61887 40695 61887 4 vdd
port 124 nsew
rlabel metal3 s 35703 61887 35703 61887 4 vdd
port 124 nsew
rlabel metal3 s 39061 61887 39061 61887 4 vdd
port 124 nsew
rlabel metal3 s 33638 63460 33638 63460 4 gnd
port 125 nsew
rlabel metal3 s 39878 63460 39878 63460 4 gnd
port 125 nsew
rlabel metal3 s 39635 67167 39635 67167 4 gnd
port 125 nsew
rlabel metal3 s 34069 61887 34069 61887 4 vdd
port 124 nsew
rlabel metal3 s 37813 61887 37813 61887 4 vdd
port 124 nsew
rlabel metal3 s 38199 61887 38199 61887 4 vdd
port 124 nsew
rlabel metal3 s 33207 61887 33207 61887 4 vdd
port 124 nsew
rlabel metal3 s 38457 65233 38457 65233 4 gnd
port 125 nsew
rlabel metal3 s 59778 49690 59778 49690 4 vdd
port 124 nsew
rlabel metal3 s 59346 50122 59346 50122 4 vdd
port 124 nsew
rlabel metal3 s 59346 46530 59346 46530 4 vdd
port 124 nsew
rlabel metal3 s 58964 47729 58964 47729 4 gnd
port 125 nsew
rlabel metal3 s 58964 47334 58964 47334 4 gnd
port 125 nsew
rlabel metal3 s 58692 48124 58692 48124 4 vdd
port 124 nsew
rlabel metal3 s 59778 48542 59778 48542 4 vdd
port 124 nsew
rlabel metal3 s 59346 49332 59346 49332 4 vdd
port 124 nsew
rlabel metal3 s 60203 50122 60203 50122 4 gnd
port 125 nsew
rlabel metal3 s 58964 46939 58964 46939 4 gnd
port 125 nsew
rlabel metal3 s 60203 46588 60203 46588 4 gnd
port 125 nsew
rlabel metal3 s 58964 49309 58964 49309 4 gnd
port 125 nsew
rlabel metal3 s 58964 49704 58964 49704 4 gnd
port 125 nsew
rlabel metal3 s 59346 49690 59346 49690 4 vdd
port 124 nsew
rlabel metal3 s 60203 48168 60203 48168 4 gnd
port 125 nsew
rlabel metal3 s 58964 46544 58964 46544 4 gnd
port 125 nsew
rlabel metal3 s 60203 49332 60203 49332 4 gnd
port 125 nsew
rlabel metal3 s 58964 48124 58964 48124 4 gnd
port 125 nsew
rlabel metal3 s 59778 46962 59778 46962 4 vdd
port 124 nsew
rlabel metal3 s 58692 50099 58692 50099 4 vdd
port 124 nsew
rlabel metal3 s 58692 46544 58692 46544 4 vdd
port 124 nsew
rlabel metal3 s 59778 47752 59778 47752 4 vdd
port 124 nsew
rlabel metal3 s 60203 48958 60203 48958 4 gnd
port 125 nsew
rlabel metal3 s 58964 48914 58964 48914 4 gnd
port 125 nsew
rlabel metal3 s 58692 49704 58692 49704 4 vdd
port 124 nsew
rlabel metal3 s 59346 48900 59346 48900 4 vdd
port 124 nsew
rlabel metal3 s 59778 46530 59778 46530 4 vdd
port 124 nsew
rlabel metal3 s 60203 47378 60203 47378 4 gnd
port 125 nsew
rlabel metal3 s 58692 47334 58692 47334 4 vdd
port 124 nsew
rlabel metal3 s 58692 48519 58692 48519 4 vdd
port 124 nsew
rlabel metal3 s 58692 49309 58692 49309 4 vdd
port 124 nsew
rlabel metal3 s 59778 47320 59778 47320 4 vdd
port 124 nsew
rlabel metal3 s 59346 48542 59346 48542 4 vdd
port 124 nsew
rlabel metal3 s 58692 47729 58692 47729 4 vdd
port 124 nsew
rlabel metal3 s 60203 47752 60203 47752 4 gnd
port 125 nsew
rlabel metal3 s 58692 46939 58692 46939 4 vdd
port 124 nsew
rlabel metal3 s 59778 50122 59778 50122 4 vdd
port 124 nsew
rlabel metal3 s 60203 48542 60203 48542 4 gnd
port 125 nsew
rlabel metal3 s 59346 47320 59346 47320 4 vdd
port 124 nsew
rlabel metal3 s 59778 49332 59778 49332 4 vdd
port 124 nsew
rlabel metal3 s 60203 46962 60203 46962 4 gnd
port 125 nsew
rlabel metal3 s 59346 48110 59346 48110 4 vdd
port 124 nsew
rlabel metal3 s 58692 48914 58692 48914 4 vdd
port 124 nsew
rlabel metal3 s 60203 49748 60203 49748 4 gnd
port 125 nsew
rlabel metal3 s 59778 48900 59778 48900 4 vdd
port 124 nsew
rlabel metal3 s 59346 46962 59346 46962 4 vdd
port 124 nsew
rlabel metal3 s 59778 48110 59778 48110 4 vdd
port 124 nsew
rlabel metal3 s 58964 48519 58964 48519 4 gnd
port 125 nsew
rlabel metal3 s 59346 47752 59346 47752 4 vdd
port 124 nsew
rlabel metal3 s 58964 50099 58964 50099 4 gnd
port 125 nsew
rlabel metal3 s 59346 45382 59346 45382 4 vdd
port 124 nsew
rlabel metal3 s 58692 42989 58692 42989 4 vdd
port 124 nsew
rlabel metal3 s 58692 44569 58692 44569 4 vdd
port 124 nsew
rlabel metal3 s 59778 45740 59778 45740 4 vdd
port 124 nsew
rlabel metal3 s 60203 42222 60203 42222 4 gnd
port 125 nsew
rlabel metal3 s 59778 43012 59778 43012 4 vdd
port 124 nsew
rlabel metal3 s 59346 44160 59346 44160 4 vdd
port 124 nsew
rlabel metal3 s 58692 46149 58692 46149 4 vdd
port 124 nsew
rlabel metal3 s 59346 45740 59346 45740 4 vdd
port 124 nsew
rlabel metal3 s 58964 44174 58964 44174 4 gnd
port 125 nsew
rlabel metal3 s 60203 45382 60203 45382 4 gnd
port 125 nsew
rlabel metal3 s 59346 44950 59346 44950 4 vdd
port 124 nsew
rlabel metal3 s 60203 43428 60203 43428 4 gnd
port 125 nsew
rlabel metal3 s 58964 44964 58964 44964 4 gnd
port 125 nsew
rlabel metal3 s 58692 42594 58692 42594 4 vdd
port 124 nsew
rlabel metal3 s 60203 43802 60203 43802 4 gnd
port 125 nsew
rlabel metal3 s 59346 42580 59346 42580 4 vdd
port 124 nsew
rlabel metal3 s 59778 44950 59778 44950 4 vdd
port 124 nsew
rlabel metal3 s 60203 43012 60203 43012 4 gnd
port 125 nsew
rlabel metal3 s 59778 45382 59778 45382 4 vdd
port 124 nsew
rlabel metal3 s 60203 45008 60203 45008 4 gnd
port 125 nsew
rlabel metal3 s 58964 43779 58964 43779 4 gnd
port 125 nsew
rlabel metal3 s 58964 45754 58964 45754 4 gnd
port 125 nsew
rlabel metal3 s 58692 44964 58692 44964 4 vdd
port 124 nsew
rlabel metal3 s 59346 44592 59346 44592 4 vdd
port 124 nsew
rlabel metal3 s 59778 43370 59778 43370 4 vdd
port 124 nsew
rlabel metal3 s 58964 43384 58964 43384 4 gnd
port 125 nsew
rlabel metal3 s 58692 44174 58692 44174 4 vdd
port 124 nsew
rlabel metal3 s 58692 42199 58692 42199 4 vdd
port 124 nsew
rlabel metal3 s 59778 42580 59778 42580 4 vdd
port 124 nsew
rlabel metal3 s 60203 45798 60203 45798 4 gnd
port 125 nsew
rlabel metal3 s 59346 43802 59346 43802 4 vdd
port 124 nsew
rlabel metal3 s 59346 46172 59346 46172 4 vdd
port 124 nsew
rlabel metal3 s 59346 42222 59346 42222 4 vdd
port 124 nsew
rlabel metal3 s 58964 44569 58964 44569 4 gnd
port 125 nsew
rlabel metal3 s 58964 45359 58964 45359 4 gnd
port 125 nsew
rlabel metal3 s 59346 43012 59346 43012 4 vdd
port 124 nsew
rlabel metal3 s 58964 42989 58964 42989 4 gnd
port 125 nsew
rlabel metal3 s 59778 46172 59778 46172 4 vdd
port 124 nsew
rlabel metal3 s 59778 44160 59778 44160 4 vdd
port 124 nsew
rlabel metal3 s 58692 43384 58692 43384 4 vdd
port 124 nsew
rlabel metal3 s 59346 43370 59346 43370 4 vdd
port 124 nsew
rlabel metal3 s 58692 45754 58692 45754 4 vdd
port 124 nsew
rlabel metal3 s 59778 43802 59778 43802 4 vdd
port 124 nsew
rlabel metal3 s 59778 44592 59778 44592 4 vdd
port 124 nsew
rlabel metal3 s 58964 46149 58964 46149 4 gnd
port 125 nsew
rlabel metal3 s 58964 42594 58964 42594 4 gnd
port 125 nsew
rlabel metal3 s 58964 42199 58964 42199 4 gnd
port 125 nsew
rlabel metal3 s 60203 46172 60203 46172 4 gnd
port 125 nsew
rlabel metal3 s 60203 44218 60203 44218 4 gnd
port 125 nsew
rlabel metal3 s 59778 42222 59778 42222 4 vdd
port 124 nsew
rlabel metal3 s 58692 43779 58692 43779 4 vdd
port 124 nsew
rlabel metal3 s 58692 45359 58692 45359 4 vdd
port 124 nsew
rlabel metal3 s 60203 42638 60203 42638 4 gnd
port 125 nsew
rlabel metal3 s 60203 44592 60203 44592 4 gnd
port 125 nsew
rlabel metal3 s 53990 44145 53990 44145 4 gnd
port 125 nsew
rlabel metal3 s 53990 48648 53990 48648 4 gnd
port 125 nsew
rlabel metal3 s 53990 45488 53990 45488 4 gnd
port 125 nsew
rlabel metal3 s 53990 44935 53990 44935 4 gnd
port 125 nsew
rlabel metal3 s 53990 49675 53990 49675 4 gnd
port 125 nsew
rlabel metal3 s 53990 49912 53990 49912 4 gnd
port 125 nsew
rlabel metal3 s 53990 46278 53990 46278 4 gnd
port 125 nsew
rlabel metal3 s 53990 43118 53990 43118 4 gnd
port 125 nsew
rlabel metal3 s 53990 50228 53990 50228 4 gnd
port 125 nsew
rlabel metal3 s 53990 44698 53990 44698 4 gnd
port 125 nsew
rlabel metal3 s 53990 46515 53990 46515 4 gnd
port 125 nsew
rlabel metal3 s 53990 43355 53990 43355 4 gnd
port 125 nsew
rlabel metal3 s 53990 42328 53990 42328 4 gnd
port 125 nsew
rlabel metal3 s 53990 48332 53990 48332 4 gnd
port 125 nsew
rlabel metal3 s 53990 45172 53990 45172 4 gnd
port 125 nsew
rlabel metal3 s 53990 49122 53990 49122 4 gnd
port 125 nsew
rlabel metal3 s 53990 45725 53990 45725 4 gnd
port 125 nsew
rlabel metal3 s 53990 42012 53990 42012 4 gnd
port 125 nsew
rlabel metal3 s 53990 42802 53990 42802 4 gnd
port 125 nsew
rlabel metal3 s 53990 46752 53990 46752 4 gnd
port 125 nsew
rlabel metal3 s 53990 42565 53990 42565 4 gnd
port 125 nsew
rlabel metal3 s 53990 43592 53990 43592 4 gnd
port 125 nsew
rlabel metal3 s 53990 47858 53990 47858 4 gnd
port 125 nsew
rlabel metal3 s 53990 48095 53990 48095 4 gnd
port 125 nsew
rlabel metal3 s 53990 48885 53990 48885 4 gnd
port 125 nsew
rlabel metal3 s 53990 44382 53990 44382 4 gnd
port 125 nsew
rlabel metal3 s 53990 47305 53990 47305 4 gnd
port 125 nsew
rlabel metal3 s 53990 49438 53990 49438 4 gnd
port 125 nsew
rlabel metal3 s 53990 45962 53990 45962 4 gnd
port 125 nsew
rlabel metal3 s 53990 47068 53990 47068 4 gnd
port 125 nsew
rlabel metal3 s 53990 43908 53990 43908 4 gnd
port 125 nsew
rlabel metal3 s 53990 47542 53990 47542 4 gnd
port 125 nsew
rlabel metal3 s 53990 41222 53990 41222 4 gnd
port 125 nsew
rlabel metal3 s 53990 34665 53990 34665 4 gnd
port 125 nsew
rlabel metal3 s 53990 35218 53990 35218 4 gnd
port 125 nsew
rlabel metal3 s 53990 36008 53990 36008 4 gnd
port 125 nsew
rlabel metal3 s 53990 39168 53990 39168 4 gnd
port 125 nsew
rlabel metal3 s 53990 34112 53990 34112 4 gnd
port 125 nsew
rlabel metal3 s 53990 38062 53990 38062 4 gnd
port 125 nsew
rlabel metal3 s 53990 38852 53990 38852 4 gnd
port 125 nsew
rlabel metal3 s 53990 37035 53990 37035 4 gnd
port 125 nsew
rlabel metal3 s 53990 40432 53990 40432 4 gnd
port 125 nsew
rlabel metal3 s 53990 34902 53990 34902 4 gnd
port 125 nsew
rlabel metal3 s 53990 39642 53990 39642 4 gnd
port 125 nsew
rlabel metal3 s 55254 35455 55254 35455 4 vdd
port 124 nsew
rlabel metal3 s 53990 35455 53990 35455 4 gnd
port 125 nsew
rlabel metal3 s 53990 33875 53990 33875 4 gnd
port 125 nsew
rlabel metal3 s 53990 39958 53990 39958 4 gnd
port 125 nsew
rlabel metal3 s 53990 39405 53990 39405 4 gnd
port 125 nsew
rlabel metal3 s 53990 34428 53990 34428 4 gnd
port 125 nsew
rlabel metal3 s 53990 37588 53990 37588 4 gnd
port 125 nsew
rlabel metal3 s 56778 35455 56778 35455 4 gnd
port 125 nsew
rlabel metal3 s 53990 40195 53990 40195 4 gnd
port 125 nsew
rlabel metal3 s 53990 38378 53990 38378 4 gnd
port 125 nsew
rlabel metal3 s 53990 36482 53990 36482 4 gnd
port 125 nsew
rlabel metal3 s 53990 38615 53990 38615 4 gnd
port 125 nsew
rlabel metal3 s 53990 40985 53990 40985 4 gnd
port 125 nsew
rlabel metal3 s 53990 35692 53990 35692 4 gnd
port 125 nsew
rlabel metal3 s 53990 40748 53990 40748 4 gnd
port 125 nsew
rlabel metal3 s 53990 41538 53990 41538 4 gnd
port 125 nsew
rlabel metal3 s 53990 36245 53990 36245 4 gnd
port 125 nsew
rlabel metal3 s 53990 33638 53990 33638 4 gnd
port 125 nsew
rlabel metal3 s 53990 37825 53990 37825 4 gnd
port 125 nsew
rlabel metal3 s 53990 41775 53990 41775 4 gnd
port 125 nsew
rlabel metal3 s 53990 36798 53990 36798 4 gnd
port 125 nsew
rlabel metal3 s 53990 37272 53990 37272 4 gnd
port 125 nsew
rlabel metal3 s 58964 40224 58964 40224 4 gnd
port 125 nsew
rlabel metal3 s 58692 39434 58692 39434 4 vdd
port 124 nsew
rlabel metal3 s 58692 37854 58692 37854 4 vdd
port 124 nsew
rlabel metal3 s 58964 40619 58964 40619 4 gnd
port 125 nsew
rlabel metal3 s 59778 41000 59778 41000 4 vdd
port 124 nsew
rlabel metal3 s 60203 39852 60203 39852 4 gnd
port 125 nsew
rlabel metal3 s 59346 39062 59346 39062 4 vdd
port 124 nsew
rlabel metal3 s 60203 40268 60203 40268 4 gnd
port 125 nsew
rlabel metal3 s 60203 37898 60203 37898 4 gnd
port 125 nsew
rlabel metal3 s 58964 41014 58964 41014 4 gnd
port 125 nsew
rlabel metal3 s 60203 39062 60203 39062 4 gnd
port 125 nsew
rlabel metal3 s 58692 38249 58692 38249 4 vdd
port 124 nsew
rlabel metal3 s 60203 38272 60203 38272 4 gnd
port 125 nsew
rlabel metal3 s 58964 39434 58964 39434 4 gnd
port 125 nsew
rlabel metal3 s 60203 38688 60203 38688 4 gnd
port 125 nsew
rlabel metal3 s 59346 41790 59346 41790 4 vdd
port 124 nsew
rlabel metal3 s 60203 40642 60203 40642 4 gnd
port 125 nsew
rlabel metal3 s 59778 39420 59778 39420 4 vdd
port 124 nsew
rlabel metal3 s 58964 39039 58964 39039 4 gnd
port 125 nsew
rlabel metal3 s 59346 37840 59346 37840 4 vdd
port 124 nsew
rlabel metal3 s 59346 41000 59346 41000 4 vdd
port 124 nsew
rlabel metal3 s 58692 41409 58692 41409 4 vdd
port 124 nsew
rlabel metal3 s 59778 38630 59778 38630 4 vdd
port 124 nsew
rlabel metal3 s 59778 40642 59778 40642 4 vdd
port 124 nsew
rlabel metal3 s 59346 38272 59346 38272 4 vdd
port 124 nsew
rlabel metal3 s 58692 38644 58692 38644 4 vdd
port 124 nsew
rlabel metal3 s 59346 40210 59346 40210 4 vdd
port 124 nsew
rlabel metal3 s 58692 39039 58692 39039 4 vdd
port 124 nsew
rlabel metal3 s 59778 40210 59778 40210 4 vdd
port 124 nsew
rlabel metal3 s 60203 41848 60203 41848 4 gnd
port 125 nsew
rlabel metal3 s 59346 39420 59346 39420 4 vdd
port 124 nsew
rlabel metal3 s 58964 41409 58964 41409 4 gnd
port 125 nsew
rlabel metal3 s 58964 38644 58964 38644 4 gnd
port 125 nsew
rlabel metal3 s 58692 39829 58692 39829 4 vdd
port 124 nsew
rlabel metal3 s 59778 38272 59778 38272 4 vdd
port 124 nsew
rlabel metal3 s 58692 40619 58692 40619 4 vdd
port 124 nsew
rlabel metal3 s 58964 38249 58964 38249 4 gnd
port 125 nsew
rlabel metal3 s 58692 41014 58692 41014 4 vdd
port 124 nsew
rlabel metal3 s 59778 39852 59778 39852 4 vdd
port 124 nsew
rlabel metal3 s 60203 41432 60203 41432 4 gnd
port 125 nsew
rlabel metal3 s 59778 41790 59778 41790 4 vdd
port 124 nsew
rlabel metal3 s 58692 40224 58692 40224 4 vdd
port 124 nsew
rlabel metal3 s 59346 40642 59346 40642 4 vdd
port 124 nsew
rlabel metal3 s 59346 39852 59346 39852 4 vdd
port 124 nsew
rlabel metal3 s 59778 37840 59778 37840 4 vdd
port 124 nsew
rlabel metal3 s 59778 41432 59778 41432 4 vdd
port 124 nsew
rlabel metal3 s 58964 37854 58964 37854 4 gnd
port 125 nsew
rlabel metal3 s 58964 41804 58964 41804 4 gnd
port 125 nsew
rlabel metal3 s 59346 41432 59346 41432 4 vdd
port 124 nsew
rlabel metal3 s 58964 39829 58964 39829 4 gnd
port 125 nsew
rlabel metal3 s 59346 38630 59346 38630 4 vdd
port 124 nsew
rlabel metal3 s 58692 41804 58692 41804 4 vdd
port 124 nsew
rlabel metal3 s 59778 39062 59778 39062 4 vdd
port 124 nsew
rlabel metal3 s 60203 39478 60203 39478 4 gnd
port 125 nsew
rlabel metal3 s 60203 41058 60203 41058 4 gnd
port 125 nsew
rlabel metal3 s 60203 34738 60203 34738 4 gnd
port 125 nsew
rlabel metal3 s 59778 35112 59778 35112 4 vdd
port 124 nsew
rlabel metal3 s 58692 35089 58692 35089 4 vdd
port 124 nsew
rlabel metal3 s 60203 35112 60203 35112 4 gnd
port 125 nsew
rlabel metal3 s 58964 37459 58964 37459 4 gnd
port 125 nsew
rlabel metal3 s 59346 34322 59346 34322 4 vdd
port 124 nsew
rlabel metal3 s 59778 34322 59778 34322 4 vdd
port 124 nsew
rlabel metal3 s 58692 35484 58692 35484 4 vdd
port 124 nsew
rlabel metal3 s 60203 35902 60203 35902 4 gnd
port 125 nsew
rlabel metal3 s 58964 35089 58964 35089 4 gnd
port 125 nsew
rlabel metal3 s 58692 34694 58692 34694 4 vdd
port 124 nsew
rlabel metal3 s 58692 36669 58692 36669 4 vdd
port 124 nsew
rlabel metal3 s 60203 33948 60203 33948 4 gnd
port 125 nsew
rlabel metal3 s 58692 33904 58692 33904 4 vdd
port 124 nsew
rlabel metal3 s 58964 35484 58964 35484 4 gnd
port 125 nsew
rlabel metal3 s 58964 34694 58964 34694 4 gnd
port 125 nsew
rlabel metal3 s 58692 35879 58692 35879 4 vdd
port 124 nsew
rlabel metal3 s 58964 35879 58964 35879 4 gnd
port 125 nsew
rlabel metal3 s 58964 34299 58964 34299 4 gnd
port 125 nsew
rlabel metal3 s 60203 36318 60203 36318 4 gnd
port 125 nsew
rlabel metal3 s 57821 35439 57821 35439 4 vdd
port 124 nsew
rlabel metal3 s 59778 35902 59778 35902 4 vdd
port 124 nsew
rlabel metal3 s 58964 33904 58964 33904 4 gnd
port 125 nsew
rlabel metal3 s 59346 36260 59346 36260 4 vdd
port 124 nsew
rlabel metal3 s 58964 36669 58964 36669 4 gnd
port 125 nsew
rlabel metal3 s 58692 34299 58692 34299 4 vdd
port 124 nsew
rlabel metal3 s 59346 37050 59346 37050 4 vdd
port 124 nsew
rlabel metal3 s 59346 33890 59346 33890 4 vdd
port 124 nsew
rlabel metal3 s 58964 36274 58964 36274 4 gnd
port 125 nsew
rlabel metal3 s 58964 37064 58964 37064 4 gnd
port 125 nsew
rlabel metal3 s 59346 37482 59346 37482 4 vdd
port 124 nsew
rlabel metal3 s 59778 34680 59778 34680 4 vdd
port 124 nsew
rlabel metal3 s 59346 35902 59346 35902 4 vdd
port 124 nsew
rlabel metal3 s 59778 37050 59778 37050 4 vdd
port 124 nsew
rlabel metal3 s 60203 37108 60203 37108 4 gnd
port 125 nsew
rlabel metal3 s 58692 37459 58692 37459 4 vdd
port 124 nsew
rlabel metal3 s 60203 37482 60203 37482 4 gnd
port 125 nsew
rlabel metal3 s 60203 36692 60203 36692 4 gnd
port 125 nsew
rlabel metal3 s 59778 35470 59778 35470 4 vdd
port 124 nsew
rlabel metal3 s 60203 35528 60203 35528 4 gnd
port 125 nsew
rlabel metal3 s 59346 35112 59346 35112 4 vdd
port 124 nsew
rlabel metal3 s 59778 36692 59778 36692 4 vdd
port 124 nsew
rlabel metal3 s 60203 34322 60203 34322 4 gnd
port 125 nsew
rlabel metal3 s 58692 36274 58692 36274 4 vdd
port 124 nsew
rlabel metal3 s 58246 35440 58246 35440 4 gnd
port 125 nsew
rlabel metal3 s 59346 35470 59346 35470 4 vdd
port 124 nsew
rlabel metal3 s 59778 37482 59778 37482 4 vdd
port 124 nsew
rlabel metal3 s 59778 33890 59778 33890 4 vdd
port 124 nsew
rlabel metal3 s 59346 34680 59346 34680 4 vdd
port 124 nsew
rlabel metal3 s 59346 36692 59346 36692 4 vdd
port 124 nsew
rlabel metal3 s 58692 37064 58692 37064 4 vdd
port 124 nsew
rlabel metal3 s 59778 36260 59778 36260 4 vdd
port 124 nsew
rlabel metal3 s 31573 61887 31573 61887 4 vdd
port 124 nsew
rlabel metal3 s 27155 66845 27155 66845 4 vdd
port 124 nsew
rlabel metal3 s 27829 61887 27829 61887 4 vdd
port 124 nsew
rlabel metal3 s 27398 63460 27398 63460 4 gnd
port 125 nsew
rlabel metal3 s 32135 66007 32135 66007 4 vdd
port 124 nsew
rlabel metal3 s 32702 61296 32702 61296 4 vdd
port 124 nsew
rlabel metal3 s 30206 61296 30206 61296 4 vdd
port 124 nsew
rlabel metal3 s 25214 61296 25214 61296 4 vdd
port 124 nsew
rlabel metal3 s 28391 66007 28391 66007 4 vdd
port 124 nsew
rlabel metal3 s 30325 61887 30325 61887 4 vdd
port 124 nsew
rlabel metal3 s 28215 61887 28215 61887 4 vdd
port 124 nsew
rlabel metal3 s 28403 66845 28403 66845 4 vdd
port 124 nsew
rlabel metal3 s 29894 63460 29894 63460 4 gnd
port 125 nsew
rlabel metal3 s 32390 63460 32390 63460 4 gnd
port 125 nsew
rlabel metal3 s 30830 61296 30830 61296 4 vdd
port 124 nsew
rlabel metal3 s 27225 65233 27225 65233 4 gnd
port 125 nsew
rlabel metal3 s 32147 66845 32147 66845 4 vdd
port 124 nsew
rlabel metal3 s 25907 67167 25907 67167 4 gnd
port 125 nsew
rlabel metal3 s 28473 65233 28473 65233 4 gnd
port 125 nsew
rlabel metal3 s 25977 65233 25977 65233 4 gnd
port 125 nsew
rlabel metal3 s 27086 61296 27086 61296 4 vdd
port 124 nsew
rlabel metal3 s 31454 61296 31454 61296 4 vdd
port 124 nsew
rlabel metal3 s 27143 66007 27143 66007 4 vdd
port 124 nsew
rlabel metal3 s 30899 67167 30899 67167 4 gnd
port 125 nsew
rlabel metal3 s 32821 61887 32821 61887 4 vdd
port 124 nsew
rlabel metal3 s 26150 63460 26150 63460 4 gnd
port 125 nsew
rlabel metal3 s 29651 67167 29651 67167 4 gnd
port 125 nsew
rlabel metal3 s 28403 67167 28403 67167 4 gnd
port 125 nsew
rlabel metal3 s 29582 61296 29582 61296 4 vdd
port 124 nsew
rlabel metal3 s 27710 61296 27710 61296 4 vdd
port 124 nsew
rlabel metal3 s 30969 65233 30969 65233 4 gnd
port 125 nsew
rlabel metal3 s 25719 61887 25719 61887 4 vdd
port 124 nsew
rlabel metal3 s 29651 66845 29651 66845 4 vdd
port 124 nsew
rlabel metal3 s 29463 61887 29463 61887 4 vdd
port 124 nsew
rlabel metal3 s 29077 61887 29077 61887 4 vdd
port 124 nsew
rlabel metal3 s 26581 61887 26581 61887 4 vdd
port 124 nsew
rlabel metal3 s 28958 61296 28958 61296 4 vdd
port 124 nsew
rlabel metal3 s 31142 63460 31142 63460 4 gnd
port 125 nsew
rlabel metal3 s 26967 61887 26967 61887 4 vdd
port 124 nsew
rlabel metal3 s 31959 61887 31959 61887 4 vdd
port 124 nsew
rlabel metal3 s 28334 61296 28334 61296 4 vdd
port 124 nsew
rlabel metal3 s 30887 66007 30887 66007 4 vdd
port 124 nsew
rlabel metal3 s 32078 61296 32078 61296 4 vdd
port 124 nsew
rlabel metal3 s 29721 65233 29721 65233 4 gnd
port 125 nsew
rlabel metal3 s 25895 66007 25895 66007 4 vdd
port 124 nsew
rlabel metal3 s 25333 61887 25333 61887 4 vdd
port 124 nsew
rlabel metal3 s 25838 61296 25838 61296 4 vdd
port 124 nsew
rlabel metal3 s 26462 61296 26462 61296 4 vdd
port 124 nsew
rlabel metal3 s 30711 61887 30711 61887 4 vdd
port 124 nsew
rlabel metal3 s 30899 66845 30899 66845 4 vdd
port 124 nsew
rlabel metal3 s 29639 66007 29639 66007 4 vdd
port 124 nsew
rlabel metal3 s 28646 63460 28646 63460 4 gnd
port 125 nsew
rlabel metal3 s 27155 67167 27155 67167 4 gnd
port 125 nsew
rlabel metal3 s 32217 65233 32217 65233 4 gnd
port 125 nsew
rlabel metal3 s 25907 66845 25907 66845 4 vdd
port 124 nsew
rlabel metal3 s 32147 67167 32147 67167 4 gnd
port 125 nsew
rlabel metal3 s 23399 66007 23399 66007 4 vdd
port 124 nsew
rlabel metal3 s 20341 61887 20341 61887 4 vdd
port 124 nsew
rlabel metal3 s 19093 61887 19093 61887 4 vdd
port 124 nsew
rlabel metal3 s 22094 61296 22094 61296 4 vdd
port 124 nsew
rlabel metal3 s 23342 61296 23342 61296 4 vdd
port 124 nsew
rlabel metal3 s 18662 63460 18662 63460 4 gnd
port 125 nsew
rlabel metal3 s 18350 61296 18350 61296 4 vdd
port 124 nsew
rlabel metal3 s 24659 66845 24659 66845 4 vdd
port 124 nsew
rlabel metal3 s 17726 61296 17726 61296 4 vdd
port 124 nsew
rlabel metal3 s 17171 67167 17171 67167 4 gnd
port 125 nsew
rlabel metal3 s 24647 66007 24647 66007 4 vdd
port 124 nsew
rlabel metal3 s 17159 66007 17159 66007 4 vdd
port 124 nsew
rlabel metal3 s 20915 66845 20915 66845 4 vdd
port 124 nsew
rlabel metal3 s 23481 65233 23481 65233 4 gnd
port 125 nsew
rlabel metal3 s 24729 65233 24729 65233 4 gnd
port 125 nsew
rlabel metal3 s 17845 61887 17845 61887 4 vdd
port 124 nsew
rlabel metal3 s 19910 63460 19910 63460 4 gnd
port 125 nsew
rlabel metal3 s 18407 66007 18407 66007 4 vdd
port 124 nsew
rlabel metal3 s 20903 66007 20903 66007 4 vdd
port 124 nsew
rlabel metal3 s 18231 61887 18231 61887 4 vdd
port 124 nsew
rlabel metal3 s 20846 61296 20846 61296 4 vdd
port 124 nsew
rlabel metal3 s 23411 67167 23411 67167 4 gnd
port 125 nsew
rlabel metal3 s 19667 67167 19667 67167 4 gnd
port 125 nsew
rlabel metal3 s 21975 61887 21975 61887 4 vdd
port 124 nsew
rlabel metal3 s 18489 65233 18489 65233 4 gnd
port 125 nsew
rlabel metal3 s 17414 63460 17414 63460 4 gnd
port 125 nsew
rlabel metal3 s 22233 65233 22233 65233 4 gnd
port 125 nsew
rlabel metal3 s 18974 61296 18974 61296 4 vdd
port 124 nsew
rlabel metal3 s 18419 66845 18419 66845 4 vdd
port 124 nsew
rlabel metal3 s 21158 63460 21158 63460 4 gnd
port 125 nsew
rlabel metal3 s 23411 66845 23411 66845 4 vdd
port 124 nsew
rlabel metal3 s 18419 67167 18419 67167 4 gnd
port 125 nsew
rlabel metal3 s 22151 66007 22151 66007 4 vdd
port 124 nsew
rlabel metal3 s 22163 66845 22163 66845 4 vdd
port 124 nsew
rlabel metal3 s 22406 63460 22406 63460 4 gnd
port 125 nsew
rlabel metal3 s 24659 67167 24659 67167 4 gnd
port 125 nsew
rlabel metal3 s 23654 63460 23654 63460 4 gnd
port 125 nsew
rlabel metal3 s 20915 67167 20915 67167 4 gnd
port 125 nsew
rlabel metal3 s 24590 61296 24590 61296 4 vdd
port 124 nsew
rlabel metal3 s 20985 65233 20985 65233 4 gnd
port 125 nsew
rlabel metal3 s 22837 61887 22837 61887 4 vdd
port 124 nsew
rlabel metal3 s 17171 66845 17171 66845 4 vdd
port 124 nsew
rlabel metal3 s 22163 67167 22163 67167 4 gnd
port 125 nsew
rlabel metal3 s 19737 65233 19737 65233 4 gnd
port 125 nsew
rlabel metal3 s 24902 63460 24902 63460 4 gnd
port 125 nsew
rlabel metal3 s 24085 61887 24085 61887 4 vdd
port 124 nsew
rlabel metal3 s 17241 65233 17241 65233 4 gnd
port 125 nsew
rlabel metal3 s 21589 61887 21589 61887 4 vdd
port 124 nsew
rlabel metal3 s 20727 61887 20727 61887 4 vdd
port 124 nsew
rlabel metal3 s 20222 61296 20222 61296 4 vdd
port 124 nsew
rlabel metal3 s 19598 61296 19598 61296 4 vdd
port 124 nsew
rlabel metal3 s 19655 66007 19655 66007 4 vdd
port 124 nsew
rlabel metal3 s 24471 61887 24471 61887 4 vdd
port 124 nsew
rlabel metal3 s 19479 61887 19479 61887 4 vdd
port 124 nsew
rlabel metal3 s 21470 61296 21470 61296 4 vdd
port 124 nsew
rlabel metal3 s 19667 66845 19667 66845 4 vdd
port 124 nsew
rlabel metal3 s 23966 61296 23966 61296 4 vdd
port 124 nsew
rlabel metal3 s 22718 61296 22718 61296 4 vdd
port 124 nsew
rlabel metal3 s 23223 61887 23223 61887 4 vdd
port 124 nsew
rlabel metal3 s 15349 61887 15349 61887 4 vdd
port 124 nsew
rlabel metal3 s 13427 67167 13427 67167 4 gnd
port 125 nsew
rlabel metal3 s 14663 66007 14663 66007 4 vdd
port 124 nsew
rlabel metal3 s 16597 61887 16597 61887 4 vdd
port 124 nsew
rlabel metal3 s 13670 63460 13670 63460 4 gnd
port 125 nsew
rlabel metal3 s 13982 61296 13982 61296 4 vdd
port 124 nsew
rlabel metal3 s 14487 61887 14487 61887 4 vdd
port 124 nsew
rlabel metal3 s 13415 66007 13415 66007 4 vdd
port 124 nsew
rlabel metal3 s 14918 63460 14918 63460 4 gnd
port 125 nsew
rlabel metal3 s 13427 66845 13427 66845 4 vdd
port 124 nsew
rlabel metal3 s 12038 59708 12038 59708 4 gnd
port 125 nsew
rlabel metal3 s 16983 61887 16983 61887 4 vdd
port 124 nsew
rlabel metal3 s 15923 67167 15923 67167 4 gnd
port 125 nsew
rlabel metal3 s 15923 66845 15923 66845 4 vdd
port 124 nsew
rlabel metal3 s 12734 61296 12734 61296 4 vdd
port 124 nsew
rlabel metal3 s 14745 65233 14745 65233 4 gnd
port 125 nsew
rlabel metal3 s 14675 66845 14675 66845 4 vdd
port 124 nsew
rlabel metal3 s 12038 60182 12038 60182 4 gnd
port 125 nsew
rlabel metal3 s 12038 59392 12038 59392 4 gnd
port 125 nsew
rlabel metal3 s 12038 60498 12038 60498 4 gnd
port 125 nsew
rlabel metal3 s 17102 61296 17102 61296 4 vdd
port 124 nsew
rlabel metal3 s 14675 67167 14675 67167 4 gnd
port 125 nsew
rlabel metal3 s 12038 59155 12038 59155 4 gnd
port 125 nsew
rlabel metal3 s 12038 60972 12038 60972 4 gnd
port 125 nsew
rlabel metal3 s 15735 61887 15735 61887 4 vdd
port 124 nsew
rlabel metal3 s 14606 61296 14606 61296 4 vdd
port 124 nsew
rlabel metal3 s 15993 65233 15993 65233 4 gnd
port 125 nsew
rlabel metal3 s 16478 61296 16478 61296 4 vdd
port 124 nsew
rlabel metal3 s 15230 61296 15230 61296 4 vdd
port 124 nsew
rlabel metal3 s 15854 61296 15854 61296 4 vdd
port 124 nsew
rlabel metal3 s 16166 63460 16166 63460 4 gnd
port 125 nsew
rlabel metal3 s 12038 58918 12038 58918 4 gnd
port 125 nsew
rlabel metal3 s 12038 59945 12038 59945 4 gnd
port 125 nsew
rlabel metal3 s 13239 61887 13239 61887 4 vdd
port 124 nsew
rlabel metal3 s 13358 61296 13358 61296 4 vdd
port 124 nsew
rlabel metal3 s 15911 66007 15911 66007 4 vdd
port 124 nsew
rlabel metal3 s 13497 65233 13497 65233 4 gnd
port 125 nsew
rlabel metal3 s 12038 60735 12038 60735 4 gnd
port 125 nsew
rlabel metal3 s 14101 61887 14101 61887 4 vdd
port 124 nsew
rlabel metal3 s 6682 59960 6682 59960 4 vdd
port 124 nsew
rlabel metal3 s 7064 58789 7064 58789 4 gnd
port 125 nsew
rlabel metal3 s 7336 60369 7336 60369 4 vdd
port 124 nsew
rlabel metal3 s 7336 59184 7336 59184 4 vdd
port 124 nsew
rlabel metal3 s 6250 59170 6250 59170 4 vdd
port 124 nsew
rlabel metal3 s 6250 58812 6250 58812 4 vdd
port 124 nsew
rlabel metal3 s 5825 59228 5825 59228 4 gnd
port 125 nsew
rlabel metal3 s 7064 60369 7064 60369 4 gnd
port 125 nsew
rlabel metal3 s 5825 58812 5825 58812 4 gnd
port 125 nsew
rlabel metal3 s 7336 59579 7336 59579 4 vdd
port 124 nsew
rlabel metal3 s 5825 59602 5825 59602 4 gnd
port 125 nsew
rlabel metal3 s 6250 60392 6250 60392 4 vdd
port 124 nsew
rlabel metal3 s 6682 59602 6682 59602 4 vdd
port 124 nsew
rlabel metal3 s 6250 59602 6250 59602 4 vdd
port 124 nsew
rlabel metal3 s 5825 60392 5825 60392 4 gnd
port 125 nsew
rlabel metal3 s 6682 58812 6682 58812 4 vdd
port 124 nsew
rlabel metal3 s 7336 59974 7336 59974 4 vdd
port 124 nsew
rlabel metal3 s 6682 60392 6682 60392 4 vdd
port 124 nsew
rlabel metal3 s 7064 59184 7064 59184 4 gnd
port 125 nsew
rlabel metal3 s 6250 59960 6250 59960 4 vdd
port 124 nsew
rlabel metal3 s 7064 59974 7064 59974 4 gnd
port 125 nsew
rlabel metal3 s 5825 60018 5825 60018 4 gnd
port 125 nsew
rlabel metal3 s 7336 58789 7336 58789 4 vdd
port 124 nsew
rlabel metal3 s 7064 59579 7064 59579 4 gnd
port 125 nsew
rlabel metal3 s 6682 59170 6682 59170 4 vdd
port 124 nsew
rlabel metal3 s 6250 56442 6250 56442 4 vdd
port 124 nsew
rlabel metal3 s 6682 56010 6682 56010 4 vdd
port 124 nsew
rlabel metal3 s 7064 57604 7064 57604 4 gnd
port 125 nsew
rlabel metal3 s 7064 58394 7064 58394 4 gnd
port 125 nsew
rlabel metal3 s 7064 57999 7064 57999 4 gnd
port 125 nsew
rlabel metal3 s 6682 58380 6682 58380 4 vdd
port 124 nsew
rlabel metal3 s 7336 57209 7336 57209 4 vdd
port 124 nsew
rlabel metal3 s 6250 55652 6250 55652 4 vdd
port 124 nsew
rlabel metal3 s 7064 54839 7064 54839 4 gnd
port 125 nsew
rlabel metal3 s 6682 56442 6682 56442 4 vdd
port 124 nsew
rlabel metal3 s 5825 56858 5825 56858 4 gnd
port 125 nsew
rlabel metal3 s 6682 57590 6682 57590 4 vdd
port 124 nsew
rlabel metal3 s 6250 54862 6250 54862 4 vdd
port 124 nsew
rlabel metal3 s 5825 56442 5825 56442 4 gnd
port 125 nsew
rlabel metal3 s 7336 56024 7336 56024 4 vdd
port 124 nsew
rlabel metal3 s 5825 55278 5825 55278 4 gnd
port 125 nsew
rlabel metal3 s 7064 55629 7064 55629 4 gnd
port 125 nsew
rlabel metal3 s 5825 57232 5825 57232 4 gnd
port 125 nsew
rlabel metal3 s 6250 56800 6250 56800 4 vdd
port 124 nsew
rlabel metal3 s 7336 56419 7336 56419 4 vdd
port 124 nsew
rlabel metal3 s 7064 57209 7064 57209 4 gnd
port 125 nsew
rlabel metal3 s 6682 56800 6682 56800 4 vdd
port 124 nsew
rlabel metal3 s 5825 56068 5825 56068 4 gnd
port 125 nsew
rlabel metal3 s 5825 55652 5825 55652 4 gnd
port 125 nsew
rlabel metal3 s 6250 55220 6250 55220 4 vdd
port 124 nsew
rlabel metal3 s 5825 57648 5825 57648 4 gnd
port 125 nsew
rlabel metal3 s 6682 55220 6682 55220 4 vdd
port 124 nsew
rlabel metal3 s 6250 57590 6250 57590 4 vdd
port 124 nsew
rlabel metal3 s 6250 56010 6250 56010 4 vdd
port 124 nsew
rlabel metal3 s 7336 56814 7336 56814 4 vdd
port 124 nsew
rlabel metal3 s 6250 57232 6250 57232 4 vdd
port 124 nsew
rlabel metal3 s 7064 56419 7064 56419 4 gnd
port 125 nsew
rlabel metal3 s 6250 58380 6250 58380 4 vdd
port 124 nsew
rlabel metal3 s 5825 54862 5825 54862 4 gnd
port 125 nsew
rlabel metal3 s 7064 56814 7064 56814 4 gnd
port 125 nsew
rlabel metal3 s 6682 55652 6682 55652 4 vdd
port 124 nsew
rlabel metal3 s 6682 54862 6682 54862 4 vdd
port 124 nsew
rlabel metal3 s 6250 58022 6250 58022 4 vdd
port 124 nsew
rlabel metal3 s 7064 56024 7064 56024 4 gnd
port 125 nsew
rlabel metal3 s 6682 57232 6682 57232 4 vdd
port 124 nsew
rlabel metal3 s 7336 55234 7336 55234 4 vdd
port 124 nsew
rlabel metal3 s 5825 58022 5825 58022 4 gnd
port 125 nsew
rlabel metal3 s 7336 57604 7336 57604 4 vdd
port 124 nsew
rlabel metal3 s 7336 54839 7336 54839 4 vdd
port 124 nsew
rlabel metal3 s 7336 57999 7336 57999 4 vdd
port 124 nsew
rlabel metal3 s 7064 55234 7064 55234 4 gnd
port 125 nsew
rlabel metal3 s 5825 58438 5825 58438 4 gnd
port 125 nsew
rlabel metal3 s 7336 58394 7336 58394 4 vdd
port 124 nsew
rlabel metal3 s 6682 58022 6682 58022 4 vdd
port 124 nsew
rlabel metal3 s 7336 55629 7336 55629 4 vdd
port 124 nsew
rlabel metal3 s 6250 54430 6250 54430 4 vdd
port 124 nsew
rlabel metal3 s 6250 52492 6250 52492 4 vdd
port 124 nsew
rlabel metal3 s 7064 50494 7064 50494 4 gnd
port 125 nsew
rlabel metal3 s 7336 54444 7336 54444 4 vdd
port 124 nsew
rlabel metal3 s 7336 50889 7336 50889 4 vdd
port 124 nsew
rlabel metal3 s 6682 52492 6682 52492 4 vdd
port 124 nsew
rlabel metal3 s 6682 52850 6682 52850 4 vdd
port 124 nsew
rlabel metal3 s 7336 52074 7336 52074 4 vdd
port 124 nsew
rlabel metal3 s 6250 50480 6250 50480 4 vdd
port 124 nsew
rlabel metal3 s 6250 50912 6250 50912 4 vdd
port 124 nsew
rlabel metal3 s 6250 54072 6250 54072 4 vdd
port 124 nsew
rlabel metal3 s 7064 52864 7064 52864 4 gnd
port 125 nsew
rlabel metal3 s 7064 54444 7064 54444 4 gnd
port 125 nsew
rlabel metal3 s 7064 51679 7064 51679 4 gnd
port 125 nsew
rlabel metal3 s 6682 51270 6682 51270 4 vdd
port 124 nsew
rlabel metal3 s 6250 52850 6250 52850 4 vdd
port 124 nsew
rlabel metal3 s 5825 52908 5825 52908 4 gnd
port 125 nsew
rlabel metal3 s 7336 52864 7336 52864 4 vdd
port 124 nsew
rlabel metal3 s 5825 54072 5825 54072 4 gnd
port 125 nsew
rlabel metal3 s 7336 51679 7336 51679 4 vdd
port 124 nsew
rlabel metal3 s 6682 54430 6682 54430 4 vdd
port 124 nsew
rlabel metal3 s 5825 53698 5825 53698 4 gnd
port 125 nsew
rlabel metal3 s 6250 53282 6250 53282 4 vdd
port 124 nsew
rlabel metal3 s 5825 50912 5825 50912 4 gnd
port 125 nsew
rlabel metal3 s 7064 51284 7064 51284 4 gnd
port 125 nsew
rlabel metal3 s 7064 53654 7064 53654 4 gnd
port 125 nsew
rlabel metal3 s 7336 52469 7336 52469 4 vdd
port 124 nsew
rlabel metal3 s 6250 53640 6250 53640 4 vdd
port 124 nsew
rlabel metal3 s 6250 52060 6250 52060 4 vdd
port 124 nsew
rlabel metal3 s 6682 50912 6682 50912 4 vdd
port 124 nsew
rlabel metal3 s 7064 54049 7064 54049 4 gnd
port 125 nsew
rlabel metal3 s 5825 52492 5825 52492 4 gnd
port 125 nsew
rlabel metal3 s 6682 53640 6682 53640 4 vdd
port 124 nsew
rlabel metal3 s 5825 51328 5825 51328 4 gnd
port 125 nsew
rlabel metal3 s 6250 51270 6250 51270 4 vdd
port 124 nsew
rlabel metal3 s 5825 54488 5825 54488 4 gnd
port 125 nsew
rlabel metal3 s 6682 53282 6682 53282 4 vdd
port 124 nsew
rlabel metal3 s 5825 53282 5825 53282 4 gnd
port 125 nsew
rlabel metal3 s 5825 51702 5825 51702 4 gnd
port 125 nsew
rlabel metal3 s 7336 50494 7336 50494 4 vdd
port 124 nsew
rlabel metal3 s 6682 52060 6682 52060 4 vdd
port 124 nsew
rlabel metal3 s 6250 51702 6250 51702 4 vdd
port 124 nsew
rlabel metal3 s 6682 51702 6682 51702 4 vdd
port 124 nsew
rlabel metal3 s 5825 50538 5825 50538 4 gnd
port 125 nsew
rlabel metal3 s 6682 50480 6682 50480 4 vdd
port 124 nsew
rlabel metal3 s 7336 53259 7336 53259 4 vdd
port 124 nsew
rlabel metal3 s 5825 52118 5825 52118 4 gnd
port 125 nsew
rlabel metal3 s 7336 54049 7336 54049 4 vdd
port 124 nsew
rlabel metal3 s 7336 53654 7336 53654 4 vdd
port 124 nsew
rlabel metal3 s 7064 50889 7064 50889 4 gnd
port 125 nsew
rlabel metal3 s 6682 54072 6682 54072 4 vdd
port 124 nsew
rlabel metal3 s 7064 52074 7064 52074 4 gnd
port 125 nsew
rlabel metal3 s 7064 52469 7064 52469 4 gnd
port 125 nsew
rlabel metal3 s 7336 51284 7336 51284 4 vdd
port 124 nsew
rlabel metal3 s 7064 53259 7064 53259 4 gnd
port 125 nsew
rlabel metal3 s 12038 53625 12038 53625 4 gnd
port 125 nsew
rlabel metal3 s 12038 58602 12038 58602 4 gnd
port 125 nsew
rlabel metal3 s 12038 55758 12038 55758 4 gnd
port 125 nsew
rlabel metal3 s 12038 58128 12038 58128 4 gnd
port 125 nsew
rlabel metal3 s 12038 50465 12038 50465 4 gnd
port 125 nsew
rlabel metal3 s 12038 54968 12038 54968 4 gnd
port 125 nsew
rlabel metal3 s 12038 52598 12038 52598 4 gnd
port 125 nsew
rlabel metal3 s 12038 56232 12038 56232 4 gnd
port 125 nsew
rlabel metal3 s 12038 55205 12038 55205 4 gnd
port 125 nsew
rlabel metal3 s 12038 50702 12038 50702 4 gnd
port 125 nsew
rlabel metal3 s 12038 54415 12038 54415 4 gnd
port 125 nsew
rlabel metal3 s 12038 53862 12038 53862 4 gnd
port 125 nsew
rlabel metal3 s 12038 56548 12038 56548 4 gnd
port 125 nsew
rlabel metal3 s 12038 56785 12038 56785 4 gnd
port 125 nsew
rlabel metal3 s 12038 57812 12038 57812 4 gnd
port 125 nsew
rlabel metal3 s 12038 51492 12038 51492 4 gnd
port 125 nsew
rlabel metal3 s 12038 57575 12038 57575 4 gnd
port 125 nsew
rlabel metal3 s 12038 52835 12038 52835 4 gnd
port 125 nsew
rlabel metal3 s 12038 54652 12038 54652 4 gnd
port 125 nsew
rlabel metal3 s 12038 53388 12038 53388 4 gnd
port 125 nsew
rlabel metal3 s 12038 53072 12038 53072 4 gnd
port 125 nsew
rlabel metal3 s 12038 52045 12038 52045 4 gnd
port 125 nsew
rlabel metal3 s 12038 57022 12038 57022 4 gnd
port 125 nsew
rlabel metal3 s 12038 54178 12038 54178 4 gnd
port 125 nsew
rlabel metal3 s 12038 55995 12038 55995 4 gnd
port 125 nsew
rlabel metal3 s 12038 55442 12038 55442 4 gnd
port 125 nsew
rlabel metal3 s 12038 51808 12038 51808 4 gnd
port 125 nsew
rlabel metal3 s 12038 51255 12038 51255 4 gnd
port 125 nsew
rlabel metal3 s 12038 57338 12038 57338 4 gnd
port 125 nsew
rlabel metal3 s 12038 58365 12038 58365 4 gnd
port 125 nsew
rlabel metal3 s 12038 52282 12038 52282 4 gnd
port 125 nsew
rlabel metal3 s 12038 51018 12038 51018 4 gnd
port 125 nsew
rlabel metal3 s 12038 45962 12038 45962 4 gnd
port 125 nsew
rlabel metal3 s 12038 47068 12038 47068 4 gnd
port 125 nsew
rlabel metal3 s 12038 50228 12038 50228 4 gnd
port 125 nsew
rlabel metal3 s 12038 42328 12038 42328 4 gnd
port 125 nsew
rlabel metal3 s 12038 47858 12038 47858 4 gnd
port 125 nsew
rlabel metal3 s 12038 47305 12038 47305 4 gnd
port 125 nsew
rlabel metal3 s 12038 44935 12038 44935 4 gnd
port 125 nsew
rlabel metal3 s 12038 47542 12038 47542 4 gnd
port 125 nsew
rlabel metal3 s 12038 48648 12038 48648 4 gnd
port 125 nsew
rlabel metal3 s 12038 46515 12038 46515 4 gnd
port 125 nsew
rlabel metal3 s 12038 42802 12038 42802 4 gnd
port 125 nsew
rlabel metal3 s 12038 45725 12038 45725 4 gnd
port 125 nsew
rlabel metal3 s 12038 49122 12038 49122 4 gnd
port 125 nsew
rlabel metal3 s 12038 49912 12038 49912 4 gnd
port 125 nsew
rlabel metal3 s 12038 43908 12038 43908 4 gnd
port 125 nsew
rlabel metal3 s 12038 48095 12038 48095 4 gnd
port 125 nsew
rlabel metal3 s 12038 44382 12038 44382 4 gnd
port 125 nsew
rlabel metal3 s 12038 43118 12038 43118 4 gnd
port 125 nsew
rlabel metal3 s 12038 46752 12038 46752 4 gnd
port 125 nsew
rlabel metal3 s 12038 42565 12038 42565 4 gnd
port 125 nsew
rlabel metal3 s 12038 49438 12038 49438 4 gnd
port 125 nsew
rlabel metal3 s 12038 49675 12038 49675 4 gnd
port 125 nsew
rlabel metal3 s 12038 45172 12038 45172 4 gnd
port 125 nsew
rlabel metal3 s 12038 45488 12038 45488 4 gnd
port 125 nsew
rlabel metal3 s 12038 43592 12038 43592 4 gnd
port 125 nsew
rlabel metal3 s 12038 46278 12038 46278 4 gnd
port 125 nsew
rlabel metal3 s 12038 44698 12038 44698 4 gnd
port 125 nsew
rlabel metal3 s 12038 48332 12038 48332 4 gnd
port 125 nsew
rlabel metal3 s 12038 44145 12038 44145 4 gnd
port 125 nsew
rlabel metal3 s 12038 43355 12038 43355 4 gnd
port 125 nsew
rlabel metal3 s 12038 48885 12038 48885 4 gnd
port 125 nsew
rlabel metal3 s 12038 42012 12038 42012 4 gnd
port 125 nsew
rlabel metal3 s 6250 47752 6250 47752 4 vdd
port 124 nsew
rlabel metal3 s 7336 48124 7336 48124 4 vdd
port 124 nsew
rlabel metal3 s 6682 47320 6682 47320 4 vdd
port 124 nsew
rlabel metal3 s 6250 48542 6250 48542 4 vdd
port 124 nsew
rlabel metal3 s 6682 48900 6682 48900 4 vdd
port 124 nsew
rlabel metal3 s 7336 49704 7336 49704 4 vdd
port 124 nsew
rlabel metal3 s 6250 46962 6250 46962 4 vdd
port 124 nsew
rlabel metal3 s 5825 49332 5825 49332 4 gnd
port 125 nsew
rlabel metal3 s 7336 46939 7336 46939 4 vdd
port 124 nsew
rlabel metal3 s 6250 46530 6250 46530 4 vdd
port 124 nsew
rlabel metal3 s 6682 48110 6682 48110 4 vdd
port 124 nsew
rlabel metal3 s 6682 46530 6682 46530 4 vdd
port 124 nsew
rlabel metal3 s 7336 46544 7336 46544 4 vdd
port 124 nsew
rlabel metal3 s 6682 49332 6682 49332 4 vdd
port 124 nsew
rlabel metal3 s 7064 50099 7064 50099 4 gnd
port 125 nsew
rlabel metal3 s 5825 47752 5825 47752 4 gnd
port 125 nsew
rlabel metal3 s 5825 49748 5825 49748 4 gnd
port 125 nsew
rlabel metal3 s 5825 46588 5825 46588 4 gnd
port 125 nsew
rlabel metal3 s 6682 47752 6682 47752 4 vdd
port 124 nsew
rlabel metal3 s 5825 50122 5825 50122 4 gnd
port 125 nsew
rlabel metal3 s 6250 49332 6250 49332 4 vdd
port 124 nsew
rlabel metal3 s 7064 48914 7064 48914 4 gnd
port 125 nsew
rlabel metal3 s 5825 48958 5825 48958 4 gnd
port 125 nsew
rlabel metal3 s 5825 48542 5825 48542 4 gnd
port 125 nsew
rlabel metal3 s 7064 46939 7064 46939 4 gnd
port 125 nsew
rlabel metal3 s 5825 47378 5825 47378 4 gnd
port 125 nsew
rlabel metal3 s 7336 47334 7336 47334 4 vdd
port 124 nsew
rlabel metal3 s 7064 47334 7064 47334 4 gnd
port 125 nsew
rlabel metal3 s 6682 46962 6682 46962 4 vdd
port 124 nsew
rlabel metal3 s 5825 46962 5825 46962 4 gnd
port 125 nsew
rlabel metal3 s 6250 50122 6250 50122 4 vdd
port 124 nsew
rlabel metal3 s 6250 48900 6250 48900 4 vdd
port 124 nsew
rlabel metal3 s 7336 47729 7336 47729 4 vdd
port 124 nsew
rlabel metal3 s 7336 49309 7336 49309 4 vdd
port 124 nsew
rlabel metal3 s 6682 49690 6682 49690 4 vdd
port 124 nsew
rlabel metal3 s 7336 48914 7336 48914 4 vdd
port 124 nsew
rlabel metal3 s 6250 47320 6250 47320 4 vdd
port 124 nsew
rlabel metal3 s 7064 47729 7064 47729 4 gnd
port 125 nsew
rlabel metal3 s 6250 48110 6250 48110 4 vdd
port 124 nsew
rlabel metal3 s 7064 46544 7064 46544 4 gnd
port 125 nsew
rlabel metal3 s 7064 49309 7064 49309 4 gnd
port 125 nsew
rlabel metal3 s 6250 49690 6250 49690 4 vdd
port 124 nsew
rlabel metal3 s 7336 48519 7336 48519 4 vdd
port 124 nsew
rlabel metal3 s 7064 48519 7064 48519 4 gnd
port 125 nsew
rlabel metal3 s 6682 50122 6682 50122 4 vdd
port 124 nsew
rlabel metal3 s 5825 48168 5825 48168 4 gnd
port 125 nsew
rlabel metal3 s 7064 49704 7064 49704 4 gnd
port 125 nsew
rlabel metal3 s 6682 48542 6682 48542 4 vdd
port 124 nsew
rlabel metal3 s 7064 48124 7064 48124 4 gnd
port 125 nsew
rlabel metal3 s 7336 50099 7336 50099 4 vdd
port 124 nsew
rlabel metal3 s 7064 43779 7064 43779 4 gnd
port 125 nsew
rlabel metal3 s 7336 45359 7336 45359 4 vdd
port 124 nsew
rlabel metal3 s 6682 44160 6682 44160 4 vdd
port 124 nsew
rlabel metal3 s 6250 43802 6250 43802 4 vdd
port 124 nsew
rlabel metal3 s 6250 44160 6250 44160 4 vdd
port 124 nsew
rlabel metal3 s 7064 42594 7064 42594 4 gnd
port 125 nsew
rlabel metal3 s 6682 46172 6682 46172 4 vdd
port 124 nsew
rlabel metal3 s 7336 42989 7336 42989 4 vdd
port 124 nsew
rlabel metal3 s 5825 44218 5825 44218 4 gnd
port 125 nsew
rlabel metal3 s 5825 46172 5825 46172 4 gnd
port 125 nsew
rlabel metal3 s 6682 43802 6682 43802 4 vdd
port 124 nsew
rlabel metal3 s 6682 44950 6682 44950 4 vdd
port 124 nsew
rlabel metal3 s 6682 42580 6682 42580 4 vdd
port 124 nsew
rlabel metal3 s 7064 44569 7064 44569 4 gnd
port 125 nsew
rlabel metal3 s 6250 43370 6250 43370 4 vdd
port 124 nsew
rlabel metal3 s 5825 42222 5825 42222 4 gnd
port 125 nsew
rlabel metal3 s 7064 45754 7064 45754 4 gnd
port 125 nsew
rlabel metal3 s 6682 45740 6682 45740 4 vdd
port 124 nsew
rlabel metal3 s 7336 42594 7336 42594 4 vdd
port 124 nsew
rlabel metal3 s 7336 43384 7336 43384 4 vdd
port 124 nsew
rlabel metal3 s 6250 45740 6250 45740 4 vdd
port 124 nsew
rlabel metal3 s 6250 44592 6250 44592 4 vdd
port 124 nsew
rlabel metal3 s 6250 42222 6250 42222 4 vdd
port 124 nsew
rlabel metal3 s 7064 45359 7064 45359 4 gnd
port 125 nsew
rlabel metal3 s 7064 46149 7064 46149 4 gnd
port 125 nsew
rlabel metal3 s 6250 45382 6250 45382 4 vdd
port 124 nsew
rlabel metal3 s 7064 44174 7064 44174 4 gnd
port 125 nsew
rlabel metal3 s 7336 46149 7336 46149 4 vdd
port 124 nsew
rlabel metal3 s 5825 42638 5825 42638 4 gnd
port 125 nsew
rlabel metal3 s 6682 42222 6682 42222 4 vdd
port 124 nsew
rlabel metal3 s 7336 44569 7336 44569 4 vdd
port 124 nsew
rlabel metal3 s 5825 43012 5825 43012 4 gnd
port 125 nsew
rlabel metal3 s 5825 45382 5825 45382 4 gnd
port 125 nsew
rlabel metal3 s 7336 44174 7336 44174 4 vdd
port 124 nsew
rlabel metal3 s 6682 44592 6682 44592 4 vdd
port 124 nsew
rlabel metal3 s 7336 42199 7336 42199 4 vdd
port 124 nsew
rlabel metal3 s 5825 45798 5825 45798 4 gnd
port 125 nsew
rlabel metal3 s 6682 43370 6682 43370 4 vdd
port 124 nsew
rlabel metal3 s 7064 43384 7064 43384 4 gnd
port 125 nsew
rlabel metal3 s 7336 44964 7336 44964 4 vdd
port 124 nsew
rlabel metal3 s 6250 44950 6250 44950 4 vdd
port 124 nsew
rlabel metal3 s 5825 43428 5825 43428 4 gnd
port 125 nsew
rlabel metal3 s 6682 43012 6682 43012 4 vdd
port 124 nsew
rlabel metal3 s 6250 43012 6250 43012 4 vdd
port 124 nsew
rlabel metal3 s 7336 43779 7336 43779 4 vdd
port 124 nsew
rlabel metal3 s 7064 42989 7064 42989 4 gnd
port 125 nsew
rlabel metal3 s 7064 44964 7064 44964 4 gnd
port 125 nsew
rlabel metal3 s 7336 45754 7336 45754 4 vdd
port 124 nsew
rlabel metal3 s 5825 45008 5825 45008 4 gnd
port 125 nsew
rlabel metal3 s 5825 43802 5825 43802 4 gnd
port 125 nsew
rlabel metal3 s 6682 45382 6682 45382 4 vdd
port 124 nsew
rlabel metal3 s 6250 42580 6250 42580 4 vdd
port 124 nsew
rlabel metal3 s 7064 42199 7064 42199 4 gnd
port 125 nsew
rlabel metal3 s 6250 46172 6250 46172 4 vdd
port 124 nsew
rlabel metal3 s 5825 44592 5825 44592 4 gnd
port 125 nsew
rlabel metal3 s 6250 41000 6250 41000 4 vdd
port 124 nsew
rlabel metal3 s 7336 41014 7336 41014 4 vdd
port 124 nsew
rlabel metal3 s 6250 40210 6250 40210 4 vdd
port 124 nsew
rlabel metal3 s 6250 39420 6250 39420 4 vdd
port 124 nsew
rlabel metal3 s 6250 39852 6250 39852 4 vdd
port 124 nsew
rlabel metal3 s 6250 37840 6250 37840 4 vdd
port 124 nsew
rlabel metal3 s 6250 38272 6250 38272 4 vdd
port 124 nsew
rlabel metal3 s 7064 40224 7064 40224 4 gnd
port 125 nsew
rlabel metal3 s 7336 41409 7336 41409 4 vdd
port 124 nsew
rlabel metal3 s 5825 37898 5825 37898 4 gnd
port 125 nsew
rlabel metal3 s 7336 39039 7336 39039 4 vdd
port 124 nsew
rlabel metal3 s 7064 38644 7064 38644 4 gnd
port 125 nsew
rlabel metal3 s 6682 40210 6682 40210 4 vdd
port 124 nsew
rlabel metal3 s 6682 41000 6682 41000 4 vdd
port 124 nsew
rlabel metal3 s 6682 39852 6682 39852 4 vdd
port 124 nsew
rlabel metal3 s 7336 37854 7336 37854 4 vdd
port 124 nsew
rlabel metal3 s 7336 38644 7336 38644 4 vdd
port 124 nsew
rlabel metal3 s 5825 41432 5825 41432 4 gnd
port 125 nsew
rlabel metal3 s 6682 38272 6682 38272 4 vdd
port 124 nsew
rlabel metal3 s 7064 40619 7064 40619 4 gnd
port 125 nsew
rlabel metal3 s 7064 39039 7064 39039 4 gnd
port 125 nsew
rlabel metal3 s 6250 39062 6250 39062 4 vdd
port 124 nsew
rlabel metal3 s 5825 39478 5825 39478 4 gnd
port 125 nsew
rlabel metal3 s 6682 39062 6682 39062 4 vdd
port 124 nsew
rlabel metal3 s 7064 41014 7064 41014 4 gnd
port 125 nsew
rlabel metal3 s 7336 39829 7336 39829 4 vdd
port 124 nsew
rlabel metal3 s 7336 39434 7336 39434 4 vdd
port 124 nsew
rlabel metal3 s 7336 40224 7336 40224 4 vdd
port 124 nsew
rlabel metal3 s 6250 41790 6250 41790 4 vdd
port 124 nsew
rlabel metal3 s 6682 40642 6682 40642 4 vdd
port 124 nsew
rlabel metal3 s 5825 41848 5825 41848 4 gnd
port 125 nsew
rlabel metal3 s 5825 41058 5825 41058 4 gnd
port 125 nsew
rlabel metal3 s 6682 37840 6682 37840 4 vdd
port 124 nsew
rlabel metal3 s 5825 39062 5825 39062 4 gnd
port 125 nsew
rlabel metal3 s 7336 40619 7336 40619 4 vdd
port 124 nsew
rlabel metal3 s 7064 39829 7064 39829 4 gnd
port 125 nsew
rlabel metal3 s 6682 38630 6682 38630 4 vdd
port 124 nsew
rlabel metal3 s 6682 39420 6682 39420 4 vdd
port 124 nsew
rlabel metal3 s 6682 41432 6682 41432 4 vdd
port 124 nsew
rlabel metal3 s 5825 40268 5825 40268 4 gnd
port 125 nsew
rlabel metal3 s 7064 41409 7064 41409 4 gnd
port 125 nsew
rlabel metal3 s 5825 38688 5825 38688 4 gnd
port 125 nsew
rlabel metal3 s 5825 38272 5825 38272 4 gnd
port 125 nsew
rlabel metal3 s 7336 38249 7336 38249 4 vdd
port 124 nsew
rlabel metal3 s 5825 39852 5825 39852 4 gnd
port 125 nsew
rlabel metal3 s 6250 38630 6250 38630 4 vdd
port 124 nsew
rlabel metal3 s 7336 41804 7336 41804 4 vdd
port 124 nsew
rlabel metal3 s 7064 38249 7064 38249 4 gnd
port 125 nsew
rlabel metal3 s 7064 37854 7064 37854 4 gnd
port 125 nsew
rlabel metal3 s 7064 41804 7064 41804 4 gnd
port 125 nsew
rlabel metal3 s 6682 41790 6682 41790 4 vdd
port 124 nsew
rlabel metal3 s 6250 41432 6250 41432 4 vdd
port 124 nsew
rlabel metal3 s 5825 40642 5825 40642 4 gnd
port 125 nsew
rlabel metal3 s 7064 39434 7064 39434 4 gnd
port 125 nsew
rlabel metal3 s 6250 40642 6250 40642 4 vdd
port 124 nsew
rlabel metal3 s 5825 35528 5825 35528 4 gnd
port 125 nsew
rlabel metal3 s 5825 34322 5825 34322 4 gnd
port 125 nsew
rlabel metal3 s 6682 35470 6682 35470 4 vdd
port 124 nsew
rlabel metal3 s 7064 33904 7064 33904 4 gnd
port 125 nsew
rlabel metal3 s 6250 36692 6250 36692 4 vdd
port 124 nsew
rlabel metal3 s 6250 35112 6250 35112 4 vdd
port 124 nsew
rlabel metal3 s 6682 36692 6682 36692 4 vdd
port 124 nsew
rlabel metal3 s 5825 34738 5825 34738 4 gnd
port 125 nsew
rlabel metal3 s 6682 36260 6682 36260 4 vdd
port 124 nsew
rlabel metal3 s 6682 37482 6682 37482 4 vdd
port 124 nsew
rlabel metal3 s 6682 34680 6682 34680 4 vdd
port 124 nsew
rlabel metal3 s 7782 35440 7782 35440 4 gnd
port 125 nsew
rlabel metal3 s 6250 36260 6250 36260 4 vdd
port 124 nsew
rlabel metal3 s 5825 35112 5825 35112 4 gnd
port 125 nsew
rlabel metal3 s 6250 34322 6250 34322 4 vdd
port 124 nsew
rlabel metal3 s 6682 34322 6682 34322 4 vdd
port 124 nsew
rlabel metal3 s 7064 35089 7064 35089 4 gnd
port 125 nsew
rlabel metal3 s 7336 36669 7336 36669 4 vdd
port 124 nsew
rlabel metal3 s 5825 36318 5825 36318 4 gnd
port 125 nsew
rlabel metal3 s 7336 34694 7336 34694 4 vdd
port 124 nsew
rlabel metal3 s 5825 37482 5825 37482 4 gnd
port 125 nsew
rlabel metal3 s 5825 33948 5825 33948 4 gnd
port 125 nsew
rlabel metal3 s 7064 37064 7064 37064 4 gnd
port 125 nsew
rlabel metal3 s 7064 34299 7064 34299 4 gnd
port 125 nsew
rlabel metal3 s 6250 37482 6250 37482 4 vdd
port 124 nsew
rlabel metal3 s 7064 34694 7064 34694 4 gnd
port 125 nsew
rlabel metal3 s 6682 35112 6682 35112 4 vdd
port 124 nsew
rlabel metal3 s 8207 35439 8207 35439 4 vdd
port 124 nsew
rlabel metal3 s 7064 36669 7064 36669 4 gnd
port 125 nsew
rlabel metal3 s 6250 35902 6250 35902 4 vdd
port 124 nsew
rlabel metal3 s 7336 34299 7336 34299 4 vdd
port 124 nsew
rlabel metal3 s 6682 35902 6682 35902 4 vdd
port 124 nsew
rlabel metal3 s 5825 37108 5825 37108 4 gnd
port 125 nsew
rlabel metal3 s 6250 33890 6250 33890 4 vdd
port 124 nsew
rlabel metal3 s 6682 37050 6682 37050 4 vdd
port 124 nsew
rlabel metal3 s 7336 36274 7336 36274 4 vdd
port 124 nsew
rlabel metal3 s 7336 37064 7336 37064 4 vdd
port 124 nsew
rlabel metal3 s 7336 35089 7336 35089 4 vdd
port 124 nsew
rlabel metal3 s 5825 35902 5825 35902 4 gnd
port 125 nsew
rlabel metal3 s 7064 37459 7064 37459 4 gnd
port 125 nsew
rlabel metal3 s 7336 35879 7336 35879 4 vdd
port 124 nsew
rlabel metal3 s 7336 37459 7336 37459 4 vdd
port 124 nsew
rlabel metal3 s 6250 35470 6250 35470 4 vdd
port 124 nsew
rlabel metal3 s 6682 33890 6682 33890 4 vdd
port 124 nsew
rlabel metal3 s 6250 37050 6250 37050 4 vdd
port 124 nsew
rlabel metal3 s 6250 34680 6250 34680 4 vdd
port 124 nsew
rlabel metal3 s 7064 36274 7064 36274 4 gnd
port 125 nsew
rlabel metal3 s 7336 35484 7336 35484 4 vdd
port 124 nsew
rlabel metal3 s 5825 36692 5825 36692 4 gnd
port 125 nsew
rlabel metal3 s 7336 33904 7336 33904 4 vdd
port 124 nsew
rlabel metal3 s 7064 35484 7064 35484 4 gnd
port 125 nsew
rlabel metal3 s 7064 35879 7064 35879 4 gnd
port 125 nsew
rlabel metal3 s 12038 41222 12038 41222 4 gnd
port 125 nsew
rlabel metal3 s 10774 35455 10774 35455 4 vdd
port 124 nsew
rlabel metal3 s 12038 34112 12038 34112 4 gnd
port 125 nsew
rlabel metal3 s 12038 36798 12038 36798 4 gnd
port 125 nsew
rlabel metal3 s 12038 40195 12038 40195 4 gnd
port 125 nsew
rlabel metal3 s 12038 33875 12038 33875 4 gnd
port 125 nsew
rlabel metal3 s 12038 38062 12038 38062 4 gnd
port 125 nsew
rlabel metal3 s 12038 34665 12038 34665 4 gnd
port 125 nsew
rlabel metal3 s 12038 34902 12038 34902 4 gnd
port 125 nsew
rlabel metal3 s 12038 40748 12038 40748 4 gnd
port 125 nsew
rlabel metal3 s 12038 36008 12038 36008 4 gnd
port 125 nsew
rlabel metal3 s 12038 38378 12038 38378 4 gnd
port 125 nsew
rlabel metal3 s 12038 40432 12038 40432 4 gnd
port 125 nsew
rlabel metal3 s 12038 39405 12038 39405 4 gnd
port 125 nsew
rlabel metal3 s 12038 35455 12038 35455 4 gnd
port 125 nsew
rlabel metal3 s 12038 41538 12038 41538 4 gnd
port 125 nsew
rlabel metal3 s 12038 37588 12038 37588 4 gnd
port 125 nsew
rlabel metal3 s 12038 38852 12038 38852 4 gnd
port 125 nsew
rlabel metal3 s 12038 39168 12038 39168 4 gnd
port 125 nsew
rlabel metal3 s 12038 36482 12038 36482 4 gnd
port 125 nsew
rlabel metal3 s 12038 34428 12038 34428 4 gnd
port 125 nsew
rlabel metal3 s 9250 35455 9250 35455 4 gnd
port 125 nsew
rlabel metal3 s 12038 37035 12038 37035 4 gnd
port 125 nsew
rlabel metal3 s 12038 36245 12038 36245 4 gnd
port 125 nsew
rlabel metal3 s 12038 38615 12038 38615 4 gnd
port 125 nsew
rlabel metal3 s 12038 40985 12038 40985 4 gnd
port 125 nsew
rlabel metal3 s 12038 33638 12038 33638 4 gnd
port 125 nsew
rlabel metal3 s 12038 37272 12038 37272 4 gnd
port 125 nsew
rlabel metal3 s 12038 41775 12038 41775 4 gnd
port 125 nsew
rlabel metal3 s 12038 35692 12038 35692 4 gnd
port 125 nsew
rlabel metal3 s 12038 39958 12038 39958 4 gnd
port 125 nsew
rlabel metal3 s 12038 35218 12038 35218 4 gnd
port 125 nsew
rlabel metal3 s 12038 37825 12038 37825 4 gnd
port 125 nsew
rlabel metal3 s 12038 39642 12038 39642 4 gnd
port 125 nsew
rlabel metal3 s 12038 30478 12038 30478 4 gnd
port 125 nsew
rlabel metal3 s 12038 32295 12038 32295 4 gnd
port 125 nsew
rlabel metal3 s 12038 28345 12038 28345 4 gnd
port 125 nsew
rlabel metal3 s 12038 25738 12038 25738 4 gnd
port 125 nsew
rlabel metal3 s 12038 31268 12038 31268 4 gnd
port 125 nsew
rlabel metal3 s 12038 27002 12038 27002 4 gnd
port 125 nsew
rlabel metal3 s 12038 30952 12038 30952 4 gnd
port 125 nsew
rlabel metal3 s 12038 27555 12038 27555 4 gnd
port 125 nsew
rlabel metal3 s 12038 32058 12038 32058 4 gnd
port 125 nsew
rlabel metal3 s 12038 33322 12038 33322 4 gnd
port 125 nsew
rlabel metal3 s 12038 31505 12038 31505 4 gnd
port 125 nsew
rlabel metal3 s 12038 25422 12038 25422 4 gnd
port 125 nsew
rlabel metal3 s 12038 29135 12038 29135 4 gnd
port 125 nsew
rlabel metal3 s 12038 30715 12038 30715 4 gnd
port 125 nsew
rlabel metal3 s 12038 26212 12038 26212 4 gnd
port 125 nsew
rlabel metal3 s 12038 30162 12038 30162 4 gnd
port 125 nsew
rlabel metal3 s 12038 29688 12038 29688 4 gnd
port 125 nsew
rlabel metal3 s 12038 32532 12038 32532 4 gnd
port 125 nsew
rlabel metal3 s 12038 28898 12038 28898 4 gnd
port 125 nsew
rlabel metal3 s 12038 27792 12038 27792 4 gnd
port 125 nsew
rlabel metal3 s 12038 29372 12038 29372 4 gnd
port 125 nsew
rlabel metal3 s 12038 29925 12038 29925 4 gnd
port 125 nsew
rlabel metal3 s 12038 33085 12038 33085 4 gnd
port 125 nsew
rlabel metal3 s 12038 26765 12038 26765 4 gnd
port 125 nsew
rlabel metal3 s 12038 26528 12038 26528 4 gnd
port 125 nsew
rlabel metal3 s 12038 28108 12038 28108 4 gnd
port 125 nsew
rlabel metal3 s 12038 31742 12038 31742 4 gnd
port 125 nsew
rlabel metal3 s 12038 28582 12038 28582 4 gnd
port 125 nsew
rlabel metal3 s 12038 25975 12038 25975 4 gnd
port 125 nsew
rlabel metal3 s 12038 32848 12038 32848 4 gnd
port 125 nsew
rlabel metal3 s 12038 27318 12038 27318 4 gnd
port 125 nsew
rlabel metal3 s 7064 31534 7064 31534 4 gnd
port 125 nsew
rlabel metal3 s 7336 31534 7336 31534 4 vdd
port 124 nsew
rlabel metal3 s 7336 31929 7336 31929 4 vdd
port 124 nsew
rlabel metal3 s 6250 31952 6250 31952 4 vdd
port 124 nsew
rlabel metal3 s 6250 32742 6250 32742 4 vdd
port 124 nsew
rlabel metal3 s 5825 32368 5825 32368 4 gnd
port 125 nsew
rlabel metal3 s 7336 30349 7336 30349 4 vdd
port 124 nsew
rlabel metal3 s 6250 33532 6250 33532 4 vdd
port 124 nsew
rlabel metal3 s 7064 31929 7064 31929 4 gnd
port 125 nsew
rlabel metal3 s 7064 29559 7064 29559 4 gnd
port 125 nsew
rlabel metal3 s 6682 29940 6682 29940 4 vdd
port 124 nsew
rlabel metal3 s 6250 29940 6250 29940 4 vdd
port 124 nsew
rlabel metal3 s 6682 31162 6682 31162 4 vdd
port 124 nsew
rlabel metal3 s 6250 30372 6250 30372 4 vdd
port 124 nsew
rlabel metal3 s 7336 32324 7336 32324 4 vdd
port 124 nsew
rlabel metal3 s 7336 29954 7336 29954 4 vdd
port 124 nsew
rlabel metal3 s 7064 33114 7064 33114 4 gnd
port 125 nsew
rlabel metal3 s 5825 31578 5825 31578 4 gnd
port 125 nsew
rlabel metal3 s 6250 32310 6250 32310 4 vdd
port 124 nsew
rlabel metal3 s 6682 31952 6682 31952 4 vdd
port 124 nsew
rlabel metal3 s 5825 33532 5825 33532 4 gnd
port 125 nsew
rlabel metal3 s 7064 30744 7064 30744 4 gnd
port 125 nsew
rlabel metal3 s 6682 33100 6682 33100 4 vdd
port 124 nsew
rlabel metal3 s 5825 33158 5825 33158 4 gnd
port 125 nsew
rlabel metal3 s 5825 31952 5825 31952 4 gnd
port 125 nsew
rlabel metal3 s 6682 32742 6682 32742 4 vdd
port 124 nsew
rlabel metal3 s 6250 31520 6250 31520 4 vdd
port 124 nsew
rlabel metal3 s 6250 29582 6250 29582 4 vdd
port 124 nsew
rlabel metal3 s 7336 29559 7336 29559 4 vdd
port 124 nsew
rlabel metal3 s 6682 32310 6682 32310 4 vdd
port 124 nsew
rlabel metal3 s 7336 32719 7336 32719 4 vdd
port 124 nsew
rlabel metal3 s 6682 31520 6682 31520 4 vdd
port 124 nsew
rlabel metal3 s 7064 33509 7064 33509 4 gnd
port 125 nsew
rlabel metal3 s 6250 30730 6250 30730 4 vdd
port 124 nsew
rlabel metal3 s 6682 33532 6682 33532 4 vdd
port 124 nsew
rlabel metal3 s 7064 29954 7064 29954 4 gnd
port 125 nsew
rlabel metal3 s 6682 30372 6682 30372 4 vdd
port 124 nsew
rlabel metal3 s 5825 29582 5825 29582 4 gnd
port 125 nsew
rlabel metal3 s 7064 32324 7064 32324 4 gnd
port 125 nsew
rlabel metal3 s 5825 29998 5825 29998 4 gnd
port 125 nsew
rlabel metal3 s 7064 30349 7064 30349 4 gnd
port 125 nsew
rlabel metal3 s 7064 32719 7064 32719 4 gnd
port 125 nsew
rlabel metal3 s 5825 31162 5825 31162 4 gnd
port 125 nsew
rlabel metal3 s 7336 33114 7336 33114 4 vdd
port 124 nsew
rlabel metal3 s 6682 30730 6682 30730 4 vdd
port 124 nsew
rlabel metal3 s 7064 31139 7064 31139 4 gnd
port 125 nsew
rlabel metal3 s 5825 30788 5825 30788 4 gnd
port 125 nsew
rlabel metal3 s 6250 33100 6250 33100 4 vdd
port 124 nsew
rlabel metal3 s 7336 33509 7336 33509 4 vdd
port 124 nsew
rlabel metal3 s 6250 31162 6250 31162 4 vdd
port 124 nsew
rlabel metal3 s 7336 30744 7336 30744 4 vdd
port 124 nsew
rlabel metal3 s 7336 31139 7336 31139 4 vdd
port 124 nsew
rlabel metal3 s 6682 29582 6682 29582 4 vdd
port 124 nsew
rlabel metal3 s 5825 32742 5825 32742 4 gnd
port 125 nsew
rlabel metal3 s 5825 30372 5825 30372 4 gnd
port 125 nsew
rlabel metal3 s 6250 28360 6250 28360 4 vdd
port 124 nsew
rlabel metal3 s 6682 28360 6682 28360 4 vdd
port 124 nsew
rlabel metal3 s 6682 27212 6682 27212 4 vdd
port 124 nsew
rlabel metal3 s 7336 26794 7336 26794 4 vdd
port 124 nsew
rlabel metal3 s 7064 27979 7064 27979 4 gnd
port 125 nsew
rlabel metal3 s 7064 28769 7064 28769 4 gnd
port 125 nsew
rlabel metal3 s 5825 28418 5825 28418 4 gnd
port 125 nsew
rlabel metal3 s 7064 26794 7064 26794 4 gnd
port 125 nsew
rlabel metal3 s 7336 25214 7336 25214 4 vdd
port 124 nsew
rlabel metal3 s 5825 26422 5825 26422 4 gnd
port 125 nsew
rlabel metal3 s 6250 27570 6250 27570 4 vdd
port 124 nsew
rlabel metal3 s 6250 25200 6250 25200 4 vdd
port 124 nsew
rlabel metal3 s 5825 28002 5825 28002 4 gnd
port 125 nsew
rlabel metal3 s 7336 27189 7336 27189 4 vdd
port 124 nsew
rlabel metal3 s 7336 27979 7336 27979 4 vdd
port 124 nsew
rlabel metal3 s 5825 27628 5825 27628 4 gnd
port 125 nsew
rlabel metal3 s 6682 25990 6682 25990 4 vdd
port 124 nsew
rlabel metal3 s 5825 26048 5825 26048 4 gnd
port 125 nsew
rlabel metal3 s 5825 25258 5825 25258 4 gnd
port 125 nsew
rlabel metal3 s 6682 28002 6682 28002 4 vdd
port 124 nsew
rlabel metal3 s 7336 25609 7336 25609 4 vdd
port 124 nsew
rlabel metal3 s 7336 27584 7336 27584 4 vdd
port 124 nsew
rlabel metal3 s 6682 25632 6682 25632 4 vdd
port 124 nsew
rlabel metal3 s 6682 26780 6682 26780 4 vdd
port 124 nsew
rlabel metal3 s 6682 26422 6682 26422 4 vdd
port 124 nsew
rlabel metal3 s 6682 29150 6682 29150 4 vdd
port 124 nsew
rlabel metal3 s 6682 28792 6682 28792 4 vdd
port 124 nsew
rlabel metal3 s 6250 25990 6250 25990 4 vdd
port 124 nsew
rlabel metal3 s 7336 28374 7336 28374 4 vdd
port 124 nsew
rlabel metal3 s 6250 26422 6250 26422 4 vdd
port 124 nsew
rlabel metal3 s 7064 25214 7064 25214 4 gnd
port 125 nsew
rlabel metal3 s 5825 27212 5825 27212 4 gnd
port 125 nsew
rlabel metal3 s 7336 29164 7336 29164 4 vdd
port 124 nsew
rlabel metal3 s 5825 28792 5825 28792 4 gnd
port 125 nsew
rlabel metal3 s 7336 28769 7336 28769 4 vdd
port 124 nsew
rlabel metal3 s 6250 25632 6250 25632 4 vdd
port 124 nsew
rlabel metal3 s 6250 28002 6250 28002 4 vdd
port 124 nsew
rlabel metal3 s 7064 25609 7064 25609 4 gnd
port 125 nsew
rlabel metal3 s 7064 27584 7064 27584 4 gnd
port 125 nsew
rlabel metal3 s 7064 27189 7064 27189 4 gnd
port 125 nsew
rlabel metal3 s 7064 26399 7064 26399 4 gnd
port 125 nsew
rlabel metal3 s 7064 29164 7064 29164 4 gnd
port 125 nsew
rlabel metal3 s 7336 26004 7336 26004 4 vdd
port 124 nsew
rlabel metal3 s 6250 28792 6250 28792 4 vdd
port 124 nsew
rlabel metal3 s 7064 26004 7064 26004 4 gnd
port 125 nsew
rlabel metal3 s 5825 29208 5825 29208 4 gnd
port 125 nsew
rlabel metal3 s 5825 25632 5825 25632 4 gnd
port 125 nsew
rlabel metal3 s 7336 26399 7336 26399 4 vdd
port 124 nsew
rlabel metal3 s 5825 26838 5825 26838 4 gnd
port 125 nsew
rlabel metal3 s 6682 27570 6682 27570 4 vdd
port 124 nsew
rlabel metal3 s 7064 28374 7064 28374 4 gnd
port 125 nsew
rlabel metal3 s 6250 27212 6250 27212 4 vdd
port 124 nsew
rlabel metal3 s 6250 26780 6250 26780 4 vdd
port 124 nsew
rlabel metal3 s 6250 29150 6250 29150 4 vdd
port 124 nsew
rlabel metal3 s 6682 25200 6682 25200 4 vdd
port 124 nsew
rlabel metal3 s 5825 24468 5825 24468 4 gnd
port 125 nsew
rlabel metal3 s 5825 22888 5825 22888 4 gnd
port 125 nsew
rlabel metal3 s 6250 24052 6250 24052 4 vdd
port 124 nsew
rlabel metal3 s 6682 21682 6682 21682 4 vdd
port 124 nsew
rlabel metal3 s 6250 22830 6250 22830 4 vdd
port 124 nsew
rlabel metal3 s 6682 22472 6682 22472 4 vdd
port 124 nsew
rlabel metal3 s 5825 21308 5825 21308 4 gnd
port 125 nsew
rlabel metal3 s 7336 21264 7336 21264 4 vdd
port 124 nsew
rlabel metal3 s 6682 21250 6682 21250 4 vdd
port 124 nsew
rlabel metal3 s 7336 21659 7336 21659 4 vdd
port 124 nsew
rlabel metal3 s 5825 22472 5825 22472 4 gnd
port 125 nsew
rlabel metal3 s 6682 22830 6682 22830 4 vdd
port 124 nsew
rlabel metal3 s 7064 24819 7064 24819 4 gnd
port 125 nsew
rlabel metal3 s 7336 24029 7336 24029 4 vdd
port 124 nsew
rlabel metal3 s 7064 23239 7064 23239 4 gnd
port 125 nsew
rlabel metal3 s 7336 23634 7336 23634 4 vdd
port 124 nsew
rlabel metal3 s 7064 24424 7064 24424 4 gnd
port 125 nsew
rlabel metal3 s 6250 23620 6250 23620 4 vdd
port 124 nsew
rlabel metal3 s 7336 23239 7336 23239 4 vdd
port 124 nsew
rlabel metal3 s 6250 21250 6250 21250 4 vdd
port 124 nsew
rlabel metal3 s 6250 22040 6250 22040 4 vdd
port 124 nsew
rlabel metal3 s 5825 24842 5825 24842 4 gnd
port 125 nsew
rlabel metal3 s 6250 24410 6250 24410 4 vdd
port 124 nsew
rlabel metal3 s 7336 22054 7336 22054 4 vdd
port 124 nsew
rlabel metal3 s 6682 24842 6682 24842 4 vdd
port 124 nsew
rlabel metal3 s 7336 22449 7336 22449 4 vdd
port 124 nsew
rlabel metal3 s 6250 23262 6250 23262 4 vdd
port 124 nsew
rlabel metal3 s 7064 22844 7064 22844 4 gnd
port 125 nsew
rlabel metal3 s 7064 22449 7064 22449 4 gnd
port 125 nsew
rlabel metal3 s 6682 24052 6682 24052 4 vdd
port 124 nsew
rlabel metal3 s 6682 24410 6682 24410 4 vdd
port 124 nsew
rlabel metal3 s 7336 24819 7336 24819 4 vdd
port 124 nsew
rlabel metal3 s 5825 22098 5825 22098 4 gnd
port 125 nsew
rlabel metal3 s 7064 23634 7064 23634 4 gnd
port 125 nsew
rlabel metal3 s 7064 21659 7064 21659 4 gnd
port 125 nsew
rlabel metal3 s 6250 22472 6250 22472 4 vdd
port 124 nsew
rlabel metal3 s 5825 21682 5825 21682 4 gnd
port 125 nsew
rlabel metal3 s 7064 21264 7064 21264 4 gnd
port 125 nsew
rlabel metal3 s 6682 23262 6682 23262 4 vdd
port 124 nsew
rlabel metal3 s 7336 22844 7336 22844 4 vdd
port 124 nsew
rlabel metal3 s 5825 23262 5825 23262 4 gnd
port 125 nsew
rlabel metal3 s 6682 22040 6682 22040 4 vdd
port 124 nsew
rlabel metal3 s 6682 23620 6682 23620 4 vdd
port 124 nsew
rlabel metal3 s 7336 24424 7336 24424 4 vdd
port 124 nsew
rlabel metal3 s 5825 23678 5825 23678 4 gnd
port 125 nsew
rlabel metal3 s 7064 22054 7064 22054 4 gnd
port 125 nsew
rlabel metal3 s 6250 21682 6250 21682 4 vdd
port 124 nsew
rlabel metal3 s 7064 24029 7064 24029 4 gnd
port 125 nsew
rlabel metal3 s 5825 24052 5825 24052 4 gnd
port 125 nsew
rlabel metal3 s 6250 24842 6250 24842 4 vdd
port 124 nsew
rlabel metal3 s 3392 16942 3392 16942 4 vdd
port 124 nsew
rlabel metal3 s 2960 16942 2960 16942 4 vdd
port 124 nsew
rlabel metal3 s 3774 16919 3774 16919 4 gnd
port 125 nsew
rlabel metal3 s 3392 17732 3392 17732 4 vdd
port 124 nsew
rlabel metal3 s 4046 17709 4046 17709 4 vdd
port 124 nsew
rlabel metal3 s 3774 17709 3774 17709 4 gnd
port 125 nsew
rlabel metal3 s 2535 16942 2535 16942 4 gnd
port 125 nsew
rlabel metal3 s 2960 17732 2960 17732 4 vdd
port 124 nsew
rlabel metal3 s 2535 17732 2535 17732 4 gnd
port 125 nsew
rlabel metal3 s 4046 16919 4046 16919 4 vdd
port 124 nsew
rlabel metal3 s 6682 18522 6682 18522 4 vdd
port 124 nsew
rlabel metal3 s 6682 19312 6682 19312 4 vdd
port 124 nsew
rlabel metal3 s 6250 18090 6250 18090 4 vdd
port 124 nsew
rlabel metal3 s 7064 18499 7064 18499 4 gnd
port 125 nsew
rlabel metal3 s 7336 18894 7336 18894 4 vdd
port 124 nsew
rlabel metal3 s 6682 17300 6682 17300 4 vdd
port 124 nsew
rlabel metal3 s 7336 20474 7336 20474 4 vdd
port 124 nsew
rlabel metal3 s 6250 18522 6250 18522 4 vdd
port 124 nsew
rlabel metal3 s 7064 17314 7064 17314 4 gnd
port 125 nsew
rlabel metal3 s 7064 16919 7064 16919 4 gnd
port 125 nsew
rlabel metal3 s 7336 18499 7336 18499 4 vdd
port 124 nsew
rlabel metal3 s 7336 16919 7336 16919 4 vdd
port 124 nsew
rlabel metal3 s 7064 19289 7064 19289 4 gnd
port 125 nsew
rlabel metal3 s 7336 19289 7336 19289 4 vdd
port 124 nsew
rlabel metal3 s 5825 20102 5825 20102 4 gnd
port 125 nsew
rlabel metal3 s 6682 19670 6682 19670 4 vdd
port 124 nsew
rlabel metal3 s 6250 19312 6250 19312 4 vdd
port 124 nsew
rlabel metal3 s 6250 17300 6250 17300 4 vdd
port 124 nsew
rlabel metal3 s 5825 20892 5825 20892 4 gnd
port 125 nsew
rlabel metal3 s 7064 18104 7064 18104 4 gnd
port 125 nsew
rlabel metal3 s 7064 19684 7064 19684 4 gnd
port 125 nsew
rlabel metal3 s 6250 20102 6250 20102 4 vdd
port 124 nsew
rlabel metal3 s 6682 18090 6682 18090 4 vdd
port 124 nsew
rlabel metal3 s 6250 20460 6250 20460 4 vdd
port 124 nsew
rlabel metal3 s 5825 19728 5825 19728 4 gnd
port 125 nsew
rlabel metal3 s 6250 16942 6250 16942 4 vdd
port 124 nsew
rlabel metal3 s 7336 19684 7336 19684 4 vdd
port 124 nsew
rlabel metal3 s 7336 17709 7336 17709 4 vdd
port 124 nsew
rlabel metal3 s 6682 20102 6682 20102 4 vdd
port 124 nsew
rlabel metal3 s 5825 18148 5825 18148 4 gnd
port 125 nsew
rlabel metal3 s 5825 17358 5825 17358 4 gnd
port 125 nsew
rlabel metal3 s 5825 19312 5825 19312 4 gnd
port 125 nsew
rlabel metal3 s 7064 20869 7064 20869 4 gnd
port 125 nsew
rlabel metal3 s 7064 17709 7064 17709 4 gnd
port 125 nsew
rlabel metal3 s 6682 16942 6682 16942 4 vdd
port 124 nsew
rlabel metal3 s 7336 20869 7336 20869 4 vdd
port 124 nsew
rlabel metal3 s 5825 20518 5825 20518 4 gnd
port 125 nsew
rlabel metal3 s 5825 18938 5825 18938 4 gnd
port 125 nsew
rlabel metal3 s 5825 17732 5825 17732 4 gnd
port 125 nsew
rlabel metal3 s 6250 19670 6250 19670 4 vdd
port 124 nsew
rlabel metal3 s 7336 17314 7336 17314 4 vdd
port 124 nsew
rlabel metal3 s 6682 20892 6682 20892 4 vdd
port 124 nsew
rlabel metal3 s 6682 18880 6682 18880 4 vdd
port 124 nsew
rlabel metal3 s 5825 16942 5825 16942 4 gnd
port 125 nsew
rlabel metal3 s 6250 18880 6250 18880 4 vdd
port 124 nsew
rlabel metal3 s 7336 20079 7336 20079 4 vdd
port 124 nsew
rlabel metal3 s 6682 17732 6682 17732 4 vdd
port 124 nsew
rlabel metal3 s 7064 18894 7064 18894 4 gnd
port 125 nsew
rlabel metal3 s 5825 18522 5825 18522 4 gnd
port 125 nsew
rlabel metal3 s 7064 20079 7064 20079 4 gnd
port 125 nsew
rlabel metal3 s 6250 20892 6250 20892 4 vdd
port 124 nsew
rlabel metal3 s 7064 20474 7064 20474 4 gnd
port 125 nsew
rlabel metal3 s 6250 17732 6250 17732 4 vdd
port 124 nsew
rlabel metal3 s 6682 20460 6682 20460 4 vdd
port 124 nsew
rlabel metal3 s 7336 18104 7336 18104 4 vdd
port 124 nsew
rlabel metal3 s 12038 24948 12038 24948 4 gnd
port 125 nsew
rlabel metal3 s 12038 22025 12038 22025 4 gnd
port 125 nsew
rlabel metal3 s 12038 21788 12038 21788 4 gnd
port 125 nsew
rlabel metal3 s 12038 20445 12038 20445 4 gnd
port 125 nsew
rlabel metal3 s 12038 17838 12038 17838 4 gnd
port 125 nsew
rlabel metal3 s 12038 21472 12038 21472 4 gnd
port 125 nsew
rlabel metal3 s 12038 24158 12038 24158 4 gnd
port 125 nsew
rlabel metal3 s 12038 18075 12038 18075 4 gnd
port 125 nsew
rlabel metal3 s 12038 24632 12038 24632 4 gnd
port 125 nsew
rlabel metal3 s 12038 25185 12038 25185 4 gnd
port 125 nsew
rlabel metal3 s 12038 23842 12038 23842 4 gnd
port 125 nsew
rlabel metal3 s 12038 18312 12038 18312 4 gnd
port 125 nsew
rlabel metal3 s 12038 23368 12038 23368 4 gnd
port 125 nsew
rlabel metal3 s 12038 17522 12038 17522 4 gnd
port 125 nsew
rlabel metal3 s 12038 23605 12038 23605 4 gnd
port 125 nsew
rlabel metal3 s 12038 17048 12038 17048 4 gnd
port 125 nsew
rlabel metal3 s 12038 20682 12038 20682 4 gnd
port 125 nsew
rlabel metal3 s 12038 18628 12038 18628 4 gnd
port 125 nsew
rlabel metal3 s 12038 19892 12038 19892 4 gnd
port 125 nsew
rlabel metal3 s 12038 20208 12038 20208 4 gnd
port 125 nsew
rlabel metal3 s 12038 22578 12038 22578 4 gnd
port 125 nsew
rlabel metal3 s 12038 19655 12038 19655 4 gnd
port 125 nsew
rlabel metal3 s 12038 19418 12038 19418 4 gnd
port 125 nsew
rlabel metal3 s 12038 17285 12038 17285 4 gnd
port 125 nsew
rlabel metal3 s 12038 19102 12038 19102 4 gnd
port 125 nsew
rlabel metal3 s 12038 23052 12038 23052 4 gnd
port 125 nsew
rlabel metal3 s 12038 20998 12038 20998 4 gnd
port 125 nsew
rlabel metal3 s 12038 22815 12038 22815 4 gnd
port 125 nsew
rlabel metal3 s 12038 21235 12038 21235 4 gnd
port 125 nsew
rlabel metal3 s 12038 22262 12038 22262 4 gnd
port 125 nsew
rlabel metal3 s 12038 18865 12038 18865 4 gnd
port 125 nsew
rlabel metal3 s 12038 24395 12038 24395 4 gnd
port 125 nsew
rlabel metal3 s 14606 9614 14606 9614 4 vdd
port 124 nsew
rlabel metal3 s 17102 9614 17102 9614 4 vdd
port 124 nsew
rlabel metal3 s 16597 9023 16597 9023 4 vdd
port 124 nsew
rlabel metal3 s 12853 9023 12853 9023 4 vdd
port 124 nsew
rlabel metal3 s 12038 10175 12038 10175 4 gnd
port 125 nsew
rlabel metal3 s 14101 9023 14101 9023 4 vdd
port 124 nsew
rlabel metal3 s 12038 14125 12038 14125 4 gnd
port 125 nsew
rlabel metal3 s 12038 15468 12038 15468 4 gnd
port 125 nsew
rlabel metal3 s 13358 9614 13358 9614 4 vdd
port 124 nsew
rlabel metal3 s 16983 9023 16983 9023 4 vdd
port 124 nsew
rlabel metal3 s 12038 15705 12038 15705 4 gnd
port 125 nsew
rlabel metal3 s 12038 13888 12038 13888 4 gnd
port 125 nsew
rlabel metal3 s 13239 9023 13239 9023 4 vdd
port 124 nsew
rlabel metal3 s 12038 10412 12038 10412 4 gnd
port 125 nsew
rlabel metal3 s 12038 15942 12038 15942 4 gnd
port 125 nsew
rlabel metal3 s 12038 14915 12038 14915 4 gnd
port 125 nsew
rlabel metal3 s 12038 11755 12038 11755 4 gnd
port 125 nsew
rlabel metal3 s 15349 9023 15349 9023 4 vdd
port 124 nsew
rlabel metal3 s 12038 10728 12038 10728 4 gnd
port 125 nsew
rlabel metal3 s 12734 9614 12734 9614 4 vdd
port 124 nsew
rlabel metal3 s 12038 16495 12038 16495 4 gnd
port 125 nsew
rlabel metal3 s 12038 10965 12038 10965 4 gnd
port 125 nsew
rlabel metal3 s 12038 11992 12038 11992 4 gnd
port 125 nsew
rlabel metal3 s 12038 14678 12038 14678 4 gnd
port 125 nsew
rlabel metal3 s 12038 15152 12038 15152 4 gnd
port 125 nsew
rlabel metal3 s 12038 12782 12038 12782 4 gnd
port 125 nsew
rlabel metal3 s 16478 9614 16478 9614 4 vdd
port 124 nsew
rlabel metal3 s 15230 9614 15230 9614 4 vdd
port 124 nsew
rlabel metal3 s 12038 16258 12038 16258 4 gnd
port 125 nsew
rlabel metal3 s 13982 9614 13982 9614 4 vdd
port 124 nsew
rlabel metal3 s 12038 11202 12038 11202 4 gnd
port 125 nsew
rlabel metal3 s 15735 9023 15735 9023 4 vdd
port 124 nsew
rlabel metal3 s 12038 9938 12038 9938 4 gnd
port 125 nsew
rlabel metal3 s 12038 13335 12038 13335 4 gnd
port 125 nsew
rlabel metal3 s 12038 13572 12038 13572 4 gnd
port 125 nsew
rlabel metal3 s 12038 13098 12038 13098 4 gnd
port 125 nsew
rlabel metal3 s 12038 16732 12038 16732 4 gnd
port 125 nsew
rlabel metal3 s 15854 9614 15854 9614 4 vdd
port 124 nsew
rlabel metal3 s 12038 12308 12038 12308 4 gnd
port 125 nsew
rlabel metal3 s 12038 14362 12038 14362 4 gnd
port 125 nsew
rlabel metal3 s 12038 12545 12038 12545 4 gnd
port 125 nsew
rlabel metal3 s 12038 11518 12038 11518 4 gnd
port 125 nsew
rlabel metal3 s 14487 9023 14487 9023 4 vdd
port 124 nsew
rlabel metal3 s 7064 15734 7064 15734 4 gnd
port 125 nsew
rlabel metal3 s 6682 14140 6682 14140 4 vdd
port 124 nsew
rlabel metal3 s 6682 14930 6682 14930 4 vdd
port 124 nsew
rlabel metal3 s 7064 13364 7064 13364 4 gnd
port 125 nsew
rlabel metal3 s 7336 13364 7336 13364 4 vdd
port 124 nsew
rlabel metal3 s 7064 14549 7064 14549 4 gnd
port 125 nsew
rlabel metal3 s 7336 14549 7336 14549 4 vdd
port 124 nsew
rlabel metal3 s 7064 12969 7064 12969 4 gnd
port 125 nsew
rlabel metal3 s 6250 16510 6250 16510 4 vdd
port 124 nsew
rlabel metal3 s 5825 12618 5825 12618 4 gnd
port 125 nsew
rlabel metal3 s 7336 13759 7336 13759 4 vdd
port 124 nsew
rlabel metal3 s 6682 16152 6682 16152 4 vdd
port 124 nsew
rlabel metal3 s 5825 16152 5825 16152 4 gnd
port 125 nsew
rlabel metal3 s 6250 14572 6250 14572 4 vdd
port 124 nsew
rlabel metal3 s 7336 14944 7336 14944 4 vdd
port 124 nsew
rlabel metal3 s 6682 15362 6682 15362 4 vdd
port 124 nsew
rlabel metal3 s 6682 16510 6682 16510 4 vdd
port 124 nsew
rlabel metal3 s 6250 15720 6250 15720 4 vdd
port 124 nsew
rlabel metal3 s 6250 14140 6250 14140 4 vdd
port 124 nsew
rlabel metal3 s 6682 15720 6682 15720 4 vdd
port 124 nsew
rlabel metal3 s 6250 13782 6250 13782 4 vdd
port 124 nsew
rlabel metal3 s 6250 13350 6250 13350 4 vdd
port 124 nsew
rlabel metal3 s 7064 13759 7064 13759 4 gnd
port 125 nsew
rlabel metal3 s 7336 12969 7336 12969 4 vdd
port 124 nsew
rlabel metal3 s 6250 15362 6250 15362 4 vdd
port 124 nsew
rlabel metal3 s 7336 15339 7336 15339 4 vdd
port 124 nsew
rlabel metal3 s 6682 13350 6682 13350 4 vdd
port 124 nsew
rlabel metal3 s 5825 15778 5825 15778 4 gnd
port 125 nsew
rlabel metal3 s 7336 16129 7336 16129 4 vdd
port 124 nsew
rlabel metal3 s 7064 16524 7064 16524 4 gnd
port 125 nsew
rlabel metal3 s 6250 12992 6250 12992 4 vdd
port 124 nsew
rlabel metal3 s 5825 13782 5825 13782 4 gnd
port 125 nsew
rlabel metal3 s 7336 16524 7336 16524 4 vdd
port 124 nsew
rlabel metal3 s 6250 16152 6250 16152 4 vdd
port 124 nsew
rlabel metal3 s 5825 12992 5825 12992 4 gnd
port 125 nsew
rlabel metal3 s 6682 12992 6682 12992 4 vdd
port 124 nsew
rlabel metal3 s 5825 13408 5825 13408 4 gnd
port 125 nsew
rlabel metal3 s 6682 13782 6682 13782 4 vdd
port 124 nsew
rlabel metal3 s 7336 14154 7336 14154 4 vdd
port 124 nsew
rlabel metal3 s 5825 14572 5825 14572 4 gnd
port 125 nsew
rlabel metal3 s 7064 14154 7064 14154 4 gnd
port 125 nsew
rlabel metal3 s 7064 15339 7064 15339 4 gnd
port 125 nsew
rlabel metal3 s 7064 14944 7064 14944 4 gnd
port 125 nsew
rlabel metal3 s 5825 15362 5825 15362 4 gnd
port 125 nsew
rlabel metal3 s 5825 14198 5825 14198 4 gnd
port 125 nsew
rlabel metal3 s 5825 16568 5825 16568 4 gnd
port 125 nsew
rlabel metal3 s 6250 14930 6250 14930 4 vdd
port 124 nsew
rlabel metal3 s 7336 15734 7336 15734 4 vdd
port 124 nsew
rlabel metal3 s 6682 14572 6682 14572 4 vdd
port 124 nsew
rlabel metal3 s 7064 16129 7064 16129 4 gnd
port 125 nsew
rlabel metal3 s 5825 14988 5825 14988 4 gnd
port 125 nsew
rlabel metal3 s 2970 12976 2970 12976 4 gnd
port 125 nsew
rlabel metal3 s 2535 15362 2535 15362 4 gnd
port 125 nsew
rlabel metal3 s 3774 15339 3774 15339 4 gnd
port 125 nsew
rlabel metal3 s 3395 13766 3395 13766 4 vdd
port 124 nsew
rlabel metal3 s 3774 13759 3774 13759 4 gnd
port 125 nsew
rlabel metal3 s 3395 12976 3395 12976 4 vdd
port 124 nsew
rlabel metal3 s 3392 15362 3392 15362 4 vdd
port 124 nsew
rlabel metal3 s 2072 12969 2072 12969 4 vdd
port 124 nsew
rlabel metal3 s 3774 16129 3774 16129 4 gnd
port 125 nsew
rlabel metal3 s 1476 15339 1476 15339 4 vdd
port 124 nsew
rlabel metal3 s 1800 12969 1800 12969 4 gnd
port 125 nsew
rlabel metal3 s 4046 13759 4046 13759 4 vdd
port 124 nsew
rlabel metal3 s 2960 16152 2960 16152 4 vdd
port 124 nsew
rlabel metal3 s 2960 15362 2960 15362 4 vdd
port 124 nsew
rlabel metal3 s 2970 13766 2970 13766 4 gnd
port 125 nsew
rlabel metal3 s 4046 16129 4046 16129 4 vdd
port 124 nsew
rlabel metal3 s 2535 16152 2535 16152 4 gnd
port 125 nsew
rlabel metal3 s 1204 15339 1204 15339 4 gnd
port 125 nsew
rlabel metal3 s 4046 12969 4046 12969 4 vdd
port 124 nsew
rlabel metal3 s 3774 12969 3774 12969 4 gnd
port 125 nsew
rlabel metal3 s 4046 15339 4046 15339 4 vdd
port 124 nsew
rlabel metal3 s 3392 16152 3392 16152 4 vdd
port 124 nsew
rlabel metal3 s 3395 11396 3395 11396 4 vdd
port 124 nsew
rlabel metal3 s 2970 11396 2970 11396 4 gnd
port 125 nsew
rlabel metal3 s 4046 11389 4046 11389 4 vdd
port 124 nsew
rlabel metal3 s 3774 11389 3774 11389 4 gnd
port 125 nsew
rlabel metal3 s 2072 10599 2072 10599 4 vdd
port 124 nsew
rlabel metal3 s 3395 10606 3395 10606 4 vdd
port 124 nsew
rlabel metal3 s 4046 10599 4046 10599 4 vdd
port 124 nsew
rlabel metal3 s 1800 10599 1800 10599 4 gnd
port 125 nsew
rlabel metal3 s 2970 10606 2970 10606 4 gnd
port 125 nsew
rlabel metal3 s 3774 10599 3774 10599 4 gnd
port 125 nsew
rlabel metal3 s 6682 11770 6682 11770 4 vdd
port 124 nsew
rlabel metal3 s 5825 12202 5825 12202 4 gnd
port 125 nsew
rlabel metal3 s 7336 12574 7336 12574 4 vdd
port 124 nsew
rlabel metal3 s 6250 12560 6250 12560 4 vdd
port 124 nsew
rlabel metal3 s 5825 11038 5825 11038 4 gnd
port 125 nsew
rlabel metal3 s 6682 11412 6682 11412 4 vdd
port 124 nsew
rlabel metal3 s 7064 11389 7064 11389 4 gnd
port 125 nsew
rlabel metal3 s 6250 10980 6250 10980 4 vdd
port 124 nsew
rlabel metal3 s 5825 10622 5825 10622 4 gnd
port 125 nsew
rlabel metal3 s 6682 10980 6682 10980 4 vdd
port 124 nsew
rlabel metal3 s 7336 11784 7336 11784 4 vdd
port 124 nsew
rlabel metal3 s 6250 10622 6250 10622 4 vdd
port 124 nsew
rlabel metal3 s 6250 12202 6250 12202 4 vdd
port 124 nsew
rlabel metal3 s 7336 12179 7336 12179 4 vdd
port 124 nsew
rlabel metal3 s 5825 11412 5825 11412 4 gnd
port 125 nsew
rlabel metal3 s 7064 10994 7064 10994 4 gnd
port 125 nsew
rlabel metal3 s 6682 12560 6682 12560 4 vdd
port 124 nsew
rlabel metal3 s 7336 10599 7336 10599 4 vdd
port 124 nsew
rlabel metal3 s 7064 12179 7064 12179 4 gnd
port 125 nsew
rlabel metal3 s 6682 12202 6682 12202 4 vdd
port 124 nsew
rlabel metal3 s 6682 10622 6682 10622 4 vdd
port 124 nsew
rlabel metal3 s 6250 11770 6250 11770 4 vdd
port 124 nsew
rlabel metal3 s 7064 11784 7064 11784 4 gnd
port 125 nsew
rlabel metal3 s 7336 10994 7336 10994 4 vdd
port 124 nsew
rlabel metal3 s 7064 10599 7064 10599 4 gnd
port 125 nsew
rlabel metal3 s 5825 11828 5825 11828 4 gnd
port 125 nsew
rlabel metal3 s 7336 11389 7336 11389 4 vdd
port 124 nsew
rlabel metal3 s 6250 11412 6250 11412 4 vdd
port 124 nsew
rlabel metal3 s 7064 12574 7064 12574 4 gnd
port 125 nsew
rlabel metal3 s 6488 6203 6488 6203 4 vdd
port 124 nsew
rlabel metal3 s 6488 7617 6488 7617 4 gnd
port 125 nsew
rlabel metal3 s 6483 8255 6483 8255 4 rbl_bl0
port 127 nsew
rlabel metal3 s 6488 4789 6488 4789 4 gnd
port 125 nsew
rlabel metal3 s 14663 4903 14663 4903 4 vdd
port 124 nsew
rlabel metal3 s 14671 2181 14671 2181 4 gnd
port 125 nsew
rlabel metal3 s 15818 1563 15818 1563 4 vdd
port 124 nsew
rlabel metal3 s 15798 2513 15798 2513 4 vdd
port 124 nsew
rlabel metal3 s 13302 2513 13302 2513 4 vdd
port 124 nsew
rlabel metal3 s 13419 1120 13419 1120 4 vdd
port 124 nsew
rlabel metal3 s 17057 2950 17057 2950 4 gnd
port 125 nsew
rlabel metal3 s 15809 2950 15809 2950 4 gnd
port 125 nsew
rlabel metal3 s 13322 1563 13322 1563 4 vdd
port 124 nsew
rlabel metal3 s 14550 2513 14550 2513 4 vdd
port 124 nsew
rlabel metal3 s 14745 5677 14745 5677 4 gnd
port 125 nsew
rlabel metal3 s 15911 4903 15911 4903 4 vdd
port 124 nsew
rlabel metal3 s 14675 4065 14675 4065 4 vdd
port 124 nsew
rlabel metal3 s 13415 4903 13415 4903 4 vdd
port 124 nsew
rlabel metal3 s 13419 0 13419 0 4 gnd
port 125 nsew
rlabel metal3 s 15923 4065 15923 4065 4 vdd
port 124 nsew
rlabel metal3 s 17046 2513 17046 2513 4 vdd
port 124 nsew
rlabel metal3 s 15919 2181 15919 2181 4 gnd
port 125 nsew
rlabel metal3 s 14918 7450 14918 7450 4 gnd
port 125 nsew
rlabel metal3 s 13670 7450 13670 7450 4 gnd
port 125 nsew
rlabel metal3 s 15804 1979 15804 1979 4 gnd
port 125 nsew
rlabel metal3 s 13313 2950 13313 2950 4 gnd
port 125 nsew
rlabel metal3 s 16166 7450 16166 7450 4 gnd
port 125 nsew
rlabel metal3 s 14570 1563 14570 1563 4 vdd
port 124 nsew
rlabel metal3 s 13308 1979 13308 1979 4 gnd
port 125 nsew
rlabel metal3 s 13427 3743 13427 3743 4 gnd
port 125 nsew
rlabel metal3 s 13427 4065 13427 4065 4 vdd
port 124 nsew
rlabel metal3 s 14561 2950 14561 2950 4 gnd
port 125 nsew
rlabel metal3 s 15923 3743 15923 3743 4 gnd
port 125 nsew
rlabel metal3 s 14675 3743 14675 3743 4 gnd
port 125 nsew
rlabel metal3 s 15993 5677 15993 5677 4 gnd
port 125 nsew
rlabel metal3 s 13497 5677 13497 5677 4 gnd
port 125 nsew
rlabel metal3 s 14556 1979 14556 1979 4 gnd
port 125 nsew
rlabel metal3 s 17066 1563 17066 1563 4 vdd
port 124 nsew
rlabel metal3 s 13423 2181 13423 2181 4 gnd
port 125 nsew
rlabel metal3 s 17052 1979 17052 1979 4 gnd
port 125 nsew
rlabel metal3 s 30325 9023 30325 9023 4 vdd
port 124 nsew
rlabel metal3 s 25719 9023 25719 9023 4 vdd
port 124 nsew
rlabel metal3 s 26967 9023 26967 9023 4 vdd
port 124 nsew
rlabel metal3 s 26581 9023 26581 9023 4 vdd
port 124 nsew
rlabel metal3 s 32078 9614 32078 9614 4 vdd
port 124 nsew
rlabel metal3 s 28958 9614 28958 9614 4 vdd
port 124 nsew
rlabel metal3 s 31959 9023 31959 9023 4 vdd
port 124 nsew
rlabel metal3 s 30830 9614 30830 9614 4 vdd
port 124 nsew
rlabel metal3 s 29582 9614 29582 9614 4 vdd
port 124 nsew
rlabel metal3 s 27086 9614 27086 9614 4 vdd
port 124 nsew
rlabel metal3 s 27710 9614 27710 9614 4 vdd
port 124 nsew
rlabel metal3 s 31454 9614 31454 9614 4 vdd
port 124 nsew
rlabel metal3 s 26462 9614 26462 9614 4 vdd
port 124 nsew
rlabel metal3 s 31573 9023 31573 9023 4 vdd
port 124 nsew
rlabel metal3 s 32702 9614 32702 9614 4 vdd
port 124 nsew
rlabel metal3 s 27829 9023 27829 9023 4 vdd
port 124 nsew
rlabel metal3 s 29463 9023 29463 9023 4 vdd
port 124 nsew
rlabel metal3 s 25214 9614 25214 9614 4 vdd
port 124 nsew
rlabel metal3 s 30711 9023 30711 9023 4 vdd
port 124 nsew
rlabel metal3 s 25333 9023 25333 9023 4 vdd
port 124 nsew
rlabel metal3 s 29077 9023 29077 9023 4 vdd
port 124 nsew
rlabel metal3 s 25838 9614 25838 9614 4 vdd
port 124 nsew
rlabel metal3 s 28215 9023 28215 9023 4 vdd
port 124 nsew
rlabel metal3 s 30206 9614 30206 9614 4 vdd
port 124 nsew
rlabel metal3 s 28334 9614 28334 9614 4 vdd
port 124 nsew
rlabel metal3 s 32821 9023 32821 9023 4 vdd
port 124 nsew
rlabel metal3 s 21975 9023 21975 9023 4 vdd
port 124 nsew
rlabel metal3 s 24471 9023 24471 9023 4 vdd
port 124 nsew
rlabel metal3 s 22094 9614 22094 9614 4 vdd
port 124 nsew
rlabel metal3 s 17726 9614 17726 9614 4 vdd
port 124 nsew
rlabel metal3 s 22837 9023 22837 9023 4 vdd
port 124 nsew
rlabel metal3 s 20727 9023 20727 9023 4 vdd
port 124 nsew
rlabel metal3 s 17845 9023 17845 9023 4 vdd
port 124 nsew
rlabel metal3 s 19598 9614 19598 9614 4 vdd
port 124 nsew
rlabel metal3 s 18974 9614 18974 9614 4 vdd
port 124 nsew
rlabel metal3 s 22718 9614 22718 9614 4 vdd
port 124 nsew
rlabel metal3 s 20846 9614 20846 9614 4 vdd
port 124 nsew
rlabel metal3 s 23342 9614 23342 9614 4 vdd
port 124 nsew
rlabel metal3 s 20222 9614 20222 9614 4 vdd
port 124 nsew
rlabel metal3 s 21589 9023 21589 9023 4 vdd
port 124 nsew
rlabel metal3 s 19093 9023 19093 9023 4 vdd
port 124 nsew
rlabel metal3 s 18350 9614 18350 9614 4 vdd
port 124 nsew
rlabel metal3 s 23223 9023 23223 9023 4 vdd
port 124 nsew
rlabel metal3 s 20341 9023 20341 9023 4 vdd
port 124 nsew
rlabel metal3 s 19479 9023 19479 9023 4 vdd
port 124 nsew
rlabel metal3 s 21470 9614 21470 9614 4 vdd
port 124 nsew
rlabel metal3 s 24085 9023 24085 9023 4 vdd
port 124 nsew
rlabel metal3 s 23966 9614 23966 9614 4 vdd
port 124 nsew
rlabel metal3 s 18231 9023 18231 9023 4 vdd
port 124 nsew
rlabel metal3 s 24590 9614 24590 9614 4 vdd
port 124 nsew
rlabel metal3 s 24729 5677 24729 5677 4 gnd
port 125 nsew
rlabel metal3 s 20810 1563 20810 1563 4 vdd
port 124 nsew
rlabel metal3 s 23654 7450 23654 7450 4 gnd
port 125 nsew
rlabel metal3 s 17414 7450 17414 7450 4 gnd
port 125 nsew
rlabel metal3 s 19667 4065 19667 4065 4 vdd
port 124 nsew
rlabel metal3 s 18489 5677 18489 5677 4 gnd
port 125 nsew
rlabel metal3 s 19737 5677 19737 5677 4 gnd
port 125 nsew
rlabel metal3 s 22151 4903 22151 4903 4 vdd
port 124 nsew
rlabel metal3 s 23292 1979 23292 1979 4 gnd
port 125 nsew
rlabel metal3 s 24902 7450 24902 7450 4 gnd
port 125 nsew
rlabel metal3 s 20915 3743 20915 3743 4 gnd
port 125 nsew
rlabel metal3 s 18419 4065 18419 4065 4 vdd
port 124 nsew
rlabel metal3 s 22049 2950 22049 2950 4 gnd
port 125 nsew
rlabel metal3 s 24554 1563 24554 1563 4 vdd
port 124 nsew
rlabel metal3 s 20790 2513 20790 2513 4 vdd
port 124 nsew
rlabel metal3 s 23411 3743 23411 3743 4 gnd
port 125 nsew
rlabel metal3 s 22058 1563 22058 1563 4 vdd
port 124 nsew
rlabel metal3 s 19553 2950 19553 2950 4 gnd
port 125 nsew
rlabel metal3 s 20796 1979 20796 1979 4 gnd
port 125 nsew
rlabel metal3 s 24655 2181 24655 2181 4 gnd
port 125 nsew
rlabel metal3 s 17167 2181 17167 2181 4 gnd
port 125 nsew
rlabel metal3 s 20985 5677 20985 5677 4 gnd
port 125 nsew
rlabel metal3 s 23399 4903 23399 4903 4 vdd
port 124 nsew
rlabel metal3 s 23411 4065 23411 4065 4 vdd
port 124 nsew
rlabel metal3 s 18407 4903 18407 4903 4 vdd
port 124 nsew
rlabel metal3 s 23407 2181 23407 2181 4 gnd
port 125 nsew
rlabel metal3 s 23297 2950 23297 2950 4 gnd
port 125 nsew
rlabel metal3 s 17241 5677 17241 5677 4 gnd
port 125 nsew
rlabel metal3 s 24540 1979 24540 1979 4 gnd
port 125 nsew
rlabel metal3 s 24659 3743 24659 3743 4 gnd
port 125 nsew
rlabel metal3 s 18314 1563 18314 1563 4 vdd
port 124 nsew
rlabel metal3 s 18419 3743 18419 3743 4 gnd
port 125 nsew
rlabel metal3 s 19655 4903 19655 4903 4 vdd
port 124 nsew
rlabel metal3 s 17171 4065 17171 4065 4 vdd
port 124 nsew
rlabel metal3 s 23286 2513 23286 2513 4 vdd
port 124 nsew
rlabel metal3 s 20903 4903 20903 4903 4 vdd
port 124 nsew
rlabel metal3 s 20911 2181 20911 2181 4 gnd
port 125 nsew
rlabel metal3 s 22233 5677 22233 5677 4 gnd
port 125 nsew
rlabel metal3 s 23403 0 23403 0 4 gnd
port 125 nsew
rlabel metal3 s 22044 1979 22044 1979 4 gnd
port 125 nsew
rlabel metal3 s 18415 2181 18415 2181 4 gnd
port 125 nsew
rlabel metal3 s 18662 7450 18662 7450 4 gnd
port 125 nsew
rlabel metal3 s 24534 2513 24534 2513 4 vdd
port 124 nsew
rlabel metal3 s 22163 4065 22163 4065 4 vdd
port 124 nsew
rlabel metal3 s 20915 4065 20915 4065 4 vdd
port 124 nsew
rlabel metal3 s 24545 2950 24545 2950 4 gnd
port 125 nsew
rlabel metal3 s 17159 4903 17159 4903 4 vdd
port 124 nsew
rlabel metal3 s 21158 7450 21158 7450 4 gnd
port 125 nsew
rlabel metal3 s 20801 2950 20801 2950 4 gnd
port 125 nsew
rlabel metal3 s 22159 2181 22159 2181 4 gnd
port 125 nsew
rlabel metal3 s 19667 3743 19667 3743 4 gnd
port 125 nsew
rlabel metal3 s 19663 2181 19663 2181 4 gnd
port 125 nsew
rlabel metal3 s 23481 5677 23481 5677 4 gnd
port 125 nsew
rlabel metal3 s 19548 1979 19548 1979 4 gnd
port 125 nsew
rlabel metal3 s 22038 2513 22038 2513 4 vdd
port 124 nsew
rlabel metal3 s 22163 3743 22163 3743 4 gnd
port 125 nsew
rlabel metal3 s 23306 1563 23306 1563 4 vdd
port 124 nsew
rlabel metal3 s 17171 3743 17171 3743 4 gnd
port 125 nsew
rlabel metal3 s 24659 4065 24659 4065 4 vdd
port 124 nsew
rlabel metal3 s 19542 2513 19542 2513 4 vdd
port 124 nsew
rlabel metal3 s 19562 1563 19562 1563 4 vdd
port 124 nsew
rlabel metal3 s 18294 2513 18294 2513 4 vdd
port 124 nsew
rlabel metal3 s 18300 1979 18300 1979 4 gnd
port 125 nsew
rlabel metal3 s 19910 7450 19910 7450 4 gnd
port 125 nsew
rlabel metal3 s 22406 7450 22406 7450 4 gnd
port 125 nsew
rlabel metal3 s 24647 4903 24647 4903 4 vdd
port 124 nsew
rlabel metal3 s 18305 2950 18305 2950 4 gnd
port 125 nsew
rlabel metal3 s 23403 1120 23403 1120 4 vdd
port 124 nsew
rlabel metal3 s 27030 2513 27030 2513 4 vdd
port 124 nsew
rlabel metal3 s 29651 3743 29651 3743 4 gnd
port 125 nsew
rlabel metal3 s 30969 5677 30969 5677 4 gnd
port 125 nsew
rlabel metal3 s 29721 5677 29721 5677 4 gnd
port 125 nsew
rlabel metal3 s 25793 2950 25793 2950 4 gnd
port 125 nsew
rlabel metal3 s 28646 7450 28646 7450 4 gnd
port 125 nsew
rlabel metal3 s 32147 4065 32147 4065 4 vdd
port 124 nsew
rlabel metal3 s 32143 2181 32143 2181 4 gnd
port 125 nsew
rlabel metal3 s 32135 4903 32135 4903 4 vdd
port 124 nsew
rlabel metal3 s 30774 2513 30774 2513 4 vdd
port 124 nsew
rlabel metal3 s 29532 1979 29532 1979 4 gnd
port 125 nsew
rlabel metal3 s 28403 4065 28403 4065 4 vdd
port 124 nsew
rlabel metal3 s 28391 4903 28391 4903 4 vdd
port 124 nsew
rlabel metal3 s 30780 1979 30780 1979 4 gnd
port 125 nsew
rlabel metal3 s 31142 7450 31142 7450 4 gnd
port 125 nsew
rlabel metal3 s 28473 5677 28473 5677 4 gnd
port 125 nsew
rlabel metal3 s 27143 4903 27143 4903 4 vdd
port 124 nsew
rlabel metal3 s 27041 2950 27041 2950 4 gnd
port 125 nsew
rlabel metal3 s 30899 3743 30899 3743 4 gnd
port 125 nsew
rlabel metal3 s 28298 1563 28298 1563 4 vdd
port 124 nsew
rlabel metal3 s 27036 1979 27036 1979 4 gnd
port 125 nsew
rlabel metal3 s 27398 7450 27398 7450 4 gnd
port 125 nsew
rlabel metal3 s 32147 3743 32147 3743 4 gnd
port 125 nsew
rlabel metal3 s 30895 2181 30895 2181 4 gnd
port 125 nsew
rlabel metal3 s 30785 2950 30785 2950 4 gnd
port 125 nsew
rlabel metal3 s 27155 4065 27155 4065 4 vdd
port 124 nsew
rlabel metal3 s 28403 3743 28403 3743 4 gnd
port 125 nsew
rlabel metal3 s 32217 5677 32217 5677 4 gnd
port 125 nsew
rlabel metal3 s 28399 2181 28399 2181 4 gnd
port 125 nsew
rlabel metal3 s 32042 1563 32042 1563 4 vdd
port 124 nsew
rlabel metal3 s 30794 1563 30794 1563 4 vdd
port 124 nsew
rlabel metal3 s 25895 4903 25895 4903 4 vdd
port 124 nsew
rlabel metal3 s 30899 4065 30899 4065 4 vdd
port 124 nsew
rlabel metal3 s 25977 5677 25977 5677 4 gnd
port 125 nsew
rlabel metal3 s 25907 3743 25907 3743 4 gnd
port 125 nsew
rlabel metal3 s 27050 1563 27050 1563 4 vdd
port 124 nsew
rlabel metal3 s 25907 4065 25907 4065 4 vdd
port 124 nsew
rlabel metal3 s 28284 1979 28284 1979 4 gnd
port 125 nsew
rlabel metal3 s 32022 2513 32022 2513 4 vdd
port 124 nsew
rlabel metal3 s 29639 4903 29639 4903 4 vdd
port 124 nsew
rlabel metal3 s 27151 2181 27151 2181 4 gnd
port 125 nsew
rlabel metal3 s 29546 1563 29546 1563 4 vdd
port 124 nsew
rlabel metal3 s 32028 1979 32028 1979 4 gnd
port 125 nsew
rlabel metal3 s 25782 2513 25782 2513 4 vdd
port 124 nsew
rlabel metal3 s 29651 4065 29651 4065 4 vdd
port 124 nsew
rlabel metal3 s 25802 1563 25802 1563 4 vdd
port 124 nsew
rlabel metal3 s 25788 1979 25788 1979 4 gnd
port 125 nsew
rlabel metal3 s 29647 2181 29647 2181 4 gnd
port 125 nsew
rlabel metal3 s 29526 2513 29526 2513 4 vdd
port 124 nsew
rlabel metal3 s 29537 2950 29537 2950 4 gnd
port 125 nsew
rlabel metal3 s 25903 2181 25903 2181 4 gnd
port 125 nsew
rlabel metal3 s 29894 7450 29894 7450 4 gnd
port 125 nsew
rlabel metal3 s 27155 3743 27155 3743 4 gnd
port 125 nsew
rlabel metal3 s 30887 4903 30887 4903 4 vdd
port 124 nsew
rlabel metal3 s 28289 2950 28289 2950 4 gnd
port 125 nsew
rlabel metal3 s 27225 5677 27225 5677 4 gnd
port 125 nsew
rlabel metal3 s 26150 7450 26150 7450 4 gnd
port 125 nsew
rlabel metal3 s 32033 2950 32033 2950 4 gnd
port 125 nsew
rlabel metal3 s 28278 2513 28278 2513 4 vdd
port 124 nsew
rlabel metal3 s 32390 7450 32390 7450 4 gnd
port 125 nsew
rlabel metal3 s 58692 31534 58692 31534 4 vdd
port 124 nsew
rlabel metal3 s 59346 32742 59346 32742 4 vdd
port 124 nsew
rlabel metal3 s 59346 31520 59346 31520 4 vdd
port 124 nsew
rlabel metal3 s 58692 31929 58692 31929 4 vdd
port 124 nsew
rlabel metal3 s 59778 31952 59778 31952 4 vdd
port 124 nsew
rlabel metal3 s 58692 29559 58692 29559 4 vdd
port 124 nsew
rlabel metal3 s 59778 33532 59778 33532 4 vdd
port 124 nsew
rlabel metal3 s 60203 33532 60203 33532 4 gnd
port 125 nsew
rlabel metal3 s 59778 32310 59778 32310 4 vdd
port 124 nsew
rlabel metal3 s 59346 30730 59346 30730 4 vdd
port 124 nsew
rlabel metal3 s 58964 30744 58964 30744 4 gnd
port 125 nsew
rlabel metal3 s 60203 31578 60203 31578 4 gnd
port 125 nsew
rlabel metal3 s 58692 29954 58692 29954 4 vdd
port 124 nsew
rlabel metal3 s 58964 30349 58964 30349 4 gnd
port 125 nsew
rlabel metal3 s 59778 29940 59778 29940 4 vdd
port 124 nsew
rlabel metal3 s 58692 30349 58692 30349 4 vdd
port 124 nsew
rlabel metal3 s 58964 32324 58964 32324 4 gnd
port 125 nsew
rlabel metal3 s 58692 30744 58692 30744 4 vdd
port 124 nsew
rlabel metal3 s 60203 32742 60203 32742 4 gnd
port 125 nsew
rlabel metal3 s 58692 33509 58692 33509 4 vdd
port 124 nsew
rlabel metal3 s 59778 31520 59778 31520 4 vdd
port 124 nsew
rlabel metal3 s 59346 33100 59346 33100 4 vdd
port 124 nsew
rlabel metal3 s 59346 32310 59346 32310 4 vdd
port 124 nsew
rlabel metal3 s 58964 33114 58964 33114 4 gnd
port 125 nsew
rlabel metal3 s 59778 33100 59778 33100 4 vdd
port 124 nsew
rlabel metal3 s 60203 31952 60203 31952 4 gnd
port 125 nsew
rlabel metal3 s 60203 33158 60203 33158 4 gnd
port 125 nsew
rlabel metal3 s 58964 31534 58964 31534 4 gnd
port 125 nsew
rlabel metal3 s 58692 33114 58692 33114 4 vdd
port 124 nsew
rlabel metal3 s 59346 31162 59346 31162 4 vdd
port 124 nsew
rlabel metal3 s 58964 29559 58964 29559 4 gnd
port 125 nsew
rlabel metal3 s 58964 33509 58964 33509 4 gnd
port 125 nsew
rlabel metal3 s 58964 31929 58964 31929 4 gnd
port 125 nsew
rlabel metal3 s 58964 31139 58964 31139 4 gnd
port 125 nsew
rlabel metal3 s 59778 30730 59778 30730 4 vdd
port 124 nsew
rlabel metal3 s 59346 33532 59346 33532 4 vdd
port 124 nsew
rlabel metal3 s 60203 31162 60203 31162 4 gnd
port 125 nsew
rlabel metal3 s 60203 29998 60203 29998 4 gnd
port 125 nsew
rlabel metal3 s 60203 32368 60203 32368 4 gnd
port 125 nsew
rlabel metal3 s 60203 30372 60203 30372 4 gnd
port 125 nsew
rlabel metal3 s 59778 31162 59778 31162 4 vdd
port 124 nsew
rlabel metal3 s 58692 32719 58692 32719 4 vdd
port 124 nsew
rlabel metal3 s 59778 30372 59778 30372 4 vdd
port 124 nsew
rlabel metal3 s 58964 32719 58964 32719 4 gnd
port 125 nsew
rlabel metal3 s 60203 30788 60203 30788 4 gnd
port 125 nsew
rlabel metal3 s 59346 30372 59346 30372 4 vdd
port 124 nsew
rlabel metal3 s 59346 29582 59346 29582 4 vdd
port 124 nsew
rlabel metal3 s 58692 32324 58692 32324 4 vdd
port 124 nsew
rlabel metal3 s 59778 29582 59778 29582 4 vdd
port 124 nsew
rlabel metal3 s 59346 29940 59346 29940 4 vdd
port 124 nsew
rlabel metal3 s 58964 29954 58964 29954 4 gnd
port 125 nsew
rlabel metal3 s 58692 31139 58692 31139 4 vdd
port 124 nsew
rlabel metal3 s 59778 32742 59778 32742 4 vdd
port 124 nsew
rlabel metal3 s 60203 29582 60203 29582 4 gnd
port 125 nsew
rlabel metal3 s 59346 31952 59346 31952 4 vdd
port 124 nsew
rlabel metal3 s 59778 28360 59778 28360 4 vdd
port 124 nsew
rlabel metal3 s 60203 26048 60203 26048 4 gnd
port 125 nsew
rlabel metal3 s 59778 27570 59778 27570 4 vdd
port 124 nsew
rlabel metal3 s 60203 29208 60203 29208 4 gnd
port 125 nsew
rlabel metal3 s 59346 29150 59346 29150 4 vdd
port 124 nsew
rlabel metal3 s 60203 28792 60203 28792 4 gnd
port 125 nsew
rlabel metal3 s 58964 29164 58964 29164 4 gnd
port 125 nsew
rlabel metal3 s 59346 25200 59346 25200 4 vdd
port 124 nsew
rlabel metal3 s 59778 25990 59778 25990 4 vdd
port 124 nsew
rlabel metal3 s 58964 26399 58964 26399 4 gnd
port 125 nsew
rlabel metal3 s 59778 26780 59778 26780 4 vdd
port 124 nsew
rlabel metal3 s 59778 27212 59778 27212 4 vdd
port 124 nsew
rlabel metal3 s 60203 25632 60203 25632 4 gnd
port 125 nsew
rlabel metal3 s 58964 25214 58964 25214 4 gnd
port 125 nsew
rlabel metal3 s 59346 28360 59346 28360 4 vdd
port 124 nsew
rlabel metal3 s 60203 27212 60203 27212 4 gnd
port 125 nsew
rlabel metal3 s 60203 26838 60203 26838 4 gnd
port 125 nsew
rlabel metal3 s 60203 25258 60203 25258 4 gnd
port 125 nsew
rlabel metal3 s 60203 28002 60203 28002 4 gnd
port 125 nsew
rlabel metal3 s 58692 26399 58692 26399 4 vdd
port 124 nsew
rlabel metal3 s 59346 28792 59346 28792 4 vdd
port 124 nsew
rlabel metal3 s 58964 27584 58964 27584 4 gnd
port 125 nsew
rlabel metal3 s 58692 26004 58692 26004 4 vdd
port 124 nsew
rlabel metal3 s 58964 28374 58964 28374 4 gnd
port 125 nsew
rlabel metal3 s 58692 26794 58692 26794 4 vdd
port 124 nsew
rlabel metal3 s 58692 27584 58692 27584 4 vdd
port 124 nsew
rlabel metal3 s 58692 27979 58692 27979 4 vdd
port 124 nsew
rlabel metal3 s 58964 28769 58964 28769 4 gnd
port 125 nsew
rlabel metal3 s 58964 26004 58964 26004 4 gnd
port 125 nsew
rlabel metal3 s 58692 28374 58692 28374 4 vdd
port 124 nsew
rlabel metal3 s 59778 25200 59778 25200 4 vdd
port 124 nsew
rlabel metal3 s 58692 25609 58692 25609 4 vdd
port 124 nsew
rlabel metal3 s 60203 28418 60203 28418 4 gnd
port 125 nsew
rlabel metal3 s 59346 26422 59346 26422 4 vdd
port 124 nsew
rlabel metal3 s 58692 27189 58692 27189 4 vdd
port 124 nsew
rlabel metal3 s 59346 25632 59346 25632 4 vdd
port 124 nsew
rlabel metal3 s 59346 26780 59346 26780 4 vdd
port 124 nsew
rlabel metal3 s 59778 28002 59778 28002 4 vdd
port 124 nsew
rlabel metal3 s 58692 29164 58692 29164 4 vdd
port 124 nsew
rlabel metal3 s 58964 25609 58964 25609 4 gnd
port 125 nsew
rlabel metal3 s 59778 28792 59778 28792 4 vdd
port 124 nsew
rlabel metal3 s 59778 26422 59778 26422 4 vdd
port 124 nsew
rlabel metal3 s 59346 28002 59346 28002 4 vdd
port 124 nsew
rlabel metal3 s 58692 28769 58692 28769 4 vdd
port 124 nsew
rlabel metal3 s 58964 27979 58964 27979 4 gnd
port 125 nsew
rlabel metal3 s 59346 27212 59346 27212 4 vdd
port 124 nsew
rlabel metal3 s 60203 26422 60203 26422 4 gnd
port 125 nsew
rlabel metal3 s 60203 27628 60203 27628 4 gnd
port 125 nsew
rlabel metal3 s 58692 25214 58692 25214 4 vdd
port 124 nsew
rlabel metal3 s 58964 26794 58964 26794 4 gnd
port 125 nsew
rlabel metal3 s 58964 27189 58964 27189 4 gnd
port 125 nsew
rlabel metal3 s 59346 27570 59346 27570 4 vdd
port 124 nsew
rlabel metal3 s 59346 25990 59346 25990 4 vdd
port 124 nsew
rlabel metal3 s 59778 29150 59778 29150 4 vdd
port 124 nsew
rlabel metal3 s 59778 25632 59778 25632 4 vdd
port 124 nsew
rlabel metal3 s 53990 25975 53990 25975 4 gnd
port 125 nsew
rlabel metal3 s 53990 28345 53990 28345 4 gnd
port 125 nsew
rlabel metal3 s 53990 27318 53990 27318 4 gnd
port 125 nsew
rlabel metal3 s 53990 28582 53990 28582 4 gnd
port 125 nsew
rlabel metal3 s 53990 31268 53990 31268 4 gnd
port 125 nsew
rlabel metal3 s 53990 32848 53990 32848 4 gnd
port 125 nsew
rlabel metal3 s 53990 29135 53990 29135 4 gnd
port 125 nsew
rlabel metal3 s 53990 30715 53990 30715 4 gnd
port 125 nsew
rlabel metal3 s 53990 32295 53990 32295 4 gnd
port 125 nsew
rlabel metal3 s 53990 27002 53990 27002 4 gnd
port 125 nsew
rlabel metal3 s 53990 26212 53990 26212 4 gnd
port 125 nsew
rlabel metal3 s 53990 30478 53990 30478 4 gnd
port 125 nsew
rlabel metal3 s 53990 33085 53990 33085 4 gnd
port 125 nsew
rlabel metal3 s 53990 33322 53990 33322 4 gnd
port 125 nsew
rlabel metal3 s 53990 29925 53990 29925 4 gnd
port 125 nsew
rlabel metal3 s 53990 27555 53990 27555 4 gnd
port 125 nsew
rlabel metal3 s 53990 32058 53990 32058 4 gnd
port 125 nsew
rlabel metal3 s 53990 25422 53990 25422 4 gnd
port 125 nsew
rlabel metal3 s 53990 27792 53990 27792 4 gnd
port 125 nsew
rlabel metal3 s 53990 31742 53990 31742 4 gnd
port 125 nsew
rlabel metal3 s 53990 25738 53990 25738 4 gnd
port 125 nsew
rlabel metal3 s 53990 32532 53990 32532 4 gnd
port 125 nsew
rlabel metal3 s 53990 30952 53990 30952 4 gnd
port 125 nsew
rlabel metal3 s 53990 29372 53990 29372 4 gnd
port 125 nsew
rlabel metal3 s 53990 26765 53990 26765 4 gnd
port 125 nsew
rlabel metal3 s 53990 28108 53990 28108 4 gnd
port 125 nsew
rlabel metal3 s 53990 30162 53990 30162 4 gnd
port 125 nsew
rlabel metal3 s 53990 26528 53990 26528 4 gnd
port 125 nsew
rlabel metal3 s 53990 28898 53990 28898 4 gnd
port 125 nsew
rlabel metal3 s 53990 31505 53990 31505 4 gnd
port 125 nsew
rlabel metal3 s 53990 29688 53990 29688 4 gnd
port 125 nsew
rlabel metal3 s 53990 22025 53990 22025 4 gnd
port 125 nsew
rlabel metal3 s 53990 21235 53990 21235 4 gnd
port 125 nsew
rlabel metal3 s 53990 20208 53990 20208 4 gnd
port 125 nsew
rlabel metal3 s 53990 22578 53990 22578 4 gnd
port 125 nsew
rlabel metal3 s 53990 23052 53990 23052 4 gnd
port 125 nsew
rlabel metal3 s 53990 20682 53990 20682 4 gnd
port 125 nsew
rlabel metal3 s 53990 17522 53990 17522 4 gnd
port 125 nsew
rlabel metal3 s 53990 22815 53990 22815 4 gnd
port 125 nsew
rlabel metal3 s 53990 20998 53990 20998 4 gnd
port 125 nsew
rlabel metal3 s 53990 23368 53990 23368 4 gnd
port 125 nsew
rlabel metal3 s 53990 19655 53990 19655 4 gnd
port 125 nsew
rlabel metal3 s 53990 25185 53990 25185 4 gnd
port 125 nsew
rlabel metal3 s 53990 21472 53990 21472 4 gnd
port 125 nsew
rlabel metal3 s 53990 19102 53990 19102 4 gnd
port 125 nsew
rlabel metal3 s 53990 19892 53990 19892 4 gnd
port 125 nsew
rlabel metal3 s 53990 20445 53990 20445 4 gnd
port 125 nsew
rlabel metal3 s 53990 17048 53990 17048 4 gnd
port 125 nsew
rlabel metal3 s 53990 21788 53990 21788 4 gnd
port 125 nsew
rlabel metal3 s 53990 17838 53990 17838 4 gnd
port 125 nsew
rlabel metal3 s 53990 18628 53990 18628 4 gnd
port 125 nsew
rlabel metal3 s 53990 24158 53990 24158 4 gnd
port 125 nsew
rlabel metal3 s 53990 24632 53990 24632 4 gnd
port 125 nsew
rlabel metal3 s 53990 24948 53990 24948 4 gnd
port 125 nsew
rlabel metal3 s 53990 23605 53990 23605 4 gnd
port 125 nsew
rlabel metal3 s 53990 17285 53990 17285 4 gnd
port 125 nsew
rlabel metal3 s 53990 18075 53990 18075 4 gnd
port 125 nsew
rlabel metal3 s 53990 24395 53990 24395 4 gnd
port 125 nsew
rlabel metal3 s 53990 22262 53990 22262 4 gnd
port 125 nsew
rlabel metal3 s 53990 23842 53990 23842 4 gnd
port 125 nsew
rlabel metal3 s 53990 18865 53990 18865 4 gnd
port 125 nsew
rlabel metal3 s 53990 19418 53990 19418 4 gnd
port 125 nsew
rlabel metal3 s 53990 18312 53990 18312 4 gnd
port 125 nsew
rlabel metal3 s 59778 21682 59778 21682 4 vdd
port 124 nsew
rlabel metal3 s 60203 24052 60203 24052 4 gnd
port 125 nsew
rlabel metal3 s 58964 23634 58964 23634 4 gnd
port 125 nsew
rlabel metal3 s 59778 22040 59778 22040 4 vdd
port 124 nsew
rlabel metal3 s 58692 24029 58692 24029 4 vdd
port 124 nsew
rlabel metal3 s 59778 23620 59778 23620 4 vdd
port 124 nsew
rlabel metal3 s 59778 21250 59778 21250 4 vdd
port 124 nsew
rlabel metal3 s 58964 22054 58964 22054 4 gnd
port 125 nsew
rlabel metal3 s 60203 22472 60203 22472 4 gnd
port 125 nsew
rlabel metal3 s 58692 21264 58692 21264 4 vdd
port 124 nsew
rlabel metal3 s 58692 22054 58692 22054 4 vdd
port 124 nsew
rlabel metal3 s 59778 22472 59778 22472 4 vdd
port 124 nsew
rlabel metal3 s 58964 24029 58964 24029 4 gnd
port 125 nsew
rlabel metal3 s 58692 21659 58692 21659 4 vdd
port 124 nsew
rlabel metal3 s 59346 22040 59346 22040 4 vdd
port 124 nsew
rlabel metal3 s 60203 22098 60203 22098 4 gnd
port 125 nsew
rlabel metal3 s 58692 23239 58692 23239 4 vdd
port 124 nsew
rlabel metal3 s 59778 24052 59778 24052 4 vdd
port 124 nsew
rlabel metal3 s 59778 24410 59778 24410 4 vdd
port 124 nsew
rlabel metal3 s 59346 24410 59346 24410 4 vdd
port 124 nsew
rlabel metal3 s 58964 23239 58964 23239 4 gnd
port 125 nsew
rlabel metal3 s 60203 23262 60203 23262 4 gnd
port 125 nsew
rlabel metal3 s 59346 24842 59346 24842 4 vdd
port 124 nsew
rlabel metal3 s 59346 23620 59346 23620 4 vdd
port 124 nsew
rlabel metal3 s 60203 24468 60203 24468 4 gnd
port 125 nsew
rlabel metal3 s 59346 24052 59346 24052 4 vdd
port 124 nsew
rlabel metal3 s 58692 22449 58692 22449 4 vdd
port 124 nsew
rlabel metal3 s 58964 21264 58964 21264 4 gnd
port 125 nsew
rlabel metal3 s 59346 23262 59346 23262 4 vdd
port 124 nsew
rlabel metal3 s 60203 24842 60203 24842 4 gnd
port 125 nsew
rlabel metal3 s 60203 22888 60203 22888 4 gnd
port 125 nsew
rlabel metal3 s 59346 21682 59346 21682 4 vdd
port 124 nsew
rlabel metal3 s 59346 22472 59346 22472 4 vdd
port 124 nsew
rlabel metal3 s 58964 21659 58964 21659 4 gnd
port 125 nsew
rlabel metal3 s 59778 22830 59778 22830 4 vdd
port 124 nsew
rlabel metal3 s 59778 24842 59778 24842 4 vdd
port 124 nsew
rlabel metal3 s 58692 24819 58692 24819 4 vdd
port 124 nsew
rlabel metal3 s 58692 24424 58692 24424 4 vdd
port 124 nsew
rlabel metal3 s 60203 21308 60203 21308 4 gnd
port 125 nsew
rlabel metal3 s 59778 23262 59778 23262 4 vdd
port 124 nsew
rlabel metal3 s 59346 21250 59346 21250 4 vdd
port 124 nsew
rlabel metal3 s 58964 24819 58964 24819 4 gnd
port 125 nsew
rlabel metal3 s 58692 23634 58692 23634 4 vdd
port 124 nsew
rlabel metal3 s 58964 22449 58964 22449 4 gnd
port 125 nsew
rlabel metal3 s 59346 22830 59346 22830 4 vdd
port 124 nsew
rlabel metal3 s 58964 22844 58964 22844 4 gnd
port 125 nsew
rlabel metal3 s 58964 24424 58964 24424 4 gnd
port 125 nsew
rlabel metal3 s 58692 22844 58692 22844 4 vdd
port 124 nsew
rlabel metal3 s 60203 21682 60203 21682 4 gnd
port 125 nsew
rlabel metal3 s 60203 23678 60203 23678 4 gnd
port 125 nsew
rlabel metal3 s 59346 18522 59346 18522 4 vdd
port 124 nsew
rlabel metal3 s 58964 16919 58964 16919 4 gnd
port 125 nsew
rlabel metal3 s 58964 19289 58964 19289 4 gnd
port 125 nsew
rlabel metal3 s 58692 20079 58692 20079 4 vdd
port 124 nsew
rlabel metal3 s 59778 20460 59778 20460 4 vdd
port 124 nsew
rlabel metal3 s 60203 17358 60203 17358 4 gnd
port 125 nsew
rlabel metal3 s 59778 17732 59778 17732 4 vdd
port 124 nsew
rlabel metal3 s 58964 17314 58964 17314 4 gnd
port 125 nsew
rlabel metal3 s 60203 18522 60203 18522 4 gnd
port 125 nsew
rlabel metal3 s 60203 19312 60203 19312 4 gnd
port 125 nsew
rlabel metal3 s 59346 19312 59346 19312 4 vdd
port 124 nsew
rlabel metal3 s 58964 18499 58964 18499 4 gnd
port 125 nsew
rlabel metal3 s 59778 19312 59778 19312 4 vdd
port 124 nsew
rlabel metal3 s 59346 18090 59346 18090 4 vdd
port 124 nsew
rlabel metal3 s 59346 16942 59346 16942 4 vdd
port 124 nsew
rlabel metal3 s 58964 19684 58964 19684 4 gnd
port 125 nsew
rlabel metal3 s 58964 18894 58964 18894 4 gnd
port 125 nsew
rlabel metal3 s 58964 20869 58964 20869 4 gnd
port 125 nsew
rlabel metal3 s 60203 20518 60203 20518 4 gnd
port 125 nsew
rlabel metal3 s 58964 20474 58964 20474 4 gnd
port 125 nsew
rlabel metal3 s 59346 19670 59346 19670 4 vdd
port 124 nsew
rlabel metal3 s 60203 16942 60203 16942 4 gnd
port 125 nsew
rlabel metal3 s 58964 17709 58964 17709 4 gnd
port 125 nsew
rlabel metal3 s 60203 17732 60203 17732 4 gnd
port 125 nsew
rlabel metal3 s 58692 17709 58692 17709 4 vdd
port 124 nsew
rlabel metal3 s 59778 17300 59778 17300 4 vdd
port 124 nsew
rlabel metal3 s 58692 19289 58692 19289 4 vdd
port 124 nsew
rlabel metal3 s 59778 20102 59778 20102 4 vdd
port 124 nsew
rlabel metal3 s 59778 18090 59778 18090 4 vdd
port 124 nsew
rlabel metal3 s 58692 18104 58692 18104 4 vdd
port 124 nsew
rlabel metal3 s 58692 20474 58692 20474 4 vdd
port 124 nsew
rlabel metal3 s 60203 20102 60203 20102 4 gnd
port 125 nsew
rlabel metal3 s 59346 20892 59346 20892 4 vdd
port 124 nsew
rlabel metal3 s 60203 18148 60203 18148 4 gnd
port 125 nsew
rlabel metal3 s 58692 18499 58692 18499 4 vdd
port 124 nsew
rlabel metal3 s 58964 20079 58964 20079 4 gnd
port 125 nsew
rlabel metal3 s 59346 17732 59346 17732 4 vdd
port 124 nsew
rlabel metal3 s 59778 18522 59778 18522 4 vdd
port 124 nsew
rlabel metal3 s 60203 18938 60203 18938 4 gnd
port 125 nsew
rlabel metal3 s 58692 19684 58692 19684 4 vdd
port 124 nsew
rlabel metal3 s 58692 18894 58692 18894 4 vdd
port 124 nsew
rlabel metal3 s 60203 19728 60203 19728 4 gnd
port 125 nsew
rlabel metal3 s 59346 18880 59346 18880 4 vdd
port 124 nsew
rlabel metal3 s 58692 17314 58692 17314 4 vdd
port 124 nsew
rlabel metal3 s 58964 18104 58964 18104 4 gnd
port 125 nsew
rlabel metal3 s 59778 18880 59778 18880 4 vdd
port 124 nsew
rlabel metal3 s 59346 20102 59346 20102 4 vdd
port 124 nsew
rlabel metal3 s 58692 20869 58692 20869 4 vdd
port 124 nsew
rlabel metal3 s 59778 19670 59778 19670 4 vdd
port 124 nsew
rlabel metal3 s 59778 20892 59778 20892 4 vdd
port 124 nsew
rlabel metal3 s 59778 16942 59778 16942 4 vdd
port 124 nsew
rlabel metal3 s 60203 20892 60203 20892 4 gnd
port 125 nsew
rlabel metal3 s 59346 17300 59346 17300 4 vdd
port 124 nsew
rlabel metal3 s 59346 20460 59346 20460 4 vdd
port 124 nsew
rlabel metal3 s 58692 16919 58692 16919 4 vdd
port 124 nsew
rlabel metal3 s 61982 16919 61982 16919 4 vdd
port 124 nsew
rlabel metal3 s 61982 17709 61982 17709 4 vdd
port 124 nsew
rlabel metal3 s 62254 17709 62254 17709 4 gnd
port 125 nsew
rlabel metal3 s 62636 16942 62636 16942 4 vdd
port 124 nsew
rlabel metal3 s 62636 17732 62636 17732 4 vdd
port 124 nsew
rlabel metal3 s 62254 16919 62254 16919 4 gnd
port 125 nsew
rlabel metal3 s 63068 16942 63068 16942 4 vdd
port 124 nsew
rlabel metal3 s 63493 16942 63493 16942 4 gnd
port 125 nsew
rlabel metal3 s 63068 17732 63068 17732 4 vdd
port 124 nsew
rlabel metal3 s 63493 17732 63493 17732 4 gnd
port 125 nsew
rlabel metal3 s 45301 9023 45301 9023 4 vdd
port 124 nsew
rlabel metal3 s 43191 9023 43191 9023 4 vdd
port 124 nsew
rlabel metal3 s 44439 9023 44439 9023 4 vdd
port 124 nsew
rlabel metal3 s 44053 9023 44053 9023 4 vdd
port 124 nsew
rlabel metal3 s 43934 9614 43934 9614 4 vdd
port 124 nsew
rlabel metal3 s 48183 9023 48183 9023 4 vdd
port 124 nsew
rlabel metal3 s 48302 9614 48302 9614 4 vdd
port 124 nsew
rlabel metal3 s 41438 9614 41438 9614 4 vdd
port 124 nsew
rlabel metal3 s 47797 9023 47797 9023 4 vdd
port 124 nsew
rlabel metal3 s 42686 9614 42686 9614 4 vdd
port 124 nsew
rlabel metal3 s 46430 9614 46430 9614 4 vdd
port 124 nsew
rlabel metal3 s 41943 9023 41943 9023 4 vdd
port 124 nsew
rlabel metal3 s 45182 9614 45182 9614 4 vdd
port 124 nsew
rlabel metal3 s 42805 9023 42805 9023 4 vdd
port 124 nsew
rlabel metal3 s 44558 9614 44558 9614 4 vdd
port 124 nsew
rlabel metal3 s 46935 9023 46935 9023 4 vdd
port 124 nsew
rlabel metal3 s 47054 9614 47054 9614 4 vdd
port 124 nsew
rlabel metal3 s 45687 9023 45687 9023 4 vdd
port 124 nsew
rlabel metal3 s 47678 9614 47678 9614 4 vdd
port 124 nsew
rlabel metal3 s 41557 9023 41557 9023 4 vdd
port 124 nsew
rlabel metal3 s 42062 9614 42062 9614 4 vdd
port 124 nsew
rlabel metal3 s 45806 9614 45806 9614 4 vdd
port 124 nsew
rlabel metal3 s 46549 9023 46549 9023 4 vdd
port 124 nsew
rlabel metal3 s 43310 9614 43310 9614 4 vdd
port 124 nsew
rlabel metal3 s 37694 9614 37694 9614 4 vdd
port 124 nsew
rlabel metal3 s 36446 9614 36446 9614 4 vdd
port 124 nsew
rlabel metal3 s 38318 9614 38318 9614 4 vdd
port 124 nsew
rlabel metal3 s 36565 9023 36565 9023 4 vdd
port 124 nsew
rlabel metal3 s 38199 9023 38199 9023 4 vdd
port 124 nsew
rlabel metal3 s 33326 9614 33326 9614 4 vdd
port 124 nsew
rlabel metal3 s 40695 9023 40695 9023 4 vdd
port 124 nsew
rlabel metal3 s 36951 9023 36951 9023 4 vdd
port 124 nsew
rlabel metal3 s 37070 9614 37070 9614 4 vdd
port 124 nsew
rlabel metal3 s 35822 9614 35822 9614 4 vdd
port 124 nsew
rlabel metal3 s 34574 9614 34574 9614 4 vdd
port 124 nsew
rlabel metal3 s 39566 9614 39566 9614 4 vdd
port 124 nsew
rlabel metal3 s 35703 9023 35703 9023 4 vdd
port 124 nsew
rlabel metal3 s 34069 9023 34069 9023 4 vdd
port 124 nsew
rlabel metal3 s 40190 9614 40190 9614 4 vdd
port 124 nsew
rlabel metal3 s 37813 9023 37813 9023 4 vdd
port 124 nsew
rlabel metal3 s 35317 9023 35317 9023 4 vdd
port 124 nsew
rlabel metal3 s 38942 9614 38942 9614 4 vdd
port 124 nsew
rlabel metal3 s 40814 9614 40814 9614 4 vdd
port 124 nsew
rlabel metal3 s 33207 9023 33207 9023 4 vdd
port 124 nsew
rlabel metal3 s 40309 9023 40309 9023 4 vdd
port 124 nsew
rlabel metal3 s 34455 9023 34455 9023 4 vdd
port 124 nsew
rlabel metal3 s 39061 9023 39061 9023 4 vdd
port 124 nsew
rlabel metal3 s 35198 9614 35198 9614 4 vdd
port 124 nsew
rlabel metal3 s 33950 9614 33950 9614 4 vdd
port 124 nsew
rlabel metal3 s 39447 9023 39447 9023 4 vdd
port 124 nsew
rlabel metal3 s 38262 2513 38262 2513 4 vdd
port 124 nsew
rlabel metal3 s 37139 3743 37139 3743 4 gnd
port 125 nsew
rlabel metal3 s 37209 5677 37209 5677 4 gnd
port 125 nsew
rlabel metal3 s 35766 2513 35766 2513 4 vdd
port 124 nsew
rlabel metal3 s 38387 3743 38387 3743 4 gnd
port 125 nsew
rlabel metal3 s 39631 2181 39631 2181 4 gnd
port 125 nsew
rlabel metal3 s 35777 2950 35777 2950 4 gnd
port 125 nsew
rlabel metal3 s 39530 1563 39530 1563 4 vdd
port 124 nsew
rlabel metal3 s 40764 1979 40764 1979 4 gnd
port 125 nsew
rlabel metal3 s 35786 1563 35786 1563 4 vdd
port 124 nsew
rlabel metal3 s 37014 2513 37014 2513 4 vdd
port 124 nsew
rlabel metal3 s 37025 2950 37025 2950 4 gnd
port 125 nsew
rlabel metal3 s 35879 4903 35879 4903 4 vdd
port 124 nsew
rlabel metal3 s 33383 4903 33383 4903 4 vdd
port 124 nsew
rlabel metal3 s 39516 1979 39516 1979 4 gnd
port 125 nsew
rlabel metal3 s 33465 5677 33465 5677 4 gnd
port 125 nsew
rlabel metal3 s 39878 7450 39878 7450 4 gnd
port 125 nsew
rlabel metal3 s 39635 4065 39635 4065 4 vdd
port 124 nsew
rlabel metal3 s 38273 2950 38273 2950 4 gnd
port 125 nsew
rlabel metal3 s 33290 1563 33290 1563 4 vdd
port 124 nsew
rlabel metal3 s 38383 2181 38383 2181 4 gnd
port 125 nsew
rlabel metal3 s 37020 1979 37020 1979 4 gnd
port 125 nsew
rlabel metal3 s 35891 3743 35891 3743 4 gnd
port 125 nsew
rlabel metal3 s 40953 5677 40953 5677 4 gnd
port 125 nsew
rlabel metal3 s 33638 7450 33638 7450 4 gnd
port 125 nsew
rlabel metal3 s 34631 4903 34631 4903 4 vdd
port 124 nsew
rlabel metal3 s 33387 0 33387 0 4 gnd
port 125 nsew
rlabel metal3 s 38387 4065 38387 4065 4 vdd
port 124 nsew
rlabel metal3 s 40769 2950 40769 2950 4 gnd
port 125 nsew
rlabel metal3 s 39623 4903 39623 4903 4 vdd
port 124 nsew
rlabel metal3 s 40778 1563 40778 1563 4 vdd
port 124 nsew
rlabel metal3 s 37135 2181 37135 2181 4 gnd
port 125 nsew
rlabel metal3 s 37034 1563 37034 1563 4 vdd
port 124 nsew
rlabel metal3 s 39635 3743 39635 3743 4 gnd
port 125 nsew
rlabel metal3 s 36134 7450 36134 7450 4 gnd
port 125 nsew
rlabel metal3 s 35961 5677 35961 5677 4 gnd
port 125 nsew
rlabel metal3 s 34643 3743 34643 3743 4 gnd
port 125 nsew
rlabel metal3 s 38282 1563 38282 1563 4 vdd
port 124 nsew
rlabel metal3 s 40758 2513 40758 2513 4 vdd
port 124 nsew
rlabel metal3 s 39521 2950 39521 2950 4 gnd
port 125 nsew
rlabel metal3 s 33395 3743 33395 3743 4 gnd
port 125 nsew
rlabel metal3 s 37382 7450 37382 7450 4 gnd
port 125 nsew
rlabel metal3 s 33281 2950 33281 2950 4 gnd
port 125 nsew
rlabel metal3 s 33276 1979 33276 1979 4 gnd
port 125 nsew
rlabel metal3 s 38268 1979 38268 1979 4 gnd
port 125 nsew
rlabel metal3 s 34886 7450 34886 7450 4 gnd
port 125 nsew
rlabel metal3 s 35891 4065 35891 4065 4 vdd
port 124 nsew
rlabel metal3 s 33387 1120 33387 1120 4 vdd
port 124 nsew
rlabel metal3 s 40883 3743 40883 3743 4 gnd
port 125 nsew
rlabel metal3 s 39510 2513 39510 2513 4 vdd
port 124 nsew
rlabel metal3 s 34643 4065 34643 4065 4 vdd
port 124 nsew
rlabel metal3 s 33270 2513 33270 2513 4 vdd
port 124 nsew
rlabel metal3 s 40883 4065 40883 4065 4 vdd
port 124 nsew
rlabel metal3 s 35772 1979 35772 1979 4 gnd
port 125 nsew
rlabel metal3 s 33395 4065 33395 4065 4 vdd
port 124 nsew
rlabel metal3 s 34524 1979 34524 1979 4 gnd
port 125 nsew
rlabel metal3 s 38630 7450 38630 7450 4 gnd
port 125 nsew
rlabel metal3 s 38375 4903 38375 4903 4 vdd
port 124 nsew
rlabel metal3 s 34518 2513 34518 2513 4 vdd
port 124 nsew
rlabel metal3 s 34538 1563 34538 1563 4 vdd
port 124 nsew
rlabel metal3 s 34639 2181 34639 2181 4 gnd
port 125 nsew
rlabel metal3 s 37127 4903 37127 4903 4 vdd
port 124 nsew
rlabel metal3 s 34529 2950 34529 2950 4 gnd
port 125 nsew
rlabel metal3 s 35887 2181 35887 2181 4 gnd
port 125 nsew
rlabel metal3 s 40879 2181 40879 2181 4 gnd
port 125 nsew
rlabel metal3 s 39705 5677 39705 5677 4 gnd
port 125 nsew
rlabel metal3 s 38457 5677 38457 5677 4 gnd
port 125 nsew
rlabel metal3 s 37139 4065 37139 4065 4 vdd
port 124 nsew
rlabel metal3 s 34713 5677 34713 5677 4 gnd
port 125 nsew
rlabel metal3 s 40871 4903 40871 4903 4 vdd
port 124 nsew
rlabel metal3 s 33391 2181 33391 2181 4 gnd
port 125 nsew
rlabel metal3 s 45875 3743 45875 3743 4 gnd
port 125 nsew
rlabel metal3 s 48367 2181 48367 2181 4 gnd
port 125 nsew
rlabel metal3 s 48246 2513 48246 2513 4 vdd
port 124 nsew
rlabel metal3 s 48266 1563 48266 1563 4 vdd
port 124 nsew
rlabel metal3 s 44513 2950 44513 2950 4 gnd
port 125 nsew
rlabel metal3 s 44615 4903 44615 4903 4 vdd
port 124 nsew
rlabel metal3 s 43379 4065 43379 4065 4 vdd
port 124 nsew
rlabel metal3 s 47119 2181 47119 2181 4 gnd
port 125 nsew
rlabel metal3 s 43260 1979 43260 1979 4 gnd
port 125 nsew
rlabel metal3 s 43274 1563 43274 1563 4 vdd
port 124 nsew
rlabel metal3 s 48371 3743 48371 3743 4 gnd
port 125 nsew
rlabel metal3 s 42017 2950 42017 2950 4 gnd
port 125 nsew
rlabel metal3 s 42026 1563 42026 1563 4 vdd
port 124 nsew
rlabel metal3 s 43371 0 43371 0 4 gnd
port 125 nsew
rlabel metal3 s 48359 4903 48359 4903 4 vdd
port 124 nsew
rlabel metal3 s 48257 2950 48257 2950 4 gnd
port 125 nsew
rlabel metal3 s 42374 7450 42374 7450 4 gnd
port 125 nsew
rlabel metal3 s 45875 4065 45875 4065 4 vdd
port 124 nsew
rlabel metal3 s 45761 2950 45761 2950 4 gnd
port 125 nsew
rlabel metal3 s 45871 2181 45871 2181 4 gnd
port 125 nsew
rlabel metal3 s 44627 4065 44627 4065 4 vdd
port 124 nsew
rlabel metal3 s 48252 1979 48252 1979 4 gnd
port 125 nsew
rlabel metal3 s 42119 4903 42119 4903 4 vdd
port 124 nsew
rlabel metal3 s 43379 3743 43379 3743 4 gnd
port 125 nsew
rlabel metal3 s 42012 1979 42012 1979 4 gnd
port 125 nsew
rlabel metal3 s 47193 5677 47193 5677 4 gnd
port 125 nsew
rlabel metal3 s 47009 2950 47009 2950 4 gnd
port 125 nsew
rlabel metal3 s 43367 4903 43367 4903 4 vdd
port 124 nsew
rlabel metal3 s 42006 2513 42006 2513 4 vdd
port 124 nsew
rlabel metal3 s 44627 3743 44627 3743 4 gnd
port 125 nsew
rlabel metal3 s 48614 7450 48614 7450 4 gnd
port 125 nsew
rlabel metal3 s 47018 1563 47018 1563 4 vdd
port 124 nsew
rlabel metal3 s 47366 7450 47366 7450 4 gnd
port 125 nsew
rlabel metal3 s 43622 7450 43622 7450 4 gnd
port 125 nsew
rlabel metal3 s 44623 2181 44623 2181 4 gnd
port 125 nsew
rlabel metal3 s 47004 1979 47004 1979 4 gnd
port 125 nsew
rlabel metal3 s 42131 4065 42131 4065 4 vdd
port 124 nsew
rlabel metal3 s 43265 2950 43265 2950 4 gnd
port 125 nsew
rlabel metal3 s 44870 7450 44870 7450 4 gnd
port 125 nsew
rlabel metal3 s 44502 2513 44502 2513 4 vdd
port 124 nsew
rlabel metal3 s 47123 3743 47123 3743 4 gnd
port 125 nsew
rlabel metal3 s 45770 1563 45770 1563 4 vdd
port 124 nsew
rlabel metal3 s 44508 1979 44508 1979 4 gnd
port 125 nsew
rlabel metal3 s 42127 2181 42127 2181 4 gnd
port 125 nsew
rlabel metal3 s 46118 7450 46118 7450 4 gnd
port 125 nsew
rlabel metal3 s 46998 2513 46998 2513 4 vdd
port 124 nsew
rlabel metal3 s 45750 2513 45750 2513 4 vdd
port 124 nsew
rlabel metal3 s 45756 1979 45756 1979 4 gnd
port 125 nsew
rlabel metal3 s 43371 1120 43371 1120 4 vdd
port 124 nsew
rlabel metal3 s 45863 4903 45863 4903 4 vdd
port 124 nsew
rlabel metal3 s 41126 7450 41126 7450 4 gnd
port 125 nsew
rlabel metal3 s 43375 2181 43375 2181 4 gnd
port 125 nsew
rlabel metal3 s 43254 2513 43254 2513 4 vdd
port 124 nsew
rlabel metal3 s 42201 5677 42201 5677 4 gnd
port 125 nsew
rlabel metal3 s 45945 5677 45945 5677 4 gnd
port 125 nsew
rlabel metal3 s 48371 4065 48371 4065 4 vdd
port 124 nsew
rlabel metal3 s 48441 5677 48441 5677 4 gnd
port 125 nsew
rlabel metal3 s 44522 1563 44522 1563 4 vdd
port 124 nsew
rlabel metal3 s 47123 4065 47123 4065 4 vdd
port 124 nsew
rlabel metal3 s 44697 5677 44697 5677 4 gnd
port 125 nsew
rlabel metal3 s 43449 5677 43449 5677 4 gnd
port 125 nsew
rlabel metal3 s 47111 4903 47111 4903 4 vdd
port 124 nsew
rlabel metal3 s 42131 3743 42131 3743 4 gnd
port 125 nsew
rlabel metal3 s 61982 13759 61982 13759 4 vdd
port 124 nsew
rlabel metal3 s 62633 13766 62633 13766 4 vdd
port 124 nsew
rlabel metal3 s 63956 12969 63956 12969 4 vdd
port 124 nsew
rlabel metal3 s 63068 15362 63068 15362 4 vdd
port 124 nsew
rlabel metal3 s 62633 12976 62633 12976 4 vdd
port 124 nsew
rlabel metal3 s 64824 15339 64824 15339 4 gnd
port 125 nsew
rlabel metal3 s 61982 15339 61982 15339 4 vdd
port 124 nsew
rlabel metal3 s 64228 12969 64228 12969 4 gnd
port 125 nsew
rlabel metal3 s 62636 15362 62636 15362 4 vdd
port 124 nsew
rlabel metal3 s 63068 16152 63068 16152 4 vdd
port 124 nsew
rlabel metal3 s 61982 16129 61982 16129 4 vdd
port 124 nsew
rlabel metal3 s 64552 15339 64552 15339 4 vdd
port 124 nsew
rlabel metal3 s 63058 13766 63058 13766 4 gnd
port 125 nsew
rlabel metal3 s 63058 12976 63058 12976 4 gnd
port 125 nsew
rlabel metal3 s 62254 15339 62254 15339 4 gnd
port 125 nsew
rlabel metal3 s 62254 16129 62254 16129 4 gnd
port 125 nsew
rlabel metal3 s 63493 16152 63493 16152 4 gnd
port 125 nsew
rlabel metal3 s 61982 12969 61982 12969 4 vdd
port 124 nsew
rlabel metal3 s 62254 13759 62254 13759 4 gnd
port 125 nsew
rlabel metal3 s 63493 15362 63493 15362 4 gnd
port 125 nsew
rlabel metal3 s 62636 16152 62636 16152 4 vdd
port 124 nsew
rlabel metal3 s 62254 12969 62254 12969 4 gnd
port 125 nsew
rlabel metal3 s 60203 12992 60203 12992 4 gnd
port 125 nsew
rlabel metal3 s 59346 16510 59346 16510 4 vdd
port 124 nsew
rlabel metal3 s 60203 15362 60203 15362 4 gnd
port 125 nsew
rlabel metal3 s 59346 15362 59346 15362 4 vdd
port 124 nsew
rlabel metal3 s 58964 13759 58964 13759 4 gnd
port 125 nsew
rlabel metal3 s 58692 14549 58692 14549 4 vdd
port 124 nsew
rlabel metal3 s 59778 13350 59778 13350 4 vdd
port 124 nsew
rlabel metal3 s 58964 14944 58964 14944 4 gnd
port 125 nsew
rlabel metal3 s 58692 14944 58692 14944 4 vdd
port 124 nsew
rlabel metal3 s 60203 14198 60203 14198 4 gnd
port 125 nsew
rlabel metal3 s 60203 13408 60203 13408 4 gnd
port 125 nsew
rlabel metal3 s 59346 16152 59346 16152 4 vdd
port 124 nsew
rlabel metal3 s 59778 14572 59778 14572 4 vdd
port 124 nsew
rlabel metal3 s 58692 16129 58692 16129 4 vdd
port 124 nsew
rlabel metal3 s 58964 14549 58964 14549 4 gnd
port 125 nsew
rlabel metal3 s 59346 14140 59346 14140 4 vdd
port 124 nsew
rlabel metal3 s 59346 14572 59346 14572 4 vdd
port 124 nsew
rlabel metal3 s 58964 15339 58964 15339 4 gnd
port 125 nsew
rlabel metal3 s 59346 13782 59346 13782 4 vdd
port 124 nsew
rlabel metal3 s 58964 15734 58964 15734 4 gnd
port 125 nsew
rlabel metal3 s 59346 13350 59346 13350 4 vdd
port 124 nsew
rlabel metal3 s 60203 14572 60203 14572 4 gnd
port 125 nsew
rlabel metal3 s 59778 16510 59778 16510 4 vdd
port 124 nsew
rlabel metal3 s 58692 12969 58692 12969 4 vdd
port 124 nsew
rlabel metal3 s 59346 15720 59346 15720 4 vdd
port 124 nsew
rlabel metal3 s 59346 12992 59346 12992 4 vdd
port 124 nsew
rlabel metal3 s 58692 13364 58692 13364 4 vdd
port 124 nsew
rlabel metal3 s 59778 14930 59778 14930 4 vdd
port 124 nsew
rlabel metal3 s 60203 16152 60203 16152 4 gnd
port 125 nsew
rlabel metal3 s 59778 15362 59778 15362 4 vdd
port 124 nsew
rlabel metal3 s 58964 12969 58964 12969 4 gnd
port 125 nsew
rlabel metal3 s 59778 12992 59778 12992 4 vdd
port 124 nsew
rlabel metal3 s 60203 12618 60203 12618 4 gnd
port 125 nsew
rlabel metal3 s 60203 15778 60203 15778 4 gnd
port 125 nsew
rlabel metal3 s 60203 13782 60203 13782 4 gnd
port 125 nsew
rlabel metal3 s 59778 13782 59778 13782 4 vdd
port 124 nsew
rlabel metal3 s 58692 15339 58692 15339 4 vdd
port 124 nsew
rlabel metal3 s 59778 15720 59778 15720 4 vdd
port 124 nsew
rlabel metal3 s 59778 14140 59778 14140 4 vdd
port 124 nsew
rlabel metal3 s 58964 16524 58964 16524 4 gnd
port 125 nsew
rlabel metal3 s 59346 14930 59346 14930 4 vdd
port 124 nsew
rlabel metal3 s 60203 14988 60203 14988 4 gnd
port 125 nsew
rlabel metal3 s 58964 13364 58964 13364 4 gnd
port 125 nsew
rlabel metal3 s 58692 14154 58692 14154 4 vdd
port 124 nsew
rlabel metal3 s 58692 13759 58692 13759 4 vdd
port 124 nsew
rlabel metal3 s 58964 14154 58964 14154 4 gnd
port 125 nsew
rlabel metal3 s 59778 16152 59778 16152 4 vdd
port 124 nsew
rlabel metal3 s 58692 16524 58692 16524 4 vdd
port 124 nsew
rlabel metal3 s 58964 16129 58964 16129 4 gnd
port 125 nsew
rlabel metal3 s 58692 15734 58692 15734 4 vdd
port 124 nsew
rlabel metal3 s 60203 16568 60203 16568 4 gnd
port 125 nsew
rlabel metal3 s 60203 12202 60203 12202 4 gnd
port 125 nsew
rlabel metal3 s 58964 10994 58964 10994 4 gnd
port 125 nsew
rlabel metal3 s 59778 12202 59778 12202 4 vdd
port 124 nsew
rlabel metal3 s 58692 12574 58692 12574 4 vdd
port 124 nsew
rlabel metal3 s 58964 12179 58964 12179 4 gnd
port 125 nsew
rlabel metal3 s 59778 10622 59778 10622 4 vdd
port 124 nsew
rlabel metal3 s 59346 10622 59346 10622 4 vdd
port 124 nsew
rlabel metal3 s 58692 11389 58692 11389 4 vdd
port 124 nsew
rlabel metal3 s 59778 10980 59778 10980 4 vdd
port 124 nsew
rlabel metal3 s 58692 12179 58692 12179 4 vdd
port 124 nsew
rlabel metal3 s 58964 11389 58964 11389 4 gnd
port 125 nsew
rlabel metal3 s 58964 12574 58964 12574 4 gnd
port 125 nsew
rlabel metal3 s 59778 11770 59778 11770 4 vdd
port 124 nsew
rlabel metal3 s 59346 12202 59346 12202 4 vdd
port 124 nsew
rlabel metal3 s 59346 11412 59346 11412 4 vdd
port 124 nsew
rlabel metal3 s 58964 10599 58964 10599 4 gnd
port 125 nsew
rlabel metal3 s 59346 10980 59346 10980 4 vdd
port 124 nsew
rlabel metal3 s 58692 11784 58692 11784 4 vdd
port 124 nsew
rlabel metal3 s 58964 11784 58964 11784 4 gnd
port 125 nsew
rlabel metal3 s 60203 11412 60203 11412 4 gnd
port 125 nsew
rlabel metal3 s 60203 10622 60203 10622 4 gnd
port 125 nsew
rlabel metal3 s 59346 11770 59346 11770 4 vdd
port 124 nsew
rlabel metal3 s 58692 10599 58692 10599 4 vdd
port 124 nsew
rlabel metal3 s 60203 11038 60203 11038 4 gnd
port 125 nsew
rlabel metal3 s 59346 12560 59346 12560 4 vdd
port 124 nsew
rlabel metal3 s 59778 11412 59778 11412 4 vdd
port 124 nsew
rlabel metal3 s 60203 11828 60203 11828 4 gnd
port 125 nsew
rlabel metal3 s 59778 12560 59778 12560 4 vdd
port 124 nsew
rlabel metal3 s 58692 10994 58692 10994 4 vdd
port 124 nsew
rlabel metal3 s 63058 10606 63058 10606 4 gnd
port 125 nsew
rlabel metal3 s 62633 11396 62633 11396 4 vdd
port 124 nsew
rlabel metal3 s 62254 11389 62254 11389 4 gnd
port 125 nsew
rlabel metal3 s 62633 10606 62633 10606 4 vdd
port 124 nsew
rlabel metal3 s 64228 10599 64228 10599 4 gnd
port 125 nsew
rlabel metal3 s 63956 10599 63956 10599 4 vdd
port 124 nsew
rlabel metal3 s 61982 11389 61982 11389 4 vdd
port 124 nsew
rlabel metal3 s 61982 10599 61982 10599 4 vdd
port 124 nsew
rlabel metal3 s 63058 11396 63058 11396 4 gnd
port 125 nsew
rlabel metal3 s 62254 10599 62254 10599 4 gnd
port 125 nsew
rlabel metal3 s 53990 14678 53990 14678 4 gnd
port 125 nsew
rlabel metal3 s 53990 13098 53990 13098 4 gnd
port 125 nsew
rlabel metal3 s 51541 9023 51541 9023 4 vdd
port 124 nsew
rlabel metal3 s 53990 16732 53990 16732 4 gnd
port 125 nsew
rlabel metal3 s 52046 9614 52046 9614 4 vdd
port 124 nsew
rlabel metal3 s 53990 11202 53990 11202 4 gnd
port 125 nsew
rlabel metal3 s 53990 13572 53990 13572 4 gnd
port 125 nsew
rlabel metal3 s 53990 16495 53990 16495 4 gnd
port 125 nsew
rlabel metal3 s 53990 12545 53990 12545 4 gnd
port 125 nsew
rlabel metal3 s 53990 10175 53990 10175 4 gnd
port 125 nsew
rlabel metal3 s 53990 14125 53990 14125 4 gnd
port 125 nsew
rlabel metal3 s 53990 12782 53990 12782 4 gnd
port 125 nsew
rlabel metal3 s 53990 11992 53990 11992 4 gnd
port 125 nsew
rlabel metal3 s 53990 10412 53990 10412 4 gnd
port 125 nsew
rlabel metal3 s 53990 12308 53990 12308 4 gnd
port 125 nsew
rlabel metal3 s 53990 9938 53990 9938 4 gnd
port 125 nsew
rlabel metal3 s 49431 9023 49431 9023 4 vdd
port 124 nsew
rlabel metal3 s 53990 15468 53990 15468 4 gnd
port 125 nsew
rlabel metal3 s 52789 9023 52789 9023 4 vdd
port 124 nsew
rlabel metal3 s 53990 16258 53990 16258 4 gnd
port 125 nsew
rlabel metal3 s 49045 9023 49045 9023 4 vdd
port 124 nsew
rlabel metal3 s 53990 10965 53990 10965 4 gnd
port 125 nsew
rlabel metal3 s 53990 10728 53990 10728 4 gnd
port 125 nsew
rlabel metal3 s 50174 9614 50174 9614 4 vdd
port 124 nsew
rlabel metal3 s 53990 13888 53990 13888 4 gnd
port 125 nsew
rlabel metal3 s 53990 15152 53990 15152 4 gnd
port 125 nsew
rlabel metal3 s 48926 9614 48926 9614 4 vdd
port 124 nsew
rlabel metal3 s 51927 9023 51927 9023 4 vdd
port 124 nsew
rlabel metal3 s 53990 13335 53990 13335 4 gnd
port 125 nsew
rlabel metal3 s 53990 14362 53990 14362 4 gnd
port 125 nsew
rlabel metal3 s 53990 14915 53990 14915 4 gnd
port 125 nsew
rlabel metal3 s 53990 15942 53990 15942 4 gnd
port 125 nsew
rlabel metal3 s 53990 11755 53990 11755 4 gnd
port 125 nsew
rlabel metal3 s 49550 9614 49550 9614 4 vdd
port 124 nsew
rlabel metal3 s 53990 15705 53990 15705 4 gnd
port 125 nsew
rlabel metal3 s 51422 9614 51422 9614 4 vdd
port 124 nsew
rlabel metal3 s 50798 9614 50798 9614 4 vdd
port 124 nsew
rlabel metal3 s 53990 11518 53990 11518 4 gnd
port 125 nsew
rlabel metal3 s 52670 9614 52670 9614 4 vdd
port 124 nsew
rlabel metal3 s 50679 9023 50679 9023 4 vdd
port 124 nsew
rlabel metal3 s 53294 9614 53294 9614 4 vdd
port 124 nsew
rlabel metal3 s 50293 9023 50293 9023 4 vdd
port 124 nsew
rlabel metal3 s 52115 3743 52115 3743 4 gnd
port 125 nsew
rlabel metal3 s 49619 3743 49619 3743 4 gnd
port 125 nsew
rlabel metal3 s 52111 2181 52111 2181 4 gnd
port 125 nsew
rlabel metal3 s 50753 2950 50753 2950 4 gnd
port 125 nsew
rlabel metal3 s 49505 2950 49505 2950 4 gnd
port 125 nsew
rlabel metal3 s 51996 1979 51996 1979 4 gnd
port 125 nsew
rlabel metal3 s 50867 4065 50867 4065 4 vdd
port 124 nsew
rlabel metal3 s 49514 1563 49514 1563 4 vdd
port 124 nsew
rlabel metal3 s 49689 5677 49689 5677 4 gnd
port 125 nsew
rlabel metal3 s 50867 3743 50867 3743 4 gnd
port 125 nsew
rlabel metal3 s 49615 2181 49615 2181 4 gnd
port 125 nsew
rlabel metal3 s 50937 5677 50937 5677 4 gnd
port 125 nsew
rlabel metal3 s 52001 2950 52001 2950 4 gnd
port 125 nsew
rlabel metal3 s 50863 2181 50863 2181 4 gnd
port 125 nsew
rlabel metal3 s 52185 5677 52185 5677 4 gnd
port 125 nsew
rlabel metal3 s 50762 1563 50762 1563 4 vdd
port 124 nsew
rlabel metal3 s 49607 4903 49607 4903 4 vdd
port 124 nsew
rlabel metal3 s 50748 1979 50748 1979 4 gnd
port 125 nsew
rlabel metal3 s 51110 7450 51110 7450 4 gnd
port 125 nsew
rlabel metal3 s 50742 2513 50742 2513 4 vdd
port 124 nsew
rlabel metal3 s 51990 2513 51990 2513 4 vdd
port 124 nsew
rlabel metal3 s 52103 4903 52103 4903 4 vdd
port 124 nsew
rlabel metal3 s 49500 1979 49500 1979 4 gnd
port 125 nsew
rlabel metal3 s 49619 4065 49619 4065 4 vdd
port 124 nsew
rlabel metal3 s 52010 1563 52010 1563 4 vdd
port 124 nsew
rlabel metal3 s 52358 7450 52358 7450 4 gnd
port 125 nsew
rlabel metal3 s 50855 4903 50855 4903 4 vdd
port 124 nsew
rlabel metal3 s 49862 7450 49862 7450 4 gnd
port 125 nsew
rlabel metal3 s 52115 4065 52115 4065 4 vdd
port 124 nsew
rlabel metal3 s 49494 2513 49494 2513 4 vdd
port 124 nsew
<< properties >>
string FIXED_BBOX 0 0 66112 67359
string GDS_END 6425618
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 5901526
<< end >>
