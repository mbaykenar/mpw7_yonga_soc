magic
tech sky130B
magscale 12 1
timestamp 1598777679
<< metal5 >>
rect 0 20 15 75
rect 30 20 45 75
rect 60 20 75 75
rect 0 10 75 20
rect 5 5 75 10
rect 10 0 30 5
rect 45 0 75 5
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
