VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO axi_node_intf_wrap
  CLASS BLOCK ;
  FOREIGN axi_node_intf_wrap ;
  ORIGIN 0.000 0.000 ;
  SIZE 2400.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 0.000 1954.910 4.000 ;
    END
  END clk
  PIN m00_ar_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END m00_ar_addr[0]
  PIN m00_ar_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 596.000 808.590 600.000 ;
    END
  END m00_ar_addr[10]
  PIN m00_ar_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END m00_ar_addr[11]
  PIN m00_ar_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 596.000 409.310 600.000 ;
    END
  END m00_ar_addr[12]
  PIN m00_ar_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 596.000 1716.630 600.000 ;
    END
  END m00_ar_addr[13]
  PIN m00_ar_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END m00_ar_addr[14]
  PIN m00_ar_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 596.000 850.450 600.000 ;
    END
  END m00_ar_addr[15]
  PIN m00_ar_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 596.000 1211.090 600.000 ;
    END
  END m00_ar_addr[16]
  PIN m00_ar_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 23.840 2400.000 24.440 ;
    END
  END m00_ar_addr[17]
  PIN m00_ar_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 0.000 2212.510 4.000 ;
    END
  END m00_ar_addr[18]
  PIN m00_ar_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 0.000 2257.590 4.000 ;
    END
  END m00_ar_addr[19]
  PIN m00_ar_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 496.440 2400.000 497.040 ;
    END
  END m00_ar_addr[1]
  PIN m00_ar_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 596.000 1030.770 600.000 ;
    END
  END m00_ar_addr[20]
  PIN m00_ar_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 0.000 2270.470 4.000 ;
    END
  END m00_ar_addr[21]
  PIN m00_ar_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 596.000 1314.130 600.000 ;
    END
  END m00_ar_addr[22]
  PIN m00_ar_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 596.000 299.830 600.000 ;
    END
  END m00_ar_addr[23]
  PIN m00_ar_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.750 0.000 1781.030 4.000 ;
    END
  END m00_ar_addr[24]
  PIN m00_ar_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.030 0.000 2341.310 4.000 ;
    END
  END m00_ar_addr[25]
  PIN m00_ar_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END m00_ar_addr[26]
  PIN m00_ar_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END m00_ar_addr[27]
  PIN m00_ar_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 596.000 1703.750 600.000 ;
    END
  END m00_ar_addr[28]
  PIN m00_ar_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 596.000 863.330 600.000 ;
    END
  END m00_ar_addr[29]
  PIN m00_ar_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.310 596.000 1774.590 600.000 ;
    END
  END m00_ar_addr[2]
  PIN m00_ar_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 596.000 84.090 600.000 ;
    END
  END m00_ar_addr[30]
  PIN m00_ar_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END m00_ar_addr[31]
  PIN m00_ar_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 129.240 2400.000 129.840 ;
    END
  END m00_ar_addr[3]
  PIN m00_ar_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END m00_ar_addr[4]
  PIN m00_ar_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 0.000 1835.770 4.000 ;
    END
  END m00_ar_addr[5]
  PIN m00_ar_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 596.000 554.210 600.000 ;
    END
  END m00_ar_addr[6]
  PIN m00_ar_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 596.000 1178.890 600.000 ;
    END
  END m00_ar_addr[7]
  PIN m00_ar_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END m00_ar_addr[8]
  PIN m00_ar_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END m00_ar_addr[9]
  PIN m00_ar_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 596.000 534.890 600.000 ;
    END
  END m00_ar_burst[0]
  PIN m00_ar_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END m00_ar_burst[1]
  PIN m00_ar_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 596.000 579.970 600.000 ;
    END
  END m00_ar_cache[0]
  PIN m00_ar_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 596.000 1790.690 600.000 ;
    END
  END m00_ar_cache[1]
  PIN m00_ar_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END m00_ar_cache[2]
  PIN m00_ar_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 596.000 1658.670 600.000 ;
    END
  END m00_ar_cache[3]
  PIN m00_ar_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END m00_ar_id[0]
  PIN m00_ar_id[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END m00_ar_id[10]
  PIN m00_ar_id[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END m00_ar_id[11]
  PIN m00_ar_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 340.040 2400.000 340.640 ;
    END
  END m00_ar_id[1]
  PIN m00_ar_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 125.840 2400.000 126.440 ;
    END
  END m00_ar_id[2]
  PIN m00_ar_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END m00_ar_id[3]
  PIN m00_ar_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 265.240 2400.000 265.840 ;
    END
  END m00_ar_id[4]
  PIN m00_ar_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 596.000 383.550 600.000 ;
    END
  END m00_ar_id[5]
  PIN m00_ar_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 550.840 2400.000 551.440 ;
    END
  END m00_ar_id[6]
  PIN m00_ar_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 0.000 1822.890 4.000 ;
    END
  END m00_ar_id[7]
  PIN m00_ar_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 596.000 1330.230 600.000 ;
    END
  END m00_ar_id[8]
  PIN m00_ar_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 493.040 2400.000 493.640 ;
    END
  END m00_ar_id[9]
  PIN m00_ar_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 596.000 901.970 600.000 ;
    END
  END m00_ar_len[0]
  PIN m00_ar_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 596.000 1111.270 600.000 ;
    END
  END m00_ar_len[1]
  PIN m00_ar_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 596.000 1317.350 600.000 ;
    END
  END m00_ar_len[2]
  PIN m00_ar_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 596.000 959.930 600.000 ;
    END
  END m00_ar_len[3]
  PIN m00_ar_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 596.000 821.470 600.000 ;
    END
  END m00_ar_len[4]
  PIN m00_ar_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END m00_ar_len[5]
  PIN m00_ar_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 596.000 1758.490 600.000 ;
    END
  END m00_ar_len[6]
  PIN m00_ar_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.790 0.000 2045.070 4.000 ;
    END
  END m00_ar_len[7]
  PIN m00_ar_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 596.000 1401.070 600.000 ;
    END
  END m00_ar_lock
  PIN m00_ar_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 596.000 2212.510 600.000 ;
    END
  END m00_ar_prot[0]
  PIN m00_ar_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.090 0.000 2093.370 4.000 ;
    END
  END m00_ar_prot[1]
  PIN m00_ar_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 596.000 847.230 600.000 ;
    END
  END m00_ar_prot[2]
  PIN m00_ar_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 61.240 2400.000 61.840 ;
    END
  END m00_ar_qos[0]
  PIN m00_ar_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 596.000 1291.590 600.000 ;
    END
  END m00_ar_qos[1]
  PIN m00_ar_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 81.640 2400.000 82.240 ;
    END
  END m00_ar_qos[2]
  PIN m00_ar_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 596.000 1127.370 600.000 ;
    END
  END m00_ar_qos[3]
  PIN m00_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END m00_ar_ready
  PIN m00_ar_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END m00_ar_region[0]
  PIN m00_ar_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END m00_ar_region[1]
  PIN m00_ar_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 596.000 1603.930 600.000 ;
    END
  END m00_ar_region[2]
  PIN m00_ar_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 596.000 35.790 600.000 ;
    END
  END m00_ar_region[3]
  PIN m00_ar_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 596.000 6.810 600.000 ;
    END
  END m00_ar_size[0]
  PIN m00_ar_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 380.840 2400.000 381.440 ;
    END
  END m00_ar_size[1]
  PIN m00_ar_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 0.000 1536.310 4.000 ;
    END
  END m00_ar_size[2]
  PIN m00_ar_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END m00_ar_user[-1]
  PIN m00_ar_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 596.000 853.670 600.000 ;
    END
  END m00_ar_user[0]
  PIN m00_ar_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 596.000 1826.110 600.000 ;
    END
  END m00_ar_valid
  PIN m00_aw_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END m00_aw_addr[0]
  PIN m00_aw_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 596.000 1932.370 600.000 ;
    END
  END m00_aw_addr[10]
  PIN m00_aw_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 596.000 509.130 600.000 ;
    END
  END m00_aw_addr[11]
  PIN m00_aw_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END m00_aw_addr[12]
  PIN m00_aw_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 503.240 2400.000 503.840 ;
    END
  END m00_aw_addr[13]
  PIN m00_aw_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 40.840 2400.000 41.440 ;
    END
  END m00_aw_addr[14]
  PIN m00_aw_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END m00_aw_addr[15]
  PIN m00_aw_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 224.440 2400.000 225.040 ;
    END
  END m00_aw_addr[16]
  PIN m00_aw_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.930 596.000 2164.210 600.000 ;
    END
  END m00_aw_addr[17]
  PIN m00_aw_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 326.440 2400.000 327.040 ;
    END
  END m00_aw_addr[18]
  PIN m00_aw_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END m00_aw_addr[19]
  PIN m00_aw_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 414.840 2400.000 415.440 ;
    END
  END m00_aw_addr[1]
  PIN m00_aw_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END m00_aw_addr[20]
  PIN m00_aw_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END m00_aw_addr[21]
  PIN m00_aw_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 596.000 1249.730 600.000 ;
    END
  END m00_aw_addr[22]
  PIN m00_aw_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 0.000 1481.570 4.000 ;
    END
  END m00_aw_addr[23]
  PIN m00_aw_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 596.000 1021.110 600.000 ;
    END
  END m00_aw_addr[24]
  PIN m00_aw_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 596.000 496.250 600.000 ;
    END
  END m00_aw_addr[25]
  PIN m00_aw_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END m00_aw_addr[26]
  PIN m00_aw_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.710 0.000 1838.990 4.000 ;
    END
  END m00_aw_addr[27]
  PIN m00_aw_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 387.640 2400.000 388.240 ;
    END
  END m00_aw_addr[28]
  PIN m00_aw_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 596.000 96.970 600.000 ;
    END
  END m00_aw_addr[29]
  PIN m00_aw_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.330 0.000 2067.610 4.000 ;
    END
  END m00_aw_addr[2]
  PIN m00_aw_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 596.000 2106.250 600.000 ;
    END
  END m00_aw_addr[30]
  PIN m00_aw_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END m00_aw_addr[31]
  PIN m00_aw_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.710 596.000 1999.990 600.000 ;
    END
  END m00_aw_addr[3]
  PIN m00_aw_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 4.000 ;
    END
  END m00_aw_addr[4]
  PIN m00_aw_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 596.000 245.090 600.000 ;
    END
  END m00_aw_addr[5]
  PIN m00_aw_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END m00_aw_addr[6]
  PIN m00_aw_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END m00_aw_addr[7]
  PIN m00_aw_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 596.000 998.570 600.000 ;
    END
  END m00_aw_addr[8]
  PIN m00_aw_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END m00_aw_addr[9]
  PIN m00_aw_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 4.000 ;
    END
  END m00_aw_burst[0]
  PIN m00_aw_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END m00_aw_burst[1]
  PIN m00_aw_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END m00_aw_cache[0]
  PIN m00_aw_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 596.000 1623.250 600.000 ;
    END
  END m00_aw_cache[1]
  PIN m00_aw_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 370.640 2400.000 371.240 ;
    END
  END m00_aw_cache[2]
  PIN m00_aw_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END m00_aw_cache[3]
  PIN m00_aw_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 596.000 567.090 600.000 ;
    END
  END m00_aw_id[0]
  PIN m00_aw_id[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 4.000 ;
    END
  END m00_aw_id[10]
  PIN m00_aw_id[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END m00_aw_id[11]
  PIN m00_aw_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 596.000 937.390 600.000 ;
    END
  END m00_aw_id[1]
  PIN m00_aw_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 596.000 1050.090 600.000 ;
    END
  END m00_aw_id[2]
  PIN m00_aw_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 596.000 180.690 600.000 ;
    END
  END m00_aw_id[3]
  PIN m00_aw_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 584.840 2400.000 585.440 ;
    END
  END m00_aw_id[4]
  PIN m00_aw_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END m00_aw_id[5]
  PIN m00_aw_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END m00_aw_id[6]
  PIN m00_aw_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 0.000 1851.870 4.000 ;
    END
  END m00_aw_id[7]
  PIN m00_aw_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 596.000 93.750 600.000 ;
    END
  END m00_aw_id[8]
  PIN m00_aw_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 596.000 531.670 600.000 ;
    END
  END m00_aw_id[9]
  PIN m00_aw_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END m00_aw_len[0]
  PIN m00_aw_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.550 596.000 2231.830 600.000 ;
    END
  END m00_aw_len[1]
  PIN m00_aw_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END m00_aw_len[2]
  PIN m00_aw_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 357.040 2400.000 357.640 ;
    END
  END m00_aw_len[3]
  PIN m00_aw_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 596.000 576.750 600.000 ;
    END
  END m00_aw_len[4]
  PIN m00_aw_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END m00_aw_len[5]
  PIN m00_aw_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 596.000 966.370 600.000 ;
    END
  END m00_aw_len[6]
  PIN m00_aw_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 596.000 927.730 600.000 ;
    END
  END m00_aw_len[7]
  PIN m00_aw_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 596.000 831.130 600.000 ;
    END
  END m00_aw_lock
  PIN m00_aw_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END m00_aw_prot[0]
  PIN m00_aw_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 596.000 1417.170 600.000 ;
    END
  END m00_aw_prot[1]
  PIN m00_aw_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END m00_aw_prot[2]
  PIN m00_aw_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 596.000 45.450 600.000 ;
    END
  END m00_aw_qos[0]
  PIN m00_aw_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 596.000 1288.370 600.000 ;
    END
  END m00_aw_qos[1]
  PIN m00_aw_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END m00_aw_qos[2]
  PIN m00_aw_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 596.000 132.390 600.000 ;
    END
  END m00_aw_qos[3]
  PIN m00_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.350 596.000 1877.630 600.000 ;
    END
  END m00_aw_ready
  PIN m00_aw_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 0.000 1314.130 4.000 ;
    END
  END m00_aw_region[0]
  PIN m00_aw_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END m00_aw_region[1]
  PIN m00_aw_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END m00_aw_region[2]
  PIN m00_aw_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END m00_aw_region[3]
  PIN m00_aw_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 596.000 1240.070 600.000 ;
    END
  END m00_aw_size[0]
  PIN m00_aw_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END m00_aw_size[1]
  PIN m00_aw_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 516.840 2400.000 517.440 ;
    END
  END m00_aw_size[2]
  PIN m00_aw_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END m00_aw_user[-1]
  PIN m00_aw_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 596.000 1858.310 600.000 ;
    END
  END m00_aw_user[0]
  PIN m00_aw_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.910 0.000 2032.190 4.000 ;
    END
  END m00_aw_valid
  PIN m00_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END m00_b_id[0]
  PIN m00_b_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END m00_b_id[10]
  PIN m00_b_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 596.000 1726.290 600.000 ;
    END
  END m00_b_id[11]
  PIN m00_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END m00_b_id[1]
  PIN m00_b_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.870 0.000 2090.150 4.000 ;
    END
  END m00_b_id[2]
  PIN m00_b_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 465.840 2400.000 466.440 ;
    END
  END m00_b_id[3]
  PIN m00_b_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END m00_b_id[4]
  PIN m00_b_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 0.000 1771.370 4.000 ;
    END
  END m00_b_id[5]
  PIN m00_b_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END m00_b_id[6]
  PIN m00_b_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 596.000 1468.690 600.000 ;
    END
  END m00_b_id[7]
  PIN m00_b_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 0.000 1880.850 4.000 ;
    END
  END m00_b_id[8]
  PIN m00_b_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END m00_b_id[9]
  PIN m00_b_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END m00_b_ready
  PIN m00_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 0.000 2012.870 4.000 ;
    END
  END m00_b_resp[0]
  PIN m00_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END m00_b_resp[1]
  PIN m00_b_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 4.000 ;
    END
  END m00_b_user[-1]
  PIN m00_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 445.440 2400.000 446.040 ;
    END
  END m00_b_user[0]
  PIN m00_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END m00_b_valid
  PIN m00_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 596.000 1391.410 600.000 ;
    END
  END m00_r_data[0]
  PIN m00_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END m00_r_data[10]
  PIN m00_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 596.000 1143.470 600.000 ;
    END
  END m00_r_data[11]
  PIN m00_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.990 0.000 2238.270 4.000 ;
    END
  END m00_r_data[12]
  PIN m00_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END m00_r_data[13]
  PIN m00_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 0.000 1339.890 4.000 ;
    END
  END m00_r_data[14]
  PIN m00_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.110 596.000 2386.390 600.000 ;
    END
  END m00_r_data[15]
  PIN m00_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 596.000 328.810 600.000 ;
    END
  END m00_r_data[16]
  PIN m00_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END m00_r_data[17]
  PIN m00_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END m00_r_data[18]
  PIN m00_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END m00_r_data[19]
  PIN m00_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END m00_r_data[1]
  PIN m00_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 596.000 55.110 600.000 ;
    END
  END m00_r_data[20]
  PIN m00_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 438.640 2400.000 439.240 ;
    END
  END m00_r_data[21]
  PIN m00_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END m00_r_data[22]
  PIN m00_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 596.000 779.610 600.000 ;
    END
  END m00_r_data[23]
  PIN m00_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 596.000 0.370 600.000 ;
    END
  END m00_r_data[24]
  PIN m00_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 51.040 2400.000 51.640 ;
    END
  END m00_r_data[25]
  PIN m00_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END m00_r_data[26]
  PIN m00_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 596.000 1082.290 600.000 ;
    END
  END m00_r_data[27]
  PIN m00_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 44.240 2400.000 44.840 ;
    END
  END m00_r_data[28]
  PIN m00_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END m00_r_data[29]
  PIN m00_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 596.000 444.730 600.000 ;
    END
  END m00_r_data[2]
  PIN m00_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 596.000 1355.990 600.000 ;
    END
  END m00_r_data[30]
  PIN m00_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 596.000 528.450 600.000 ;
    END
  END m00_r_data[31]
  PIN m00_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 596.000 177.470 600.000 ;
    END
  END m00_r_data[3]
  PIN m00_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 596.000 212.890 600.000 ;
    END
  END m00_r_data[4]
  PIN m00_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 596.000 650.810 600.000 ;
    END
  END m00_r_data[5]
  PIN m00_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 596.000 618.610 600.000 ;
    END
  END m00_r_data[6]
  PIN m00_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 0.000 1681.210 4.000 ;
    END
  END m00_r_data[7]
  PIN m00_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 596.000 1874.410 600.000 ;
    END
  END m00_r_data[8]
  PIN m00_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END m00_r_data[9]
  PIN m00_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 596.000 934.170 600.000 ;
    END
  END m00_r_id[0]
  PIN m00_r_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 510.040 2400.000 510.640 ;
    END
  END m00_r_id[10]
  PIN m00_r_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END m00_r_id[11]
  PIN m00_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 596.000 486.590 600.000 ;
    END
  END m00_r_id[1]
  PIN m00_r_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 596.000 1855.090 600.000 ;
    END
  END m00_r_id[2]
  PIN m00_r_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END m00_r_id[3]
  PIN m00_r_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 596.000 1723.070 600.000 ;
    END
  END m00_r_id[4]
  PIN m00_r_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 596.000 119.510 600.000 ;
    END
  END m00_r_id[5]
  PIN m00_r_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 596.000 1642.570 600.000 ;
    END
  END m00_r_id[6]
  PIN m00_r_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 596.000 1793.910 600.000 ;
    END
  END m00_r_id[7]
  PIN m00_r_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END m00_r_id[8]
  PIN m00_r_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END m00_r_id[9]
  PIN m00_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END m00_r_last
  PIN m00_r_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END m00_r_ready
  PIN m00_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END m00_r_resp[0]
  PIN m00_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.710 0.000 1999.990 4.000 ;
    END
  END m00_r_resp[1]
  PIN m00_r_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END m00_r_user[-1]
  PIN m00_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END m00_r_user[0]
  PIN m00_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 0.000 2396.050 4.000 ;
    END
  END m00_r_valid
  PIN m00_w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END m00_w_data[0]
  PIN m00_w_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 596.000 1961.350 600.000 ;
    END
  END m00_w_data[10]
  PIN m00_w_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.030 596.000 2341.310 600.000 ;
    END
  END m00_w_data[11]
  PIN m00_w_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END m00_w_data[12]
  PIN m00_w_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 596.000 203.230 600.000 ;
    END
  END m00_w_data[13]
  PIN m00_w_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END m00_w_data[14]
  PIN m00_w_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END m00_w_data[15]
  PIN m00_w_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END m00_w_data[16]
  PIN m00_w_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 596.000 1600.710 600.000 ;
    END
  END m00_w_data[17]
  PIN m00_w_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END m00_w_data[18]
  PIN m00_w_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 596.000 1806.790 600.000 ;
    END
  END m00_w_data[19]
  PIN m00_w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END m00_w_data[1]
  PIN m00_w_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END m00_w_data[20]
  PIN m00_w_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 0.000 2177.090 4.000 ;
    END
  END m00_w_data[21]
  PIN m00_w_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 596.000 367.450 600.000 ;
    END
  END m00_w_data[22]
  PIN m00_w_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END m00_w_data[23]
  PIN m00_w_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 0.040 2400.000 0.640 ;
    END
  END m00_w_data[24]
  PIN m00_w_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 377.440 2400.000 378.040 ;
    END
  END m00_w_data[25]
  PIN m00_w_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.370 596.000 2009.650 600.000 ;
    END
  END m00_w_data[26]
  PIN m00_w_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 595.040 2400.000 595.640 ;
    END
  END m00_w_data[27]
  PIN m00_w_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 596.000 1677.990 600.000 ;
    END
  END m00_w_data[28]
  PIN m00_w_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END m00_w_data[29]
  PIN m00_w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END m00_w_data[2]
  PIN m00_w_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END m00_w_data[30]
  PIN m00_w_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END m00_w_data[31]
  PIN m00_w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.170 596.000 1977.450 600.000 ;
    END
  END m00_w_data[3]
  PIN m00_w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 596.000 1542.750 600.000 ;
    END
  END m00_w_data[4]
  PIN m00_w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END m00_w_data[5]
  PIN m00_w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.410 596.000 2273.690 600.000 ;
    END
  END m00_w_data[6]
  PIN m00_w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END m00_w_data[7]
  PIN m00_w_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.350 596.000 2038.630 600.000 ;
    END
  END m00_w_data[8]
  PIN m00_w_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END m00_w_data[9]
  PIN m00_w_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 30.640 2400.000 31.240 ;
    END
  END m00_w_last
  PIN m00_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 540.640 2400.000 541.240 ;
    END
  END m00_w_ready
  PIN m00_w_strb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 353.640 2400.000 354.240 ;
    END
  END m00_w_strb[0]
  PIN m00_w_strb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 17.040 2400.000 17.640 ;
    END
  END m00_w_strb[1]
  PIN m00_w_strb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.670 0.000 2379.950 4.000 ;
    END
  END m00_w_strb[2]
  PIN m00_w_strb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 596.000 422.190 600.000 ;
    END
  END m00_w_strb[3]
  PIN m00_w_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 0.000 1797.130 4.000 ;
    END
  END m00_w_user[-1]
  PIN m00_w_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.670 596.000 2057.950 600.000 ;
    END
  END m00_w_user[0]
  PIN m00_w_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 596.000 776.390 600.000 ;
    END
  END m00_w_valid
  PIN m01_ar_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 596.000 1810.010 600.000 ;
    END
  END m01_ar_addr[0]
  PIN m01_ar_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END m01_ar_addr[10]
  PIN m01_ar_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END m01_ar_addr[11]
  PIN m01_ar_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 596.000 77.650 600.000 ;
    END
  END m01_ar_addr[12]
  PIN m01_ar_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.490 0.000 1996.770 4.000 ;
    END
  END m01_ar_addr[13]
  PIN m01_ar_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.130 0.000 2196.410 4.000 ;
    END
  END m01_ar_addr[14]
  PIN m01_ar_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END m01_ar_addr[15]
  PIN m01_ar_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.590 0.000 2334.870 4.000 ;
    END
  END m01_ar_addr[16]
  PIN m01_ar_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 596.000 670.130 600.000 ;
    END
  END m01_ar_addr[17]
  PIN m01_ar_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 4.000 ;
    END
  END m01_ar_addr[18]
  PIN m01_ar_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 596.000 2109.470 600.000 ;
    END
  END m01_ar_addr[19]
  PIN m01_ar_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END m01_ar_addr[1]
  PIN m01_ar_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.870 0.000 2251.150 4.000 ;
    END
  END m01_ar_addr[20]
  PIN m01_ar_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 596.000 2186.750 600.000 ;
    END
  END m01_ar_addr[21]
  PIN m01_ar_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 596.000 1800.350 600.000 ;
    END
  END m01_ar_addr[22]
  PIN m01_ar_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END m01_ar_addr[23]
  PIN m01_ar_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 596.000 1903.390 600.000 ;
    END
  END m01_ar_addr[24]
  PIN m01_ar_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END m01_ar_addr[25]
  PIN m01_ar_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END m01_ar_addr[26]
  PIN m01_ar_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 596.000 2183.530 600.000 ;
    END
  END m01_ar_addr[27]
  PIN m01_ar_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 596.000 1652.230 600.000 ;
    END
  END m01_ar_addr[28]
  PIN m01_ar_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.530 596.000 2260.810 600.000 ;
    END
  END m01_ar_addr[29]
  PIN m01_ar_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END m01_ar_addr[2]
  PIN m01_ar_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END m01_ar_addr[30]
  PIN m01_ar_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 0.000 1690.870 4.000 ;
    END
  END m01_ar_addr[31]
  PIN m01_ar_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 0.000 1745.610 4.000 ;
    END
  END m01_ar_addr[3]
  PIN m01_ar_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 596.000 261.190 600.000 ;
    END
  END m01_ar_addr[4]
  PIN m01_ar_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END m01_ar_addr[5]
  PIN m01_ar_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 596.000 1764.930 600.000 ;
    END
  END m01_ar_addr[6]
  PIN m01_ar_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END m01_ar_addr[7]
  PIN m01_ar_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 596.000 406.090 600.000 ;
    END
  END m01_ar_addr[8]
  PIN m01_ar_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END m01_ar_addr[9]
  PIN m01_ar_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END m01_ar_burst[0]
  PIN m01_ar_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 159.840 2400.000 160.440 ;
    END
  END m01_ar_burst[1]
  PIN m01_ar_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 596.000 1304.470 600.000 ;
    END
  END m01_ar_cache[0]
  PIN m01_ar_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 596.000 451.170 600.000 ;
    END
  END m01_ar_cache[1]
  PIN m01_ar_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END m01_ar_cache[2]
  PIN m01_ar_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 0.000 1706.970 4.000 ;
    END
  END m01_ar_cache[3]
  PIN m01_ar_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END m01_ar_id[0]
  PIN m01_ar_id[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 47.640 2400.000 48.240 ;
    END
  END m01_ar_id[10]
  PIN m01_ar_id[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 333.240 2400.000 333.840 ;
    END
  END m01_ar_id[11]
  PIN m01_ar_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END m01_ar_id[1]
  PIN m01_ar_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END m01_ar_id[2]
  PIN m01_ar_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 251.640 2400.000 252.240 ;
    END
  END m01_ar_id[3]
  PIN m01_ar_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2366.790 596.000 2367.070 600.000 ;
    END
  END m01_ar_id[4]
  PIN m01_ar_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 596.000 1349.550 600.000 ;
    END
  END m01_ar_id[5]
  PIN m01_ar_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 596.000 1880.850 600.000 ;
    END
  END m01_ar_id[6]
  PIN m01_ar_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END m01_ar_id[7]
  PIN m01_ar_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 0.000 2354.190 4.000 ;
    END
  END m01_ar_id[8]
  PIN m01_ar_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 0.000 2199.630 4.000 ;
    END
  END m01_ar_id[9]
  PIN m01_ar_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END m01_ar_len[0]
  PIN m01_ar_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 506.640 2400.000 507.240 ;
    END
  END m01_ar_len[1]
  PIN m01_ar_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END m01_ar_len[2]
  PIN m01_ar_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END m01_ar_len[3]
  PIN m01_ar_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.930 596.000 2325.210 600.000 ;
    END
  END m01_ar_len[4]
  PIN m01_ar_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 397.840 2400.000 398.440 ;
    END
  END m01_ar_len[5]
  PIN m01_ar_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END m01_ar_len[6]
  PIN m01_ar_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END m01_ar_len[7]
  PIN m01_ar_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END m01_ar_lock
  PIN m01_ar_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END m01_ar_prot[0]
  PIN m01_ar_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.670 0.000 1896.950 4.000 ;
    END
  END m01_ar_prot[1]
  PIN m01_ar_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END m01_ar_prot[2]
  PIN m01_ar_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END m01_ar_qos[0]
  PIN m01_ar_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END m01_ar_qos[1]
  PIN m01_ar_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 596.000 386.770 600.000 ;
    END
  END m01_ar_qos[2]
  PIN m01_ar_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 596.000 1062.970 600.000 ;
    END
  END m01_ar_qos[3]
  PIN m01_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 204.040 2400.000 204.640 ;
    END
  END m01_ar_ready
  PIN m01_ar_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 596.000 1768.150 600.000 ;
    END
  END m01_ar_region[0]
  PIN m01_ar_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 306.040 2400.000 306.640 ;
    END
  END m01_ar_region[1]
  PIN m01_ar_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 596.000 724.870 600.000 ;
    END
  END m01_ar_region[2]
  PIN m01_ar_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.270 596.000 1993.550 600.000 ;
    END
  END m01_ar_region[3]
  PIN m01_ar_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 596.000 644.370 600.000 ;
    END
  END m01_ar_size[0]
  PIN m01_ar_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 596.000 753.850 600.000 ;
    END
  END m01_ar_size[1]
  PIN m01_ar_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END m01_ar_size[2]
  PIN m01_ar_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.510 596.000 2128.790 600.000 ;
    END
  END m01_ar_user[-1]
  PIN m01_ar_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.410 0.000 2273.690 4.000 ;
    END
  END m01_ar_user[0]
  PIN m01_ar_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 596.000 1848.650 600.000 ;
    END
  END m01_ar_valid
  PIN m01_aw_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.430 596.000 2083.710 600.000 ;
    END
  END m01_aw_addr[0]
  PIN m01_aw_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 596.000 876.210 600.000 ;
    END
  END m01_aw_addr[10]
  PIN m01_aw_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 596.000 67.990 600.000 ;
    END
  END m01_aw_addr[11]
  PIN m01_aw_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END m01_aw_addr[12]
  PIN m01_aw_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END m01_aw_addr[13]
  PIN m01_aw_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.050 596.000 2151.330 600.000 ;
    END
  END m01_aw_addr[14]
  PIN m01_aw_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END m01_aw_addr[15]
  PIN m01_aw_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END m01_aw_addr[16]
  PIN m01_aw_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 596.000 109.850 600.000 ;
    END
  END m01_aw_addr[17]
  PIN m01_aw_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 596.000 1439.710 600.000 ;
    END
  END m01_aw_addr[18]
  PIN m01_aw_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 596.000 32.570 600.000 ;
    END
  END m01_aw_addr[19]
  PIN m01_aw_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END m01_aw_addr[1]
  PIN m01_aw_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.670 596.000 1896.950 600.000 ;
    END
  END m01_aw_addr[20]
  PIN m01_aw_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END m01_aw_addr[21]
  PIN m01_aw_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690 596.000 2350.970 600.000 ;
    END
  END m01_aw_addr[22]
  PIN m01_aw_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END m01_aw_addr[23]
  PIN m01_aw_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END m01_aw_addr[24]
  PIN m01_aw_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END m01_aw_addr[25]
  PIN m01_aw_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 578.040 2400.000 578.640 ;
    END
  END m01_aw_addr[26]
  PIN m01_aw_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END m01_aw_addr[27]
  PIN m01_aw_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END m01_aw_addr[28]
  PIN m01_aw_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 596.000 377.110 600.000 ;
    END
  END m01_aw_addr[29]
  PIN m01_aw_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.250 0.000 2022.530 4.000 ;
    END
  END m01_aw_addr[2]
  PIN m01_aw_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 596.000 138.830 600.000 ;
    END
  END m01_aw_addr[30]
  PIN m01_aw_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END m01_aw_addr[31]
  PIN m01_aw_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 0.000 1871.190 4.000 ;
    END
  END m01_aw_addr[3]
  PIN m01_aw_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END m01_aw_addr[4]
  PIN m01_aw_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END m01_aw_addr[5]
  PIN m01_aw_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 596.000 322.370 600.000 ;
    END
  END m01_aw_addr[6]
  PIN m01_aw_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END m01_aw_addr[7]
  PIN m01_aw_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 596.000 1909.830 600.000 ;
    END
  END m01_aw_addr[8]
  PIN m01_aw_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 596.000 493.030 600.000 ;
    END
  END m01_aw_addr[9]
  PIN m01_aw_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END m01_aw_burst[0]
  PIN m01_aw_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 193.840 2400.000 194.440 ;
    END
  END m01_aw_burst[1]
  PIN m01_aw_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 596.000 467.270 600.000 ;
    END
  END m01_aw_cache[0]
  PIN m01_aw_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END m01_aw_cache[1]
  PIN m01_aw_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.130 0.000 2357.410 4.000 ;
    END
  END m01_aw_cache[2]
  PIN m01_aw_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 0.000 1935.590 4.000 ;
    END
  END m01_aw_cache[3]
  PIN m01_aw_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END m01_aw_id[0]
  PIN m01_aw_id[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 482.840 2400.000 483.440 ;
    END
  END m01_aw_id[10]
  PIN m01_aw_id[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 596.000 357.790 600.000 ;
    END
  END m01_aw_id[11]
  PIN m01_aw_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 596.000 1610.370 600.000 ;
    END
  END m01_aw_id[1]
  PIN m01_aw_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 248.240 2400.000 248.840 ;
    END
  END m01_aw_id[2]
  PIN m01_aw_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END m01_aw_id[3]
  PIN m01_aw_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 596.000 1713.410 600.000 ;
    END
  END m01_aw_id[4]
  PIN m01_aw_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 596.000 1365.650 600.000 ;
    END
  END m01_aw_id[5]
  PIN m01_aw_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 596.000 216.110 600.000 ;
    END
  END m01_aw_id[6]
  PIN m01_aw_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 596.000 1690.870 600.000 ;
    END
  END m01_aw_id[7]
  PIN m01_aw_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 596.000 1639.350 600.000 ;
    END
  END m01_aw_id[8]
  PIN m01_aw_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 596.000 61.550 600.000 ;
    END
  END m01_aw_id[9]
  PIN m01_aw_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END m01_aw_len[0]
  PIN m01_aw_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.090 0.000 2254.370 4.000 ;
    END
  END m01_aw_len[1]
  PIN m01_aw_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 596.000 1732.730 600.000 ;
    END
  END m01_aw_len[2]
  PIN m01_aw_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 289.040 2400.000 289.640 ;
    END
  END m01_aw_len[3]
  PIN m01_aw_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.070 0.000 2283.350 4.000 ;
    END
  END m01_aw_len[4]
  PIN m01_aw_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END m01_aw_len[5]
  PIN m01_aw_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 596.000 676.570 600.000 ;
    END
  END m01_aw_len[6]
  PIN m01_aw_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 596.000 1545.970 600.000 ;
    END
  END m01_aw_len[7]
  PIN m01_aw_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 596.000 113.070 600.000 ;
    END
  END m01_aw_lock
  PIN m01_aw_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 596.000 1938.810 600.000 ;
    END
  END m01_aw_prot[0]
  PIN m01_aw_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 0.000 1858.310 4.000 ;
    END
  END m01_aw_prot[1]
  PIN m01_aw_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 596.000 2199.630 600.000 ;
    END
  END m01_aw_prot[2]
  PIN m01_aw_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.290 596.000 1964.570 600.000 ;
    END
  END m01_aw_qos[0]
  PIN m01_aw_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 596.000 1710.190 600.000 ;
    END
  END m01_aw_qos[1]
  PIN m01_aw_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END m01_aw_qos[2]
  PIN m01_aw_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END m01_aw_qos[3]
  PIN m01_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END m01_aw_ready
  PIN m01_aw_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END m01_aw_region[0]
  PIN m01_aw_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.990 596.000 2399.270 600.000 ;
    END
  END m01_aw_region[1]
  PIN m01_aw_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 596.000 399.650 600.000 ;
    END
  END m01_aw_region[2]
  PIN m01_aw_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 596.000 1156.350 600.000 ;
    END
  END m01_aw_region[3]
  PIN m01_aw_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 596.000 428.630 600.000 ;
    END
  END m01_aw_size[0]
  PIN m01_aw_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END m01_aw_size[1]
  PIN m01_aw_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 596.000 1117.710 600.000 ;
    END
  END m01_aw_size[2]
  PIN m01_aw_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.070 596.000 2283.350 600.000 ;
    END
  END m01_aw_user[-1]
  PIN m01_aw_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END m01_aw_user[0]
  PIN m01_aw_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END m01_aw_valid
  PIN m01_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END m01_b_id[0]
  PIN m01_b_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 547.440 2400.000 548.040 ;
    END
  END m01_b_id[10]
  PIN m01_b_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END m01_b_id[11]
  PIN m01_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END m01_b_id[1]
  PIN m01_b_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END m01_b_id[2]
  PIN m01_b_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END m01_b_id[3]
  PIN m01_b_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 596.000 866.550 600.000 ;
    END
  END m01_b_id[4]
  PIN m01_b_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 302.640 2400.000 303.240 ;
    END
  END m01_b_id[5]
  PIN m01_b_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 596.000 235.430 600.000 ;
    END
  END m01_b_id[6]
  PIN m01_b_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 596.000 969.590 600.000 ;
    END
  END m01_b_id[7]
  PIN m01_b_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END m01_b_id[8]
  PIN m01_b_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END m01_b_id[9]
  PIN m01_b_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 596.000 789.270 600.000 ;
    END
  END m01_b_ready
  PIN m01_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.550 0.000 2231.830 4.000 ;
    END
  END m01_b_resp[0]
  PIN m01_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END m01_b_resp[1]
  PIN m01_b_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.130 596.000 2035.410 600.000 ;
    END
  END m01_b_user[-1]
  PIN m01_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 596.000 209.670 600.000 ;
    END
  END m01_b_user[0]
  PIN m01_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.650 0.000 1925.930 4.000 ;
    END
  END m01_b_valid
  PIN m01_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END m01_r_data[0]
  PIN m01_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END m01_r_data[10]
  PIN m01_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 0.000 1507.330 4.000 ;
    END
  END m01_r_data[11]
  PIN m01_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 596.000 389.990 600.000 ;
    END
  END m01_r_data[12]
  PIN m01_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END m01_r_data[13]
  PIN m01_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END m01_r_data[14]
  PIN m01_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END m01_r_data[15]
  PIN m01_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 4.000 ;
    END
  END m01_r_data[16]
  PIN m01_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 596.000 1027.550 600.000 ;
    END
  END m01_r_data[17]
  PIN m01_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.930 0.000 2325.210 4.000 ;
    END
  END m01_r_data[18]
  PIN m01_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 596.000 525.230 600.000 ;
    END
  END m01_r_data[19]
  PIN m01_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 596.000 1958.130 600.000 ;
    END
  END m01_r_data[1]
  PIN m01_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 596.000 1539.530 600.000 ;
    END
  END m01_r_data[20]
  PIN m01_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 596.000 705.550 600.000 ;
    END
  END m01_r_data[21]
  PIN m01_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.030 0.000 2180.310 4.000 ;
    END
  END m01_r_data[22]
  PIN m01_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END m01_r_data[23]
  PIN m01_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 596.000 1201.430 600.000 ;
    END
  END m01_r_data[24]
  PIN m01_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.490 596.000 2318.770 600.000 ;
    END
  END m01_r_data[25]
  PIN m01_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 469.240 2400.000 469.840 ;
    END
  END m01_r_data[26]
  PIN m01_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 596.000 1890.510 600.000 ;
    END
  END m01_r_data[27]
  PIN m01_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END m01_r_data[28]
  PIN m01_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 596.000 2122.350 600.000 ;
    END
  END m01_r_data[29]
  PIN m01_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 596.000 1578.170 600.000 ;
    END
  END m01_r_data[2]
  PIN m01_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 596.000 1368.870 600.000 ;
    END
  END m01_r_data[30]
  PIN m01_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END m01_r_data[31]
  PIN m01_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 596.000 1359.210 600.000 ;
    END
  END m01_r_data[3]
  PIN m01_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 596.000 1185.330 600.000 ;
    END
  END m01_r_data[4]
  PIN m01_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 0.000 1365.650 4.000 ;
    END
  END m01_r_data[5]
  PIN m01_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 596.000 1861.530 600.000 ;
    END
  END m01_r_data[6]
  PIN m01_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END m01_r_data[7]
  PIN m01_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 596.000 1597.490 600.000 ;
    END
  END m01_r_data[8]
  PIN m01_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END m01_r_data[9]
  PIN m01_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 596.000 992.130 600.000 ;
    END
  END m01_r_id[0]
  PIN m01_r_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END m01_r_id[10]
  PIN m01_r_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 596.000 1748.830 600.000 ;
    END
  END m01_r_id[11]
  PIN m01_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END m01_r_id[1]
  PIN m01_r_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 596.000 924.510 600.000 ;
    END
  END m01_r_id[2]
  PIN m01_r_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.730 596.000 2132.010 600.000 ;
    END
  END m01_r_id[3]
  PIN m01_r_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.790 0.000 2206.070 4.000 ;
    END
  END m01_r_id[4]
  PIN m01_r_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END m01_r_id[5]
  PIN m01_r_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 596.000 361.010 600.000 ;
    END
  END m01_r_id[6]
  PIN m01_r_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END m01_r_id[7]
  PIN m01_r_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 513.440 2400.000 514.040 ;
    END
  END m01_r_id[8]
  PIN m01_r_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END m01_r_id[9]
  PIN m01_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 596.000 1098.390 600.000 ;
    END
  END m01_r_last
  PIN m01_r_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 0.000 1748.830 4.000 ;
    END
  END m01_r_ready
  PIN m01_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END m01_r_resp[0]
  PIN m01_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 596.000 125.950 600.000 ;
    END
  END m01_r_resp[1]
  PIN m01_r_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 591.640 2400.000 592.240 ;
    END
  END m01_r_user[-1]
  PIN m01_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END m01_r_user[0]
  PIN m01_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END m01_r_valid
  PIN m01_w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END m01_w_data[0]
  PIN m01_w_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END m01_w_data[10]
  PIN m01_w_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.470 596.000 2025.750 600.000 ;
    END
  END m01_w_data[11]
  PIN m01_w_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.570 596.000 2363.850 600.000 ;
    END
  END m01_w_data[12]
  PIN m01_w_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 596.000 306.270 600.000 ;
    END
  END m01_w_data[13]
  PIN m01_w_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 596.000 370.670 600.000 ;
    END
  END m01_w_data[14]
  PIN m01_w_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 596.000 882.650 600.000 ;
    END
  END m01_w_data[15]
  PIN m01_w_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 596.000 319.150 600.000 ;
    END
  END m01_w_data[16]
  PIN m01_w_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END m01_w_data[17]
  PIN m01_w_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END m01_w_data[18]
  PIN m01_w_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 596.000 2148.110 600.000 ;
    END
  END m01_w_data[19]
  PIN m01_w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 596.000 1394.630 600.000 ;
    END
  END m01_w_data[1]
  PIN m01_w_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 596.000 1230.410 600.000 ;
    END
  END m01_w_data[20]
  PIN m01_w_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END m01_w_data[21]
  PIN m01_w_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 596.000 148.490 600.000 ;
    END
  END m01_w_data[22]
  PIN m01_w_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 596.000 2048.290 600.000 ;
    END
  END m01_w_data[23]
  PIN m01_w_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 596.000 315.930 600.000 ;
    END
  END m01_w_data[24]
  PIN m01_w_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 596.000 1207.870 600.000 ;
    END
  END m01_w_data[25]
  PIN m01_w_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END m01_w_data[26]
  PIN m01_w_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END m01_w_data[27]
  PIN m01_w_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.450 596.000 2376.730 600.000 ;
    END
  END m01_w_data[28]
  PIN m01_w_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 448.840 2400.000 449.440 ;
    END
  END m01_w_data[29]
  PIN m01_w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 596.000 763.510 600.000 ;
    END
  END m01_w_data[2]
  PIN m01_w_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END m01_w_data[30]
  PIN m01_w_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END m01_w_data[31]
  PIN m01_w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END m01_w_data[3]
  PIN m01_w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 596.000 2099.810 600.000 ;
    END
  END m01_w_data[4]
  PIN m01_w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END m01_w_data[5]
  PIN m01_w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 596.000 818.250 600.000 ;
    END
  END m01_w_data[6]
  PIN m01_w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END m01_w_data[7]
  PIN m01_w_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 0.000 1913.050 4.000 ;
    END
  END m01_w_data[8]
  PIN m01_w_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 221.040 2400.000 221.640 ;
    END
  END m01_w_data[9]
  PIN m01_w_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END m01_w_last
  PIN m01_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 319.640 2400.000 320.240 ;
    END
  END m01_w_ready
  PIN m01_w_strb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END m01_w_strb[0]
  PIN m01_w_strb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END m01_w_strb[1]
  PIN m01_w_strb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 596.000 1987.110 600.000 ;
    END
  END m01_w_strb[2]
  PIN m01_w_strb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 596.000 1729.510 600.000 ;
    END
  END m01_w_strb[3]
  PIN m01_w_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 596.000 2354.190 600.000 ;
    END
  END m01_w_user[-1]
  PIN m01_w_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 596.000 663.690 600.000 ;
    END
  END m01_w_user[0]
  PIN m01_w_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 596.000 995.350 600.000 ;
    END
  END m01_w_valid
  PIN m02_ar_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END m02_ar_addr[0]
  PIN m02_ar_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.250 0.000 2344.530 4.000 ;
    END
  END m02_ar_addr[10]
  PIN m02_ar_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 596.000 1407.510 600.000 ;
    END
  END m02_ar_addr[11]
  PIN m02_ar_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 596.000 335.250 600.000 ;
    END
  END m02_ar_addr[12]
  PIN m02_ar_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 596.000 64.770 600.000 ;
    END
  END m02_ar_addr[13]
  PIN m02_ar_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END m02_ar_addr[14]
  PIN m02_ar_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 596.000 1745.610 600.000 ;
    END
  END m02_ar_addr[15]
  PIN m02_ar_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END m02_ar_addr[16]
  PIN m02_ar_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 132.640 2400.000 133.240 ;
    END
  END m02_ar_addr[17]
  PIN m02_ar_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.450 596.000 2215.730 600.000 ;
    END
  END m02_ar_addr[18]
  PIN m02_ar_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 596.000 573.530 600.000 ;
    END
  END m02_ar_addr[19]
  PIN m02_ar_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 596.000 380.330 600.000 ;
    END
  END m02_ar_addr[1]
  PIN m02_ar_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 292.440 2400.000 293.040 ;
    END
  END m02_ar_addr[20]
  PIN m02_ar_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.150 0.000 2167.430 4.000 ;
    END
  END m02_ar_addr[21]
  PIN m02_ar_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.950 0.000 2296.230 4.000 ;
    END
  END m02_ar_addr[22]
  PIN m02_ar_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 596.000 1095.170 600.000 ;
    END
  END m02_ar_addr[23]
  PIN m02_ar_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END m02_ar_addr[24]
  PIN m02_ar_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 596.000 87.310 600.000 ;
    END
  END m02_ar_addr[25]
  PIN m02_ar_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 596.000 1922.710 600.000 ;
    END
  END m02_ar_addr[26]
  PIN m02_ar_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END m02_ar_addr[27]
  PIN m02_ar_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 596.000 338.470 600.000 ;
    END
  END m02_ar_addr[28]
  PIN m02_ar_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 0.000 1903.390 4.000 ;
    END
  END m02_ar_addr[29]
  PIN m02_ar_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 596.000 1797.130 600.000 ;
    END
  END m02_ar_addr[2]
  PIN m02_ar_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END m02_ar_addr[30]
  PIN m02_ar_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END m02_ar_addr[31]
  PIN m02_ar_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 596.000 1182.110 600.000 ;
    END
  END m02_ar_addr[3]
  PIN m02_ar_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END m02_ar_addr[4]
  PIN m02_ar_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 0.000 1723.070 4.000 ;
    END
  END m02_ar_addr[5]
  PIN m02_ar_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 596.000 702.330 600.000 ;
    END
  END m02_ar_addr[6]
  PIN m02_ar_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END m02_ar_addr[7]
  PIN m02_ar_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END m02_ar_addr[8]
  PIN m02_ar_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 596.000 1478.350 600.000 ;
    END
  END m02_ar_addr[9]
  PIN m02_ar_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 596.000 1059.750 600.000 ;
    END
  END m02_ar_burst[0]
  PIN m02_ar_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END m02_ar_burst[1]
  PIN m02_ar_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.970 596.000 1784.250 600.000 ;
    END
  END m02_ar_cache[0]
  PIN m02_ar_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.790 596.000 1884.070 600.000 ;
    END
  END m02_ar_cache[1]
  PIN m02_ar_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 596.000 187.130 600.000 ;
    END
  END m02_ar_cache[2]
  PIN m02_ar_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.950 596.000 2296.230 600.000 ;
    END
  END m02_ar_cache[3]
  PIN m02_ar_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END m02_ar_id[0]
  PIN m02_ar_id[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END m02_ar_id[10]
  PIN m02_ar_id[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 596.000 1526.650 600.000 ;
    END
  END m02_ar_id[11]
  PIN m02_ar_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END m02_ar_id[1]
  PIN m02_ar_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END m02_ar_id[2]
  PIN m02_ar_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 596.000 885.870 600.000 ;
    END
  END m02_ar_id[3]
  PIN m02_ar_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END m02_ar_id[4]
  PIN m02_ar_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END m02_ar_id[5]
  PIN m02_ar_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 596.000 976.030 600.000 ;
    END
  END m02_ar_id[6]
  PIN m02_ar_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 596.000 1954.910 600.000 ;
    END
  END m02_ar_id[7]
  PIN m02_ar_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END m02_ar_id[8]
  PIN m02_ar_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 596.000 1510.550 600.000 ;
    END
  END m02_ar_id[9]
  PIN m02_ar_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 596.000 106.630 600.000 ;
    END
  END m02_ar_len[0]
  PIN m02_ar_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END m02_ar_len[1]
  PIN m02_ar_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END m02_ar_len[2]
  PIN m02_ar_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END m02_ar_len[3]
  PIN m02_ar_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END m02_ar_len[4]
  PIN m02_ar_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 596.000 476.930 600.000 ;
    END
  END m02_ar_len[5]
  PIN m02_ar_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END m02_ar_len[6]
  PIN m02_ar_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 0.000 2115.910 4.000 ;
    END
  END m02_ar_len[7]
  PIN m02_ar_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 0.000 2138.450 4.000 ;
    END
  END m02_ar_lock
  PIN m02_ar_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 74.840 2400.000 75.440 ;
    END
  END m02_ar_prot[0]
  PIN m02_ar_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 596.000 2218.950 600.000 ;
    END
  END m02_ar_prot[1]
  PIN m02_ar_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 596.000 596.070 600.000 ;
    END
  END m02_ar_prot[2]
  PIN m02_ar_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.550 596.000 1587.830 600.000 ;
    END
  END m02_ar_qos[0]
  PIN m02_ar_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.690 0.000 2028.970 4.000 ;
    END
  END m02_ar_qos[1]
  PIN m02_ar_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END m02_ar_qos[2]
  PIN m02_ar_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END m02_ar_qos[3]
  PIN m02_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 596.000 1375.310 600.000 ;
    END
  END m02_ar_ready
  PIN m02_ar_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END m02_ar_region[0]
  PIN m02_ar_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END m02_ar_region[1]
  PIN m02_ar_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 596.000 834.350 600.000 ;
    END
  END m02_ar_region[2]
  PIN m02_ar_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 596.000 2241.490 600.000 ;
    END
  END m02_ar_region[3]
  PIN m02_ar_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.550 0.000 1587.830 4.000 ;
    END
  END m02_ar_size[0]
  PIN m02_ar_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END m02_ar_size[1]
  PIN m02_ar_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END m02_ar_size[2]
  PIN m02_ar_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 596.000 718.430 600.000 ;
    END
  END m02_ar_user[-1]
  PIN m02_ar_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END m02_ar_user[0]
  PIN m02_ar_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END m02_ar_valid
  PIN m02_aw_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.770 0.000 2235.050 4.000 ;
    END
  END m02_aw_addr[0]
  PIN m02_aw_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 418.240 2400.000 418.840 ;
    END
  END m02_aw_addr[10]
  PIN m02_aw_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 596.000 232.210 600.000 ;
    END
  END m02_aw_addr[11]
  PIN m02_aw_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 238.040 2400.000 238.640 ;
    END
  END m02_aw_addr[12]
  PIN m02_aw_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END m02_aw_addr[13]
  PIN m02_aw_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 596.000 599.290 600.000 ;
    END
  END m02_aw_addr[14]
  PIN m02_aw_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.350 0.000 2360.630 4.000 ;
    END
  END m02_aw_addr[15]
  PIN m02_aw_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 596.000 1475.130 600.000 ;
    END
  END m02_aw_addr[16]
  PIN m02_aw_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 596.000 200.010 600.000 ;
    END
  END m02_aw_addr[17]
  PIN m02_aw_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.470 0.000 2347.750 4.000 ;
    END
  END m02_aw_addr[18]
  PIN m02_aw_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 0.000 2086.930 4.000 ;
    END
  END m02_aw_addr[19]
  PIN m02_aw_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 596.000 1056.530 600.000 ;
    END
  END m02_aw_addr[1]
  PIN m02_aw_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 596.000 10.030 600.000 ;
    END
  END m02_aw_addr[20]
  PIN m02_aw_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END m02_aw_addr[21]
  PIN m02_aw_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 596.000 740.970 600.000 ;
    END
  END m02_aw_addr[22]
  PIN m02_aw_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 596.000 312.710 600.000 ;
    END
  END m02_aw_addr[23]
  PIN m02_aw_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 71.440 2400.000 72.040 ;
    END
  END m02_aw_addr[24]
  PIN m02_aw_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 428.440 2400.000 429.040 ;
    END
  END m02_aw_addr[25]
  PIN m02_aw_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 596.000 1700.530 600.000 ;
    END
  END m02_aw_addr[26]
  PIN m02_aw_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 227.840 2400.000 228.440 ;
    END
  END m02_aw_addr[27]
  PIN m02_aw_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 596.000 686.230 600.000 ;
    END
  END m02_aw_addr[28]
  PIN m02_aw_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.130 596.000 2357.410 600.000 ;
    END
  END m02_aw_addr[29]
  PIN m02_aw_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.770 0.000 2074.050 4.000 ;
    END
  END m02_aw_addr[2]
  PIN m02_aw_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END m02_aw_addr[30]
  PIN m02_aw_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END m02_aw_addr[31]
  PIN m02_aw_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 596.000 1269.050 600.000 ;
    END
  END m02_aw_addr[3]
  PIN m02_aw_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 596.000 1043.650 600.000 ;
    END
  END m02_aw_addr[4]
  PIN m02_aw_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END m02_aw_addr[5]
  PIN m02_aw_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 596.000 1735.950 600.000 ;
    END
  END m02_aw_addr[6]
  PIN m02_aw_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 596.000 174.250 600.000 ;
    END
  END m02_aw_addr[7]
  PIN m02_aw_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END m02_aw_addr[8]
  PIN m02_aw_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.090 596.000 2093.370 600.000 ;
    END
  END m02_aw_addr[9]
  PIN m02_aw_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 27.240 2400.000 27.840 ;
    END
  END m02_aw_burst[0]
  PIN m02_aw_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 0.000 1810.010 4.000 ;
    END
  END m02_aw_burst[1]
  PIN m02_aw_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END m02_aw_cache[0]
  PIN m02_aw_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.150 0.000 2006.430 4.000 ;
    END
  END m02_aw_cache[1]
  PIN m02_aw_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 476.040 2400.000 476.640 ;
    END
  END m02_aw_cache[2]
  PIN m02_aw_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.350 0.000 1877.630 4.000 ;
    END
  END m02_aw_cache[3]
  PIN m02_aw_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END m02_aw_id[0]
  PIN m02_aw_id[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END m02_aw_id[10]
  PIN m02_aw_id[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 596.000 1169.230 600.000 ;
    END
  END m02_aw_id[11]
  PIN m02_aw_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END m02_aw_id[1]
  PIN m02_aw_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.690 596.000 2028.970 600.000 ;
    END
  END m02_aw_id[2]
  PIN m02_aw_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 596.000 1687.650 600.000 ;
    END
  END m02_aw_id[3]
  PIN m02_aw_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END m02_aw_id[4]
  PIN m02_aw_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 596.000 795.710 600.000 ;
    END
  END m02_aw_id[5]
  PIN m02_aw_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 596.000 364.230 600.000 ;
    END
  END m02_aw_id[6]
  PIN m02_aw_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END m02_aw_id[7]
  PIN m02_aw_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END m02_aw_id[8]
  PIN m02_aw_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 596.000 277.290 600.000 ;
    END
  END m02_aw_id[9]
  PIN m02_aw_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END m02_aw_len[0]
  PIN m02_aw_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END m02_aw_len[1]
  PIN m02_aw_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 596.000 1140.250 600.000 ;
    END
  END m02_aw_len[2]
  PIN m02_aw_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END m02_aw_len[3]
  PIN m02_aw_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 596.000 1471.910 600.000 ;
    END
  END m02_aw_len[4]
  PIN m02_aw_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 596.000 22.910 600.000 ;
    END
  END m02_aw_len[5]
  PIN m02_aw_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 0.000 1958.130 4.000 ;
    END
  END m02_aw_len[6]
  PIN m02_aw_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END m02_aw_len[7]
  PIN m02_aw_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 207.440 2400.000 208.040 ;
    END
  END m02_aw_lock
  PIN m02_aw_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 596.000 943.830 600.000 ;
    END
  END m02_aw_prot[0]
  PIN m02_aw_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 596.000 953.490 600.000 ;
    END
  END m02_aw_prot[1]
  PIN m02_aw_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END m02_aw_prot[2]
  PIN m02_aw_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END m02_aw_qos[0]
  PIN m02_aw_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 596.000 972.810 600.000 ;
    END
  END m02_aw_qos[1]
  PIN m02_aw_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 554.240 2400.000 554.840 ;
    END
  END m02_aw_qos[2]
  PIN m02_aw_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 4.000 ;
    END
  END m02_aw_qos[3]
  PIN m02_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.350 596.000 2360.630 600.000 ;
    END
  END m02_aw_ready
  PIN m02_aw_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 431.840 2400.000 432.440 ;
    END
  END m02_aw_region[0]
  PIN m02_aw_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.430 0.000 2083.710 4.000 ;
    END
  END m02_aw_region[1]
  PIN m02_aw_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.530 0.000 2260.810 4.000 ;
    END
  END m02_aw_region[2]
  PIN m02_aw_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 596.000 811.810 600.000 ;
    END
  END m02_aw_region[3]
  PIN m02_aw_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 596.000 824.690 600.000 ;
    END
  END m02_aw_size[0]
  PIN m02_aw_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 596.000 1053.310 600.000 ;
    END
  END m02_aw_size[1]
  PIN m02_aw_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END m02_aw_size[2]
  PIN m02_aw_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END m02_aw_user[-1]
  PIN m02_aw_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END m02_aw_user[0]
  PIN m02_aw_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.990 596.000 2238.270 600.000 ;
    END
  END m02_aw_valid
  PIN m02_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 596.000 1661.890 600.000 ;
    END
  END m02_b_id[0]
  PIN m02_b_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 596.000 158.150 600.000 ;
    END
  END m02_b_id[10]
  PIN m02_b_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 596.000 1104.830 600.000 ;
    END
  END m02_b_id[11]
  PIN m02_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END m02_b_id[1]
  PIN m02_b_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END m02_b_id[2]
  PIN m02_b_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 596.000 1449.370 600.000 ;
    END
  END m02_b_id[3]
  PIN m02_b_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 596.000 251.530 600.000 ;
    END
  END m02_b_id[4]
  PIN m02_b_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 596.000 1558.850 600.000 ;
    END
  END m02_b_id[5]
  PIN m02_b_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 374.040 2400.000 374.640 ;
    END
  END m02_b_id[6]
  PIN m02_b_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 0.000 1842.210 4.000 ;
    END
  END m02_b_id[7]
  PIN m02_b_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 596.000 1137.030 600.000 ;
    END
  END m02_b_id[8]
  PIN m02_b_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.630 596.000 2276.910 600.000 ;
    END
  END m02_b_id[9]
  PIN m02_b_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.450 0.000 2215.730 4.000 ;
    END
  END m02_b_ready
  PIN m02_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END m02_b_resp[0]
  PIN m02_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.170 0.000 2299.450 4.000 ;
    END
  END m02_b_resp[1]
  PIN m02_b_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 596.000 1220.750 600.000 ;
    END
  END m02_b_user[-1]
  PIN m02_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 596.000 171.030 600.000 ;
    END
  END m02_b_user[0]
  PIN m02_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 596.000 798.930 600.000 ;
    END
  END m02_b_valid
  PIN m02_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END m02_r_data[0]
  PIN m02_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END m02_r_data[10]
  PIN m02_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 197.240 2400.000 197.840 ;
    END
  END m02_r_data[11]
  PIN m02_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 596.000 2247.930 600.000 ;
    END
  END m02_r_data[12]
  PIN m02_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 0.000 1893.730 4.000 ;
    END
  END m02_r_data[13]
  PIN m02_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END m02_r_data[14]
  PIN m02_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END m02_r_data[15]
  PIN m02_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 596.000 51.890 600.000 ;
    END
  END m02_r_data[16]
  PIN m02_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 4.000 ;
    END
  END m02_r_data[17]
  PIN m02_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END m02_r_data[18]
  PIN m02_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 596.000 2070.830 600.000 ;
    END
  END m02_r_data[19]
  PIN m02_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END m02_r_data[1]
  PIN m02_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.250 596.000 2022.530 600.000 ;
    END
  END m02_r_data[20]
  PIN m02_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.950 596.000 1974.230 600.000 ;
    END
  END m02_r_data[21]
  PIN m02_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 596.000 1175.670 600.000 ;
    END
  END m02_r_data[22]
  PIN m02_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 596.000 1301.250 600.000 ;
    END
  END m02_r_data[23]
  PIN m02_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 142.840 2400.000 143.440 ;
    END
  END m02_r_data[24]
  PIN m02_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 596.000 557.430 600.000 ;
    END
  END m02_r_data[25]
  PIN m02_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END m02_r_data[26]
  PIN m02_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 596.000 293.390 600.000 ;
    END
  END m02_r_data[27]
  PIN m02_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.610 0.000 2144.890 4.000 ;
    END
  END m02_r_data[28]
  PIN m02_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 596.000 1694.090 600.000 ;
    END
  END m02_r_data[29]
  PIN m02_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 596.000 1101.610 600.000 ;
    END
  END m02_r_data[2]
  PIN m02_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 596.000 1223.970 600.000 ;
    END
  END m02_r_data[30]
  PIN m02_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END m02_r_data[31]
  PIN m02_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END m02_r_data[3]
  PIN m02_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END m02_r_data[4]
  PIN m02_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END m02_r_data[5]
  PIN m02_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END m02_r_data[6]
  PIN m02_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END m02_r_data[7]
  PIN m02_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END m02_r_data[8]
  PIN m02_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 0.000 1246.510 4.000 ;
    END
  END m02_r_data[9]
  PIN m02_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END m02_r_id[0]
  PIN m02_r_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 0.000 1764.930 4.000 ;
    END
  END m02_r_id[10]
  PIN m02_r_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END m02_r_id[11]
  PIN m02_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END m02_r_id[1]
  PIN m02_r_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END m02_r_id[2]
  PIN m02_r_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END m02_r_id[3]
  PIN m02_r_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 0.000 1900.170 4.000 ;
    END
  END m02_r_id[4]
  PIN m02_r_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 285.640 2400.000 286.240 ;
    END
  END m02_r_id[5]
  PIN m02_r_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 596.000 1194.990 600.000 ;
    END
  END m02_r_id[6]
  PIN m02_r_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END m02_r_id[7]
  PIN m02_r_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 596.000 544.550 600.000 ;
    END
  END m02_r_id[8]
  PIN m02_r_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END m02_r_id[9]
  PIN m02_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 596.000 425.410 600.000 ;
    END
  END m02_r_last
  PIN m02_r_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 176.840 2400.000 177.440 ;
    END
  END m02_r_ready
  PIN m02_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END m02_r_resp[0]
  PIN m02_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END m02_r_resp[1]
  PIN m02_r_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END m02_r_user[-1]
  PIN m02_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END m02_r_user[0]
  PIN m02_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END m02_r_valid
  PIN m02_w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 596.000 1259.390 600.000 ;
    END
  END m02_w_data[0]
  PIN m02_w_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END m02_w_data[10]
  PIN m02_w_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END m02_w_data[11]
  PIN m02_w_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END m02_w_data[12]
  PIN m02_w_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 596.000 1565.290 600.000 ;
    END
  END m02_w_data[13]
  PIN m02_w_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END m02_w_data[14]
  PIN m02_w_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END m02_w_data[15]
  PIN m02_w_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 0.000 1542.750 4.000 ;
    END
  END m02_w_data[16]
  PIN m02_w_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 596.000 286.950 600.000 ;
    END
  END m02_w_data[17]
  PIN m02_w_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END m02_w_data[18]
  PIN m02_w_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END m02_w_data[19]
  PIN m02_w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 596.000 589.630 600.000 ;
    END
  END m02_w_data[1]
  PIN m02_w_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 596.000 1581.390 600.000 ;
    END
  END m02_w_data[20]
  PIN m02_w_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.050 0.000 2151.330 4.000 ;
    END
  END m02_w_data[21]
  PIN m02_w_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 596.000 135.610 600.000 ;
    END
  END m02_w_data[22]
  PIN m02_w_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.790 596.000 2206.070 600.000 ;
    END
  END m02_w_data[23]
  PIN m02_w_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END m02_w_data[24]
  PIN m02_w_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END m02_w_data[25]
  PIN m02_w_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 115.640 2400.000 116.240 ;
    END
  END m02_w_data[26]
  PIN m02_w_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 596.000 71.210 600.000 ;
    END
  END m02_w_data[27]
  PIN m02_w_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 596.000 470.490 600.000 ;
    END
  END m02_w_data[28]
  PIN m02_w_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 156.440 2400.000 157.040 ;
    END
  END m02_w_data[29]
  PIN m02_w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END m02_w_data[2]
  PIN m02_w_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 0.000 1710.190 4.000 ;
    END
  END m02_w_data[30]
  PIN m02_w_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 0.000 2293.010 4.000 ;
    END
  END m02_w_data[31]
  PIN m02_w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END m02_w_data[3]
  PIN m02_w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END m02_w_data[4]
  PIN m02_w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END m02_w_data[5]
  PIN m02_w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 596.000 505.910 600.000 ;
    END
  END m02_w_data[6]
  PIN m02_w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.590 0.000 2173.870 4.000 ;
    END
  END m02_w_data[7]
  PIN m02_w_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END m02_w_data[8]
  PIN m02_w_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 0.000 1713.410 4.000 ;
    END
  END m02_w_data[9]
  PIN m02_w_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 3.440 2400.000 4.040 ;
    END
  END m02_w_last
  PIN m02_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END m02_w_ready
  PIN m02_w_strb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 0.000 2241.490 4.000 ;
    END
  END m02_w_strb[0]
  PIN m02_w_strb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 596.000 344.910 600.000 ;
    END
  END m02_w_strb[1]
  PIN m02_w_strb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 596.000 2119.130 600.000 ;
    END
  END m02_w_strb[2]
  PIN m02_w_strb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END m02_w_strb[3]
  PIN m02_w_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END m02_w_user[-1]
  PIN m02_w_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 537.240 2400.000 537.840 ;
    END
  END m02_w_user[0]
  PIN m02_w_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 596.000 1114.490 600.000 ;
    END
  END m02_w_valid
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END rst_n
  PIN s00_ar_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 596.000 29.350 600.000 ;
    END
  END s00_ar_addr[0]
  PIN s00_ar_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 596.000 2257.590 600.000 ;
    END
  END s00_ar_addr[10]
  PIN s00_ar_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 596.000 1413.950 600.000 ;
    END
  END s00_ar_addr[11]
  PIN s00_ar_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 596.000 1252.950 600.000 ;
    END
  END s00_ar_addr[12]
  PIN s00_ar_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.330 0.000 1906.610 4.000 ;
    END
  END s00_ar_addr[13]
  PIN s00_ar_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END s00_ar_addr[14]
  PIN s00_ar_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 596.000 2270.470 600.000 ;
    END
  END s00_ar_addr[15]
  PIN s00_ar_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END s00_ar_addr[16]
  PIN s00_ar_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END s00_ar_addr[17]
  PIN s00_ar_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 596.000 1281.930 600.000 ;
    END
  END s00_ar_addr[18]
  PIN s00_ar_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.770 596.000 2235.050 600.000 ;
    END
  END s00_ar_addr[19]
  PIN s00_ar_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END s00_ar_addr[1]
  PIN s00_ar_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 98.640 2400.000 99.240 ;
    END
  END s00_ar_addr[20]
  PIN s00_ar_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 596.000 747.410 600.000 ;
    END
  END s00_ar_addr[21]
  PIN s00_ar_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END s00_ar_addr[22]
  PIN s00_ar_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.310 0.000 2096.590 4.000 ;
    END
  END s00_ar_addr[23]
  PIN s00_ar_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 214.240 2400.000 214.840 ;
    END
  END s00_ar_addr[24]
  PIN s00_ar_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 596.000 1333.450 600.000 ;
    END
  END s00_ar_addr[25]
  PIN s00_ar_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END s00_ar_addr[26]
  PIN s00_ar_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.470 0.000 2025.750 4.000 ;
    END
  END s00_ar_addr[27]
  PIN s00_ar_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END s00_ar_addr[28]
  PIN s00_ar_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END s00_ar_addr[29]
  PIN s00_ar_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 4.000 ;
    END
  END s00_ar_addr[2]
  PIN s00_ar_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 596.000 515.570 600.000 ;
    END
  END s00_ar_addr[30]
  PIN s00_ar_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END s00_ar_addr[31]
  PIN s00_ar_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END s00_ar_addr[3]
  PIN s00_ar_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END s00_ar_addr[4]
  PIN s00_ar_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END s00_ar_addr[5]
  PIN s00_ar_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.510 596.000 1967.790 600.000 ;
    END
  END s00_ar_addr[6]
  PIN s00_ar_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END s00_ar_addr[7]
  PIN s00_ar_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END s00_ar_addr[8]
  PIN s00_ar_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 596.000 660.470 600.000 ;
    END
  END s00_ar_addr[9]
  PIN s00_ar_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 596.000 348.130 600.000 ;
    END
  END s00_ar_burst[0]
  PIN s00_ar_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END s00_ar_burst[1]
  PIN s00_ar_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 472.640 2400.000 473.240 ;
    END
  END s00_ar_cache[0]
  PIN s00_ar_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 596.000 1204.650 600.000 ;
    END
  END s00_ar_cache[1]
  PIN s00_ar_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.810 596.000 2338.090 600.000 ;
    END
  END s00_ar_cache[2]
  PIN s00_ar_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 596.000 431.850 600.000 ;
    END
  END s00_ar_cache[3]
  PIN s00_ar_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 596.000 1813.230 600.000 ;
    END
  END s00_ar_id[0]
  PIN s00_ar_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 0.000 1983.890 4.000 ;
    END
  END s00_ar_id[1]
  PIN s00_ar_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.890 596.000 2383.170 600.000 ;
    END
  END s00_ar_id[2]
  PIN s00_ar_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 217.640 2400.000 218.240 ;
    END
  END s00_ar_id[3]
  PIN s00_ar_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END s00_ar_id[4]
  PIN s00_ar_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 187.040 2400.000 187.640 ;
    END
  END s00_ar_id[5]
  PIN s00_ar_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 596.000 518.790 600.000 ;
    END
  END s00_ar_id[6]
  PIN s00_ar_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END s00_ar_id[7]
  PIN s00_ar_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 596.000 2086.930 600.000 ;
    END
  END s00_ar_id[8]
  PIN s00_ar_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 0.000 1832.550 4.000 ;
    END
  END s00_ar_id[9]
  PIN s00_ar_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 596.000 911.630 600.000 ;
    END
  END s00_ar_len[0]
  PIN s00_ar_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.370 0.000 2170.650 4.000 ;
    END
  END s00_ar_len[1]
  PIN s00_ar_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END s00_ar_len[2]
  PIN s00_ar_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 596.000 154.930 600.000 ;
    END
  END s00_ar_len[3]
  PIN s00_ar_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.250 596.000 2344.530 600.000 ;
    END
  END s00_ar_len[4]
  PIN s00_ar_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 596.000 1162.790 600.000 ;
    END
  END s00_ar_len[5]
  PIN s00_ar_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 0.000 1887.290 4.000 ;
    END
  END s00_ar_len[6]
  PIN s00_ar_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 596.000 2103.030 600.000 ;
    END
  END s00_ar_len[7]
  PIN s00_ar_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END s00_ar_lock
  PIN s00_ar_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 596.000 1681.210 600.000 ;
    END
  END s00_ar_prot[0]
  PIN s00_ar_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 0.000 2080.490 4.000 ;
    END
  END s00_ar_prot[1]
  PIN s00_ar_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.870 596.000 2090.150 600.000 ;
    END
  END s00_ar_prot[2]
  PIN s00_ar_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END s00_ar_qos[0]
  PIN s00_ar_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.930 0.000 2003.210 4.000 ;
    END
  END s00_ar_qos[1]
  PIN s00_ar_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END s00_ar_qos[2]
  PIN s00_ar_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 596.000 715.210 600.000 ;
    END
  END s00_ar_qos[3]
  PIN s00_ar_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 0.000 2148.110 4.000 ;
    END
  END s00_ar_ready
  PIN s00_ar_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END s00_ar_region[0]
  PIN s00_ar_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 421.640 2400.000 422.240 ;
    END
  END s00_ar_region[1]
  PIN s00_ar_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 0.000 1639.350 4.000 ;
    END
  END s00_ar_region[2]
  PIN s00_ar_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 596.000 2019.310 600.000 ;
    END
  END s00_ar_region[3]
  PIN s00_ar_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.830 596.000 2309.110 600.000 ;
    END
  END s00_ar_size[0]
  PIN s00_ar_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.450 0.000 2054.730 4.000 ;
    END
  END s00_ar_size[1]
  PIN s00_ar_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END s00_ar_size[2]
  PIN s00_ar_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 596.000 892.310 600.000 ;
    END
  END s00_ar_user[-1]
  PIN s00_ar_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END s00_ar_user[0]
  PIN s00_ar_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END s00_ar_valid
  PIN s00_aw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 557.640 2400.000 558.240 ;
    END
  END s00_aw_addr[0]
  PIN s00_aw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 596.000 1188.550 600.000 ;
    END
  END s00_aw_addr[10]
  PIN s00_aw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 596.000 744.190 600.000 ;
    END
  END s00_aw_addr[11]
  PIN s00_aw_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 596.000 1433.270 600.000 ;
    END
  END s00_aw_addr[12]
  PIN s00_aw_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 596.000 193.570 600.000 ;
    END
  END s00_aw_addr[13]
  PIN s00_aw_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END s00_aw_addr[14]
  PIN s00_aw_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.930 0.000 2164.210 4.000 ;
    END
  END s00_aw_addr[15]
  PIN s00_aw_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 596.000 283.730 600.000 ;
    END
  END s00_aw_addr[16]
  PIN s00_aw_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 4.000 ;
    END
  END s00_aw_addr[17]
  PIN s00_aw_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END s00_aw_addr[18]
  PIN s00_aw_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END s00_aw_addr[19]
  PIN s00_aw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 596.000 460.830 600.000 ;
    END
  END s00_aw_addr[1]
  PIN s00_aw_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END s00_aw_addr[20]
  PIN s00_aw_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END s00_aw_addr[21]
  PIN s00_aw_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 170.040 2400.000 170.640 ;
    END
  END s00_aw_addr[22]
  PIN s00_aw_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 596.000 1871.190 600.000 ;
    END
  END s00_aw_addr[23]
  PIN s00_aw_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END s00_aw_addr[24]
  PIN s00_aw_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 4.000 ;
    END
  END s00_aw_addr[25]
  PIN s00_aw_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 596.000 435.070 600.000 ;
    END
  END s00_aw_addr[26]
  PIN s00_aw_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 596.000 782.830 600.000 ;
    END
  END s00_aw_addr[27]
  PIN s00_aw_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.890 596.000 2061.170 600.000 ;
    END
  END s00_aw_addr[28]
  PIN s00_aw_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 596.000 1008.230 600.000 ;
    END
  END s00_aw_addr[29]
  PIN s00_aw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END s00_aw_addr[2]
  PIN s00_aw_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 596.000 1645.790 600.000 ;
    END
  END s00_aw_addr[30]
  PIN s00_aw_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END s00_aw_addr[31]
  PIN s00_aw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 596.000 560.650 600.000 ;
    END
  END s00_aw_addr[3]
  PIN s00_aw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 596.000 1706.970 600.000 ;
    END
  END s00_aw_addr[4]
  PIN s00_aw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 596.000 1120.930 600.000 ;
    END
  END s00_aw_addr[5]
  PIN s00_aw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END s00_aw_addr[6]
  PIN s00_aw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END s00_aw_addr[7]
  PIN s00_aw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END s00_aw_addr[8]
  PIN s00_aw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 200.640 2400.000 201.240 ;
    END
  END s00_aw_addr[9]
  PIN s00_aw_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END s00_aw_burst[0]
  PIN s00_aw_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END s00_aw_burst[1]
  PIN s00_aw_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 596.000 766.730 600.000 ;
    END
  END s00_aw_cache[0]
  PIN s00_aw_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END s00_aw_cache[1]
  PIN s00_aw_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END s00_aw_cache[2]
  PIN s00_aw_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 596.000 1835.770 600.000 ;
    END
  END s00_aw_cache[3]
  PIN s00_aw_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 596.000 602.510 600.000 ;
    END
  END s00_aw_id[0]
  PIN s00_aw_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 0.000 2112.690 4.000 ;
    END
  END s00_aw_id[1]
  PIN s00_aw_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END s00_aw_id[2]
  PIN s00_aw_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 0.000 1919.490 4.000 ;
    END
  END s00_aw_id[3]
  PIN s00_aw_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.630 0.000 2276.910 4.000 ;
    END
  END s00_aw_id[4]
  PIN s00_aw_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 163.240 2400.000 163.840 ;
    END
  END s00_aw_id[5]
  PIN s00_aw_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 0.000 1793.910 4.000 ;
    END
  END s00_aw_id[6]
  PIN s00_aw_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 596.000 48.670 600.000 ;
    END
  END s00_aw_id[7]
  PIN s00_aw_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 596.000 654.030 600.000 ;
    END
  END s00_aw_id[8]
  PIN s00_aw_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END s00_aw_id[9]
  PIN s00_aw_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 596.000 586.410 600.000 ;
    END
  END s00_aw_len[0]
  PIN s00_aw_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.390 0.000 2302.670 4.000 ;
    END
  END s00_aw_len[1]
  PIN s00_aw_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END s00_aw_len[2]
  PIN s00_aw_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 596.000 351.350 600.000 ;
    END
  END s00_aw_len[3]
  PIN s00_aw_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END s00_aw_len[4]
  PIN s00_aw_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 0.000 1922.710 4.000 ;
    END
  END s00_aw_len[5]
  PIN s00_aw_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 596.000 905.190 600.000 ;
    END
  END s00_aw_len[6]
  PIN s00_aw_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END s00_aw_len[7]
  PIN s00_aw_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 596.000 219.330 600.000 ;
    END
  END s00_aw_lock
  PIN s00_aw_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 596.000 1426.830 600.000 ;
    END
  END s00_aw_prot[0]
  PIN s00_aw_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.610 596.000 2144.890 600.000 ;
    END
  END s00_aw_prot[1]
  PIN s00_aw_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END s00_aw_prot[2]
  PIN s00_aw_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END s00_aw_qos[0]
  PIN s00_aw_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END s00_aw_qos[1]
  PIN s00_aw_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 596.000 1410.730 600.000 ;
    END
  END s00_aw_qos[2]
  PIN s00_aw_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 68.040 2400.000 68.640 ;
    END
  END s00_aw_qos[3]
  PIN s00_aw_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END s00_aw_ready
  PIN s00_aw_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 598.440 2400.000 599.040 ;
    END
  END s00_aw_region[0]
  PIN s00_aw_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END s00_aw_region[1]
  PIN s00_aw_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 596.000 1942.030 600.000 ;
    END
  END s00_aw_region[2]
  PIN s00_aw_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END s00_aw_region[3]
  PIN s00_aw_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END s00_aw_size[0]
  PIN s00_aw_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END s00_aw_size[1]
  PIN s00_aw_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 596.000 1323.790 600.000 ;
    END
  END s00_aw_size[2]
  PIN s00_aw_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 596.000 985.690 600.000 ;
    END
  END s00_aw_user[-1]
  PIN s00_aw_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 596.000 1085.510 600.000 ;
    END
  END s00_aw_user[0]
  PIN s00_aw_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 596.000 914.850 600.000 ;
    END
  END s00_aw_valid
  PIN s00_b_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END s00_b_id[0]
  PIN s00_b_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 0.000 1433.270 4.000 ;
    END
  END s00_b_id[1]
  PIN s00_b_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 486.240 2400.000 486.840 ;
    END
  END s00_b_id[2]
  PIN s00_b_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 596.000 1649.010 600.000 ;
    END
  END s00_b_id[3]
  PIN s00_b_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 596.000 1227.190 600.000 ;
    END
  END s00_b_id[4]
  PIN s00_b_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 183.640 2400.000 184.240 ;
    END
  END s00_b_id[5]
  PIN s00_b_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 0.000 1864.750 4.000 ;
    END
  END s00_b_id[6]
  PIN s00_b_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 596.000 1867.970 600.000 ;
    END
  END s00_b_id[7]
  PIN s00_b_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END s00_b_id[8]
  PIN s00_b_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END s00_b_id[9]
  PIN s00_b_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 596.000 608.950 600.000 ;
    END
  END s00_b_ready
  PIN s00_b_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END s00_b_resp[0]
  PIN s00_b_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.490 0.000 2318.770 4.000 ;
    END
  END s00_b_resp[1]
  PIN s00_b_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 596.000 988.910 600.000 ;
    END
  END s00_b_user[-1]
  PIN s00_b_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.510 0.000 1967.790 4.000 ;
    END
  END s00_b_user[0]
  PIN s00_b_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END s00_b_valid
  PIN s00_r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END s00_r_data[0]
  PIN s00_r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END s00_r_data[10]
  PIN s00_r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END s00_r_data[11]
  PIN s00_r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.510 596.000 2289.790 600.000 ;
    END
  END s00_r_data[12]
  PIN s00_r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 596.000 1513.770 600.000 ;
    END
  END s00_r_data[13]
  PIN s00_r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END s00_r_data[14]
  PIN s00_r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END s00_r_data[15]
  PIN s00_r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END s00_r_data[16]
  PIN s00_r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END s00_r_data[17]
  PIN s00_r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 596.000 1430.050 600.000 ;
    END
  END s00_r_data[18]
  PIN s00_r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 462.440 2400.000 463.040 ;
    END
  END s00_r_data[19]
  PIN s00_r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 596.000 1285.150 600.000 ;
    END
  END s00_r_data[1]
  PIN s00_r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 596.000 1523.430 600.000 ;
    END
  END s00_r_data[20]
  PIN s00_r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END s00_r_data[21]
  PIN s00_r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END s00_r_data[22]
  PIN s00_r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END s00_r_data[23]
  PIN s00_r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 596.000 151.710 600.000 ;
    END
  END s00_r_data[24]
  PIN s00_r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 596.000 634.710 600.000 ;
    END
  END s00_r_data[25]
  PIN s00_r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 596.000 2312.330 600.000 ;
    END
  END s00_r_data[26]
  PIN s00_r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END s00_r_data[27]
  PIN s00_r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END s00_r_data[28]
  PIN s00_r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END s00_r_data[29]
  PIN s00_r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END s00_r_data[2]
  PIN s00_r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.270 596.000 2154.550 600.000 ;
    END
  END s00_r_data[30]
  PIN s00_r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.010 0.000 2209.290 4.000 ;
    END
  END s00_r_data[31]
  PIN s00_r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 596.000 1494.450 600.000 ;
    END
  END s00_r_data[3]
  PIN s00_r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 596.000 464.050 600.000 ;
    END
  END s00_r_data[4]
  PIN s00_r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 596.000 1684.430 600.000 ;
    END
  END s00_r_data[5]
  PIN s00_r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.350 0.000 2038.630 4.000 ;
    END
  END s00_r_data[6]
  PIN s00_r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END s00_r_data[7]
  PIN s00_r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 596.000 631.490 600.000 ;
    END
  END s00_r_data[8]
  PIN s00_r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 596.000 1017.890 600.000 ;
    END
  END s00_r_data[9]
  PIN s00_r_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END s00_r_id[0]
  PIN s00_r_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 596.000 592.850 600.000 ;
    END
  END s00_r_id[1]
  PIN s00_r_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END s00_r_id[2]
  PIN s00_r_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 596.000 570.310 600.000 ;
    END
  END s00_r_id[3]
  PIN s00_r_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END s00_r_id[4]
  PIN s00_r_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END s00_r_id[5]
  PIN s00_r_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 0.000 1423.610 4.000 ;
    END
  END s00_r_id[6]
  PIN s00_r_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END s00_r_id[7]
  PIN s00_r_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 0.000 1285.150 4.000 ;
    END
  END s00_r_id[8]
  PIN s00_r_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.490 596.000 1996.770 600.000 ;
    END
  END s00_r_id[9]
  PIN s00_r_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END s00_r_last
  PIN s00_r_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 596.000 711.990 600.000 ;
    END
  END s00_r_ready
  PIN s00_r_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END s00_r_resp[0]
  PIN s00_r_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 0.000 1516.990 4.000 ;
    END
  END s00_r_resp[1]
  PIN s00_r_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 295.840 2400.000 296.440 ;
    END
  END s00_r_user[-1]
  PIN s00_r_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END s00_r_user[0]
  PIN s00_r_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END s00_r_valid
  PIN s00_w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END s00_w_data[0]
  PIN s00_w_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.390 596.000 2302.670 600.000 ;
    END
  END s00_w_data[10]
  PIN s00_w_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 596.000 512.350 600.000 ;
    END
  END s00_w_data[11]
  PIN s00_w_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 596.000 1153.130 600.000 ;
    END
  END s00_w_data[12]
  PIN s00_w_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END s00_w_data[13]
  PIN s00_w_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.730 0.000 1971.010 4.000 ;
    END
  END s00_w_data[14]
  PIN s00_w_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END s00_w_data[15]
  PIN s00_w_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END s00_w_data[16]
  PIN s00_w_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.570 0.000 2363.850 4.000 ;
    END
  END s00_w_data[17]
  PIN s00_w_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 596.000 805.370 600.000 ;
    END
  END s00_w_data[18]
  PIN s00_w_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END s00_w_data[19]
  PIN s00_w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 596.000 1484.790 600.000 ;
    END
  END s00_w_data[1]
  PIN s00_w_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 596.000 341.690 600.000 ;
    END
  END s00_w_data[20]
  PIN s00_w_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END s00_w_data[21]
  PIN s00_w_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 596.000 612.170 600.000 ;
    END
  END s00_w_data[22]
  PIN s00_w_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END s00_w_data[23]
  PIN s00_w_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.270 0.000 2154.550 4.000 ;
    END
  END s00_w_data[24]
  PIN s00_w_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 0.000 1401.070 4.000 ;
    END
  END s00_w_data[25]
  PIN s00_w_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END s00_w_data[26]
  PIN s00_w_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 360.440 2400.000 361.040 ;
    END
  END s00_w_data[27]
  PIN s00_w_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 596.000 303.050 600.000 ;
    END
  END s00_w_data[28]
  PIN s00_w_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 346.840 2400.000 347.440 ;
    END
  END s00_w_data[29]
  PIN s00_w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.790 596.000 2045.070 600.000 ;
    END
  END s00_w_data[2]
  PIN s00_w_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 533.840 2400.000 534.440 ;
    END
  END s00_w_data[30]
  PIN s00_w_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END s00_w_data[31]
  PIN s00_w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 596.000 1327.010 600.000 ;
    END
  END s00_w_data[3]
  PIN s00_w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END s00_w_data[4]
  PIN s00_w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.570 0.000 2041.850 4.000 ;
    END
  END s00_w_data[5]
  PIN s00_w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END s00_w_data[6]
  PIN s00_w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END s00_w_data[7]
  PIN s00_w_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END s00_w_data[8]
  PIN s00_w_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 596.000 3.590 600.000 ;
    END
  END s00_w_data[9]
  PIN s00_w_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 268.640 2400.000 269.240 ;
    END
  END s00_w_last
  PIN s00_w_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 37.440 2400.000 38.040 ;
    END
  END s00_w_ready
  PIN s00_w_strb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END s00_w_strb[0]
  PIN s00_w_strb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 596.000 621.830 600.000 ;
    END
  END s00_w_strb[1]
  PIN s00_w_strb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END s00_w_strb[2]
  PIN s00_w_strb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.750 0.000 2264.030 4.000 ;
    END
  END s00_w_strb[3]
  PIN s00_w_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 596.000 1668.330 600.000 ;
    END
  END s00_w_user[-1]
  PIN s00_w_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 394.440 2400.000 395.040 ;
    END
  END s00_w_user[0]
  PIN s00_w_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.930 596.000 2003.210 600.000 ;
    END
  END s00_w_valid
  PIN s01_ar_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 596.000 1636.130 600.000 ;
    END
  END s01_ar_addr[0]
  PIN s01_ar_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 0.000 1578.170 4.000 ;
    END
  END s01_ar_addr[10]
  PIN s01_ar_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.330 0.000 2228.610 4.000 ;
    END
  END s01_ar_addr[11]
  PIN s01_ar_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 4.000 ;
    END
  END s01_ar_addr[12]
  PIN s01_ar_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END s01_ar_addr[13]
  PIN s01_ar_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END s01_ar_addr[14]
  PIN s01_ar_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END s01_ar_addr[15]
  PIN s01_ar_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END s01_ar_addr[16]
  PIN s01_ar_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.970 596.000 1945.250 600.000 ;
    END
  END s01_ar_addr[17]
  PIN s01_ar_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 596.000 1079.070 600.000 ;
    END
  END s01_ar_addr[18]
  PIN s01_ar_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 0.000 1549.190 4.000 ;
    END
  END s01_ar_addr[19]
  PIN s01_ar_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 596.000 145.270 600.000 ;
    END
  END s01_ar_addr[1]
  PIN s01_ar_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END s01_ar_addr[20]
  PIN s01_ar_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END s01_ar_addr[21]
  PIN s01_ar_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 596.000 947.050 600.000 ;
    END
  END s01_ar_addr[22]
  PIN s01_ar_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 596.000 1397.850 600.000 ;
    END
  END s01_ar_addr[23]
  PIN s01_ar_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 596.000 1462.250 600.000 ;
    END
  END s01_ar_addr[24]
  PIN s01_ar_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.710 0.000 2321.990 4.000 ;
    END
  END s01_ar_addr[25]
  PIN s01_ar_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 596.000 950.270 600.000 ;
    END
  END s01_ar_addr[26]
  PIN s01_ar_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 0.000 2247.930 4.000 ;
    END
  END s01_ar_addr[27]
  PIN s01_ar_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END s01_ar_addr[28]
  PIN s01_ar_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END s01_ar_addr[29]
  PIN s01_ar_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 596.000 1584.610 600.000 ;
    END
  END s01_ar_addr[2]
  PIN s01_ar_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 596.000 1481.570 600.000 ;
    END
  END s01_ar_addr[30]
  PIN s01_ar_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END s01_ar_addr[31]
  PIN s01_ar_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END s01_ar_addr[3]
  PIN s01_ar_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 596.000 908.410 600.000 ;
    END
  END s01_ar_addr[4]
  PIN s01_ar_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 596.000 1752.050 600.000 ;
    END
  END s01_ar_addr[5]
  PIN s01_ar_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 596.000 1166.010 600.000 ;
    END
  END s01_ar_addr[6]
  PIN s01_ar_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 596.000 637.930 600.000 ;
    END
  END s01_ar_addr[7]
  PIN s01_ar_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 596.000 1452.590 600.000 ;
    END
  END s01_ar_addr[8]
  PIN s01_ar_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END s01_ar_addr[9]
  PIN s01_ar_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 596.000 1500.890 600.000 ;
    END
  END s01_ar_burst[0]
  PIN s01_ar_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 596.000 1272.270 600.000 ;
    END
  END s01_ar_burst[1]
  PIN s01_ar_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END s01_ar_cache[0]
  PIN s01_ar_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END s01_ar_cache[1]
  PIN s01_ar_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 275.440 2400.000 276.040 ;
    END
  END s01_ar_cache[2]
  PIN s01_ar_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 596.000 42.230 600.000 ;
    END
  END s01_ar_cache[3]
  PIN s01_ar_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END s01_ar_id[0]
  PIN s01_ar_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2366.790 0.000 2367.070 4.000 ;
    END
  END s01_ar_id[1]
  PIN s01_ar_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END s01_ar_id[2]
  PIN s01_ar_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 0.000 2070.830 4.000 ;
    END
  END s01_ar_id[3]
  PIN s01_ar_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 596.000 1037.210 600.000 ;
    END
  END s01_ar_id[4]
  PIN s01_ar_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END s01_ar_id[5]
  PIN s01_ar_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END s01_ar_id[6]
  PIN s01_ar_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 596.000 1771.370 600.000 ;
    END
  END s01_ar_id[7]
  PIN s01_ar_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.230 0.000 2051.510 4.000 ;
    END
  END s01_ar_id[8]
  PIN s01_ar_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 408.040 2400.000 408.640 ;
    END
  END s01_ar_id[9]
  PIN s01_ar_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 6.840 2400.000 7.440 ;
    END
  END s01_ar_len[0]
  PIN s01_ar_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 309.440 2400.000 310.040 ;
    END
  END s01_ar_len[1]
  PIN s01_ar_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 596.000 325.590 600.000 ;
    END
  END s01_ar_len[2]
  PIN s01_ar_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END s01_ar_len[3]
  PIN s01_ar_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.570 596.000 2041.850 600.000 ;
    END
  END s01_ar_len[4]
  PIN s01_ar_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.390 0.000 1819.670 4.000 ;
    END
  END s01_ar_len[5]
  PIN s01_ar_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 261.840 2400.000 262.440 ;
    END
  END s01_ar_len[6]
  PIN s01_ar_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 596.000 1562.070 600.000 ;
    END
  END s01_ar_len[7]
  PIN s01_ar_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 596.000 1620.030 600.000 ;
    END
  END s01_ar_lock
  PIN s01_ar_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 0.000 2048.290 4.000 ;
    END
  END s01_ar_prot[0]
  PIN s01_ar_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 0.000 1652.230 4.000 ;
    END
  END s01_ar_prot[1]
  PIN s01_ar_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 596.000 1243.290 600.000 ;
    END
  END s01_ar_prot[2]
  PIN s01_ar_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 596.000 1001.790 600.000 ;
    END
  END s01_ar_qos[0]
  PIN s01_ar_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 91.840 2400.000 92.440 ;
    END
  END s01_ar_qos[1]
  PIN s01_ar_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END s01_ar_qos[2]
  PIN s01_ar_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END s01_ar_qos[3]
  PIN s01_ar_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END s01_ar_ready
  PIN s01_ar_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 312.840 2400.000 313.440 ;
    END
  END s01_ar_region[0]
  PIN s01_ar_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 596.000 802.150 600.000 ;
    END
  END s01_ar_region[1]
  PIN s01_ar_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.490 0.000 2157.770 4.000 ;
    END
  END s01_ar_region[2]
  PIN s01_ar_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 596.000 19.690 600.000 ;
    END
  END s01_ar_region[3]
  PIN s01_ar_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2305.610 0.000 2305.890 4.000 ;
    END
  END s01_ar_size[0]
  PIN s01_ar_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 596.000 550.990 600.000 ;
    END
  END s01_ar_size[1]
  PIN s01_ar_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END s01_ar_size[2]
  PIN s01_ar_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 425.040 2400.000 425.640 ;
    END
  END s01_ar_user[-1]
  PIN s01_ar_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 596.000 2293.010 600.000 ;
    END
  END s01_ar_user[0]
  PIN s01_ar_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 596.000 1742.390 600.000 ;
    END
  END s01_ar_valid
  PIN s01_aw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.690 596.000 2189.970 600.000 ;
    END
  END s01_aw_addr[0]
  PIN s01_aw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 401.240 2400.000 401.840 ;
    END
  END s01_aw_addr[10]
  PIN s01_aw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 0.000 1568.510 4.000 ;
    END
  END s01_aw_addr[11]
  PIN s01_aw_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.370 596.000 2170.650 600.000 ;
    END
  END s01_aw_addr[12]
  PIN s01_aw_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END s01_aw_addr[13]
  PIN s01_aw_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END s01_aw_addr[14]
  PIN s01_aw_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 0.000 2125.570 4.000 ;
    END
  END s01_aw_addr[15]
  PIN s01_aw_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END s01_aw_addr[16]
  PIN s01_aw_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 596.000 196.790 600.000 ;
    END
  END s01_aw_addr[17]
  PIN s01_aw_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.170 596.000 2299.450 600.000 ;
    END
  END s01_aw_addr[18]
  PIN s01_aw_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END s01_aw_addr[19]
  PIN s01_aw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END s01_aw_addr[1]
  PIN s01_aw_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 596.000 1072.630 600.000 ;
    END
  END s01_aw_addr[20]
  PIN s01_aw_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 596.000 615.390 600.000 ;
    END
  END s01_aw_addr[21]
  PIN s01_aw_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 0.000 1942.030 4.000 ;
    END
  END s01_aw_addr[22]
  PIN s01_aw_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.230 596.000 2373.510 600.000 ;
    END
  END s01_aw_addr[23]
  PIN s01_aw_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 596.000 238.650 600.000 ;
    END
  END s01_aw_addr[24]
  PIN s01_aw_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.890 0.000 2383.170 4.000 ;
    END
  END s01_aw_addr[25]
  PIN s01_aw_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 596.000 441.510 600.000 ;
    END
  END s01_aw_addr[26]
  PIN s01_aw_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END s01_aw_addr[27]
  PIN s01_aw_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 4.000 ;
    END
  END s01_aw_addr[28]
  PIN s01_aw_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END s01_aw_addr[29]
  PIN s01_aw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 596.000 1124.150 600.000 ;
    END
  END s01_aw_addr[2]
  PIN s01_aw_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 520.240 2400.000 520.840 ;
    END
  END s01_aw_addr[30]
  PIN s01_aw_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 596.000 1262.610 600.000 ;
    END
  END s01_aw_addr[31]
  PIN s01_aw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 596.000 760.290 600.000 ;
    END
  END s01_aw_addr[3]
  PIN s01_aw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.190 0.000 1626.470 4.000 ;
    END
  END s01_aw_addr[4]
  PIN s01_aw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END s01_aw_addr[5]
  PIN s01_aw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 153.040 2400.000 153.640 ;
    END
  END s01_aw_addr[6]
  PIN s01_aw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 272.040 2400.000 272.640 ;
    END
  END s01_aw_addr[7]
  PIN s01_aw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 564.440 2400.000 565.040 ;
    END
  END s01_aw_addr[8]
  PIN s01_aw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 596.000 895.530 600.000 ;
    END
  END s01_aw_addr[9]
  PIN s01_aw_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 596.000 1916.270 600.000 ;
    END
  END s01_aw_burst[0]
  PIN s01_aw_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END s01_aw_burst[1]
  PIN s01_aw_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 596.000 1246.510 600.000 ;
    END
  END s01_aw_cache[0]
  PIN s01_aw_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END s01_aw_cache[1]
  PIN s01_aw_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 596.000 1616.810 600.000 ;
    END
  END s01_aw_cache[2]
  PIN s01_aw_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 459.040 2400.000 459.640 ;
    END
  END s01_aw_cache[3]
  PIN s01_aw_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 596.000 1442.930 600.000 ;
    END
  END s01_aw_id[0]
  PIN s01_aw_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 596.000 1919.490 600.000 ;
    END
  END s01_aw_id[1]
  PIN s01_aw_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END s01_aw_id[2]
  PIN s01_aw_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 596.000 1436.490 600.000 ;
    END
  END s01_aw_id[3]
  PIN s01_aw_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END s01_aw_id[4]
  PIN s01_aw_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 596.000 1388.190 600.000 ;
    END
  END s01_aw_id[5]
  PIN s01_aw_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 596.000 1607.150 600.000 ;
    END
  END s01_aw_id[6]
  PIN s01_aw_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 596.000 2141.670 600.000 ;
    END
  END s01_aw_id[7]
  PIN s01_aw_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.090 596.000 2254.370 600.000 ;
    END
  END s01_aw_id[8]
  PIN s01_aw_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END s01_aw_id[9]
  PIN s01_aw_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END s01_aw_len[0]
  PIN s01_aw_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 596.000 721.650 600.000 ;
    END
  END s01_aw_len[1]
  PIN s01_aw_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END s01_aw_len[2]
  PIN s01_aw_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 452.240 2400.000 452.840 ;
    END
  END s01_aw_len[3]
  PIN s01_aw_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 596.000 1420.390 600.000 ;
    END
  END s01_aw_len[4]
  PIN s01_aw_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 596.000 1336.670 600.000 ;
    END
  END s01_aw_len[5]
  PIN s01_aw_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 105.440 2400.000 106.040 ;
    END
  END s01_aw_len[6]
  PIN s01_aw_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 596.000 1346.330 600.000 ;
    END
  END s01_aw_len[7]
  PIN s01_aw_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END s01_aw_lock
  PIN s01_aw_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END s01_aw_prot[0]
  PIN s01_aw_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END s01_aw_prot[1]
  PIN s01_aw_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END s01_aw_prot[2]
  PIN s01_aw_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END s01_aw_qos[0]
  PIN s01_aw_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.110 0.000 2386.390 4.000 ;
    END
  END s01_aw_qos[1]
  PIN s01_aw_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 0.000 2328.430 4.000 ;
    END
  END s01_aw_qos[2]
  PIN s01_aw_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 112.240 2400.000 112.840 ;
    END
  END s01_aw_qos[3]
  PIN s01_aw_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 596.000 930.950 600.000 ;
    END
  END s01_aw_ready
  PIN s01_aw_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 596.000 167.810 600.000 ;
    END
  END s01_aw_region[0]
  PIN s01_aw_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END s01_aw_region[1]
  PIN s01_aw_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.670 596.000 2379.950 600.000 ;
    END
  END s01_aw_region[2]
  PIN s01_aw_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END s01_aw_region[3]
  PIN s01_aw_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 596.000 254.750 600.000 ;
    END
  END s01_aw_size[0]
  PIN s01_aw_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END s01_aw_size[1]
  PIN s01_aw_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 596.000 1378.530 600.000 ;
    END
  END s01_aw_size[2]
  PIN s01_aw_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 64.640 2400.000 65.240 ;
    END
  END s01_aw_user[-1]
  PIN s01_aw_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 596.000 1159.570 600.000 ;
    END
  END s01_aw_user[0]
  PIN s01_aw_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END s01_aw_valid
  PIN s01_b_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END s01_b_id[0]
  PIN s01_b_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.810 596.000 2016.090 600.000 ;
    END
  END s01_b_id[1]
  PIN s01_b_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END s01_b_id[2]
  PIN s01_b_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.850 596.000 2280.130 600.000 ;
    END
  END s01_b_id[3]
  PIN s01_b_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 596.000 116.290 600.000 ;
    END
  END s01_b_id[4]
  PIN s01_b_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 596.000 1533.090 600.000 ;
    END
  END s01_b_id[5]
  PIN s01_b_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 596.000 1075.850 600.000 ;
    END
  END s01_b_id[6]
  PIN s01_b_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 596.000 222.550 600.000 ;
    END
  END s01_b_id[7]
  PIN s01_b_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 596.000 483.370 600.000 ;
    END
  END s01_b_id[8]
  PIN s01_b_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 0.000 1829.330 4.000 ;
    END
  END s01_b_id[9]
  PIN s01_b_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.910 596.000 2193.190 600.000 ;
    END
  END s01_b_ready
  PIN s01_b_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 596.000 1040.430 600.000 ;
    END
  END s01_b_resp[0]
  PIN s01_b_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END s01_b_resp[1]
  PIN s01_b_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END s01_b_user[-1]
  PIN s01_b_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 596.000 2396.050 600.000 ;
    END
  END s01_b_user[0]
  PIN s01_b_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END s01_b_valid
  PIN s01_r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 596.000 190.350 600.000 ;
    END
  END s01_r_data[0]
  PIN s01_r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END s01_r_data[10]
  PIN s01_r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END s01_r_data[11]
  PIN s01_r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 596.000 2077.270 600.000 ;
    END
  END s01_r_data[12]
  PIN s01_r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END s01_r_data[13]
  PIN s01_r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END s01_r_data[14]
  PIN s01_r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 596.000 2225.390 600.000 ;
    END
  END s01_r_data[15]
  PIN s01_r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 596.000 402.870 600.000 ;
    END
  END s01_r_data[16]
  PIN s01_r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 363.840 2400.000 364.440 ;
    END
  END s01_r_data[17]
  PIN s01_r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 596.000 1372.090 600.000 ;
    END
  END s01_r_data[18]
  PIN s01_r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END s01_r_data[19]
  PIN s01_r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END s01_r_data[1]
  PIN s01_r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END s01_r_data[20]
  PIN s01_r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.450 0.000 2376.730 4.000 ;
    END
  END s01_r_data[21]
  PIN s01_r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 596.000 296.610 600.000 ;
    END
  END s01_r_data[22]
  PIN s01_r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END s01_r_data[23]
  PIN s01_r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 596.000 1459.030 600.000 ;
    END
  END s01_r_data[24]
  PIN s01_r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.190 596.000 1626.470 600.000 ;
    END
  END s01_r_data[25]
  PIN s01_r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END s01_r_data[26]
  PIN s01_r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 596.000 1536.310 600.000 ;
    END
  END s01_r_data[27]
  PIN s01_r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 119.040 2400.000 119.640 ;
    END
  END s01_r_data[28]
  PIN s01_r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 0.000 1874.410 4.000 ;
    END
  END s01_r_data[29]
  PIN s01_r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 596.000 257.970 600.000 ;
    END
  END s01_r_data[2]
  PIN s01_r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END s01_r_data[30]
  PIN s01_r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 596.000 2392.830 600.000 ;
    END
  END s01_r_data[31]
  PIN s01_r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END s01_r_data[3]
  PIN s01_r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 0.000 1735.950 4.000 ;
    END
  END s01_r_data[4]
  PIN s01_r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 596.000 1574.950 600.000 ;
    END
  END s01_r_data[5]
  PIN s01_r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 596.000 473.710 600.000 ;
    END
  END s01_r_data[6]
  PIN s01_r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END s01_r_data[7]
  PIN s01_r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END s01_r_data[8]
  PIN s01_r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 596.000 393.210 600.000 ;
    END
  END s01_r_data[9]
  PIN s01_r_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 596.000 1755.270 600.000 ;
    END
  END s01_r_id[0]
  PIN s01_r_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END s01_r_id[1]
  PIN s01_r_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 596.000 2177.090 600.000 ;
    END
  END s01_r_id[2]
  PIN s01_r_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 442.040 2400.000 442.640 ;
    END
  END s01_r_id[3]
  PIN s01_r_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END s01_r_id[4]
  PIN s01_r_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 244.840 2400.000 245.440 ;
    END
  END s01_r_id[5]
  PIN s01_r_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 596.000 673.350 600.000 ;
    END
  END s01_r_id[6]
  PIN s01_r_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 0.000 2135.230 4.000 ;
    END
  END s01_r_id[7]
  PIN s01_r_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.810 0.000 2338.090 4.000 ;
    END
  END s01_r_id[8]
  PIN s01_r_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 139.440 2400.000 140.040 ;
    END
  END s01_r_id[9]
  PIN s01_r_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END s01_r_last
  PIN s01_r_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 596.000 2112.690 600.000 ;
    END
  END s01_r_ready
  PIN s01_r_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END s01_r_resp[0]
  PIN s01_r_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.370 596.000 2331.650 600.000 ;
    END
  END s01_r_resp[1]
  PIN s01_r_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 596.000 1011.450 600.000 ;
    END
  END s01_r_user[-1]
  PIN s01_r_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 0.000 1655.450 4.000 ;
    END
  END s01_r_user[0]
  PIN s01_r_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END s01_r_valid
  PIN s01_w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END s01_w_data[0]
  PIN s01_w_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END s01_w_data[10]
  PIN s01_w_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 0.000 1980.670 4.000 ;
    END
  END s01_w_data[11]
  PIN s01_w_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 20.440 2400.000 21.040 ;
    END
  END s01_w_data[12]
  PIN s01_w_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 596.000 657.250 600.000 ;
    END
  END s01_w_data[13]
  PIN s01_w_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 571.240 2400.000 571.840 ;
    END
  END s01_w_data[14]
  PIN s01_w_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END s01_w_data[15]
  PIN s01_w_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END s01_w_data[16]
  PIN s01_w_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 596.000 538.110 600.000 ;
    END
  END s01_w_data[17]
  PIN s01_w_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END s01_w_data[18]
  PIN s01_w_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 596.000 228.990 600.000 ;
    END
  END s01_w_data[19]
  PIN s01_w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 0.000 1459.030 4.000 ;
    END
  END s01_w_data[1]
  PIN s01_w_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 596.000 1913.050 600.000 ;
    END
  END s01_w_data[20]
  PIN s01_w_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 10.240 2400.000 10.840 ;
    END
  END s01_w_data[21]
  PIN s01_w_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 596.000 1983.890 600.000 ;
    END
  END s01_w_data[22]
  PIN s01_w_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END s01_w_data[23]
  PIN s01_w_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 596.000 447.950 600.000 ;
    END
  END s01_w_data[24]
  PIN s01_w_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 596.000 679.790 600.000 ;
    END
  END s01_w_data[25]
  PIN s01_w_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END s01_w_data[26]
  PIN s01_w_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 596.000 628.270 600.000 ;
    END
  END s01_w_data[27]
  PIN s01_w_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END s01_w_data[28]
  PIN s01_w_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.310 0.000 1774.590 4.000 ;
    END
  END s01_w_data[29]
  PIN s01_w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.170 0.000 1977.450 4.000 ;
    END
  END s01_w_data[2]
  PIN s01_w_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.650 596.000 1925.930 600.000 ;
    END
  END s01_w_data[30]
  PIN s01_w_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 350.240 2400.000 350.840 ;
    END
  END s01_w_data[31]
  PIN s01_w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 149.640 2400.000 150.240 ;
    END
  END s01_w_data[3]
  PIN s01_w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END s01_w_data[4]
  PIN s01_w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END s01_w_data[5]
  PIN s01_w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END s01_w_data[6]
  PIN s01_w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 596.000 728.090 600.000 ;
    END
  END s01_w_data[7]
  PIN s01_w_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END s01_w_data[8]
  PIN s01_w_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END s01_w_data[9]
  PIN s01_w_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END s01_w_last
  PIN s01_w_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END s01_w_ready
  PIN s01_w_strb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.410 596.000 1951.690 600.000 ;
    END
  END s01_w_strb[0]
  PIN s01_w_strb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END s01_w_strb[1]
  PIN s01_w_strb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.990 0.000 2399.270 4.000 ;
    END
  END s01_w_strb[2]
  PIN s01_w_strb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END s01_w_strb[3]
  PIN s01_w_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 258.440 2400.000 259.040 ;
    END
  END s01_w_user[-1]
  PIN s01_w_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 136.040 2400.000 136.640 ;
    END
  END s01_w_user[0]
  PIN s01_w_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END s01_w_valid
  PIN s02_ar_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END s02_ar_addr[0]
  PIN s02_ar_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END s02_ar_addr[10]
  PIN s02_ar_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 596.000 1091.950 600.000 ;
    END
  END s02_ar_addr[11]
  PIN s02_ar_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END s02_ar_addr[12]
  PIN s02_ar_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 596.000 1294.810 600.000 ;
    END
  END s02_ar_addr[13]
  PIN s02_ar_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END s02_ar_addr[14]
  PIN s02_ar_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END s02_ar_addr[15]
  PIN s02_ar_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 596.000 2135.230 600.000 ;
    END
  END s02_ar_addr[16]
  PIN s02_ar_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END s02_ar_addr[17]
  PIN s02_ar_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END s02_ar_addr[18]
  PIN s02_ar_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END s02_ar_addr[19]
  PIN s02_ar_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 596.000 827.910 600.000 ;
    END
  END s02_ar_addr[1]
  PIN s02_ar_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 0.000 1591.050 4.000 ;
    END
  END s02_ar_addr[20]
  PIN s02_ar_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END s02_ar_addr[21]
  PIN s02_ar_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 596.000 872.990 600.000 ;
    END
  END s02_ar_addr[22]
  PIN s02_ar_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END s02_ar_addr[23]
  PIN s02_ar_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 596.000 1310.910 600.000 ;
    END
  END s02_ar_addr[24]
  PIN s02_ar_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 0.000 1629.690 4.000 ;
    END
  END s02_ar_addr[25]
  PIN s02_ar_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 329.840 2400.000 330.440 ;
    END
  END s02_ar_addr[26]
  PIN s02_ar_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 596.000 129.170 600.000 ;
    END
  END s02_ar_addr[27]
  PIN s02_ar_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 596.000 869.770 600.000 ;
    END
  END s02_ar_addr[28]
  PIN s02_ar_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 0.000 2103.030 4.000 ;
    END
  END s02_ar_addr[29]
  PIN s02_ar_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END s02_ar_addr[2]
  PIN s02_ar_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END s02_ar_addr[30]
  PIN s02_ar_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 596.000 1307.690 600.000 ;
    END
  END s02_ar_addr[31]
  PIN s02_ar_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END s02_ar_addr[3]
  PIN s02_ar_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 596.000 956.710 600.000 ;
    END
  END s02_ar_addr[4]
  PIN s02_ar_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END s02_ar_addr[5]
  PIN s02_ar_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 596.000 2160.990 600.000 ;
    END
  END s02_ar_addr[6]
  PIN s02_ar_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END s02_ar_addr[7]
  PIN s02_ar_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 596.000 1265.830 600.000 ;
    END
  END s02_ar_addr[8]
  PIN s02_ar_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.130 596.000 2196.410 600.000 ;
    END
  END s02_ar_addr[9]
  PIN s02_ar_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END s02_ar_burst[0]
  PIN s02_ar_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 596.000 889.090 600.000 ;
    END
  END s02_ar_burst[1]
  PIN s02_ar_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END s02_ar_cache[0]
  PIN s02_ar_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 596.000 74.430 600.000 ;
    END
  END s02_ar_cache[1]
  PIN s02_ar_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END s02_ar_cache[2]
  PIN s02_ar_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.270 596.000 2315.550 600.000 ;
    END
  END s02_ar_cache[3]
  PIN s02_ar_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END s02_ar_id[0]
  PIN s02_ar_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 596.000 547.770 600.000 ;
    END
  END s02_ar_id[1]
  PIN s02_ar_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 0.000 1169.230 4.000 ;
    END
  END s02_ar_id[2]
  PIN s02_ar_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END s02_ar_id[3]
  PIN s02_ar_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 596.000 1497.670 600.000 ;
    END
  END s02_ar_id[4]
  PIN s02_ar_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 384.240 2400.000 384.840 ;
    END
  END s02_ar_id[5]
  PIN s02_ar_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END s02_ar_id[6]
  PIN s02_ar_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.970 596.000 2267.250 600.000 ;
    END
  END s02_ar_id[7]
  PIN s02_ar_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 4.000 ;
    END
  END s02_ar_id[8]
  PIN s02_ar_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END s02_ar_id[9]
  PIN s02_ar_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 596.000 699.110 600.000 ;
    END
  END s02_ar_len[0]
  PIN s02_ar_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 596.000 1787.470 600.000 ;
    END
  END s02_ar_len[1]
  PIN s02_ar_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END s02_ar_len[2]
  PIN s02_ar_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 530.440 2400.000 531.040 ;
    END
  END s02_ar_len[3]
  PIN s02_ar_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 0.000 1623.250 4.000 ;
    END
  END s02_ar_len[4]
  PIN s02_ar_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 54.440 2400.000 55.040 ;
    END
  END s02_ar_len[5]
  PIN s02_ar_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 596.000 2080.490 600.000 ;
    END
  END s02_ar_len[6]
  PIN s02_ar_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 596.000 734.530 600.000 ;
    END
  END s02_ar_len[7]
  PIN s02_ar_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END s02_ar_lock
  PIN s02_ar_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END s02_ar_prot[0]
  PIN s02_ar_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END s02_ar_prot[1]
  PIN s02_ar_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.850 0.000 2280.130 4.000 ;
    END
  END s02_ar_prot[2]
  PIN s02_ar_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END s02_ar_qos[0]
  PIN s02_ar_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END s02_ar_qos[1]
  PIN s02_ar_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END s02_ar_qos[2]
  PIN s02_ar_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 596.000 1671.550 600.000 ;
    END
  END s02_ar_qos[3]
  PIN s02_ar_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 336.640 2400.000 337.240 ;
    END
  END s02_ar_ready
  PIN s02_ar_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END s02_ar_region[0]
  PIN s02_ar_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 180.240 2400.000 180.840 ;
    END
  END s02_ar_region[1]
  PIN s02_ar_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END s02_ar_region[2]
  PIN s02_ar_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 596.000 1343.110 600.000 ;
    END
  END s02_ar_region[3]
  PIN s02_ar_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 0.000 1230.410 4.000 ;
    END
  END s02_ar_size[0]
  PIN s02_ar_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 561.040 2400.000 561.640 ;
    END
  END s02_ar_size[1]
  PIN s02_ar_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 596.000 1594.270 600.000 ;
    END
  END s02_ar_size[2]
  PIN s02_ar_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 596.000 1384.970 600.000 ;
    END
  END s02_ar_user[-1]
  PIN s02_ar_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 596.000 918.070 600.000 ;
    END
  END s02_ar_user[0]
  PIN s02_ar_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 596.000 1629.690 600.000 ;
    END
  END s02_ar_valid
  PIN s02_aw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 596.000 270.850 600.000 ;
    END
  END s02_aw_addr[0]
  PIN s02_aw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END s02_aw_addr[10]
  PIN s02_aw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.370 0.000 2009.650 4.000 ;
    END
  END s02_aw_addr[11]
  PIN s02_aw_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 88.440 2400.000 89.040 ;
    END
  END s02_aw_addr[12]
  PIN s02_aw_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END s02_aw_addr[13]
  PIN s02_aw_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 596.000 695.890 600.000 ;
    END
  END s02_aw_addr[14]
  PIN s02_aw_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END s02_aw_addr[15]
  PIN s02_aw_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.150 596.000 2006.430 600.000 ;
    END
  END s02_aw_addr[16]
  PIN s02_aw_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.870 596.000 2251.150 600.000 ;
    END
  END s02_aw_addr[17]
  PIN s02_aw_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 596.000 1516.990 600.000 ;
    END
  END s02_aw_addr[18]
  PIN s02_aw_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 596.000 1851.870 600.000 ;
    END
  END s02_aw_addr[19]
  PIN s02_aw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 4.000 ;
    END
  END s02_aw_addr[1]
  PIN s02_aw_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END s02_aw_addr[20]
  PIN s02_aw_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END s02_aw_addr[21]
  PIN s02_aw_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.290 0.000 1964.570 4.000 ;
    END
  END s02_aw_addr[22]
  PIN s02_aw_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END s02_aw_addr[23]
  PIN s02_aw_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END s02_aw_addr[24]
  PIN s02_aw_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END s02_aw_addr[25]
  PIN s02_aw_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.330 0.000 2389.610 4.000 ;
    END
  END s02_aw_addr[26]
  PIN s02_aw_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.230 596.000 2051.510 600.000 ;
    END
  END s02_aw_addr[27]
  PIN s02_aw_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 596.000 844.010 600.000 ;
    END
  END s02_aw_addr[28]
  PIN s02_aw_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 596.000 769.950 600.000 ;
    END
  END s02_aw_addr[29]
  PIN s02_aw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 596.000 489.810 600.000 ;
    END
  END s02_aw_addr[2]
  PIN s02_aw_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END s02_aw_addr[30]
  PIN s02_aw_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 596.000 1893.730 600.000 ;
    END
  END s02_aw_addr[31]
  PIN s02_aw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 4.000 ;
    END
  END s02_aw_addr[3]
  PIN s02_aw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 596.000 412.530 600.000 ;
    END
  END s02_aw_addr[4]
  PIN s02_aw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END s02_aw_addr[5]
  PIN s02_aw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 596.000 2125.570 600.000 ;
    END
  END s02_aw_addr[6]
  PIN s02_aw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 596.000 1236.850 600.000 ;
    END
  END s02_aw_addr[7]
  PIN s02_aw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 596.000 1133.810 600.000 ;
    END
  END s02_aw_addr[8]
  PIN s02_aw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 596.000 1455.810 600.000 ;
    END
  END s02_aw_addr[9]
  PIN s02_aw_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 596.000 1552.410 600.000 ;
    END
  END s02_aw_burst[0]
  PIN s02_aw_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 596.000 1568.510 600.000 ;
    END
  END s02_aw_burst[1]
  PIN s02_aw_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END s02_aw_cache[0]
  PIN s02_aw_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 596.000 979.250 600.000 ;
    END
  END s02_aw_cache[1]
  PIN s02_aw_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END s02_aw_cache[2]
  PIN s02_aw_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END s02_aw_cache[3]
  PIN s02_aw_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 0.000 1581.390 4.000 ;
    END
  END s02_aw_id[0]
  PIN s02_aw_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END s02_aw_id[1]
  PIN s02_aw_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.730 0.000 2132.010 4.000 ;
    END
  END s02_aw_id[2]
  PIN s02_aw_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 596.000 1198.210 600.000 ;
    END
  END s02_aw_id[3]
  PIN s02_aw_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.290 0.000 2286.570 4.000 ;
    END
  END s02_aw_id[4]
  PIN s02_aw_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 596.000 26.130 600.000 ;
    END
  END s02_aw_id[5]
  PIN s02_aw_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END s02_aw_id[6]
  PIN s02_aw_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END s02_aw_id[7]
  PIN s02_aw_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END s02_aw_id[8]
  PIN s02_aw_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 596.000 1014.670 600.000 ;
    END
  END s02_aw_id[9]
  PIN s02_aw_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 4.000 ;
    END
  END s02_aw_len[0]
  PIN s02_aw_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END s02_aw_len[1]
  PIN s02_aw_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END s02_aw_len[2]
  PIN s02_aw_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END s02_aw_len[3]
  PIN s02_aw_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 596.000 2064.390 600.000 ;
    END
  END s02_aw_len[4]
  PIN s02_aw_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END s02_aw_len[5]
  PIN s02_aw_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 596.000 103.410 600.000 ;
    END
  END s02_aw_len[6]
  PIN s02_aw_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.970 0.000 1945.250 4.000 ;
    END
  END s02_aw_len[7]
  PIN s02_aw_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.150 596.000 2167.430 600.000 ;
    END
  END s02_aw_lock
  PIN s02_aw_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 596.000 840.790 600.000 ;
    END
  END s02_aw_prot[0]
  PIN s02_aw_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 581.440 2400.000 582.040 ;
    END
  END s02_aw_prot[1]
  PIN s02_aw_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END s02_aw_prot[2]
  PIN s02_aw_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 596.000 1275.490 600.000 ;
    END
  END s02_aw_qos[0]
  PIN s02_aw_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.510 0.000 2128.790 4.000 ;
    END
  END s02_aw_qos[1]
  PIN s02_aw_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 596.000 737.750 600.000 ;
    END
  END s02_aw_qos[2]
  PIN s02_aw_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END s02_aw_qos[3]
  PIN s02_aw_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 596.000 90.530 600.000 ;
    END
  END s02_aw_ready
  PIN s02_aw_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END s02_aw_region[0]
  PIN s02_aw_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 489.640 2400.000 490.240 ;
    END
  END s02_aw_region[1]
  PIN s02_aw_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END s02_aw_region[2]
  PIN s02_aw_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.330 596.000 2228.610 600.000 ;
    END
  END s02_aw_region[3]
  PIN s02_aw_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END s02_aw_size[0]
  PIN s02_aw_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 0.000 1800.350 4.000 ;
    END
  END s02_aw_size[1]
  PIN s02_aw_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 596.000 280.510 600.000 ;
    END
  END s02_aw_size[2]
  PIN s02_aw_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 596.000 1352.770 600.000 ;
    END
  END s02_aw_user[-1]
  PIN s02_aw_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.330 596.000 2067.610 600.000 ;
    END
  END s02_aw_user[0]
  PIN s02_aw_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 596.000 241.870 600.000 ;
    END
  END s02_aw_valid
  PIN s02_b_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 596.000 418.970 600.000 ;
    END
  END s02_b_id[0]
  PIN s02_b_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.690 0.000 2189.970 4.000 ;
    END
  END s02_b_id[1]
  PIN s02_b_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 596.000 161.370 600.000 ;
    END
  END s02_b_id[2]
  PIN s02_b_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 95.240 2400.000 95.840 ;
    END
  END s02_b_id[3]
  PIN s02_b_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 596.000 1069.410 600.000 ;
    END
  END s02_b_id[4]
  PIN s02_b_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 596.000 692.670 600.000 ;
    END
  END s02_b_id[5]
  PIN s02_b_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END s02_b_id[6]
  PIN s02_b_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END s02_b_id[7]
  PIN s02_b_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END s02_b_id[8]
  PIN s02_b_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.010 596.000 2209.290 600.000 ;
    END
  END s02_b_id[9]
  PIN s02_b_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END s02_b_ready
  PIN s02_b_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END s02_b_resp[0]
  PIN s02_b_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 527.040 2400.000 527.640 ;
    END
  END s02_b_resp[1]
  PIN s02_b_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.010 0.000 2370.290 4.000 ;
    END
  END s02_b_user[-1]
  PIN s02_b_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 4.000 ;
    END
  END s02_b_user[0]
  PIN s02_b_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END s02_b_valid
  PIN s02_r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 596.000 1665.110 600.000 ;
    END
  END s02_r_data[0]
  PIN s02_r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END s02_r_data[10]
  PIN s02_r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END s02_r_data[11]
  PIN s02_r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END s02_r_data[12]
  PIN s02_r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 596.000 264.410 600.000 ;
    END
  END s02_r_data[13]
  PIN s02_r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END s02_r_data[14]
  PIN s02_r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END s02_r_data[15]
  PIN s02_r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 596.000 683.010 600.000 ;
    END
  END s02_r_data[16]
  PIN s02_r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 404.640 2400.000 405.240 ;
    END
  END s02_r_data[17]
  PIN s02_r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 596.000 1935.590 600.000 ;
    END
  END s02_r_data[18]
  PIN s02_r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END s02_r_data[19]
  PIN s02_r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 596.000 1520.210 600.000 ;
    END
  END s02_r_data[1]
  PIN s02_r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 85.040 2400.000 85.640 ;
    END
  END s02_r_data[20]
  PIN s02_r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END s02_r_data[21]
  PIN s02_r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 596.000 1504.110 600.000 ;
    END
  END s02_r_data[22]
  PIN s02_r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END s02_r_data[23]
  PIN s02_r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END s02_r_data[24]
  PIN s02_r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END s02_r_data[25]
  PIN s02_r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END s02_r_data[26]
  PIN s02_r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 0.000 2186.750 4.000 ;
    END
  END s02_r_data[27]
  PIN s02_r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 596.000 786.050 600.000 ;
    END
  END s02_r_data[28]
  PIN s02_r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.590 596.000 2173.870 600.000 ;
    END
  END s02_r_data[29]
  PIN s02_r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END s02_r_data[2]
  PIN s02_r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 596.000 13.250 600.000 ;
    END
  END s02_r_data[30]
  PIN s02_r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END s02_r_data[31]
  PIN s02_r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END s02_r_data[3]
  PIN s02_r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END s02_r_data[4]
  PIN s02_r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 173.440 2400.000 174.040 ;
    END
  END s02_r_data[5]
  PIN s02_r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END s02_r_data[6]
  PIN s02_r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 596.000 1491.230 600.000 ;
    END
  END s02_r_data[7]
  PIN s02_r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 596.000 1900.170 600.000 ;
    END
  END s02_r_data[8]
  PIN s02_r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 596.000 454.390 600.000 ;
    END
  END s02_r_data[9]
  PIN s02_r_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END s02_r_id[0]
  PIN s02_r_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 282.240 2400.000 282.840 ;
    END
  END s02_r_id[1]
  PIN s02_r_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 596.000 1980.670 600.000 ;
    END
  END s02_r_id[2]
  PIN s02_r_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END s02_r_id[3]
  PIN s02_r_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 574.640 2400.000 575.240 ;
    END
  END s02_r_id[4]
  PIN s02_r_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.910 0.000 2193.190 4.000 ;
    END
  END s02_r_id[5]
  PIN s02_r_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END s02_r_id[6]
  PIN s02_r_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.390 596.000 1819.670 600.000 ;
    END
  END s02_r_id[7]
  PIN s02_r_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 596.000 860.110 600.000 ;
    END
  END s02_r_id[8]
  PIN s02_r_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END s02_r_id[9]
  PIN s02_r_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 231.240 2400.000 231.840 ;
    END
  END s02_r_last
  PIN s02_r_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END s02_r_ready
  PIN s02_r_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 0.000 2109.470 4.000 ;
    END
  END s02_r_resp[0]
  PIN s02_r_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END s02_r_resp[1]
  PIN s02_r_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 0.000 1684.430 4.000 ;
    END
  END s02_r_user[-1]
  PIN s02_r_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END s02_r_user[0]
  PIN s02_r_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END s02_r_valid
  PIN s02_w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 0.000 2312.330 4.000 ;
    END
  END s02_w_data[0]
  PIN s02_w_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 596.000 1832.550 600.000 ;
    END
  END s02_w_data[10]
  PIN s02_w_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.590 596.000 2334.870 600.000 ;
    END
  END s02_w_data[11]
  PIN s02_w_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 0.000 1687.650 4.000 ;
    END
  END s02_w_data[12]
  PIN s02_w_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END s02_w_data[13]
  PIN s02_w_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 108.840 2400.000 109.440 ;
    END
  END s02_w_data[14]
  PIN s02_w_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END s02_w_data[15]
  PIN s02_w_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.710 596.000 2321.990 600.000 ;
    END
  END s02_w_data[16]
  PIN s02_w_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 596.000 1816.450 600.000 ;
    END
  END s02_w_data[17]
  PIN s02_w_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END s02_w_data[18]
  PIN s02_w_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 596.000 1777.810 600.000 ;
    END
  END s02_w_data[19]
  PIN s02_w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END s02_w_data[1]
  PIN s02_w_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END s02_w_data[20]
  PIN s02_w_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END s02_w_data[21]
  PIN s02_w_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END s02_w_data[22]
  PIN s02_w_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END s02_w_data[23]
  PIN s02_w_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END s02_w_data[24]
  PIN s02_w_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 596.000 502.690 600.000 ;
    END
  END s02_w_data[25]
  PIN s02_w_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 596.000 1146.690 600.000 ;
    END
  END s02_w_data[26]
  PIN s02_w_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END s02_w_data[27]
  PIN s02_w_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END s02_w_data[28]
  PIN s02_w_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END s02_w_data[29]
  PIN s02_w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 596.000 1555.630 600.000 ;
    END
  END s02_w_data[2]
  PIN s02_w_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 596.000 1217.530 600.000 ;
    END
  END s02_w_data[30]
  PIN s02_w_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END s02_w_data[31]
  PIN s02_w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.710 596.000 1838.990 600.000 ;
    END
  END s02_w_data[3]
  PIN s02_w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 0.000 1961.350 4.000 ;
    END
  END s02_w_data[4]
  PIN s02_w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 596.000 274.070 600.000 ;
    END
  END s02_w_data[5]
  PIN s02_w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 316.240 2400.000 316.840 ;
    END
  END s02_w_data[6]
  PIN s02_w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END s02_w_data[7]
  PIN s02_w_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END s02_w_data[8]
  PIN s02_w_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END s02_w_data[9]
  PIN s02_w_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2396.000 241.440 2400.000 242.040 ;
    END
  END s02_w_last
  PIN s02_w_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END s02_w_ready
  PIN s02_w_strb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 596.000 1842.210 600.000 ;
    END
  END s02_w_strb[0]
  PIN s02_w_strb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 596.000 1829.330 600.000 ;
    END
  END s02_w_strb[1]
  PIN s02_w_strb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 596.000 757.070 600.000 ;
    END
  END s02_w_strb[2]
  PIN s02_w_strb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 596.000 1033.990 600.000 ;
    END
  END s02_w_strb[3]
  PIN s02_w_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END s02_w_user[-1]
  PIN s02_w_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END s02_w_user[0]
  PIN s02_w_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 596.000 641.150 600.000 ;
    END
  END s02_w_valid
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.890 0.000 2222.170 4.000 ;
    END
  END test_en_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2394.300 587.605 ;
      LAYER met1 ;
        RECT 0.070 4.120 2399.290 593.600 ;
      LAYER met2 ;
        RECT 0.650 595.720 3.030 598.925 ;
        RECT 3.870 595.720 6.250 598.925 ;
        RECT 7.090 595.720 9.470 598.925 ;
        RECT 10.310 595.720 12.690 598.925 ;
        RECT 13.530 595.720 19.130 598.925 ;
        RECT 19.970 595.720 22.350 598.925 ;
        RECT 23.190 595.720 25.570 598.925 ;
        RECT 26.410 595.720 28.790 598.925 ;
        RECT 29.630 595.720 32.010 598.925 ;
        RECT 32.850 595.720 35.230 598.925 ;
        RECT 36.070 595.720 41.670 598.925 ;
        RECT 42.510 595.720 44.890 598.925 ;
        RECT 45.730 595.720 48.110 598.925 ;
        RECT 48.950 595.720 51.330 598.925 ;
        RECT 52.170 595.720 54.550 598.925 ;
        RECT 55.390 595.720 60.990 598.925 ;
        RECT 61.830 595.720 64.210 598.925 ;
        RECT 65.050 595.720 67.430 598.925 ;
        RECT 68.270 595.720 70.650 598.925 ;
        RECT 71.490 595.720 73.870 598.925 ;
        RECT 74.710 595.720 77.090 598.925 ;
        RECT 77.930 595.720 83.530 598.925 ;
        RECT 84.370 595.720 86.750 598.925 ;
        RECT 87.590 595.720 89.970 598.925 ;
        RECT 90.810 595.720 93.190 598.925 ;
        RECT 94.030 595.720 96.410 598.925 ;
        RECT 97.250 595.720 102.850 598.925 ;
        RECT 103.690 595.720 106.070 598.925 ;
        RECT 106.910 595.720 109.290 598.925 ;
        RECT 110.130 595.720 112.510 598.925 ;
        RECT 113.350 595.720 115.730 598.925 ;
        RECT 116.570 595.720 118.950 598.925 ;
        RECT 119.790 595.720 125.390 598.925 ;
        RECT 126.230 595.720 128.610 598.925 ;
        RECT 129.450 595.720 131.830 598.925 ;
        RECT 132.670 595.720 135.050 598.925 ;
        RECT 135.890 595.720 138.270 598.925 ;
        RECT 139.110 595.720 144.710 598.925 ;
        RECT 145.550 595.720 147.930 598.925 ;
        RECT 148.770 595.720 151.150 598.925 ;
        RECT 151.990 595.720 154.370 598.925 ;
        RECT 155.210 595.720 157.590 598.925 ;
        RECT 158.430 595.720 160.810 598.925 ;
        RECT 161.650 595.720 167.250 598.925 ;
        RECT 168.090 595.720 170.470 598.925 ;
        RECT 171.310 595.720 173.690 598.925 ;
        RECT 174.530 595.720 176.910 598.925 ;
        RECT 177.750 595.720 180.130 598.925 ;
        RECT 180.970 595.720 186.570 598.925 ;
        RECT 187.410 595.720 189.790 598.925 ;
        RECT 190.630 595.720 193.010 598.925 ;
        RECT 193.850 595.720 196.230 598.925 ;
        RECT 197.070 595.720 199.450 598.925 ;
        RECT 200.290 595.720 202.670 598.925 ;
        RECT 203.510 595.720 209.110 598.925 ;
        RECT 209.950 595.720 212.330 598.925 ;
        RECT 213.170 595.720 215.550 598.925 ;
        RECT 216.390 595.720 218.770 598.925 ;
        RECT 219.610 595.720 221.990 598.925 ;
        RECT 222.830 595.720 228.430 598.925 ;
        RECT 229.270 595.720 231.650 598.925 ;
        RECT 232.490 595.720 234.870 598.925 ;
        RECT 235.710 595.720 238.090 598.925 ;
        RECT 238.930 595.720 241.310 598.925 ;
        RECT 242.150 595.720 244.530 598.925 ;
        RECT 245.370 595.720 250.970 598.925 ;
        RECT 251.810 595.720 254.190 598.925 ;
        RECT 255.030 595.720 257.410 598.925 ;
        RECT 258.250 595.720 260.630 598.925 ;
        RECT 261.470 595.720 263.850 598.925 ;
        RECT 264.690 595.720 270.290 598.925 ;
        RECT 271.130 595.720 273.510 598.925 ;
        RECT 274.350 595.720 276.730 598.925 ;
        RECT 277.570 595.720 279.950 598.925 ;
        RECT 280.790 595.720 283.170 598.925 ;
        RECT 284.010 595.720 286.390 598.925 ;
        RECT 287.230 595.720 292.830 598.925 ;
        RECT 293.670 595.720 296.050 598.925 ;
        RECT 296.890 595.720 299.270 598.925 ;
        RECT 300.110 595.720 302.490 598.925 ;
        RECT 303.330 595.720 305.710 598.925 ;
        RECT 306.550 595.720 312.150 598.925 ;
        RECT 312.990 595.720 315.370 598.925 ;
        RECT 316.210 595.720 318.590 598.925 ;
        RECT 319.430 595.720 321.810 598.925 ;
        RECT 322.650 595.720 325.030 598.925 ;
        RECT 325.870 595.720 328.250 598.925 ;
        RECT 329.090 595.720 334.690 598.925 ;
        RECT 335.530 595.720 337.910 598.925 ;
        RECT 338.750 595.720 341.130 598.925 ;
        RECT 341.970 595.720 344.350 598.925 ;
        RECT 345.190 595.720 347.570 598.925 ;
        RECT 348.410 595.720 350.790 598.925 ;
        RECT 351.630 595.720 357.230 598.925 ;
        RECT 358.070 595.720 360.450 598.925 ;
        RECT 361.290 595.720 363.670 598.925 ;
        RECT 364.510 595.720 366.890 598.925 ;
        RECT 367.730 595.720 370.110 598.925 ;
        RECT 370.950 595.720 376.550 598.925 ;
        RECT 377.390 595.720 379.770 598.925 ;
        RECT 380.610 595.720 382.990 598.925 ;
        RECT 383.830 595.720 386.210 598.925 ;
        RECT 387.050 595.720 389.430 598.925 ;
        RECT 390.270 595.720 392.650 598.925 ;
        RECT 393.490 595.720 399.090 598.925 ;
        RECT 399.930 595.720 402.310 598.925 ;
        RECT 403.150 595.720 405.530 598.925 ;
        RECT 406.370 595.720 408.750 598.925 ;
        RECT 409.590 595.720 411.970 598.925 ;
        RECT 412.810 595.720 418.410 598.925 ;
        RECT 419.250 595.720 421.630 598.925 ;
        RECT 422.470 595.720 424.850 598.925 ;
        RECT 425.690 595.720 428.070 598.925 ;
        RECT 428.910 595.720 431.290 598.925 ;
        RECT 432.130 595.720 434.510 598.925 ;
        RECT 435.350 595.720 440.950 598.925 ;
        RECT 441.790 595.720 444.170 598.925 ;
        RECT 445.010 595.720 447.390 598.925 ;
        RECT 448.230 595.720 450.610 598.925 ;
        RECT 451.450 595.720 453.830 598.925 ;
        RECT 454.670 595.720 460.270 598.925 ;
        RECT 461.110 595.720 463.490 598.925 ;
        RECT 464.330 595.720 466.710 598.925 ;
        RECT 467.550 595.720 469.930 598.925 ;
        RECT 470.770 595.720 473.150 598.925 ;
        RECT 473.990 595.720 476.370 598.925 ;
        RECT 477.210 595.720 482.810 598.925 ;
        RECT 483.650 595.720 486.030 598.925 ;
        RECT 486.870 595.720 489.250 598.925 ;
        RECT 490.090 595.720 492.470 598.925 ;
        RECT 493.310 595.720 495.690 598.925 ;
        RECT 496.530 595.720 502.130 598.925 ;
        RECT 502.970 595.720 505.350 598.925 ;
        RECT 506.190 595.720 508.570 598.925 ;
        RECT 509.410 595.720 511.790 598.925 ;
        RECT 512.630 595.720 515.010 598.925 ;
        RECT 515.850 595.720 518.230 598.925 ;
        RECT 519.070 595.720 524.670 598.925 ;
        RECT 525.510 595.720 527.890 598.925 ;
        RECT 528.730 595.720 531.110 598.925 ;
        RECT 531.950 595.720 534.330 598.925 ;
        RECT 535.170 595.720 537.550 598.925 ;
        RECT 538.390 595.720 543.990 598.925 ;
        RECT 544.830 595.720 547.210 598.925 ;
        RECT 548.050 595.720 550.430 598.925 ;
        RECT 551.270 595.720 553.650 598.925 ;
        RECT 554.490 595.720 556.870 598.925 ;
        RECT 557.710 595.720 560.090 598.925 ;
        RECT 560.930 595.720 566.530 598.925 ;
        RECT 567.370 595.720 569.750 598.925 ;
        RECT 570.590 595.720 572.970 598.925 ;
        RECT 573.810 595.720 576.190 598.925 ;
        RECT 577.030 595.720 579.410 598.925 ;
        RECT 580.250 595.720 585.850 598.925 ;
        RECT 586.690 595.720 589.070 598.925 ;
        RECT 589.910 595.720 592.290 598.925 ;
        RECT 593.130 595.720 595.510 598.925 ;
        RECT 596.350 595.720 598.730 598.925 ;
        RECT 599.570 595.720 601.950 598.925 ;
        RECT 602.790 595.720 608.390 598.925 ;
        RECT 609.230 595.720 611.610 598.925 ;
        RECT 612.450 595.720 614.830 598.925 ;
        RECT 615.670 595.720 618.050 598.925 ;
        RECT 618.890 595.720 621.270 598.925 ;
        RECT 622.110 595.720 627.710 598.925 ;
        RECT 628.550 595.720 630.930 598.925 ;
        RECT 631.770 595.720 634.150 598.925 ;
        RECT 634.990 595.720 637.370 598.925 ;
        RECT 638.210 595.720 640.590 598.925 ;
        RECT 641.430 595.720 643.810 598.925 ;
        RECT 644.650 595.720 650.250 598.925 ;
        RECT 651.090 595.720 653.470 598.925 ;
        RECT 654.310 595.720 656.690 598.925 ;
        RECT 657.530 595.720 659.910 598.925 ;
        RECT 660.750 595.720 663.130 598.925 ;
        RECT 663.970 595.720 669.570 598.925 ;
        RECT 670.410 595.720 672.790 598.925 ;
        RECT 673.630 595.720 676.010 598.925 ;
        RECT 676.850 595.720 679.230 598.925 ;
        RECT 680.070 595.720 682.450 598.925 ;
        RECT 683.290 595.720 685.670 598.925 ;
        RECT 686.510 595.720 692.110 598.925 ;
        RECT 692.950 595.720 695.330 598.925 ;
        RECT 696.170 595.720 698.550 598.925 ;
        RECT 699.390 595.720 701.770 598.925 ;
        RECT 702.610 595.720 704.990 598.925 ;
        RECT 705.830 595.720 711.430 598.925 ;
        RECT 712.270 595.720 714.650 598.925 ;
        RECT 715.490 595.720 717.870 598.925 ;
        RECT 718.710 595.720 721.090 598.925 ;
        RECT 721.930 595.720 724.310 598.925 ;
        RECT 725.150 595.720 727.530 598.925 ;
        RECT 728.370 595.720 733.970 598.925 ;
        RECT 734.810 595.720 737.190 598.925 ;
        RECT 738.030 595.720 740.410 598.925 ;
        RECT 741.250 595.720 743.630 598.925 ;
        RECT 744.470 595.720 746.850 598.925 ;
        RECT 747.690 595.720 753.290 598.925 ;
        RECT 754.130 595.720 756.510 598.925 ;
        RECT 757.350 595.720 759.730 598.925 ;
        RECT 760.570 595.720 762.950 598.925 ;
        RECT 763.790 595.720 766.170 598.925 ;
        RECT 767.010 595.720 769.390 598.925 ;
        RECT 770.230 595.720 775.830 598.925 ;
        RECT 776.670 595.720 779.050 598.925 ;
        RECT 779.890 595.720 782.270 598.925 ;
        RECT 783.110 595.720 785.490 598.925 ;
        RECT 786.330 595.720 788.710 598.925 ;
        RECT 789.550 595.720 795.150 598.925 ;
        RECT 795.990 595.720 798.370 598.925 ;
        RECT 799.210 595.720 801.590 598.925 ;
        RECT 802.430 595.720 804.810 598.925 ;
        RECT 805.650 595.720 808.030 598.925 ;
        RECT 808.870 595.720 811.250 598.925 ;
        RECT 812.090 595.720 817.690 598.925 ;
        RECT 818.530 595.720 820.910 598.925 ;
        RECT 821.750 595.720 824.130 598.925 ;
        RECT 824.970 595.720 827.350 598.925 ;
        RECT 828.190 595.720 830.570 598.925 ;
        RECT 831.410 595.720 833.790 598.925 ;
        RECT 834.630 595.720 840.230 598.925 ;
        RECT 841.070 595.720 843.450 598.925 ;
        RECT 844.290 595.720 846.670 598.925 ;
        RECT 847.510 595.720 849.890 598.925 ;
        RECT 850.730 595.720 853.110 598.925 ;
        RECT 853.950 595.720 859.550 598.925 ;
        RECT 860.390 595.720 862.770 598.925 ;
        RECT 863.610 595.720 865.990 598.925 ;
        RECT 866.830 595.720 869.210 598.925 ;
        RECT 870.050 595.720 872.430 598.925 ;
        RECT 873.270 595.720 875.650 598.925 ;
        RECT 876.490 595.720 882.090 598.925 ;
        RECT 882.930 595.720 885.310 598.925 ;
        RECT 886.150 595.720 888.530 598.925 ;
        RECT 889.370 595.720 891.750 598.925 ;
        RECT 892.590 595.720 894.970 598.925 ;
        RECT 895.810 595.720 901.410 598.925 ;
        RECT 902.250 595.720 904.630 598.925 ;
        RECT 905.470 595.720 907.850 598.925 ;
        RECT 908.690 595.720 911.070 598.925 ;
        RECT 911.910 595.720 914.290 598.925 ;
        RECT 915.130 595.720 917.510 598.925 ;
        RECT 918.350 595.720 923.950 598.925 ;
        RECT 924.790 595.720 927.170 598.925 ;
        RECT 928.010 595.720 930.390 598.925 ;
        RECT 931.230 595.720 933.610 598.925 ;
        RECT 934.450 595.720 936.830 598.925 ;
        RECT 937.670 595.720 943.270 598.925 ;
        RECT 944.110 595.720 946.490 598.925 ;
        RECT 947.330 595.720 949.710 598.925 ;
        RECT 950.550 595.720 952.930 598.925 ;
        RECT 953.770 595.720 956.150 598.925 ;
        RECT 956.990 595.720 959.370 598.925 ;
        RECT 960.210 595.720 965.810 598.925 ;
        RECT 966.650 595.720 969.030 598.925 ;
        RECT 969.870 595.720 972.250 598.925 ;
        RECT 973.090 595.720 975.470 598.925 ;
        RECT 976.310 595.720 978.690 598.925 ;
        RECT 979.530 595.720 985.130 598.925 ;
        RECT 985.970 595.720 988.350 598.925 ;
        RECT 989.190 595.720 991.570 598.925 ;
        RECT 992.410 595.720 994.790 598.925 ;
        RECT 995.630 595.720 998.010 598.925 ;
        RECT 998.850 595.720 1001.230 598.925 ;
        RECT 1002.070 595.720 1007.670 598.925 ;
        RECT 1008.510 595.720 1010.890 598.925 ;
        RECT 1011.730 595.720 1014.110 598.925 ;
        RECT 1014.950 595.720 1017.330 598.925 ;
        RECT 1018.170 595.720 1020.550 598.925 ;
        RECT 1021.390 595.720 1026.990 598.925 ;
        RECT 1027.830 595.720 1030.210 598.925 ;
        RECT 1031.050 595.720 1033.430 598.925 ;
        RECT 1034.270 595.720 1036.650 598.925 ;
        RECT 1037.490 595.720 1039.870 598.925 ;
        RECT 1040.710 595.720 1043.090 598.925 ;
        RECT 1043.930 595.720 1049.530 598.925 ;
        RECT 1050.370 595.720 1052.750 598.925 ;
        RECT 1053.590 595.720 1055.970 598.925 ;
        RECT 1056.810 595.720 1059.190 598.925 ;
        RECT 1060.030 595.720 1062.410 598.925 ;
        RECT 1063.250 595.720 1068.850 598.925 ;
        RECT 1069.690 595.720 1072.070 598.925 ;
        RECT 1072.910 595.720 1075.290 598.925 ;
        RECT 1076.130 595.720 1078.510 598.925 ;
        RECT 1079.350 595.720 1081.730 598.925 ;
        RECT 1082.570 595.720 1084.950 598.925 ;
        RECT 1085.790 595.720 1091.390 598.925 ;
        RECT 1092.230 595.720 1094.610 598.925 ;
        RECT 1095.450 595.720 1097.830 598.925 ;
        RECT 1098.670 595.720 1101.050 598.925 ;
        RECT 1101.890 595.720 1104.270 598.925 ;
        RECT 1105.110 595.720 1110.710 598.925 ;
        RECT 1111.550 595.720 1113.930 598.925 ;
        RECT 1114.770 595.720 1117.150 598.925 ;
        RECT 1117.990 595.720 1120.370 598.925 ;
        RECT 1121.210 595.720 1123.590 598.925 ;
        RECT 1124.430 595.720 1126.810 598.925 ;
        RECT 1127.650 595.720 1133.250 598.925 ;
        RECT 1134.090 595.720 1136.470 598.925 ;
        RECT 1137.310 595.720 1139.690 598.925 ;
        RECT 1140.530 595.720 1142.910 598.925 ;
        RECT 1143.750 595.720 1146.130 598.925 ;
        RECT 1146.970 595.720 1152.570 598.925 ;
        RECT 1153.410 595.720 1155.790 598.925 ;
        RECT 1156.630 595.720 1159.010 598.925 ;
        RECT 1159.850 595.720 1162.230 598.925 ;
        RECT 1163.070 595.720 1165.450 598.925 ;
        RECT 1166.290 595.720 1168.670 598.925 ;
        RECT 1169.510 595.720 1175.110 598.925 ;
        RECT 1175.950 595.720 1178.330 598.925 ;
        RECT 1179.170 595.720 1181.550 598.925 ;
        RECT 1182.390 595.720 1184.770 598.925 ;
        RECT 1185.610 595.720 1187.990 598.925 ;
        RECT 1188.830 595.720 1194.430 598.925 ;
        RECT 1195.270 595.720 1197.650 598.925 ;
        RECT 1198.490 595.720 1200.870 598.925 ;
        RECT 1201.710 595.720 1204.090 598.925 ;
        RECT 1204.930 595.720 1207.310 598.925 ;
        RECT 1208.150 595.720 1210.530 598.925 ;
        RECT 1211.370 595.720 1216.970 598.925 ;
        RECT 1217.810 595.720 1220.190 598.925 ;
        RECT 1221.030 595.720 1223.410 598.925 ;
        RECT 1224.250 595.720 1226.630 598.925 ;
        RECT 1227.470 595.720 1229.850 598.925 ;
        RECT 1230.690 595.720 1236.290 598.925 ;
        RECT 1237.130 595.720 1239.510 598.925 ;
        RECT 1240.350 595.720 1242.730 598.925 ;
        RECT 1243.570 595.720 1245.950 598.925 ;
        RECT 1246.790 595.720 1249.170 598.925 ;
        RECT 1250.010 595.720 1252.390 598.925 ;
        RECT 1253.230 595.720 1258.830 598.925 ;
        RECT 1259.670 595.720 1262.050 598.925 ;
        RECT 1262.890 595.720 1265.270 598.925 ;
        RECT 1266.110 595.720 1268.490 598.925 ;
        RECT 1269.330 595.720 1271.710 598.925 ;
        RECT 1272.550 595.720 1274.930 598.925 ;
        RECT 1275.770 595.720 1281.370 598.925 ;
        RECT 1282.210 595.720 1284.590 598.925 ;
        RECT 1285.430 595.720 1287.810 598.925 ;
        RECT 1288.650 595.720 1291.030 598.925 ;
        RECT 1291.870 595.720 1294.250 598.925 ;
        RECT 1295.090 595.720 1300.690 598.925 ;
        RECT 1301.530 595.720 1303.910 598.925 ;
        RECT 1304.750 595.720 1307.130 598.925 ;
        RECT 1307.970 595.720 1310.350 598.925 ;
        RECT 1311.190 595.720 1313.570 598.925 ;
        RECT 1314.410 595.720 1316.790 598.925 ;
        RECT 1317.630 595.720 1323.230 598.925 ;
        RECT 1324.070 595.720 1326.450 598.925 ;
        RECT 1327.290 595.720 1329.670 598.925 ;
        RECT 1330.510 595.720 1332.890 598.925 ;
        RECT 1333.730 595.720 1336.110 598.925 ;
        RECT 1336.950 595.720 1342.550 598.925 ;
        RECT 1343.390 595.720 1345.770 598.925 ;
        RECT 1346.610 595.720 1348.990 598.925 ;
        RECT 1349.830 595.720 1352.210 598.925 ;
        RECT 1353.050 595.720 1355.430 598.925 ;
        RECT 1356.270 595.720 1358.650 598.925 ;
        RECT 1359.490 595.720 1365.090 598.925 ;
        RECT 1365.930 595.720 1368.310 598.925 ;
        RECT 1369.150 595.720 1371.530 598.925 ;
        RECT 1372.370 595.720 1374.750 598.925 ;
        RECT 1375.590 595.720 1377.970 598.925 ;
        RECT 1378.810 595.720 1384.410 598.925 ;
        RECT 1385.250 595.720 1387.630 598.925 ;
        RECT 1388.470 595.720 1390.850 598.925 ;
        RECT 1391.690 595.720 1394.070 598.925 ;
        RECT 1394.910 595.720 1397.290 598.925 ;
        RECT 1398.130 595.720 1400.510 598.925 ;
        RECT 1401.350 595.720 1406.950 598.925 ;
        RECT 1407.790 595.720 1410.170 598.925 ;
        RECT 1411.010 595.720 1413.390 598.925 ;
        RECT 1414.230 595.720 1416.610 598.925 ;
        RECT 1417.450 595.720 1419.830 598.925 ;
        RECT 1420.670 595.720 1426.270 598.925 ;
        RECT 1427.110 595.720 1429.490 598.925 ;
        RECT 1430.330 595.720 1432.710 598.925 ;
        RECT 1433.550 595.720 1435.930 598.925 ;
        RECT 1436.770 595.720 1439.150 598.925 ;
        RECT 1439.990 595.720 1442.370 598.925 ;
        RECT 1443.210 595.720 1448.810 598.925 ;
        RECT 1449.650 595.720 1452.030 598.925 ;
        RECT 1452.870 595.720 1455.250 598.925 ;
        RECT 1456.090 595.720 1458.470 598.925 ;
        RECT 1459.310 595.720 1461.690 598.925 ;
        RECT 1462.530 595.720 1468.130 598.925 ;
        RECT 1468.970 595.720 1471.350 598.925 ;
        RECT 1472.190 595.720 1474.570 598.925 ;
        RECT 1475.410 595.720 1477.790 598.925 ;
        RECT 1478.630 595.720 1481.010 598.925 ;
        RECT 1481.850 595.720 1484.230 598.925 ;
        RECT 1485.070 595.720 1490.670 598.925 ;
        RECT 1491.510 595.720 1493.890 598.925 ;
        RECT 1494.730 595.720 1497.110 598.925 ;
        RECT 1497.950 595.720 1500.330 598.925 ;
        RECT 1501.170 595.720 1503.550 598.925 ;
        RECT 1504.390 595.720 1509.990 598.925 ;
        RECT 1510.830 595.720 1513.210 598.925 ;
        RECT 1514.050 595.720 1516.430 598.925 ;
        RECT 1517.270 595.720 1519.650 598.925 ;
        RECT 1520.490 595.720 1522.870 598.925 ;
        RECT 1523.710 595.720 1526.090 598.925 ;
        RECT 1526.930 595.720 1532.530 598.925 ;
        RECT 1533.370 595.720 1535.750 598.925 ;
        RECT 1536.590 595.720 1538.970 598.925 ;
        RECT 1539.810 595.720 1542.190 598.925 ;
        RECT 1543.030 595.720 1545.410 598.925 ;
        RECT 1546.250 595.720 1551.850 598.925 ;
        RECT 1552.690 595.720 1555.070 598.925 ;
        RECT 1555.910 595.720 1558.290 598.925 ;
        RECT 1559.130 595.720 1561.510 598.925 ;
        RECT 1562.350 595.720 1564.730 598.925 ;
        RECT 1565.570 595.720 1567.950 598.925 ;
        RECT 1568.790 595.720 1574.390 598.925 ;
        RECT 1575.230 595.720 1577.610 598.925 ;
        RECT 1578.450 595.720 1580.830 598.925 ;
        RECT 1581.670 595.720 1584.050 598.925 ;
        RECT 1584.890 595.720 1587.270 598.925 ;
        RECT 1588.110 595.720 1593.710 598.925 ;
        RECT 1594.550 595.720 1596.930 598.925 ;
        RECT 1597.770 595.720 1600.150 598.925 ;
        RECT 1600.990 595.720 1603.370 598.925 ;
        RECT 1604.210 595.720 1606.590 598.925 ;
        RECT 1607.430 595.720 1609.810 598.925 ;
        RECT 1610.650 595.720 1616.250 598.925 ;
        RECT 1617.090 595.720 1619.470 598.925 ;
        RECT 1620.310 595.720 1622.690 598.925 ;
        RECT 1623.530 595.720 1625.910 598.925 ;
        RECT 1626.750 595.720 1629.130 598.925 ;
        RECT 1629.970 595.720 1635.570 598.925 ;
        RECT 1636.410 595.720 1638.790 598.925 ;
        RECT 1639.630 595.720 1642.010 598.925 ;
        RECT 1642.850 595.720 1645.230 598.925 ;
        RECT 1646.070 595.720 1648.450 598.925 ;
        RECT 1649.290 595.720 1651.670 598.925 ;
        RECT 1652.510 595.720 1658.110 598.925 ;
        RECT 1658.950 595.720 1661.330 598.925 ;
        RECT 1662.170 595.720 1664.550 598.925 ;
        RECT 1665.390 595.720 1667.770 598.925 ;
        RECT 1668.610 595.720 1670.990 598.925 ;
        RECT 1671.830 595.720 1677.430 598.925 ;
        RECT 1678.270 595.720 1680.650 598.925 ;
        RECT 1681.490 595.720 1683.870 598.925 ;
        RECT 1684.710 595.720 1687.090 598.925 ;
        RECT 1687.930 595.720 1690.310 598.925 ;
        RECT 1691.150 595.720 1693.530 598.925 ;
        RECT 1694.370 595.720 1699.970 598.925 ;
        RECT 1700.810 595.720 1703.190 598.925 ;
        RECT 1704.030 595.720 1706.410 598.925 ;
        RECT 1707.250 595.720 1709.630 598.925 ;
        RECT 1710.470 595.720 1712.850 598.925 ;
        RECT 1713.690 595.720 1716.070 598.925 ;
        RECT 1716.910 595.720 1722.510 598.925 ;
        RECT 1723.350 595.720 1725.730 598.925 ;
        RECT 1726.570 595.720 1728.950 598.925 ;
        RECT 1729.790 595.720 1732.170 598.925 ;
        RECT 1733.010 595.720 1735.390 598.925 ;
        RECT 1736.230 595.720 1741.830 598.925 ;
        RECT 1742.670 595.720 1745.050 598.925 ;
        RECT 1745.890 595.720 1748.270 598.925 ;
        RECT 1749.110 595.720 1751.490 598.925 ;
        RECT 1752.330 595.720 1754.710 598.925 ;
        RECT 1755.550 595.720 1757.930 598.925 ;
        RECT 1758.770 595.720 1764.370 598.925 ;
        RECT 1765.210 595.720 1767.590 598.925 ;
        RECT 1768.430 595.720 1770.810 598.925 ;
        RECT 1771.650 595.720 1774.030 598.925 ;
        RECT 1774.870 595.720 1777.250 598.925 ;
        RECT 1778.090 595.720 1783.690 598.925 ;
        RECT 1784.530 595.720 1786.910 598.925 ;
        RECT 1787.750 595.720 1790.130 598.925 ;
        RECT 1790.970 595.720 1793.350 598.925 ;
        RECT 1794.190 595.720 1796.570 598.925 ;
        RECT 1797.410 595.720 1799.790 598.925 ;
        RECT 1800.630 595.720 1806.230 598.925 ;
        RECT 1807.070 595.720 1809.450 598.925 ;
        RECT 1810.290 595.720 1812.670 598.925 ;
        RECT 1813.510 595.720 1815.890 598.925 ;
        RECT 1816.730 595.720 1819.110 598.925 ;
        RECT 1819.950 595.720 1825.550 598.925 ;
        RECT 1826.390 595.720 1828.770 598.925 ;
        RECT 1829.610 595.720 1831.990 598.925 ;
        RECT 1832.830 595.720 1835.210 598.925 ;
        RECT 1836.050 595.720 1838.430 598.925 ;
        RECT 1839.270 595.720 1841.650 598.925 ;
        RECT 1842.490 595.720 1848.090 598.925 ;
        RECT 1848.930 595.720 1851.310 598.925 ;
        RECT 1852.150 595.720 1854.530 598.925 ;
        RECT 1855.370 595.720 1857.750 598.925 ;
        RECT 1858.590 595.720 1860.970 598.925 ;
        RECT 1861.810 595.720 1867.410 598.925 ;
        RECT 1868.250 595.720 1870.630 598.925 ;
        RECT 1871.470 595.720 1873.850 598.925 ;
        RECT 1874.690 595.720 1877.070 598.925 ;
        RECT 1877.910 595.720 1880.290 598.925 ;
        RECT 1881.130 595.720 1883.510 598.925 ;
        RECT 1884.350 595.720 1889.950 598.925 ;
        RECT 1890.790 595.720 1893.170 598.925 ;
        RECT 1894.010 595.720 1896.390 598.925 ;
        RECT 1897.230 595.720 1899.610 598.925 ;
        RECT 1900.450 595.720 1902.830 598.925 ;
        RECT 1903.670 595.720 1909.270 598.925 ;
        RECT 1910.110 595.720 1912.490 598.925 ;
        RECT 1913.330 595.720 1915.710 598.925 ;
        RECT 1916.550 595.720 1918.930 598.925 ;
        RECT 1919.770 595.720 1922.150 598.925 ;
        RECT 1922.990 595.720 1925.370 598.925 ;
        RECT 1926.210 595.720 1931.810 598.925 ;
        RECT 1932.650 595.720 1935.030 598.925 ;
        RECT 1935.870 595.720 1938.250 598.925 ;
        RECT 1939.090 595.720 1941.470 598.925 ;
        RECT 1942.310 595.720 1944.690 598.925 ;
        RECT 1945.530 595.720 1951.130 598.925 ;
        RECT 1951.970 595.720 1954.350 598.925 ;
        RECT 1955.190 595.720 1957.570 598.925 ;
        RECT 1958.410 595.720 1960.790 598.925 ;
        RECT 1961.630 595.720 1964.010 598.925 ;
        RECT 1964.850 595.720 1967.230 598.925 ;
        RECT 1968.070 595.720 1973.670 598.925 ;
        RECT 1974.510 595.720 1976.890 598.925 ;
        RECT 1977.730 595.720 1980.110 598.925 ;
        RECT 1980.950 595.720 1983.330 598.925 ;
        RECT 1984.170 595.720 1986.550 598.925 ;
        RECT 1987.390 595.720 1992.990 598.925 ;
        RECT 1993.830 595.720 1996.210 598.925 ;
        RECT 1997.050 595.720 1999.430 598.925 ;
        RECT 2000.270 595.720 2002.650 598.925 ;
        RECT 2003.490 595.720 2005.870 598.925 ;
        RECT 2006.710 595.720 2009.090 598.925 ;
        RECT 2009.930 595.720 2015.530 598.925 ;
        RECT 2016.370 595.720 2018.750 598.925 ;
        RECT 2019.590 595.720 2021.970 598.925 ;
        RECT 2022.810 595.720 2025.190 598.925 ;
        RECT 2026.030 595.720 2028.410 598.925 ;
        RECT 2029.250 595.720 2034.850 598.925 ;
        RECT 2035.690 595.720 2038.070 598.925 ;
        RECT 2038.910 595.720 2041.290 598.925 ;
        RECT 2042.130 595.720 2044.510 598.925 ;
        RECT 2045.350 595.720 2047.730 598.925 ;
        RECT 2048.570 595.720 2050.950 598.925 ;
        RECT 2051.790 595.720 2057.390 598.925 ;
        RECT 2058.230 595.720 2060.610 598.925 ;
        RECT 2061.450 595.720 2063.830 598.925 ;
        RECT 2064.670 595.720 2067.050 598.925 ;
        RECT 2067.890 595.720 2070.270 598.925 ;
        RECT 2071.110 595.720 2076.710 598.925 ;
        RECT 2077.550 595.720 2079.930 598.925 ;
        RECT 2080.770 595.720 2083.150 598.925 ;
        RECT 2083.990 595.720 2086.370 598.925 ;
        RECT 2087.210 595.720 2089.590 598.925 ;
        RECT 2090.430 595.720 2092.810 598.925 ;
        RECT 2093.650 595.720 2099.250 598.925 ;
        RECT 2100.090 595.720 2102.470 598.925 ;
        RECT 2103.310 595.720 2105.690 598.925 ;
        RECT 2106.530 595.720 2108.910 598.925 ;
        RECT 2109.750 595.720 2112.130 598.925 ;
        RECT 2112.970 595.720 2118.570 598.925 ;
        RECT 2119.410 595.720 2121.790 598.925 ;
        RECT 2122.630 595.720 2125.010 598.925 ;
        RECT 2125.850 595.720 2128.230 598.925 ;
        RECT 2129.070 595.720 2131.450 598.925 ;
        RECT 2132.290 595.720 2134.670 598.925 ;
        RECT 2135.510 595.720 2141.110 598.925 ;
        RECT 2141.950 595.720 2144.330 598.925 ;
        RECT 2145.170 595.720 2147.550 598.925 ;
        RECT 2148.390 595.720 2150.770 598.925 ;
        RECT 2151.610 595.720 2153.990 598.925 ;
        RECT 2154.830 595.720 2160.430 598.925 ;
        RECT 2161.270 595.720 2163.650 598.925 ;
        RECT 2164.490 595.720 2166.870 598.925 ;
        RECT 2167.710 595.720 2170.090 598.925 ;
        RECT 2170.930 595.720 2173.310 598.925 ;
        RECT 2174.150 595.720 2176.530 598.925 ;
        RECT 2177.370 595.720 2182.970 598.925 ;
        RECT 2183.810 595.720 2186.190 598.925 ;
        RECT 2187.030 595.720 2189.410 598.925 ;
        RECT 2190.250 595.720 2192.630 598.925 ;
        RECT 2193.470 595.720 2195.850 598.925 ;
        RECT 2196.690 595.720 2199.070 598.925 ;
        RECT 2199.910 595.720 2205.510 598.925 ;
        RECT 2206.350 595.720 2208.730 598.925 ;
        RECT 2209.570 595.720 2211.950 598.925 ;
        RECT 2212.790 595.720 2215.170 598.925 ;
        RECT 2216.010 595.720 2218.390 598.925 ;
        RECT 2219.230 595.720 2224.830 598.925 ;
        RECT 2225.670 595.720 2228.050 598.925 ;
        RECT 2228.890 595.720 2231.270 598.925 ;
        RECT 2232.110 595.720 2234.490 598.925 ;
        RECT 2235.330 595.720 2237.710 598.925 ;
        RECT 2238.550 595.720 2240.930 598.925 ;
        RECT 2241.770 595.720 2247.370 598.925 ;
        RECT 2248.210 595.720 2250.590 598.925 ;
        RECT 2251.430 595.720 2253.810 598.925 ;
        RECT 2254.650 595.720 2257.030 598.925 ;
        RECT 2257.870 595.720 2260.250 598.925 ;
        RECT 2261.090 595.720 2266.690 598.925 ;
        RECT 2267.530 595.720 2269.910 598.925 ;
        RECT 2270.750 595.720 2273.130 598.925 ;
        RECT 2273.970 595.720 2276.350 598.925 ;
        RECT 2277.190 595.720 2279.570 598.925 ;
        RECT 2280.410 595.720 2282.790 598.925 ;
        RECT 2283.630 595.720 2289.230 598.925 ;
        RECT 2290.070 595.720 2292.450 598.925 ;
        RECT 2293.290 595.720 2295.670 598.925 ;
        RECT 2296.510 595.720 2298.890 598.925 ;
        RECT 2299.730 595.720 2302.110 598.925 ;
        RECT 2302.950 595.720 2308.550 598.925 ;
        RECT 2309.390 595.720 2311.770 598.925 ;
        RECT 2312.610 595.720 2314.990 598.925 ;
        RECT 2315.830 595.720 2318.210 598.925 ;
        RECT 2319.050 595.720 2321.430 598.925 ;
        RECT 2322.270 595.720 2324.650 598.925 ;
        RECT 2325.490 595.720 2331.090 598.925 ;
        RECT 2331.930 595.720 2334.310 598.925 ;
        RECT 2335.150 595.720 2337.530 598.925 ;
        RECT 2338.370 595.720 2340.750 598.925 ;
        RECT 2341.590 595.720 2343.970 598.925 ;
        RECT 2344.810 595.720 2350.410 598.925 ;
        RECT 2351.250 595.720 2353.630 598.925 ;
        RECT 2354.470 595.720 2356.850 598.925 ;
        RECT 2357.690 595.720 2360.070 598.925 ;
        RECT 2360.910 595.720 2363.290 598.925 ;
        RECT 2364.130 595.720 2366.510 598.925 ;
        RECT 2367.350 595.720 2372.950 598.925 ;
        RECT 2373.790 595.720 2376.170 598.925 ;
        RECT 2377.010 595.720 2379.390 598.925 ;
        RECT 2380.230 595.720 2382.610 598.925 ;
        RECT 2383.450 595.720 2385.830 598.925 ;
        RECT 2386.670 595.720 2392.270 598.925 ;
        RECT 2393.110 595.720 2395.490 598.925 ;
        RECT 2396.330 595.720 2398.710 598.925 ;
        RECT 0.100 4.280 2399.260 595.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
        RECT 248.590 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 305.710 4.280 ;
        RECT 306.550 0.155 308.930 4.280 ;
        RECT 309.770 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 357.230 4.280 ;
        RECT 358.070 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 379.770 4.280 ;
        RECT 380.610 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 399.090 4.280 ;
        RECT 399.930 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 408.750 4.280 ;
        RECT 409.590 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 421.630 4.280 ;
        RECT 422.470 0.155 424.850 4.280 ;
        RECT 425.690 0.155 428.070 4.280 ;
        RECT 428.910 0.155 431.290 4.280 ;
        RECT 432.130 0.155 434.510 4.280 ;
        RECT 435.350 0.155 440.950 4.280 ;
        RECT 441.790 0.155 444.170 4.280 ;
        RECT 445.010 0.155 447.390 4.280 ;
        RECT 448.230 0.155 450.610 4.280 ;
        RECT 451.450 0.155 453.830 4.280 ;
        RECT 454.670 0.155 457.050 4.280 ;
        RECT 457.890 0.155 463.490 4.280 ;
        RECT 464.330 0.155 466.710 4.280 ;
        RECT 467.550 0.155 469.930 4.280 ;
        RECT 470.770 0.155 473.150 4.280 ;
        RECT 473.990 0.155 476.370 4.280 ;
        RECT 477.210 0.155 479.590 4.280 ;
        RECT 480.430 0.155 486.030 4.280 ;
        RECT 486.870 0.155 489.250 4.280 ;
        RECT 490.090 0.155 492.470 4.280 ;
        RECT 493.310 0.155 495.690 4.280 ;
        RECT 496.530 0.155 498.910 4.280 ;
        RECT 499.750 0.155 505.350 4.280 ;
        RECT 506.190 0.155 508.570 4.280 ;
        RECT 509.410 0.155 511.790 4.280 ;
        RECT 512.630 0.155 515.010 4.280 ;
        RECT 515.850 0.155 518.230 4.280 ;
        RECT 519.070 0.155 521.450 4.280 ;
        RECT 522.290 0.155 527.890 4.280 ;
        RECT 528.730 0.155 531.110 4.280 ;
        RECT 531.950 0.155 534.330 4.280 ;
        RECT 535.170 0.155 537.550 4.280 ;
        RECT 538.390 0.155 540.770 4.280 ;
        RECT 541.610 0.155 547.210 4.280 ;
        RECT 548.050 0.155 550.430 4.280 ;
        RECT 551.270 0.155 553.650 4.280 ;
        RECT 554.490 0.155 556.870 4.280 ;
        RECT 557.710 0.155 560.090 4.280 ;
        RECT 560.930 0.155 563.310 4.280 ;
        RECT 564.150 0.155 569.750 4.280 ;
        RECT 570.590 0.155 572.970 4.280 ;
        RECT 573.810 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 582.630 4.280 ;
        RECT 583.470 0.155 589.070 4.280 ;
        RECT 589.910 0.155 592.290 4.280 ;
        RECT 593.130 0.155 595.510 4.280 ;
        RECT 596.350 0.155 598.730 4.280 ;
        RECT 599.570 0.155 601.950 4.280 ;
        RECT 602.790 0.155 605.170 4.280 ;
        RECT 606.010 0.155 611.610 4.280 ;
        RECT 612.450 0.155 614.830 4.280 ;
        RECT 615.670 0.155 618.050 4.280 ;
        RECT 618.890 0.155 621.270 4.280 ;
        RECT 622.110 0.155 624.490 4.280 ;
        RECT 625.330 0.155 630.930 4.280 ;
        RECT 631.770 0.155 634.150 4.280 ;
        RECT 634.990 0.155 637.370 4.280 ;
        RECT 638.210 0.155 640.590 4.280 ;
        RECT 641.430 0.155 643.810 4.280 ;
        RECT 644.650 0.155 647.030 4.280 ;
        RECT 647.870 0.155 653.470 4.280 ;
        RECT 654.310 0.155 656.690 4.280 ;
        RECT 657.530 0.155 659.910 4.280 ;
        RECT 660.750 0.155 663.130 4.280 ;
        RECT 663.970 0.155 666.350 4.280 ;
        RECT 667.190 0.155 672.790 4.280 ;
        RECT 673.630 0.155 676.010 4.280 ;
        RECT 676.850 0.155 679.230 4.280 ;
        RECT 680.070 0.155 682.450 4.280 ;
        RECT 683.290 0.155 685.670 4.280 ;
        RECT 686.510 0.155 688.890 4.280 ;
        RECT 689.730 0.155 695.330 4.280 ;
        RECT 696.170 0.155 698.550 4.280 ;
        RECT 699.390 0.155 701.770 4.280 ;
        RECT 702.610 0.155 704.990 4.280 ;
        RECT 705.830 0.155 708.210 4.280 ;
        RECT 709.050 0.155 714.650 4.280 ;
        RECT 715.490 0.155 717.870 4.280 ;
        RECT 718.710 0.155 721.090 4.280 ;
        RECT 721.930 0.155 724.310 4.280 ;
        RECT 725.150 0.155 727.530 4.280 ;
        RECT 728.370 0.155 730.750 4.280 ;
        RECT 731.590 0.155 737.190 4.280 ;
        RECT 738.030 0.155 740.410 4.280 ;
        RECT 741.250 0.155 743.630 4.280 ;
        RECT 744.470 0.155 746.850 4.280 ;
        RECT 747.690 0.155 750.070 4.280 ;
        RECT 750.910 0.155 756.510 4.280 ;
        RECT 757.350 0.155 759.730 4.280 ;
        RECT 760.570 0.155 762.950 4.280 ;
        RECT 763.790 0.155 766.170 4.280 ;
        RECT 767.010 0.155 769.390 4.280 ;
        RECT 770.230 0.155 772.610 4.280 ;
        RECT 773.450 0.155 779.050 4.280 ;
        RECT 779.890 0.155 782.270 4.280 ;
        RECT 783.110 0.155 785.490 4.280 ;
        RECT 786.330 0.155 788.710 4.280 ;
        RECT 789.550 0.155 791.930 4.280 ;
        RECT 792.770 0.155 798.370 4.280 ;
        RECT 799.210 0.155 801.590 4.280 ;
        RECT 802.430 0.155 804.810 4.280 ;
        RECT 805.650 0.155 808.030 4.280 ;
        RECT 808.870 0.155 811.250 4.280 ;
        RECT 812.090 0.155 814.470 4.280 ;
        RECT 815.310 0.155 820.910 4.280 ;
        RECT 821.750 0.155 824.130 4.280 ;
        RECT 824.970 0.155 827.350 4.280 ;
        RECT 828.190 0.155 830.570 4.280 ;
        RECT 831.410 0.155 833.790 4.280 ;
        RECT 834.630 0.155 840.230 4.280 ;
        RECT 841.070 0.155 843.450 4.280 ;
        RECT 844.290 0.155 846.670 4.280 ;
        RECT 847.510 0.155 849.890 4.280 ;
        RECT 850.730 0.155 853.110 4.280 ;
        RECT 853.950 0.155 856.330 4.280 ;
        RECT 857.170 0.155 862.770 4.280 ;
        RECT 863.610 0.155 865.990 4.280 ;
        RECT 866.830 0.155 869.210 4.280 ;
        RECT 870.050 0.155 872.430 4.280 ;
        RECT 873.270 0.155 875.650 4.280 ;
        RECT 876.490 0.155 882.090 4.280 ;
        RECT 882.930 0.155 885.310 4.280 ;
        RECT 886.150 0.155 888.530 4.280 ;
        RECT 889.370 0.155 891.750 4.280 ;
        RECT 892.590 0.155 894.970 4.280 ;
        RECT 895.810 0.155 898.190 4.280 ;
        RECT 899.030 0.155 904.630 4.280 ;
        RECT 905.470 0.155 907.850 4.280 ;
        RECT 908.690 0.155 911.070 4.280 ;
        RECT 911.910 0.155 914.290 4.280 ;
        RECT 915.130 0.155 917.510 4.280 ;
        RECT 918.350 0.155 920.730 4.280 ;
        RECT 921.570 0.155 927.170 4.280 ;
        RECT 928.010 0.155 930.390 4.280 ;
        RECT 931.230 0.155 933.610 4.280 ;
        RECT 934.450 0.155 936.830 4.280 ;
        RECT 937.670 0.155 940.050 4.280 ;
        RECT 940.890 0.155 946.490 4.280 ;
        RECT 947.330 0.155 949.710 4.280 ;
        RECT 950.550 0.155 952.930 4.280 ;
        RECT 953.770 0.155 956.150 4.280 ;
        RECT 956.990 0.155 959.370 4.280 ;
        RECT 960.210 0.155 962.590 4.280 ;
        RECT 963.430 0.155 969.030 4.280 ;
        RECT 969.870 0.155 972.250 4.280 ;
        RECT 973.090 0.155 975.470 4.280 ;
        RECT 976.310 0.155 978.690 4.280 ;
        RECT 979.530 0.155 981.910 4.280 ;
        RECT 982.750 0.155 988.350 4.280 ;
        RECT 989.190 0.155 991.570 4.280 ;
        RECT 992.410 0.155 994.790 4.280 ;
        RECT 995.630 0.155 998.010 4.280 ;
        RECT 998.850 0.155 1001.230 4.280 ;
        RECT 1002.070 0.155 1004.450 4.280 ;
        RECT 1005.290 0.155 1010.890 4.280 ;
        RECT 1011.730 0.155 1014.110 4.280 ;
        RECT 1014.950 0.155 1017.330 4.280 ;
        RECT 1018.170 0.155 1020.550 4.280 ;
        RECT 1021.390 0.155 1023.770 4.280 ;
        RECT 1024.610 0.155 1030.210 4.280 ;
        RECT 1031.050 0.155 1033.430 4.280 ;
        RECT 1034.270 0.155 1036.650 4.280 ;
        RECT 1037.490 0.155 1039.870 4.280 ;
        RECT 1040.710 0.155 1043.090 4.280 ;
        RECT 1043.930 0.155 1046.310 4.280 ;
        RECT 1047.150 0.155 1052.750 4.280 ;
        RECT 1053.590 0.155 1055.970 4.280 ;
        RECT 1056.810 0.155 1059.190 4.280 ;
        RECT 1060.030 0.155 1062.410 4.280 ;
        RECT 1063.250 0.155 1065.630 4.280 ;
        RECT 1066.470 0.155 1072.070 4.280 ;
        RECT 1072.910 0.155 1075.290 4.280 ;
        RECT 1076.130 0.155 1078.510 4.280 ;
        RECT 1079.350 0.155 1081.730 4.280 ;
        RECT 1082.570 0.155 1084.950 4.280 ;
        RECT 1085.790 0.155 1088.170 4.280 ;
        RECT 1089.010 0.155 1094.610 4.280 ;
        RECT 1095.450 0.155 1097.830 4.280 ;
        RECT 1098.670 0.155 1101.050 4.280 ;
        RECT 1101.890 0.155 1104.270 4.280 ;
        RECT 1105.110 0.155 1107.490 4.280 ;
        RECT 1108.330 0.155 1113.930 4.280 ;
        RECT 1114.770 0.155 1117.150 4.280 ;
        RECT 1117.990 0.155 1120.370 4.280 ;
        RECT 1121.210 0.155 1123.590 4.280 ;
        RECT 1124.430 0.155 1126.810 4.280 ;
        RECT 1127.650 0.155 1130.030 4.280 ;
        RECT 1130.870 0.155 1136.470 4.280 ;
        RECT 1137.310 0.155 1139.690 4.280 ;
        RECT 1140.530 0.155 1142.910 4.280 ;
        RECT 1143.750 0.155 1146.130 4.280 ;
        RECT 1146.970 0.155 1149.350 4.280 ;
        RECT 1150.190 0.155 1155.790 4.280 ;
        RECT 1156.630 0.155 1159.010 4.280 ;
        RECT 1159.850 0.155 1162.230 4.280 ;
        RECT 1163.070 0.155 1165.450 4.280 ;
        RECT 1166.290 0.155 1168.670 4.280 ;
        RECT 1169.510 0.155 1171.890 4.280 ;
        RECT 1172.730 0.155 1178.330 4.280 ;
        RECT 1179.170 0.155 1181.550 4.280 ;
        RECT 1182.390 0.155 1184.770 4.280 ;
        RECT 1185.610 0.155 1187.990 4.280 ;
        RECT 1188.830 0.155 1191.210 4.280 ;
        RECT 1192.050 0.155 1197.650 4.280 ;
        RECT 1198.490 0.155 1200.870 4.280 ;
        RECT 1201.710 0.155 1204.090 4.280 ;
        RECT 1204.930 0.155 1207.310 4.280 ;
        RECT 1208.150 0.155 1210.530 4.280 ;
        RECT 1211.370 0.155 1213.750 4.280 ;
        RECT 1214.590 0.155 1220.190 4.280 ;
        RECT 1221.030 0.155 1223.410 4.280 ;
        RECT 1224.250 0.155 1226.630 4.280 ;
        RECT 1227.470 0.155 1229.850 4.280 ;
        RECT 1230.690 0.155 1233.070 4.280 ;
        RECT 1233.910 0.155 1239.510 4.280 ;
        RECT 1240.350 0.155 1242.730 4.280 ;
        RECT 1243.570 0.155 1245.950 4.280 ;
        RECT 1246.790 0.155 1249.170 4.280 ;
        RECT 1250.010 0.155 1252.390 4.280 ;
        RECT 1253.230 0.155 1255.610 4.280 ;
        RECT 1256.450 0.155 1262.050 4.280 ;
        RECT 1262.890 0.155 1265.270 4.280 ;
        RECT 1266.110 0.155 1268.490 4.280 ;
        RECT 1269.330 0.155 1271.710 4.280 ;
        RECT 1272.550 0.155 1274.930 4.280 ;
        RECT 1275.770 0.155 1281.370 4.280 ;
        RECT 1282.210 0.155 1284.590 4.280 ;
        RECT 1285.430 0.155 1287.810 4.280 ;
        RECT 1288.650 0.155 1291.030 4.280 ;
        RECT 1291.870 0.155 1294.250 4.280 ;
        RECT 1295.090 0.155 1297.470 4.280 ;
        RECT 1298.310 0.155 1303.910 4.280 ;
        RECT 1304.750 0.155 1307.130 4.280 ;
        RECT 1307.970 0.155 1310.350 4.280 ;
        RECT 1311.190 0.155 1313.570 4.280 ;
        RECT 1314.410 0.155 1316.790 4.280 ;
        RECT 1317.630 0.155 1323.230 4.280 ;
        RECT 1324.070 0.155 1326.450 4.280 ;
        RECT 1327.290 0.155 1329.670 4.280 ;
        RECT 1330.510 0.155 1332.890 4.280 ;
        RECT 1333.730 0.155 1336.110 4.280 ;
        RECT 1336.950 0.155 1339.330 4.280 ;
        RECT 1340.170 0.155 1345.770 4.280 ;
        RECT 1346.610 0.155 1348.990 4.280 ;
        RECT 1349.830 0.155 1352.210 4.280 ;
        RECT 1353.050 0.155 1355.430 4.280 ;
        RECT 1356.270 0.155 1358.650 4.280 ;
        RECT 1359.490 0.155 1365.090 4.280 ;
        RECT 1365.930 0.155 1368.310 4.280 ;
        RECT 1369.150 0.155 1371.530 4.280 ;
        RECT 1372.370 0.155 1374.750 4.280 ;
        RECT 1375.590 0.155 1377.970 4.280 ;
        RECT 1378.810 0.155 1381.190 4.280 ;
        RECT 1382.030 0.155 1387.630 4.280 ;
        RECT 1388.470 0.155 1390.850 4.280 ;
        RECT 1391.690 0.155 1394.070 4.280 ;
        RECT 1394.910 0.155 1397.290 4.280 ;
        RECT 1398.130 0.155 1400.510 4.280 ;
        RECT 1401.350 0.155 1403.730 4.280 ;
        RECT 1404.570 0.155 1410.170 4.280 ;
        RECT 1411.010 0.155 1413.390 4.280 ;
        RECT 1414.230 0.155 1416.610 4.280 ;
        RECT 1417.450 0.155 1419.830 4.280 ;
        RECT 1420.670 0.155 1423.050 4.280 ;
        RECT 1423.890 0.155 1429.490 4.280 ;
        RECT 1430.330 0.155 1432.710 4.280 ;
        RECT 1433.550 0.155 1435.930 4.280 ;
        RECT 1436.770 0.155 1439.150 4.280 ;
        RECT 1439.990 0.155 1442.370 4.280 ;
        RECT 1443.210 0.155 1445.590 4.280 ;
        RECT 1446.430 0.155 1452.030 4.280 ;
        RECT 1452.870 0.155 1455.250 4.280 ;
        RECT 1456.090 0.155 1458.470 4.280 ;
        RECT 1459.310 0.155 1461.690 4.280 ;
        RECT 1462.530 0.155 1464.910 4.280 ;
        RECT 1465.750 0.155 1471.350 4.280 ;
        RECT 1472.190 0.155 1474.570 4.280 ;
        RECT 1475.410 0.155 1477.790 4.280 ;
        RECT 1478.630 0.155 1481.010 4.280 ;
        RECT 1481.850 0.155 1484.230 4.280 ;
        RECT 1485.070 0.155 1487.450 4.280 ;
        RECT 1488.290 0.155 1493.890 4.280 ;
        RECT 1494.730 0.155 1497.110 4.280 ;
        RECT 1497.950 0.155 1500.330 4.280 ;
        RECT 1501.170 0.155 1503.550 4.280 ;
        RECT 1504.390 0.155 1506.770 4.280 ;
        RECT 1507.610 0.155 1513.210 4.280 ;
        RECT 1514.050 0.155 1516.430 4.280 ;
        RECT 1517.270 0.155 1519.650 4.280 ;
        RECT 1520.490 0.155 1522.870 4.280 ;
        RECT 1523.710 0.155 1526.090 4.280 ;
        RECT 1526.930 0.155 1529.310 4.280 ;
        RECT 1530.150 0.155 1535.750 4.280 ;
        RECT 1536.590 0.155 1538.970 4.280 ;
        RECT 1539.810 0.155 1542.190 4.280 ;
        RECT 1543.030 0.155 1545.410 4.280 ;
        RECT 1546.250 0.155 1548.630 4.280 ;
        RECT 1549.470 0.155 1555.070 4.280 ;
        RECT 1555.910 0.155 1558.290 4.280 ;
        RECT 1559.130 0.155 1561.510 4.280 ;
        RECT 1562.350 0.155 1564.730 4.280 ;
        RECT 1565.570 0.155 1567.950 4.280 ;
        RECT 1568.790 0.155 1571.170 4.280 ;
        RECT 1572.010 0.155 1577.610 4.280 ;
        RECT 1578.450 0.155 1580.830 4.280 ;
        RECT 1581.670 0.155 1584.050 4.280 ;
        RECT 1584.890 0.155 1587.270 4.280 ;
        RECT 1588.110 0.155 1590.490 4.280 ;
        RECT 1591.330 0.155 1596.930 4.280 ;
        RECT 1597.770 0.155 1600.150 4.280 ;
        RECT 1600.990 0.155 1603.370 4.280 ;
        RECT 1604.210 0.155 1606.590 4.280 ;
        RECT 1607.430 0.155 1609.810 4.280 ;
        RECT 1610.650 0.155 1613.030 4.280 ;
        RECT 1613.870 0.155 1619.470 4.280 ;
        RECT 1620.310 0.155 1622.690 4.280 ;
        RECT 1623.530 0.155 1625.910 4.280 ;
        RECT 1626.750 0.155 1629.130 4.280 ;
        RECT 1629.970 0.155 1632.350 4.280 ;
        RECT 1633.190 0.155 1638.790 4.280 ;
        RECT 1639.630 0.155 1642.010 4.280 ;
        RECT 1642.850 0.155 1645.230 4.280 ;
        RECT 1646.070 0.155 1648.450 4.280 ;
        RECT 1649.290 0.155 1651.670 4.280 ;
        RECT 1652.510 0.155 1654.890 4.280 ;
        RECT 1655.730 0.155 1661.330 4.280 ;
        RECT 1662.170 0.155 1664.550 4.280 ;
        RECT 1665.390 0.155 1667.770 4.280 ;
        RECT 1668.610 0.155 1670.990 4.280 ;
        RECT 1671.830 0.155 1674.210 4.280 ;
        RECT 1675.050 0.155 1680.650 4.280 ;
        RECT 1681.490 0.155 1683.870 4.280 ;
        RECT 1684.710 0.155 1687.090 4.280 ;
        RECT 1687.930 0.155 1690.310 4.280 ;
        RECT 1691.150 0.155 1693.530 4.280 ;
        RECT 1694.370 0.155 1696.750 4.280 ;
        RECT 1697.590 0.155 1703.190 4.280 ;
        RECT 1704.030 0.155 1706.410 4.280 ;
        RECT 1707.250 0.155 1709.630 4.280 ;
        RECT 1710.470 0.155 1712.850 4.280 ;
        RECT 1713.690 0.155 1716.070 4.280 ;
        RECT 1716.910 0.155 1722.510 4.280 ;
        RECT 1723.350 0.155 1725.730 4.280 ;
        RECT 1726.570 0.155 1728.950 4.280 ;
        RECT 1729.790 0.155 1732.170 4.280 ;
        RECT 1733.010 0.155 1735.390 4.280 ;
        RECT 1736.230 0.155 1738.610 4.280 ;
        RECT 1739.450 0.155 1745.050 4.280 ;
        RECT 1745.890 0.155 1748.270 4.280 ;
        RECT 1749.110 0.155 1751.490 4.280 ;
        RECT 1752.330 0.155 1754.710 4.280 ;
        RECT 1755.550 0.155 1757.930 4.280 ;
        RECT 1758.770 0.155 1764.370 4.280 ;
        RECT 1765.210 0.155 1767.590 4.280 ;
        RECT 1768.430 0.155 1770.810 4.280 ;
        RECT 1771.650 0.155 1774.030 4.280 ;
        RECT 1774.870 0.155 1777.250 4.280 ;
        RECT 1778.090 0.155 1780.470 4.280 ;
        RECT 1781.310 0.155 1786.910 4.280 ;
        RECT 1787.750 0.155 1790.130 4.280 ;
        RECT 1790.970 0.155 1793.350 4.280 ;
        RECT 1794.190 0.155 1796.570 4.280 ;
        RECT 1797.410 0.155 1799.790 4.280 ;
        RECT 1800.630 0.155 1806.230 4.280 ;
        RECT 1807.070 0.155 1809.450 4.280 ;
        RECT 1810.290 0.155 1812.670 4.280 ;
        RECT 1813.510 0.155 1815.890 4.280 ;
        RECT 1816.730 0.155 1819.110 4.280 ;
        RECT 1819.950 0.155 1822.330 4.280 ;
        RECT 1823.170 0.155 1828.770 4.280 ;
        RECT 1829.610 0.155 1831.990 4.280 ;
        RECT 1832.830 0.155 1835.210 4.280 ;
        RECT 1836.050 0.155 1838.430 4.280 ;
        RECT 1839.270 0.155 1841.650 4.280 ;
        RECT 1842.490 0.155 1844.870 4.280 ;
        RECT 1845.710 0.155 1851.310 4.280 ;
        RECT 1852.150 0.155 1854.530 4.280 ;
        RECT 1855.370 0.155 1857.750 4.280 ;
        RECT 1858.590 0.155 1860.970 4.280 ;
        RECT 1861.810 0.155 1864.190 4.280 ;
        RECT 1865.030 0.155 1870.630 4.280 ;
        RECT 1871.470 0.155 1873.850 4.280 ;
        RECT 1874.690 0.155 1877.070 4.280 ;
        RECT 1877.910 0.155 1880.290 4.280 ;
        RECT 1881.130 0.155 1883.510 4.280 ;
        RECT 1884.350 0.155 1886.730 4.280 ;
        RECT 1887.570 0.155 1893.170 4.280 ;
        RECT 1894.010 0.155 1896.390 4.280 ;
        RECT 1897.230 0.155 1899.610 4.280 ;
        RECT 1900.450 0.155 1902.830 4.280 ;
        RECT 1903.670 0.155 1906.050 4.280 ;
        RECT 1906.890 0.155 1912.490 4.280 ;
        RECT 1913.330 0.155 1915.710 4.280 ;
        RECT 1916.550 0.155 1918.930 4.280 ;
        RECT 1919.770 0.155 1922.150 4.280 ;
        RECT 1922.990 0.155 1925.370 4.280 ;
        RECT 1926.210 0.155 1928.590 4.280 ;
        RECT 1929.430 0.155 1935.030 4.280 ;
        RECT 1935.870 0.155 1938.250 4.280 ;
        RECT 1939.090 0.155 1941.470 4.280 ;
        RECT 1942.310 0.155 1944.690 4.280 ;
        RECT 1945.530 0.155 1947.910 4.280 ;
        RECT 1948.750 0.155 1954.350 4.280 ;
        RECT 1955.190 0.155 1957.570 4.280 ;
        RECT 1958.410 0.155 1960.790 4.280 ;
        RECT 1961.630 0.155 1964.010 4.280 ;
        RECT 1964.850 0.155 1967.230 4.280 ;
        RECT 1968.070 0.155 1970.450 4.280 ;
        RECT 1971.290 0.155 1976.890 4.280 ;
        RECT 1977.730 0.155 1980.110 4.280 ;
        RECT 1980.950 0.155 1983.330 4.280 ;
        RECT 1984.170 0.155 1986.550 4.280 ;
        RECT 1987.390 0.155 1989.770 4.280 ;
        RECT 1990.610 0.155 1996.210 4.280 ;
        RECT 1997.050 0.155 1999.430 4.280 ;
        RECT 2000.270 0.155 2002.650 4.280 ;
        RECT 2003.490 0.155 2005.870 4.280 ;
        RECT 2006.710 0.155 2009.090 4.280 ;
        RECT 2009.930 0.155 2012.310 4.280 ;
        RECT 2013.150 0.155 2018.750 4.280 ;
        RECT 2019.590 0.155 2021.970 4.280 ;
        RECT 2022.810 0.155 2025.190 4.280 ;
        RECT 2026.030 0.155 2028.410 4.280 ;
        RECT 2029.250 0.155 2031.630 4.280 ;
        RECT 2032.470 0.155 2038.070 4.280 ;
        RECT 2038.910 0.155 2041.290 4.280 ;
        RECT 2042.130 0.155 2044.510 4.280 ;
        RECT 2045.350 0.155 2047.730 4.280 ;
        RECT 2048.570 0.155 2050.950 4.280 ;
        RECT 2051.790 0.155 2054.170 4.280 ;
        RECT 2055.010 0.155 2060.610 4.280 ;
        RECT 2061.450 0.155 2063.830 4.280 ;
        RECT 2064.670 0.155 2067.050 4.280 ;
        RECT 2067.890 0.155 2070.270 4.280 ;
        RECT 2071.110 0.155 2073.490 4.280 ;
        RECT 2074.330 0.155 2079.930 4.280 ;
        RECT 2080.770 0.155 2083.150 4.280 ;
        RECT 2083.990 0.155 2086.370 4.280 ;
        RECT 2087.210 0.155 2089.590 4.280 ;
        RECT 2090.430 0.155 2092.810 4.280 ;
        RECT 2093.650 0.155 2096.030 4.280 ;
        RECT 2096.870 0.155 2102.470 4.280 ;
        RECT 2103.310 0.155 2105.690 4.280 ;
        RECT 2106.530 0.155 2108.910 4.280 ;
        RECT 2109.750 0.155 2112.130 4.280 ;
        RECT 2112.970 0.155 2115.350 4.280 ;
        RECT 2116.190 0.155 2121.790 4.280 ;
        RECT 2122.630 0.155 2125.010 4.280 ;
        RECT 2125.850 0.155 2128.230 4.280 ;
        RECT 2129.070 0.155 2131.450 4.280 ;
        RECT 2132.290 0.155 2134.670 4.280 ;
        RECT 2135.510 0.155 2137.890 4.280 ;
        RECT 2138.730 0.155 2144.330 4.280 ;
        RECT 2145.170 0.155 2147.550 4.280 ;
        RECT 2148.390 0.155 2150.770 4.280 ;
        RECT 2151.610 0.155 2153.990 4.280 ;
        RECT 2154.830 0.155 2157.210 4.280 ;
        RECT 2158.050 0.155 2163.650 4.280 ;
        RECT 2164.490 0.155 2166.870 4.280 ;
        RECT 2167.710 0.155 2170.090 4.280 ;
        RECT 2170.930 0.155 2173.310 4.280 ;
        RECT 2174.150 0.155 2176.530 4.280 ;
        RECT 2177.370 0.155 2179.750 4.280 ;
        RECT 2180.590 0.155 2186.190 4.280 ;
        RECT 2187.030 0.155 2189.410 4.280 ;
        RECT 2190.250 0.155 2192.630 4.280 ;
        RECT 2193.470 0.155 2195.850 4.280 ;
        RECT 2196.690 0.155 2199.070 4.280 ;
        RECT 2199.910 0.155 2205.510 4.280 ;
        RECT 2206.350 0.155 2208.730 4.280 ;
        RECT 2209.570 0.155 2211.950 4.280 ;
        RECT 2212.790 0.155 2215.170 4.280 ;
        RECT 2216.010 0.155 2218.390 4.280 ;
        RECT 2219.230 0.155 2221.610 4.280 ;
        RECT 2222.450 0.155 2228.050 4.280 ;
        RECT 2228.890 0.155 2231.270 4.280 ;
        RECT 2232.110 0.155 2234.490 4.280 ;
        RECT 2235.330 0.155 2237.710 4.280 ;
        RECT 2238.550 0.155 2240.930 4.280 ;
        RECT 2241.770 0.155 2247.370 4.280 ;
        RECT 2248.210 0.155 2250.590 4.280 ;
        RECT 2251.430 0.155 2253.810 4.280 ;
        RECT 2254.650 0.155 2257.030 4.280 ;
        RECT 2257.870 0.155 2260.250 4.280 ;
        RECT 2261.090 0.155 2263.470 4.280 ;
        RECT 2264.310 0.155 2269.910 4.280 ;
        RECT 2270.750 0.155 2273.130 4.280 ;
        RECT 2273.970 0.155 2276.350 4.280 ;
        RECT 2277.190 0.155 2279.570 4.280 ;
        RECT 2280.410 0.155 2282.790 4.280 ;
        RECT 2283.630 0.155 2286.010 4.280 ;
        RECT 2286.850 0.155 2292.450 4.280 ;
        RECT 2293.290 0.155 2295.670 4.280 ;
        RECT 2296.510 0.155 2298.890 4.280 ;
        RECT 2299.730 0.155 2302.110 4.280 ;
        RECT 2302.950 0.155 2305.330 4.280 ;
        RECT 2306.170 0.155 2311.770 4.280 ;
        RECT 2312.610 0.155 2314.990 4.280 ;
        RECT 2315.830 0.155 2318.210 4.280 ;
        RECT 2319.050 0.155 2321.430 4.280 ;
        RECT 2322.270 0.155 2324.650 4.280 ;
        RECT 2325.490 0.155 2327.870 4.280 ;
        RECT 2328.710 0.155 2334.310 4.280 ;
        RECT 2335.150 0.155 2337.530 4.280 ;
        RECT 2338.370 0.155 2340.750 4.280 ;
        RECT 2341.590 0.155 2343.970 4.280 ;
        RECT 2344.810 0.155 2347.190 4.280 ;
        RECT 2348.030 0.155 2353.630 4.280 ;
        RECT 2354.470 0.155 2356.850 4.280 ;
        RECT 2357.690 0.155 2360.070 4.280 ;
        RECT 2360.910 0.155 2363.290 4.280 ;
        RECT 2364.130 0.155 2366.510 4.280 ;
        RECT 2367.350 0.155 2369.730 4.280 ;
        RECT 2370.570 0.155 2376.170 4.280 ;
        RECT 2377.010 0.155 2379.390 4.280 ;
        RECT 2380.230 0.155 2382.610 4.280 ;
        RECT 2383.450 0.155 2385.830 4.280 ;
        RECT 2386.670 0.155 2389.050 4.280 ;
        RECT 2389.890 0.155 2395.490 4.280 ;
        RECT 2396.330 0.155 2398.710 4.280 ;
      LAYER met3 ;
        RECT 4.000 598.040 2395.600 598.905 ;
        RECT 4.000 596.040 2396.000 598.040 ;
        RECT 4.400 594.640 2395.600 596.040 ;
        RECT 4.000 592.640 2396.000 594.640 ;
        RECT 4.400 591.240 2395.600 592.640 ;
        RECT 4.000 589.240 2396.000 591.240 ;
        RECT 4.400 587.840 2396.000 589.240 ;
        RECT 4.000 585.840 2396.000 587.840 ;
        RECT 4.400 584.440 2395.600 585.840 ;
        RECT 4.000 582.440 2396.000 584.440 ;
        RECT 4.400 581.040 2395.600 582.440 ;
        RECT 4.000 579.040 2396.000 581.040 ;
        RECT 4.400 577.640 2395.600 579.040 ;
        RECT 4.000 575.640 2396.000 577.640 ;
        RECT 4.000 574.240 2395.600 575.640 ;
        RECT 4.000 572.240 2396.000 574.240 ;
        RECT 4.400 570.840 2395.600 572.240 ;
        RECT 4.000 568.840 2396.000 570.840 ;
        RECT 4.400 567.440 2396.000 568.840 ;
        RECT 4.000 565.440 2396.000 567.440 ;
        RECT 4.400 564.040 2395.600 565.440 ;
        RECT 4.000 562.040 2396.000 564.040 ;
        RECT 4.400 560.640 2395.600 562.040 ;
        RECT 4.000 558.640 2396.000 560.640 ;
        RECT 4.400 557.240 2395.600 558.640 ;
        RECT 4.000 555.240 2396.000 557.240 ;
        RECT 4.000 553.840 2395.600 555.240 ;
        RECT 4.000 551.840 2396.000 553.840 ;
        RECT 4.400 550.440 2395.600 551.840 ;
        RECT 4.000 548.440 2396.000 550.440 ;
        RECT 4.400 547.040 2395.600 548.440 ;
        RECT 4.000 545.040 2396.000 547.040 ;
        RECT 4.400 543.640 2396.000 545.040 ;
        RECT 4.000 541.640 2396.000 543.640 ;
        RECT 4.400 540.240 2395.600 541.640 ;
        RECT 4.000 538.240 2396.000 540.240 ;
        RECT 4.400 536.840 2395.600 538.240 ;
        RECT 4.000 534.840 2396.000 536.840 ;
        RECT 4.400 533.440 2395.600 534.840 ;
        RECT 4.000 531.440 2396.000 533.440 ;
        RECT 4.000 530.040 2395.600 531.440 ;
        RECT 4.000 528.040 2396.000 530.040 ;
        RECT 4.400 526.640 2395.600 528.040 ;
        RECT 4.000 524.640 2396.000 526.640 ;
        RECT 4.400 523.240 2396.000 524.640 ;
        RECT 4.000 521.240 2396.000 523.240 ;
        RECT 4.400 519.840 2395.600 521.240 ;
        RECT 4.000 517.840 2396.000 519.840 ;
        RECT 4.400 516.440 2395.600 517.840 ;
        RECT 4.000 514.440 2396.000 516.440 ;
        RECT 4.400 513.040 2395.600 514.440 ;
        RECT 4.000 511.040 2396.000 513.040 ;
        RECT 4.000 509.640 2395.600 511.040 ;
        RECT 4.000 507.640 2396.000 509.640 ;
        RECT 4.400 506.240 2395.600 507.640 ;
        RECT 4.000 504.240 2396.000 506.240 ;
        RECT 4.400 502.840 2395.600 504.240 ;
        RECT 4.000 500.840 2396.000 502.840 ;
        RECT 4.400 499.440 2396.000 500.840 ;
        RECT 4.000 497.440 2396.000 499.440 ;
        RECT 4.400 496.040 2395.600 497.440 ;
        RECT 4.000 494.040 2396.000 496.040 ;
        RECT 4.400 492.640 2395.600 494.040 ;
        RECT 4.000 490.640 2396.000 492.640 ;
        RECT 4.400 489.240 2395.600 490.640 ;
        RECT 4.000 487.240 2396.000 489.240 ;
        RECT 4.000 485.840 2395.600 487.240 ;
        RECT 4.000 483.840 2396.000 485.840 ;
        RECT 4.400 482.440 2395.600 483.840 ;
        RECT 4.000 480.440 2396.000 482.440 ;
        RECT 4.400 479.040 2396.000 480.440 ;
        RECT 4.000 477.040 2396.000 479.040 ;
        RECT 4.400 475.640 2395.600 477.040 ;
        RECT 4.000 473.640 2396.000 475.640 ;
        RECT 4.400 472.240 2395.600 473.640 ;
        RECT 4.000 470.240 2396.000 472.240 ;
        RECT 4.400 468.840 2395.600 470.240 ;
        RECT 4.000 466.840 2396.000 468.840 ;
        RECT 4.400 465.440 2395.600 466.840 ;
        RECT 4.000 463.440 2396.000 465.440 ;
        RECT 4.000 462.040 2395.600 463.440 ;
        RECT 4.000 460.040 2396.000 462.040 ;
        RECT 4.400 458.640 2395.600 460.040 ;
        RECT 4.000 456.640 2396.000 458.640 ;
        RECT 4.400 455.240 2396.000 456.640 ;
        RECT 4.000 453.240 2396.000 455.240 ;
        RECT 4.400 451.840 2395.600 453.240 ;
        RECT 4.000 449.840 2396.000 451.840 ;
        RECT 4.400 448.440 2395.600 449.840 ;
        RECT 4.000 446.440 2396.000 448.440 ;
        RECT 4.400 445.040 2395.600 446.440 ;
        RECT 4.000 443.040 2396.000 445.040 ;
        RECT 4.000 441.640 2395.600 443.040 ;
        RECT 4.000 439.640 2396.000 441.640 ;
        RECT 4.400 438.240 2395.600 439.640 ;
        RECT 4.000 436.240 2396.000 438.240 ;
        RECT 4.400 434.840 2396.000 436.240 ;
        RECT 4.000 432.840 2396.000 434.840 ;
        RECT 4.400 431.440 2395.600 432.840 ;
        RECT 4.000 429.440 2396.000 431.440 ;
        RECT 4.400 428.040 2395.600 429.440 ;
        RECT 4.000 426.040 2396.000 428.040 ;
        RECT 4.400 424.640 2395.600 426.040 ;
        RECT 4.000 422.640 2396.000 424.640 ;
        RECT 4.400 421.240 2395.600 422.640 ;
        RECT 4.000 419.240 2396.000 421.240 ;
        RECT 4.000 417.840 2395.600 419.240 ;
        RECT 4.000 415.840 2396.000 417.840 ;
        RECT 4.400 414.440 2395.600 415.840 ;
        RECT 4.000 412.440 2396.000 414.440 ;
        RECT 4.400 411.040 2396.000 412.440 ;
        RECT 4.000 409.040 2396.000 411.040 ;
        RECT 4.400 407.640 2395.600 409.040 ;
        RECT 4.000 405.640 2396.000 407.640 ;
        RECT 4.400 404.240 2395.600 405.640 ;
        RECT 4.000 402.240 2396.000 404.240 ;
        RECT 4.400 400.840 2395.600 402.240 ;
        RECT 4.000 398.840 2396.000 400.840 ;
        RECT 4.000 397.440 2395.600 398.840 ;
        RECT 4.000 395.440 2396.000 397.440 ;
        RECT 4.400 394.040 2395.600 395.440 ;
        RECT 4.000 392.040 2396.000 394.040 ;
        RECT 4.400 390.640 2396.000 392.040 ;
        RECT 4.000 388.640 2396.000 390.640 ;
        RECT 4.400 387.240 2395.600 388.640 ;
        RECT 4.000 385.240 2396.000 387.240 ;
        RECT 4.400 383.840 2395.600 385.240 ;
        RECT 4.000 381.840 2396.000 383.840 ;
        RECT 4.400 380.440 2395.600 381.840 ;
        RECT 4.000 378.440 2396.000 380.440 ;
        RECT 4.400 377.040 2395.600 378.440 ;
        RECT 4.000 375.040 2396.000 377.040 ;
        RECT 4.000 373.640 2395.600 375.040 ;
        RECT 4.000 371.640 2396.000 373.640 ;
        RECT 4.400 370.240 2395.600 371.640 ;
        RECT 4.000 368.240 2396.000 370.240 ;
        RECT 4.400 366.840 2396.000 368.240 ;
        RECT 4.000 364.840 2396.000 366.840 ;
        RECT 4.400 363.440 2395.600 364.840 ;
        RECT 4.000 361.440 2396.000 363.440 ;
        RECT 4.400 360.040 2395.600 361.440 ;
        RECT 4.000 358.040 2396.000 360.040 ;
        RECT 4.400 356.640 2395.600 358.040 ;
        RECT 4.000 354.640 2396.000 356.640 ;
        RECT 4.000 353.240 2395.600 354.640 ;
        RECT 4.000 351.240 2396.000 353.240 ;
        RECT 4.400 349.840 2395.600 351.240 ;
        RECT 4.000 347.840 2396.000 349.840 ;
        RECT 4.400 346.440 2395.600 347.840 ;
        RECT 4.000 344.440 2396.000 346.440 ;
        RECT 4.400 343.040 2396.000 344.440 ;
        RECT 4.000 341.040 2396.000 343.040 ;
        RECT 4.400 339.640 2395.600 341.040 ;
        RECT 4.000 337.640 2396.000 339.640 ;
        RECT 4.400 336.240 2395.600 337.640 ;
        RECT 4.000 334.240 2396.000 336.240 ;
        RECT 4.400 332.840 2395.600 334.240 ;
        RECT 4.000 330.840 2396.000 332.840 ;
        RECT 4.000 329.440 2395.600 330.840 ;
        RECT 4.000 327.440 2396.000 329.440 ;
        RECT 4.400 326.040 2395.600 327.440 ;
        RECT 4.000 324.040 2396.000 326.040 ;
        RECT 4.400 322.640 2396.000 324.040 ;
        RECT 4.000 320.640 2396.000 322.640 ;
        RECT 4.400 319.240 2395.600 320.640 ;
        RECT 4.000 317.240 2396.000 319.240 ;
        RECT 4.400 315.840 2395.600 317.240 ;
        RECT 4.000 313.840 2396.000 315.840 ;
        RECT 4.400 312.440 2395.600 313.840 ;
        RECT 4.000 310.440 2396.000 312.440 ;
        RECT 4.000 309.040 2395.600 310.440 ;
        RECT 4.000 307.040 2396.000 309.040 ;
        RECT 4.400 305.640 2395.600 307.040 ;
        RECT 4.000 303.640 2396.000 305.640 ;
        RECT 4.400 302.240 2395.600 303.640 ;
        RECT 4.000 300.240 2396.000 302.240 ;
        RECT 4.400 298.840 2396.000 300.240 ;
        RECT 4.000 296.840 2396.000 298.840 ;
        RECT 4.400 295.440 2395.600 296.840 ;
        RECT 4.000 293.440 2396.000 295.440 ;
        RECT 4.400 292.040 2395.600 293.440 ;
        RECT 4.000 290.040 2396.000 292.040 ;
        RECT 4.400 288.640 2395.600 290.040 ;
        RECT 4.000 286.640 2396.000 288.640 ;
        RECT 4.000 285.240 2395.600 286.640 ;
        RECT 4.000 283.240 2396.000 285.240 ;
        RECT 4.400 281.840 2395.600 283.240 ;
        RECT 4.000 279.840 2396.000 281.840 ;
        RECT 4.400 278.440 2396.000 279.840 ;
        RECT 4.000 276.440 2396.000 278.440 ;
        RECT 4.400 275.040 2395.600 276.440 ;
        RECT 4.000 273.040 2396.000 275.040 ;
        RECT 4.400 271.640 2395.600 273.040 ;
        RECT 4.000 269.640 2396.000 271.640 ;
        RECT 4.400 268.240 2395.600 269.640 ;
        RECT 4.000 266.240 2396.000 268.240 ;
        RECT 4.000 264.840 2395.600 266.240 ;
        RECT 4.000 262.840 2396.000 264.840 ;
        RECT 4.400 261.440 2395.600 262.840 ;
        RECT 4.000 259.440 2396.000 261.440 ;
        RECT 4.400 258.040 2395.600 259.440 ;
        RECT 4.000 256.040 2396.000 258.040 ;
        RECT 4.400 254.640 2396.000 256.040 ;
        RECT 4.000 252.640 2396.000 254.640 ;
        RECT 4.400 251.240 2395.600 252.640 ;
        RECT 4.000 249.240 2396.000 251.240 ;
        RECT 4.400 247.840 2395.600 249.240 ;
        RECT 4.000 245.840 2396.000 247.840 ;
        RECT 4.400 244.440 2395.600 245.840 ;
        RECT 4.000 242.440 2396.000 244.440 ;
        RECT 4.000 241.040 2395.600 242.440 ;
        RECT 4.000 239.040 2396.000 241.040 ;
        RECT 4.400 237.640 2395.600 239.040 ;
        RECT 4.000 235.640 2396.000 237.640 ;
        RECT 4.400 234.240 2396.000 235.640 ;
        RECT 4.000 232.240 2396.000 234.240 ;
        RECT 4.400 230.840 2395.600 232.240 ;
        RECT 4.000 228.840 2396.000 230.840 ;
        RECT 4.400 227.440 2395.600 228.840 ;
        RECT 4.000 225.440 2396.000 227.440 ;
        RECT 4.400 224.040 2395.600 225.440 ;
        RECT 4.000 222.040 2396.000 224.040 ;
        RECT 4.000 220.640 2395.600 222.040 ;
        RECT 4.000 218.640 2396.000 220.640 ;
        RECT 4.400 217.240 2395.600 218.640 ;
        RECT 4.000 215.240 2396.000 217.240 ;
        RECT 4.400 213.840 2395.600 215.240 ;
        RECT 4.000 211.840 2396.000 213.840 ;
        RECT 4.400 210.440 2396.000 211.840 ;
        RECT 4.000 208.440 2396.000 210.440 ;
        RECT 4.400 207.040 2395.600 208.440 ;
        RECT 4.000 205.040 2396.000 207.040 ;
        RECT 4.400 203.640 2395.600 205.040 ;
        RECT 4.000 201.640 2396.000 203.640 ;
        RECT 4.400 200.240 2395.600 201.640 ;
        RECT 4.000 198.240 2396.000 200.240 ;
        RECT 4.000 196.840 2395.600 198.240 ;
        RECT 4.000 194.840 2396.000 196.840 ;
        RECT 4.400 193.440 2395.600 194.840 ;
        RECT 4.000 191.440 2396.000 193.440 ;
        RECT 4.400 190.040 2396.000 191.440 ;
        RECT 4.000 188.040 2396.000 190.040 ;
        RECT 4.400 186.640 2395.600 188.040 ;
        RECT 4.000 184.640 2396.000 186.640 ;
        RECT 4.400 183.240 2395.600 184.640 ;
        RECT 4.000 181.240 2396.000 183.240 ;
        RECT 4.400 179.840 2395.600 181.240 ;
        RECT 4.000 177.840 2396.000 179.840 ;
        RECT 4.000 176.440 2395.600 177.840 ;
        RECT 4.000 174.440 2396.000 176.440 ;
        RECT 4.400 173.040 2395.600 174.440 ;
        RECT 4.000 171.040 2396.000 173.040 ;
        RECT 4.400 169.640 2395.600 171.040 ;
        RECT 4.000 167.640 2396.000 169.640 ;
        RECT 4.400 166.240 2396.000 167.640 ;
        RECT 4.000 164.240 2396.000 166.240 ;
        RECT 4.400 162.840 2395.600 164.240 ;
        RECT 4.000 160.840 2396.000 162.840 ;
        RECT 4.400 159.440 2395.600 160.840 ;
        RECT 4.000 157.440 2396.000 159.440 ;
        RECT 4.400 156.040 2395.600 157.440 ;
        RECT 4.000 154.040 2396.000 156.040 ;
        RECT 4.000 152.640 2395.600 154.040 ;
        RECT 4.000 150.640 2396.000 152.640 ;
        RECT 4.400 149.240 2395.600 150.640 ;
        RECT 4.000 147.240 2396.000 149.240 ;
        RECT 4.400 145.840 2396.000 147.240 ;
        RECT 4.000 143.840 2396.000 145.840 ;
        RECT 4.400 142.440 2395.600 143.840 ;
        RECT 4.000 140.440 2396.000 142.440 ;
        RECT 4.400 139.040 2395.600 140.440 ;
        RECT 4.000 137.040 2396.000 139.040 ;
        RECT 4.400 135.640 2395.600 137.040 ;
        RECT 4.000 133.640 2396.000 135.640 ;
        RECT 4.000 132.240 2395.600 133.640 ;
        RECT 4.000 130.240 2396.000 132.240 ;
        RECT 4.400 128.840 2395.600 130.240 ;
        RECT 4.000 126.840 2396.000 128.840 ;
        RECT 4.400 125.440 2395.600 126.840 ;
        RECT 4.000 123.440 2396.000 125.440 ;
        RECT 4.400 122.040 2396.000 123.440 ;
        RECT 4.000 120.040 2396.000 122.040 ;
        RECT 4.400 118.640 2395.600 120.040 ;
        RECT 4.000 116.640 2396.000 118.640 ;
        RECT 4.400 115.240 2395.600 116.640 ;
        RECT 4.000 113.240 2396.000 115.240 ;
        RECT 4.400 111.840 2395.600 113.240 ;
        RECT 4.000 109.840 2396.000 111.840 ;
        RECT 4.000 108.440 2395.600 109.840 ;
        RECT 4.000 106.440 2396.000 108.440 ;
        RECT 4.400 105.040 2395.600 106.440 ;
        RECT 4.000 103.040 2396.000 105.040 ;
        RECT 4.400 101.640 2396.000 103.040 ;
        RECT 4.000 99.640 2396.000 101.640 ;
        RECT 4.400 98.240 2395.600 99.640 ;
        RECT 4.000 96.240 2396.000 98.240 ;
        RECT 4.400 94.840 2395.600 96.240 ;
        RECT 4.000 92.840 2396.000 94.840 ;
        RECT 4.400 91.440 2395.600 92.840 ;
        RECT 4.000 89.440 2396.000 91.440 ;
        RECT 4.000 88.040 2395.600 89.440 ;
        RECT 4.000 86.040 2396.000 88.040 ;
        RECT 4.400 84.640 2395.600 86.040 ;
        RECT 4.000 82.640 2396.000 84.640 ;
        RECT 4.400 81.240 2395.600 82.640 ;
        RECT 4.000 79.240 2396.000 81.240 ;
        RECT 4.400 77.840 2396.000 79.240 ;
        RECT 4.000 75.840 2396.000 77.840 ;
        RECT 4.400 74.440 2395.600 75.840 ;
        RECT 4.000 72.440 2396.000 74.440 ;
        RECT 4.400 71.040 2395.600 72.440 ;
        RECT 4.000 69.040 2396.000 71.040 ;
        RECT 4.400 67.640 2395.600 69.040 ;
        RECT 4.000 65.640 2396.000 67.640 ;
        RECT 4.000 64.240 2395.600 65.640 ;
        RECT 4.000 62.240 2396.000 64.240 ;
        RECT 4.400 60.840 2395.600 62.240 ;
        RECT 4.000 58.840 2396.000 60.840 ;
        RECT 4.400 57.440 2396.000 58.840 ;
        RECT 4.000 55.440 2396.000 57.440 ;
        RECT 4.400 54.040 2395.600 55.440 ;
        RECT 4.000 52.040 2396.000 54.040 ;
        RECT 4.400 50.640 2395.600 52.040 ;
        RECT 4.000 48.640 2396.000 50.640 ;
        RECT 4.400 47.240 2395.600 48.640 ;
        RECT 4.000 45.240 2396.000 47.240 ;
        RECT 4.000 43.840 2395.600 45.240 ;
        RECT 4.000 41.840 2396.000 43.840 ;
        RECT 4.400 40.440 2395.600 41.840 ;
        RECT 4.000 38.440 2396.000 40.440 ;
        RECT 4.400 37.040 2395.600 38.440 ;
        RECT 4.000 35.040 2396.000 37.040 ;
        RECT 4.400 33.640 2396.000 35.040 ;
        RECT 4.000 31.640 2396.000 33.640 ;
        RECT 4.400 30.240 2395.600 31.640 ;
        RECT 4.000 28.240 2396.000 30.240 ;
        RECT 4.400 26.840 2395.600 28.240 ;
        RECT 4.000 24.840 2396.000 26.840 ;
        RECT 4.400 23.440 2395.600 24.840 ;
        RECT 4.000 21.440 2396.000 23.440 ;
        RECT 4.000 20.040 2395.600 21.440 ;
        RECT 4.000 18.040 2396.000 20.040 ;
        RECT 4.400 16.640 2395.600 18.040 ;
        RECT 4.000 14.640 2396.000 16.640 ;
        RECT 4.400 13.240 2396.000 14.640 ;
        RECT 4.000 11.240 2396.000 13.240 ;
        RECT 4.400 9.840 2395.600 11.240 ;
        RECT 4.000 7.840 2396.000 9.840 ;
        RECT 4.400 6.440 2395.600 7.840 ;
        RECT 4.000 4.440 2396.000 6.440 ;
        RECT 4.400 3.040 2395.600 4.440 ;
        RECT 4.000 1.040 2396.000 3.040 ;
        RECT 4.000 0.175 2395.600 1.040 ;
      LAYER met4 ;
        RECT 849.455 10.240 865.440 586.665 ;
        RECT 867.840 10.240 942.240 586.665 ;
        RECT 944.640 10.240 1019.040 586.665 ;
        RECT 1021.440 10.240 1095.840 586.665 ;
        RECT 1098.240 10.240 1172.640 586.665 ;
        RECT 1175.040 10.240 1249.440 586.665 ;
        RECT 1251.840 10.240 1326.240 586.665 ;
        RECT 1328.640 10.240 1403.040 586.665 ;
        RECT 1405.440 10.240 1479.840 586.665 ;
        RECT 1482.240 10.240 1556.640 586.665 ;
        RECT 1559.040 10.240 1632.705 586.665 ;
        RECT 849.455 8.335 1632.705 10.240 ;
  END
END axi_node_intf_wrap
END LIBRARY

