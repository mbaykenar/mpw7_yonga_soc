magic
tech sky130B
magscale 12 1
timestamp 1598777896
<< metal5 >>
rect 0 60 45 75
rect 20 45 45 60
rect 15 40 40 45
rect 10 35 35 40
rect 5 30 30 35
rect 0 15 25 30
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
