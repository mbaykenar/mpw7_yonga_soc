module boot_code (
	CLK,
	RSTN,
	CSN,
	A,
	Q
);
	input wire CLK;
	input wire RSTN;
	input wire CSN;
	input wire [9:0] A;
	output wire [31:0] Q;
	reg [17535:0] mem = 17536'h130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130100006f0100006f0080006f0040006f0000006f0000009300008113000081930000821300008293000083130000839300008413000084930000851300008593000086130000869300008713000087930000881300008893000089130000899300008a1300008a9300008b1300008b9300008c1300008c9300008d1300008d9300008e1300008e9300008f1300008f9300100117ef41011300000d177f8d0d1300000d977f0d8d9301bd5863000d2023004d0d13ffaddce30000051300000593072000ef000000000000000000000000000000004681110145a1460109f0051300efce060513362000ef040045813b6000ef45014581396000ef450100283de004000593420000ef55134722157d0187de8717b32190071300a0353300e788630761670937b38f99953e00f0610540f2715d8082c6864505c2a6c4a2de4ec0cada56dc52d65ed85ad266d46200efd06a458525a000ef450167854460bb8787930037c0fb0001000127b74711c3d81a10f65ff0ef8537c911059300000513024000ef7185a001476000008537051345c500ef740545a146604601468100ef451945012a602fc000ef4505458132c000ef358000ef10055433fe143ce380000637069345a1061302000513348600ef0710450127602cc000ef852245812fc000ef328000ef10055533fe153ce345214581298000ef0200069345a146010eb00513244000ef10000513298000ef450945812c8000ef1000059300ef850a853730a045d500007545051349024cb244c24c124b724ad23c4000ef4521458124c000ef07905e6349816421412c0c3300008bb77b04041300008a3716136d050693008945a102000eb005131dc000ef00ef65214581232000ef45090533262065a1012c2a4000ef8513459900ef76cbd51336e04585004900ef9522b53336204585f64900ef9522098535600513459900ef774a996a34a0388000effb3c91e324c000ef10055533fe153ce300008537051345b500ef77c500ef32604581366000ef45215e631aa064210760409a89b38bb74901041300008a377b046a8500000084961302000693051345a100ef0eb0652113a0190000ef450945811c0000ef0099853300ef65a14599202076cb85132cc000ef00495513952245852c0000eff6493533952245852b4000ef45990905774a05132a8000ef00ef94d611e32e608537fb2b059300000513022000ef78c500ef28e077b72ce0a4231a1007930007806708000001000700010001450140b64496442659f249065ad25a625bb25b425c925c2261615d0200008082ff01011300812423000005930005041300f0051300112623294000ef0000059300e00513288000ef0000059300d0051327c000ef0000059300c00513270000ef048056630000059301000513260000ef02142e630000059300b00513250000ef022426630000059300000513240000ef00342e6300c12083008124030000059300100513010101132240006f00c1208300812403010101130000806700004837f008081300869693020007131a1027b740b707330106f6b3f265b5b300e515330087881300c7871300b6e5b30107879300a8202300c7202300b7a02300008067010595931005553300a5e5b31a1027b700b7aa23000080671a1027370107071300072783ff01011300f1262300c127831007d7b30105151300f5653300a1262300c1278300f720230101011300008067001007930085859300b795b300a79533000017b7f007879300f5f5b3ee85353300a5e5331a1027b700a7a023000080671a1027b70007a783ff01011300f1262300c125030101011300008067d45597b3ff010113f455b5b300f1242300058863008127830017879300f124230001262300c126831a102737008127830207081302f6de6300072783cf0797b3fe078ce300c127830008258300c126830016869300d126230101061300279793ffc626030081268300b567a3fcd646e301010113000080671a10773700470713000726031a1007b7c016463300c720230047869300c785130085d813083007130ff5f59300e520230106a0230a70071300b7a42b00e7a0230030079300f520230006a7830f07f793c017c7b300f6a023000080671a100737014707130205886304000693000727830207f793fe078ce30015460b1a1007b7fff5859300c7a023fff6869300069663fc059ce300008067fc059ae3000080671a10073701470713000727830407f793fe078ce3000080671a1076b70006a783ff01011300f126230010079300a797b300c12703fff7c79300e7f7b300f1262300c1278300a595b300f5e53300a1262300c1278300f6a02301010113000080674f52524553203a52736e6170206e6f692049505373616c666f6e20686f6620740a646e750000000064616f4c20676e696d6f7266495053200000000a79706f4320676e6974736e4974637572736e6f690000000a636f6c420000206b6e6f642000000a6579706f4320676e69617461440000000a656e6f44756a202c6e69706d6f742067736e4920637572746e6f69744d41522000000a2e33323130373635344241393846454443000000100000000000527a010101040100020d1b0000001400000018fffff9740000005e200e42007f01114c0000003800000030fffff9ba00000274500e42007f01115a117e081112117d097b13117c117a14111611791577171178117618111a11751900000074000000180000006cfffffbf40000009c100e44007e0811487f01114c0000001000000088fffffc740000004400000000000000100000009cfffffca4000000180000000000000010000000b0fffffca800000038100e500000000010000000c4fffffccc00000030;
	reg [9:0] A_Q;
	always @(posedge CLK or negedge RSTN)
		if (~RSTN)
			A_Q <= 1'sb0;
		else if (~CSN)
			A_Q <= A;
	assign Q = mem[(547 - A_Q) * 32+:32];
endmodule
