magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -42 452 316 1184
<< pwell >>
rect -2 -6 276 246
<< mvnmos >>
rect 77 20 197 220
<< mvpmos >>
rect 77 518 197 1118
<< mvndiff >>
rect 24 208 77 220
rect 24 174 32 208
rect 66 174 77 208
rect 24 140 77 174
rect 24 106 32 140
rect 66 106 77 140
rect 24 72 77 106
rect 24 38 32 72
rect 66 38 77 72
rect 24 20 77 38
rect 197 208 250 220
rect 197 174 208 208
rect 242 174 250 208
rect 197 140 250 174
rect 197 106 208 140
rect 242 106 250 140
rect 197 72 250 106
rect 197 38 208 72
rect 242 38 250 72
rect 197 20 250 38
<< mvpdiff >>
rect 24 1106 77 1118
rect 24 1072 32 1106
rect 66 1072 77 1106
rect 24 1038 77 1072
rect 24 1004 32 1038
rect 66 1004 77 1038
rect 24 970 77 1004
rect 24 936 32 970
rect 66 936 77 970
rect 24 902 77 936
rect 24 868 32 902
rect 66 868 77 902
rect 24 834 77 868
rect 24 800 32 834
rect 66 800 77 834
rect 24 766 77 800
rect 24 732 32 766
rect 66 732 77 766
rect 24 698 77 732
rect 24 664 32 698
rect 66 664 77 698
rect 24 630 77 664
rect 24 596 32 630
rect 66 596 77 630
rect 24 518 77 596
rect 197 1106 250 1118
rect 197 1072 208 1106
rect 242 1072 250 1106
rect 197 1038 250 1072
rect 197 1004 208 1038
rect 242 1004 250 1038
rect 197 970 250 1004
rect 197 936 208 970
rect 242 936 250 970
rect 197 902 250 936
rect 197 868 208 902
rect 242 868 250 902
rect 197 834 250 868
rect 197 800 208 834
rect 242 800 250 834
rect 197 766 250 800
rect 197 732 208 766
rect 242 732 250 766
rect 197 698 250 732
rect 197 664 208 698
rect 242 664 250 698
rect 197 630 250 664
rect 197 596 208 630
rect 242 596 250 630
rect 197 518 250 596
<< mvndiffc >>
rect 32 174 66 208
rect 32 106 66 140
rect 32 38 66 72
rect 208 174 242 208
rect 208 106 242 140
rect 208 38 242 72
<< mvpdiffc >>
rect 32 1072 66 1106
rect 32 1004 66 1038
rect 32 936 66 970
rect 32 868 66 902
rect 32 800 66 834
rect 32 732 66 766
rect 32 664 66 698
rect 32 596 66 630
rect 208 1072 242 1106
rect 208 1004 242 1038
rect 208 936 242 970
rect 208 868 242 902
rect 208 800 242 834
rect 208 732 242 766
rect 208 664 242 698
rect 208 596 242 630
<< poly >>
rect 77 1118 197 1144
rect 77 418 197 518
rect 77 384 116 418
rect 150 384 197 418
rect 77 350 197 384
rect 77 316 116 350
rect 150 316 197 350
rect 77 220 197 316
rect 77 -6 197 20
<< polycont >>
rect 116 384 150 418
rect 116 316 150 350
<< locali >>
rect 32 1152 66 1192
rect 32 1106 66 1118
rect 32 1038 66 1046
rect 32 970 66 1004
rect 32 902 66 936
rect 32 834 66 868
rect 32 766 66 800
rect 32 698 66 732
rect 32 630 66 664
rect 32 580 66 596
rect 208 1106 270 1122
rect 242 1072 270 1106
rect 208 1038 270 1072
rect 242 1004 270 1038
rect 208 970 270 1004
rect 242 936 270 970
rect 208 902 270 936
rect 242 868 270 902
rect 208 834 270 868
rect 242 800 270 834
rect 208 766 270 800
rect 242 732 270 766
rect 208 698 270 732
rect 242 664 270 698
rect 208 630 270 664
rect 242 596 270 630
rect 100 384 116 418
rect 150 384 166 418
rect 100 350 166 384
rect 100 316 116 350
rect 150 316 166 350
rect 32 208 66 224
rect 32 140 66 174
rect 32 75 66 106
rect 32 3 66 38
rect 208 208 270 596
rect 242 174 270 208
rect 208 140 270 174
rect 242 106 270 140
rect 208 72 270 106
rect 242 38 270 72
rect 208 22 270 38
rect 32 -69 66 -31
<< viali >>
rect 32 1118 66 1152
rect 32 1072 66 1080
rect 32 1046 66 1072
rect 32 72 66 75
rect 32 41 66 72
rect 32 -31 66 3
rect 32 -103 66 -69
<< metal1 >>
rect -47 1152 314 1292
rect -47 1118 32 1152
rect 66 1118 314 1152
rect -47 1080 314 1118
rect -47 1046 32 1080
rect 66 1046 314 1080
rect -47 1034 314 1046
rect -47 75 314 87
rect -47 41 32 75
rect 66 41 314 75
rect -47 3 314 41
rect -47 -31 32 3
rect 66 -31 314 3
rect -47 -69 314 -31
rect -47 -103 32 -69
rect 66 -103 314 -69
rect -47 -115 314 -103
use sky130_fd_pr__model__nfet_highvoltage__example_5595914180899  sky130_fd_pr__model__nfet_highvoltage__example_5595914180899_0
timestamp 1649977179
transform 1 0 77 0 -1 220
box -28 0 148 97
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808101  sky130_fd_pr__model__pfet_highvoltage__example_55959141808101_0
timestamp 1649977179
transform 1 0 77 0 -1 1118
box -28 0 148 267
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1649977179
transform 0 -1 66 -1 0 1152
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1649977179
transform 0 -1 66 -1 0 75
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1649977179
transform 0 -1 166 1 0 300
box 0 0 1 1
<< properties >>
string GDS_END 37315268
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37314438
<< end >>
