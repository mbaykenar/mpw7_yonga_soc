magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< locali >>
rect 159 752 171 786
rect 205 752 243 786
rect 277 752 315 786
rect 349 752 387 786
rect 421 752 459 786
rect 493 752 505 786
rect 48 672 82 674
rect 48 600 82 638
rect 48 528 82 566
rect 48 456 82 494
rect 48 384 82 422
rect 48 312 82 350
rect 48 240 82 278
rect 48 168 82 206
rect 48 132 82 134
rect 582 672 616 674
rect 582 600 616 638
rect 582 528 616 566
rect 582 456 616 494
rect 582 384 616 422
rect 582 312 616 350
rect 582 240 616 278
rect 582 168 616 206
rect 582 132 616 134
rect 159 20 171 54
rect 205 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 505 54
<< viali >>
rect 171 752 205 786
rect 243 752 277 786
rect 315 752 349 786
rect 387 752 421 786
rect 459 752 493 786
rect 48 638 82 672
rect 48 566 82 600
rect 48 494 82 528
rect 48 422 82 456
rect 48 350 82 384
rect 48 278 82 312
rect 48 206 82 240
rect 48 134 82 168
rect 582 638 616 672
rect 582 566 616 600
rect 582 494 616 528
rect 582 422 616 456
rect 582 350 616 384
rect 582 278 616 312
rect 582 206 616 240
rect 582 134 616 168
rect 171 20 205 54
rect 243 20 277 54
rect 315 20 349 54
rect 387 20 421 54
rect 459 20 493 54
<< obsli1 >>
rect 159 98 193 708
rect 315 98 349 708
rect 471 98 505 708
<< metal1 >>
rect 159 786 505 806
rect 159 752 171 786
rect 205 752 243 786
rect 277 752 315 786
rect 349 752 387 786
rect 421 752 459 786
rect 493 752 505 786
rect 159 740 505 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 570 672 628 684
rect 570 638 582 672
rect 616 638 628 672
rect 570 600 628 638
rect 570 566 582 600
rect 616 566 628 600
rect 570 528 628 566
rect 570 494 582 528
rect 616 494 628 528
rect 570 456 628 494
rect 570 422 582 456
rect 616 422 628 456
rect 570 384 628 422
rect 570 350 582 384
rect 616 350 628 384
rect 570 312 628 350
rect 570 278 582 312
rect 616 278 628 312
rect 570 240 628 278
rect 570 206 582 240
rect 616 206 628 240
rect 570 168 628 206
rect 570 134 582 168
rect 616 134 628 168
rect 570 122 628 134
rect 159 54 505 66
rect 159 20 171 54
rect 205 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 505 54
rect 159 0 505 20
<< obsm1 >>
rect 150 122 202 684
rect 306 122 358 684
rect 462 122 514 684
<< metal2 >>
rect 10 428 654 684
rect 10 122 654 378
<< labels >>
rlabel viali s 582 638 616 672 6 BULK
port 1 nsew
rlabel viali s 582 566 616 600 6 BULK
port 1 nsew
rlabel viali s 582 494 616 528 6 BULK
port 1 nsew
rlabel viali s 582 422 616 456 6 BULK
port 1 nsew
rlabel viali s 582 350 616 384 6 BULK
port 1 nsew
rlabel viali s 582 278 616 312 6 BULK
port 1 nsew
rlabel viali s 582 206 616 240 6 BULK
port 1 nsew
rlabel viali s 582 134 616 168 6 BULK
port 1 nsew
rlabel viali s 48 638 82 672 6 BULK
port 1 nsew
rlabel viali s 48 566 82 600 6 BULK
port 1 nsew
rlabel viali s 48 494 82 528 6 BULK
port 1 nsew
rlabel viali s 48 422 82 456 6 BULK
port 1 nsew
rlabel viali s 48 350 82 384 6 BULK
port 1 nsew
rlabel viali s 48 278 82 312 6 BULK
port 1 nsew
rlabel viali s 48 206 82 240 6 BULK
port 1 nsew
rlabel viali s 48 134 82 168 6 BULK
port 1 nsew
rlabel locali s 582 132 616 674 6 BULK
port 1 nsew
rlabel locali s 48 132 82 674 6 BULK
port 1 nsew
rlabel metal1 s 570 122 628 684 6 BULK
port 1 nsew
rlabel metal1 s 36 122 94 684 6 BULK
port 1 nsew
rlabel metal2 s 10 428 654 684 6 DRAIN
port 2 nsew
rlabel viali s 459 752 493 786 6 GATE
port 3 nsew
rlabel viali s 459 20 493 54 6 GATE
port 3 nsew
rlabel viali s 387 752 421 786 6 GATE
port 3 nsew
rlabel viali s 387 20 421 54 6 GATE
port 3 nsew
rlabel viali s 315 752 349 786 6 GATE
port 3 nsew
rlabel viali s 315 20 349 54 6 GATE
port 3 nsew
rlabel viali s 243 752 277 786 6 GATE
port 3 nsew
rlabel viali s 243 20 277 54 6 GATE
port 3 nsew
rlabel viali s 171 752 205 786 6 GATE
port 3 nsew
rlabel viali s 171 20 205 54 6 GATE
port 3 nsew
rlabel locali s 159 752 505 786 6 GATE
port 3 nsew
rlabel locali s 159 20 505 54 6 GATE
port 3 nsew
rlabel metal1 s 159 740 505 806 6 GATE
port 3 nsew
rlabel metal1 s 159 0 505 66 6 GATE
port 3 nsew
rlabel metal2 s 10 122 654 378 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 664 806
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9894844
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9883352
<< end >>
