magic
tech sky130B
magscale 12 1
timestamp 1598769117
<< metal5 >>
rect 0 55 15 105
rect 30 55 45 105
rect 0 45 45 55
rect 5 30 40 45
rect 10 15 35 30
rect 15 0 30 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
