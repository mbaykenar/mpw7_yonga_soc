magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 16 49 661 263
rect 0 0 672 49
<< scnmos >>
rect 95 69 125 237
rect 181 69 211 237
rect 267 69 297 237
rect 345 69 375 237
rect 491 69 521 237
<< scpmoshvt >>
rect 95 367 125 619
rect 173 367 203 619
rect 263 367 293 619
rect 349 367 379 619
rect 562 367 592 619
<< ndiff >>
rect 42 192 95 237
rect 42 158 50 192
rect 84 158 95 192
rect 42 115 95 158
rect 42 81 50 115
rect 84 81 95 115
rect 42 69 95 81
rect 125 208 181 237
rect 125 174 136 208
rect 170 174 181 208
rect 125 117 181 174
rect 125 83 136 117
rect 170 83 181 117
rect 125 69 181 83
rect 211 132 267 237
rect 211 98 222 132
rect 256 98 267 132
rect 211 69 267 98
rect 297 69 345 237
rect 375 229 491 237
rect 375 195 424 229
rect 458 195 491 229
rect 375 153 491 195
rect 375 119 424 153
rect 458 119 491 153
rect 375 69 491 119
rect 521 196 635 237
rect 521 162 593 196
rect 627 162 635 196
rect 521 115 635 162
rect 521 81 593 115
rect 627 81 635 115
rect 521 69 635 81
<< pdiff >>
rect 401 621 451 639
rect 401 619 409 621
rect 42 599 95 619
rect 42 565 50 599
rect 84 565 95 599
rect 42 525 95 565
rect 42 491 50 525
rect 84 491 95 525
rect 42 447 95 491
rect 42 413 50 447
rect 84 413 95 447
rect 42 367 95 413
rect 125 367 173 619
rect 203 607 263 619
rect 203 573 214 607
rect 248 573 263 607
rect 203 531 263 573
rect 203 497 214 531
rect 248 497 263 531
rect 203 367 263 497
rect 293 607 349 619
rect 293 573 304 607
rect 338 573 349 607
rect 293 515 349 573
rect 293 481 304 515
rect 338 481 349 515
rect 293 367 349 481
rect 379 587 409 619
rect 443 587 451 621
rect 379 367 451 587
rect 505 409 562 619
rect 505 375 517 409
rect 551 375 562 409
rect 505 367 562 375
rect 592 569 645 619
rect 592 535 603 569
rect 637 535 645 569
rect 592 367 645 535
<< ndiffc >>
rect 50 158 84 192
rect 50 81 84 115
rect 136 174 170 208
rect 136 83 170 117
rect 222 98 256 132
rect 424 195 458 229
rect 424 119 458 153
rect 593 162 627 196
rect 593 81 627 115
<< pdiffc >>
rect 50 565 84 599
rect 50 491 84 525
rect 50 413 84 447
rect 214 573 248 607
rect 214 497 248 531
rect 304 573 338 607
rect 304 481 338 515
rect 409 587 443 621
rect 517 375 551 409
rect 603 535 637 569
<< poly >>
rect 95 619 125 645
rect 173 619 203 645
rect 263 619 293 645
rect 349 619 379 645
rect 562 619 592 645
rect 95 325 125 367
rect 173 325 203 367
rect 263 325 293 367
rect 349 335 379 367
rect 25 309 125 325
rect 25 275 41 309
rect 75 275 125 309
rect 25 259 125 275
rect 167 309 301 325
rect 167 275 183 309
rect 217 275 251 309
rect 285 275 301 309
rect 167 259 301 275
rect 345 319 439 335
rect 345 285 389 319
rect 423 285 439 319
rect 562 325 592 367
rect 562 309 647 325
rect 562 289 597 309
rect 345 269 439 285
rect 491 275 597 289
rect 631 275 647 309
rect 95 237 125 259
rect 181 237 211 259
rect 267 237 297 259
rect 345 237 375 269
rect 491 259 647 275
rect 491 237 521 259
rect 95 43 125 69
rect 181 43 211 69
rect 267 43 297 69
rect 345 43 375 69
rect 491 43 521 69
<< polycont >>
rect 41 275 75 309
rect 183 275 217 309
rect 251 275 285 309
rect 389 285 423 319
rect 597 275 631 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 34 599 100 615
rect 34 565 50 599
rect 84 565 100 599
rect 34 525 100 565
rect 34 491 50 525
rect 84 491 100 525
rect 34 447 100 491
rect 198 607 254 649
rect 393 621 459 649
rect 198 573 214 607
rect 248 573 254 607
rect 198 531 254 573
rect 198 497 214 531
rect 248 497 254 531
rect 198 481 254 497
rect 288 607 354 615
rect 288 573 304 607
rect 338 573 354 607
rect 393 587 409 621
rect 443 587 459 621
rect 393 583 459 587
rect 288 549 354 573
rect 587 569 653 585
rect 587 549 603 569
rect 288 535 603 549
rect 637 535 653 569
rect 288 515 653 535
rect 288 481 304 515
rect 338 481 354 515
rect 388 447 647 481
rect 34 413 50 447
rect 84 413 422 447
rect 501 409 567 413
rect 17 345 423 379
rect 501 375 517 409
rect 551 375 567 409
rect 501 359 567 375
rect 501 350 547 359
rect 17 309 91 345
rect 387 319 423 345
rect 17 275 41 309
rect 75 275 91 309
rect 17 242 91 275
rect 125 309 353 311
rect 125 275 183 309
rect 217 275 251 309
rect 285 275 353 309
rect 125 242 353 275
rect 387 285 389 319
rect 387 269 423 285
rect 457 314 547 350
rect 613 325 647 447
rect 457 233 491 314
rect 581 309 647 325
rect 581 280 597 309
rect 408 229 491 233
rect 34 192 86 208
rect 34 158 50 192
rect 84 158 86 192
rect 34 115 86 158
rect 34 81 50 115
rect 84 81 86 115
rect 34 17 86 81
rect 120 174 136 208
rect 170 174 374 208
rect 120 117 172 174
rect 120 83 136 117
rect 170 83 172 117
rect 120 67 172 83
rect 206 132 272 140
rect 206 98 222 132
rect 256 98 272 132
rect 206 17 272 98
rect 340 85 374 174
rect 408 195 424 229
rect 458 195 491 229
rect 408 153 491 195
rect 408 119 424 153
rect 458 119 491 153
rect 525 275 597 280
rect 631 275 647 309
rect 525 246 647 275
rect 525 85 559 246
rect 340 51 559 85
rect 593 196 643 212
rect 627 162 643 196
rect 593 115 643 162
rect 627 81 643 115
rect 593 17 643 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 1 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 2 nsew
rlabel comment s 0 0 0 0 4 SKY130_FD_IO__XOR2_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 3 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 5 nsew
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 5 nsew
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 5 nsew
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 6 nsew
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 6 nsew
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_END 8529162
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8523180
<< end >>
