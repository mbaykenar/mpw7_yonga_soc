magic
tech sky130B
magscale 12 1
timestamp 1598776997
<< metal5 >>
rect 0 70 35 75
rect 0 65 40 70
rect 0 55 45 65
rect 0 0 15 55
rect 30 0 45 55
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
