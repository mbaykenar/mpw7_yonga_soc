magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -66 377 1986 897
<< pwell >>
rect 1650 217 1916 283
rect 6 43 1916 217
rect -26 -43 1946 43
<< mvnmos >>
rect 89 107 189 191
rect 245 107 345 191
rect 519 107 619 191
rect 675 107 775 191
rect 817 107 917 191
rect 996 107 1096 191
rect 1138 107 1238 191
rect 1412 107 1512 191
rect 1554 107 1654 191
rect 1733 107 1833 257
<< mvpmos >>
rect 89 564 189 714
rect 245 564 345 714
rect 519 491 619 641
rect 675 491 775 641
rect 817 491 917 641
rect 996 491 1096 575
rect 1138 491 1238 575
rect 1317 443 1417 593
rect 1473 443 1573 593
rect 1652 443 1752 743
<< mvndiff >>
rect 1676 249 1733 257
rect 1676 215 1688 249
rect 1722 215 1733 249
rect 1676 191 1733 215
rect 32 166 89 191
rect 32 132 44 166
rect 78 132 89 166
rect 32 107 89 132
rect 189 166 245 191
rect 189 132 200 166
rect 234 132 245 166
rect 189 107 245 132
rect 345 166 402 191
rect 345 132 356 166
rect 390 132 402 166
rect 345 107 402 132
rect 462 166 519 191
rect 462 132 474 166
rect 508 132 519 166
rect 462 107 519 132
rect 619 154 675 191
rect 619 120 630 154
rect 664 120 675 154
rect 619 107 675 120
rect 775 107 817 191
rect 917 166 996 191
rect 917 132 951 166
rect 985 132 996 166
rect 917 107 996 132
rect 1096 107 1138 191
rect 1238 166 1295 191
rect 1238 132 1249 166
rect 1283 132 1295 166
rect 1238 107 1295 132
rect 1355 166 1412 191
rect 1355 132 1367 166
rect 1401 132 1412 166
rect 1355 107 1412 132
rect 1512 107 1554 191
rect 1654 149 1733 191
rect 1654 115 1688 149
rect 1722 115 1733 149
rect 1654 107 1733 115
rect 1833 249 1890 257
rect 1833 215 1844 249
rect 1878 215 1890 249
rect 1833 149 1890 215
rect 1833 115 1844 149
rect 1878 115 1890 149
rect 1833 107 1890 115
<< mvpdiff >>
rect 1595 735 1652 743
rect 32 706 89 714
rect 32 672 44 706
rect 78 672 89 706
rect 32 606 89 672
rect 32 572 44 606
rect 78 572 89 606
rect 32 564 89 572
rect 189 706 245 714
rect 189 672 200 706
rect 234 672 245 706
rect 189 606 245 672
rect 189 572 200 606
rect 234 572 245 606
rect 189 564 245 572
rect 345 706 402 714
rect 345 672 356 706
rect 390 672 402 706
rect 345 606 402 672
rect 1595 701 1607 735
rect 1641 701 1652 735
rect 1595 661 1652 701
rect 345 572 356 606
rect 390 572 402 606
rect 345 564 402 572
rect 462 633 519 641
rect 462 599 474 633
rect 508 599 519 633
rect 462 533 519 599
rect 462 499 474 533
rect 508 499 519 533
rect 462 491 519 499
rect 619 606 675 641
rect 619 572 630 606
rect 664 572 675 606
rect 619 491 675 572
rect 775 491 817 641
rect 917 606 974 641
rect 1595 627 1607 661
rect 1641 627 1652 661
rect 917 572 928 606
rect 962 575 974 606
rect 1595 593 1652 627
rect 1260 585 1317 593
rect 1260 575 1272 585
rect 962 572 996 575
rect 917 491 996 572
rect 1096 491 1138 575
rect 1238 551 1272 575
rect 1306 551 1317 585
rect 1238 491 1317 551
rect 1260 485 1317 491
rect 1260 451 1272 485
rect 1306 451 1317 485
rect 1260 443 1317 451
rect 1417 585 1473 593
rect 1417 551 1428 585
rect 1462 551 1473 585
rect 1417 485 1473 551
rect 1417 451 1428 485
rect 1462 451 1473 485
rect 1417 443 1473 451
rect 1573 585 1652 593
rect 1573 551 1607 585
rect 1641 551 1652 585
rect 1573 511 1652 551
rect 1573 477 1607 511
rect 1641 477 1652 511
rect 1573 443 1652 477
rect 1752 735 1809 743
rect 1752 701 1763 735
rect 1797 701 1809 735
rect 1752 652 1809 701
rect 1752 618 1763 652
rect 1797 618 1809 652
rect 1752 568 1809 618
rect 1752 534 1763 568
rect 1797 534 1809 568
rect 1752 485 1809 534
rect 1752 451 1763 485
rect 1797 451 1809 485
rect 1752 443 1809 451
<< mvndiffc >>
rect 1688 215 1722 249
rect 44 132 78 166
rect 200 132 234 166
rect 356 132 390 166
rect 474 132 508 166
rect 630 120 664 154
rect 951 132 985 166
rect 1249 132 1283 166
rect 1367 132 1401 166
rect 1688 115 1722 149
rect 1844 215 1878 249
rect 1844 115 1878 149
<< mvpdiffc >>
rect 44 672 78 706
rect 44 572 78 606
rect 200 672 234 706
rect 200 572 234 606
rect 356 672 390 706
rect 1607 701 1641 735
rect 356 572 390 606
rect 474 599 508 633
rect 474 499 508 533
rect 630 572 664 606
rect 1607 627 1641 661
rect 928 572 962 606
rect 1272 551 1306 585
rect 1272 451 1306 485
rect 1428 551 1462 585
rect 1428 451 1462 485
rect 1607 551 1641 585
rect 1607 477 1641 511
rect 1763 701 1797 735
rect 1763 618 1797 652
rect 1763 534 1797 568
rect 1763 451 1797 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
<< poly >>
rect 1652 743 1752 769
rect 89 714 189 740
rect 245 714 345 740
rect 519 641 619 667
rect 675 641 775 667
rect 817 641 917 667
rect 89 504 189 564
rect 89 470 130 504
rect 164 470 189 504
rect 89 436 189 470
rect 89 402 130 436
rect 164 402 189 436
rect 89 191 189 402
rect 245 275 345 564
rect 996 575 1096 601
rect 1138 575 1238 601
rect 1317 593 1417 619
rect 1473 593 1573 619
rect 245 241 265 275
rect 299 241 345 275
rect 245 191 345 241
rect 519 439 619 491
rect 519 405 539 439
rect 573 405 619 439
rect 519 191 619 405
rect 675 389 775 491
rect 661 369 775 389
rect 661 335 681 369
rect 715 335 775 369
rect 661 289 775 335
rect 817 439 917 491
rect 996 469 1096 491
rect 817 405 837 439
rect 871 405 917 439
rect 817 371 917 405
rect 965 443 1096 469
rect 965 409 985 443
rect 1019 409 1096 443
rect 965 393 1096 409
rect 1138 411 1238 491
rect 817 337 837 371
rect 871 351 917 371
rect 1138 377 1178 411
rect 1212 377 1238 411
rect 871 337 1096 351
rect 817 321 1096 337
rect 675 191 775 289
rect 817 263 917 279
rect 817 229 851 263
rect 885 229 917 263
rect 817 191 917 229
rect 996 191 1096 321
rect 1138 343 1238 377
rect 1317 361 1417 443
rect 1138 309 1178 343
rect 1212 309 1238 343
rect 1138 191 1238 309
rect 1286 341 1417 361
rect 1286 307 1306 341
rect 1340 307 1417 341
rect 1473 371 1573 443
rect 1473 337 1519 371
rect 1553 337 1573 371
rect 1473 321 1573 337
rect 1652 421 1752 443
rect 1652 383 1833 421
rect 1652 349 1676 383
rect 1710 349 1833 383
rect 1652 321 1833 349
rect 1286 279 1417 307
rect 1286 273 1512 279
rect 1286 239 1306 273
rect 1340 239 1512 273
rect 1286 213 1512 239
rect 1412 191 1512 213
rect 1554 263 1654 279
rect 1554 229 1574 263
rect 1608 229 1654 263
rect 1733 257 1833 321
rect 1554 191 1654 229
rect 89 81 189 107
rect 245 81 345 107
rect 519 81 619 107
rect 675 81 775 107
rect 817 81 917 107
rect 996 81 1096 107
rect 1138 81 1238 107
rect 1412 81 1512 107
rect 1554 81 1654 107
rect 1733 81 1833 107
<< polycont >>
rect 130 470 164 504
rect 130 402 164 436
rect 265 241 299 275
rect 539 405 573 439
rect 681 335 715 369
rect 837 405 871 439
rect 985 409 1019 443
rect 837 337 871 371
rect 1178 377 1212 411
rect 851 229 885 263
rect 1178 309 1212 343
rect 1306 307 1340 341
rect 1519 337 1553 371
rect 1676 349 1710 383
rect 1306 239 1340 273
rect 1574 229 1608 263
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 114 735 304 741
rect 28 706 78 722
rect 28 672 44 706
rect 28 606 78 672
rect 28 572 44 606
rect 28 350 78 572
rect 114 701 120 735
rect 154 701 192 735
rect 226 706 264 735
rect 234 701 264 706
rect 298 701 304 735
rect 560 735 750 741
rect 114 672 200 701
rect 234 672 304 701
rect 114 606 304 672
rect 114 572 200 606
rect 234 572 304 606
rect 114 556 304 572
rect 340 706 406 722
rect 340 672 356 706
rect 390 672 406 706
rect 340 606 406 672
rect 560 701 566 735
rect 600 701 638 735
rect 672 701 710 735
rect 744 701 750 735
rect 340 572 356 606
rect 390 572 406 606
rect 114 504 180 520
rect 114 470 130 504
rect 164 470 180 504
rect 114 436 180 470
rect 114 402 130 436
rect 164 402 180 436
rect 340 439 406 572
rect 458 633 524 649
rect 458 599 474 633
rect 508 599 524 633
rect 458 533 524 599
rect 560 606 750 701
rect 1141 735 1331 741
rect 1141 701 1147 735
rect 1181 701 1219 735
rect 1253 701 1291 735
rect 1325 701 1331 735
rect 560 572 630 606
rect 664 572 750 606
rect 560 545 750 572
rect 912 606 978 649
rect 912 572 928 606
rect 962 579 978 606
rect 1141 585 1331 701
rect 1514 735 1704 751
rect 1514 701 1520 735
rect 1554 701 1592 735
rect 1641 701 1664 735
rect 1698 701 1704 735
rect 1514 661 1704 701
rect 1514 627 1607 661
rect 1641 627 1704 661
rect 962 572 1105 579
rect 912 545 1105 572
rect 458 499 474 533
rect 508 509 524 533
rect 508 499 957 509
rect 458 475 957 499
rect 923 459 957 475
rect 923 443 1035 459
rect 340 405 539 439
rect 573 405 837 439
rect 871 405 887 439
rect 114 386 180 402
rect 767 371 887 405
rect 325 350 681 369
rect 28 335 681 350
rect 715 335 731 369
rect 767 337 837 371
rect 871 337 887 371
rect 28 316 359 335
rect 767 321 887 337
rect 923 409 985 443
rect 1019 409 1035 443
rect 923 393 1035 409
rect 28 166 78 316
rect 767 299 801 321
rect 121 275 359 280
rect 121 241 265 275
rect 299 241 359 275
rect 121 235 359 241
rect 395 265 801 299
rect 923 279 957 393
rect 395 199 429 265
rect 837 263 957 279
rect 1071 269 1105 545
rect 1141 551 1272 585
rect 1306 551 1331 585
rect 1141 485 1331 551
rect 1141 451 1272 485
rect 1306 451 1331 485
rect 1392 585 1478 601
rect 1392 551 1428 585
rect 1462 551 1478 585
rect 1392 485 1478 551
rect 1392 451 1428 485
rect 1462 451 1478 485
rect 1514 585 1704 627
rect 1514 551 1607 585
rect 1641 551 1704 585
rect 1514 511 1704 551
rect 1514 477 1607 511
rect 1641 477 1704 511
rect 1747 735 1895 751
rect 1747 701 1763 735
rect 1797 701 1895 735
rect 1747 652 1895 701
rect 1747 618 1763 652
rect 1797 618 1895 652
rect 1747 568 1895 618
rect 1747 534 1763 568
rect 1797 534 1895 568
rect 1747 485 1895 534
rect 1392 441 1478 451
rect 1747 451 1763 485
rect 1797 451 1895 485
rect 1392 415 1694 441
rect 1747 435 1895 451
rect 1162 411 1694 415
rect 1162 377 1178 411
rect 1212 407 1694 411
rect 1212 381 1426 407
rect 1212 377 1228 381
rect 1162 343 1228 377
rect 1162 309 1178 343
rect 1212 309 1228 343
rect 1162 305 1228 309
rect 1290 341 1356 345
rect 1290 307 1306 341
rect 1340 307 1356 341
rect 1290 273 1356 307
rect 1290 269 1306 273
rect 837 229 851 263
rect 885 245 957 263
rect 885 229 899 245
rect 28 132 44 166
rect 28 99 78 132
rect 114 166 304 199
rect 114 132 200 166
rect 234 132 304 166
rect 114 113 304 132
rect 114 79 120 113
rect 154 79 192 113
rect 226 79 264 113
rect 298 79 304 113
rect 340 166 429 199
rect 340 132 356 166
rect 390 132 429 166
rect 340 99 429 132
rect 474 195 899 229
rect 993 239 1306 269
rect 1340 239 1356 273
rect 993 235 1356 239
rect 993 199 1027 235
rect 1392 199 1426 381
rect 1660 399 1694 407
rect 1660 383 1726 399
rect 474 166 524 195
rect 508 132 524 166
rect 935 166 1027 199
rect 474 99 524 132
rect 560 154 750 159
rect 560 120 630 154
rect 664 120 750 154
rect 560 113 750 120
rect 114 73 304 79
rect 560 79 566 113
rect 600 79 638 113
rect 672 79 710 113
rect 744 79 750 113
rect 935 132 951 166
rect 985 132 1027 166
rect 935 99 1027 132
rect 1109 166 1299 199
rect 1109 132 1249 166
rect 1283 132 1299 166
rect 1109 113 1299 132
rect 560 73 750 79
rect 1109 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1259 113
rect 1293 79 1299 113
rect 1351 166 1426 199
rect 1351 132 1367 166
rect 1401 132 1426 166
rect 1503 337 1519 371
rect 1553 356 1569 371
rect 1553 337 1624 356
rect 1503 263 1624 337
rect 1660 349 1676 383
rect 1710 349 1726 383
rect 1660 333 1726 349
rect 1503 229 1574 263
rect 1608 229 1624 263
rect 1503 162 1624 229
rect 1660 249 1778 265
rect 1660 215 1688 249
rect 1722 215 1778 249
rect 1351 99 1426 132
rect 1660 149 1778 215
rect 1660 115 1688 149
rect 1722 115 1778 149
rect 1660 113 1778 115
rect 1109 73 1299 79
rect 1660 79 1666 113
rect 1700 79 1738 113
rect 1772 79 1778 113
rect 1828 249 1895 435
rect 1828 215 1844 249
rect 1878 215 1895 249
rect 1828 149 1895 215
rect 1828 115 1844 149
rect 1878 115 1895 149
rect 1828 99 1895 115
rect 1660 73 1778 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 120 701 154 735
rect 192 706 226 735
rect 192 701 200 706
rect 200 701 226 706
rect 264 701 298 735
rect 566 701 600 735
rect 638 701 672 735
rect 710 701 744 735
rect 1147 701 1181 735
rect 1219 701 1253 735
rect 1291 701 1325 735
rect 1520 701 1554 735
rect 1592 701 1607 735
rect 1607 701 1626 735
rect 1664 701 1698 735
rect 120 79 154 113
rect 192 79 226 113
rect 264 79 298 113
rect 566 79 600 113
rect 638 79 672 113
rect 710 79 744 113
rect 1115 79 1149 113
rect 1187 79 1221 113
rect 1259 79 1293 113
rect 1666 79 1700 113
rect 1738 79 1772 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 831 1920 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 0 791 1920 797
rect 0 735 1920 763
rect 0 701 120 735
rect 154 701 192 735
rect 226 701 264 735
rect 298 701 566 735
rect 600 701 638 735
rect 672 701 710 735
rect 744 701 1147 735
rect 1181 701 1219 735
rect 1253 701 1291 735
rect 1325 701 1520 735
rect 1554 701 1592 735
rect 1626 701 1664 735
rect 1698 701 1920 735
rect 0 689 1920 701
rect 0 113 1920 125
rect 0 79 120 113
rect 154 79 192 113
rect 226 79 264 113
rect 298 79 566 113
rect 600 79 638 113
rect 672 79 710 113
rect 744 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1259 113
rect 1293 79 1666 113
rect 1700 79 1738 113
rect 1772 79 1920 113
rect 0 51 1920 79
rect 0 17 1920 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -23 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrtp_1
flabel metal1 s 0 51 1920 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 1920 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 1920 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 1920 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 464 1889 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 538 1889 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 612 1889 646 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
rlabel locali s 560 73 750 159 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1109 73 1299 199 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1660 73 1778 265 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 51 1920 125 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 1920 23 1 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 1920 837 1 VPB
port 6 nsew power bidirectional
rlabel locali s 560 545 750 741 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 1141 451 1331 741 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 1514 477 1704 751 1 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 689 1920 763 1 VPWR
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 1920 814
string GDS_END 1203658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1183922
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
