magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< pwell >>
rect 370 486 386 503
<< metal1 >>
rect -88 912 788 918
rect -88 860 -12 912
rect 40 860 52 912
rect 104 860 116 912
rect 168 860 180 912
rect 232 860 244 912
rect 296 860 308 912
rect 360 860 372 912
rect 424 860 436 912
rect 488 860 500 912
rect 552 860 564 912
rect 616 860 628 912
rect 680 860 788 912
rect -88 854 788 860
rect -88 809 -34 826
rect -88 757 -87 809
rect -35 757 -34 809
rect -88 745 -34 757
rect -88 693 -87 745
rect -35 693 -34 745
rect -88 681 -34 693
rect -88 629 -87 681
rect -35 629 -34 681
rect -88 617 -34 629
rect -88 565 -87 617
rect -35 565 -34 617
rect -88 553 -34 565
rect -88 501 -87 553
rect -35 501 -34 553
rect -88 489 -34 501
rect -88 437 -87 489
rect -35 437 -34 489
rect -88 425 -34 437
rect -88 373 -87 425
rect -35 373 -34 425
rect -88 361 -34 373
rect -88 309 -87 361
rect -35 309 -34 361
rect -88 297 -34 309
rect -88 245 -87 297
rect -35 245 -34 297
rect -88 233 -34 245
rect -88 181 -87 233
rect -35 181 -34 233
rect -88 169 -34 181
rect -88 117 -87 169
rect -35 117 -34 169
rect -88 105 -34 117
rect -88 53 -87 105
rect -35 64 -34 105
rect 0 64 28 826
rect 56 92 84 854
rect 112 64 140 826
rect 168 92 196 854
rect 224 64 252 826
rect 280 92 308 854
rect 336 64 364 826
rect 392 92 420 854
rect 448 64 476 826
rect 504 92 532 854
rect 560 64 588 826
rect 616 92 644 854
rect 672 64 700 826
rect 734 790 788 854
rect 734 738 735 790
rect 787 738 788 790
rect 734 726 788 738
rect 734 674 735 726
rect 787 674 788 726
rect 734 662 788 674
rect 734 610 735 662
rect 787 610 788 662
rect 734 598 788 610
rect 734 546 735 598
rect 787 546 788 598
rect 734 534 788 546
rect 734 482 735 534
rect 787 482 788 534
rect 734 470 788 482
rect 734 418 735 470
rect 787 418 788 470
rect 734 406 788 418
rect 734 354 735 406
rect 787 354 788 406
rect 734 342 788 354
rect 734 290 735 342
rect 787 290 788 342
rect 734 278 788 290
rect 734 226 735 278
rect 787 226 788 278
rect 734 214 788 226
rect 734 162 735 214
rect 787 162 788 214
rect 734 150 788 162
rect 734 98 735 150
rect 787 98 788 150
rect 734 92 788 98
rect -35 58 788 64
rect -35 53 -12 58
rect -88 6 -12 53
rect 40 6 52 58
rect 104 6 116 58
rect 168 6 180 58
rect 232 6 244 58
rect 296 6 308 58
rect 360 6 372 58
rect 424 6 436 58
rect 488 6 500 58
rect 552 6 564 58
rect 616 6 628 58
rect 680 6 788 58
rect -88 0 788 6
<< via1 >>
rect -12 860 40 912
rect 52 860 104 912
rect 116 860 168 912
rect 180 860 232 912
rect 244 860 296 912
rect 308 860 360 912
rect 372 860 424 912
rect 436 860 488 912
rect 500 860 552 912
rect 564 860 616 912
rect 628 860 680 912
rect -87 757 -35 809
rect -87 693 -35 745
rect -87 629 -35 681
rect -87 565 -35 617
rect -87 501 -35 553
rect -87 437 -35 489
rect -87 373 -35 425
rect -87 309 -35 361
rect -87 245 -35 297
rect -87 181 -35 233
rect -87 117 -35 169
rect -87 53 -35 105
rect 735 738 787 790
rect 735 674 787 726
rect 735 610 787 662
rect 735 546 787 598
rect 735 482 787 534
rect 735 418 787 470
rect 735 354 787 406
rect 735 290 787 342
rect 735 226 787 278
rect 735 162 787 214
rect 735 98 787 150
rect -12 6 40 58
rect 52 6 104 58
rect 116 6 168 58
rect 180 6 232 58
rect 244 6 296 58
rect 308 6 360 58
rect 372 6 424 58
rect 436 6 488 58
rect 500 6 552 58
rect 564 6 616 58
rect 628 6 680 58
<< metal2 >>
rect -88 912 788 918
rect -88 860 -12 912
rect 40 860 52 912
rect 104 860 116 912
rect 168 860 180 912
rect 232 860 244 912
rect 296 860 308 912
rect 360 860 372 912
rect 424 860 436 912
rect 488 860 500 912
rect 552 860 564 912
rect 616 860 628 912
rect 680 860 788 912
rect -88 854 788 860
rect -88 809 -34 826
rect -88 757 -87 809
rect -35 757 -34 809
rect -88 745 -34 757
rect -88 693 -87 745
rect -35 693 -34 745
rect -88 681 -34 693
rect -88 629 -87 681
rect -35 629 -34 681
rect -88 617 -34 629
rect -88 565 -87 617
rect -35 565 -34 617
rect -88 553 -34 565
rect -88 501 -87 553
rect -35 501 -34 553
rect -88 489 -34 501
rect -88 437 -87 489
rect -35 437 -34 489
rect -88 425 -34 437
rect -88 373 -87 425
rect -35 373 -34 425
rect -88 361 -34 373
rect -88 309 -87 361
rect -35 309 -34 361
rect -88 297 -34 309
rect -88 245 -87 297
rect -35 245 -34 297
rect -88 233 -34 245
rect -88 181 -87 233
rect -35 181 -34 233
rect -88 169 -34 181
rect -88 117 -87 169
rect -35 117 -34 169
rect -88 105 -34 117
rect -88 53 -87 105
rect -35 64 -34 105
rect 0 92 28 854
rect 56 64 84 826
rect 112 92 140 854
rect 168 64 196 826
rect 224 92 252 854
rect 280 64 308 826
rect 336 92 364 854
rect 392 64 420 826
rect 448 92 476 854
rect 504 64 532 826
rect 560 92 588 854
rect 616 64 644 826
rect 672 92 700 854
rect 734 790 788 854
rect 734 738 735 790
rect 787 738 788 790
rect 734 726 788 738
rect 734 674 735 726
rect 787 674 788 726
rect 734 662 788 674
rect 734 610 735 662
rect 787 610 788 662
rect 734 598 788 610
rect 734 546 735 598
rect 787 546 788 598
rect 734 534 788 546
rect 734 482 735 534
rect 787 482 788 534
rect 734 470 788 482
rect 734 418 735 470
rect 787 418 788 470
rect 734 406 788 418
rect 734 354 735 406
rect 787 354 788 406
rect 734 342 788 354
rect 734 290 735 342
rect 787 290 788 342
rect 734 278 788 290
rect 734 226 735 278
rect 787 226 788 278
rect 734 214 788 226
rect 734 162 735 214
rect 787 162 788 214
rect 734 150 788 162
rect 734 98 735 150
rect 787 98 788 150
rect 734 92 788 98
rect -35 58 788 64
rect -35 53 -12 58
rect -88 6 -12 53
rect 40 6 52 58
rect 104 6 116 58
rect 168 6 180 58
rect 232 6 244 58
rect 296 6 308 58
rect 360 6 372 58
rect 424 6 436 58
rect 488 6 500 58
rect 552 6 564 58
rect 616 6 628 58
rect 680 6 788 58
rect -88 0 788 6
<< labels >>
flabel comment s 355 29 355 29 0 FreeSans 200 0 0 0 For future design recommend using caps in MTM-378
flabel metal2 s 283 165 305 192 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 338 745 359 771 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 370 486 386 503 0 FreeSans 200 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 90738
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 84420
<< end >>
