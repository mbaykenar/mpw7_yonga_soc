magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< metal4 >>
rect 0 13600 200 18593
rect 0 12410 200 13300
rect 0 11240 200 12130
rect 0 10874 200 10940
rect 0 10218 200 10814
rect 0 9266 200 9862
rect 0 9140 200 9206
rect 0 7910 200 8840
rect 0 6940 200 7630
rect 0 5970 200 6660
rect 0 4760 200 5690
rect 0 3550 200 4480
rect 0 2580 200 3270
rect 0 1370 200 2300
rect 0 0 200 1090
<< obsm4 >>
rect 0 34750 200 39593
rect 0 13380 200 13520
rect 0 12210 200 12330
rect 0 11020 200 11160
rect 0 9922 200 10158
<< metal5 >>
rect 0 34750 200 39593
rect 0 13600 200 18590
rect 0 12430 200 13280
rect 0 11260 200 12110
rect 0 9140 200 10940
rect 0 7930 200 8820
rect 0 6960 200 7610
rect 0 5990 200 6640
rect 0 4780 200 5670
rect 0 3570 200 4460
rect 0 2600 200 3250
rect 0 1390 200 2280
rect 0 20 200 1070
<< labels >>
rlabel metal4 s 0 10218 200 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 200 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 9140 200 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 200 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 200 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6960 200 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6940 200 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 2600 200 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2580 200 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 5990 200 6640 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 5970 200 6660 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 0 12430 200 13280 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 12410 200 13300 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 20 200 1070 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 0 0 200 1090 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 13600 200 18590 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 13600 200 18593 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3570 200 4460 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 3550 200 4480 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 1390 200 2280 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1370 200 2300 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 4780 200 5670 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4760 200 5690 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34750 200 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 7930 200 8820 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 0 7910 200 8840 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 0 11260 200 12110 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 0 11240 200 12130 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 200 39593
string LEFclass PAD SPACER
string LEFview TRUE
string GDS_END 2305334
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2299708
<< end >>
