magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< metal1 >>
rect 13910 1399 13916 1451
rect 13968 1399 13974 1451
rect 16406 1399 16412 1451
rect 16464 1399 16470 1451
rect 18902 1399 18908 1451
rect 18960 1399 18966 1451
rect 21398 1399 21404 1451
rect 21456 1399 21462 1451
rect 23894 1399 23900 1451
rect 23952 1399 23958 1451
rect 26390 1399 26396 1451
rect 26448 1399 26454 1451
rect 28886 1399 28892 1451
rect 28944 1399 28950 1451
rect 31382 1399 31388 1451
rect 31440 1399 31446 1451
rect 33878 1399 33884 1451
rect 33936 1399 33942 1451
rect 36374 1399 36380 1451
rect 36432 1399 36438 1451
rect 38870 1399 38876 1451
rect 38928 1399 38934 1451
rect 41366 1399 41372 1451
rect 41424 1399 41430 1451
rect 43862 1399 43868 1451
rect 43920 1399 43926 1451
rect 46358 1399 46364 1451
rect 46416 1399 46422 1451
rect 48854 1399 48860 1451
rect 48912 1399 48918 1451
rect 51350 1399 51356 1451
rect 51408 1399 51414 1451
rect 53846 1399 53852 1451
rect 53904 1399 53910 1451
rect 56342 1399 56348 1451
rect 56400 1399 56406 1451
rect 58838 1399 58844 1451
rect 58896 1399 58902 1451
rect 61334 1399 61340 1451
rect 61392 1399 61398 1451
rect 63830 1399 63836 1451
rect 63888 1399 63894 1451
rect 66326 1399 66332 1451
rect 66384 1399 66390 1451
rect 68822 1399 68828 1451
rect 68880 1399 68886 1451
rect 71318 1399 71324 1451
rect 71376 1399 71382 1451
rect 73814 1399 73820 1451
rect 73872 1399 73878 1451
rect 76310 1399 76316 1451
rect 76368 1399 76374 1451
rect 78806 1399 78812 1451
rect 78864 1399 78870 1451
rect 81302 1399 81308 1451
rect 81360 1399 81366 1451
rect 83798 1399 83804 1451
rect 83856 1399 83862 1451
rect 86294 1399 86300 1451
rect 86352 1399 86358 1451
rect 88790 1399 88796 1451
rect 88848 1399 88854 1451
rect 91286 1399 91292 1451
rect 91344 1399 91350 1451
<< via1 >>
rect 13916 1399 13968 1451
rect 16412 1399 16464 1451
rect 18908 1399 18960 1451
rect 21404 1399 21456 1451
rect 23900 1399 23952 1451
rect 26396 1399 26448 1451
rect 28892 1399 28944 1451
rect 31388 1399 31440 1451
rect 33884 1399 33936 1451
rect 36380 1399 36432 1451
rect 38876 1399 38928 1451
rect 41372 1399 41424 1451
rect 43868 1399 43920 1451
rect 46364 1399 46416 1451
rect 48860 1399 48912 1451
rect 51356 1399 51408 1451
rect 53852 1399 53904 1451
rect 56348 1399 56400 1451
rect 58844 1399 58896 1451
rect 61340 1399 61392 1451
rect 63836 1399 63888 1451
rect 66332 1399 66384 1451
rect 68828 1399 68880 1451
rect 71324 1399 71376 1451
rect 73820 1399 73872 1451
rect 76316 1399 76368 1451
rect 78812 1399 78864 1451
rect 81308 1399 81360 1451
rect 83804 1399 83856 1451
rect 86300 1399 86352 1451
rect 88796 1399 88848 1451
rect 91292 1399 91344 1451
<< metal2 >>
rect 13914 1453 13970 1462
rect 13914 1388 13970 1397
rect 16410 1453 16466 1462
rect 16410 1388 16466 1397
rect 18906 1453 18962 1462
rect 18906 1388 18962 1397
rect 21402 1453 21458 1462
rect 21402 1388 21458 1397
rect 23898 1453 23954 1462
rect 23898 1388 23954 1397
rect 26394 1453 26450 1462
rect 26394 1388 26450 1397
rect 28890 1453 28946 1462
rect 28890 1388 28946 1397
rect 31386 1453 31442 1462
rect 31386 1388 31442 1397
rect 33882 1453 33938 1462
rect 33882 1388 33938 1397
rect 36378 1453 36434 1462
rect 36378 1388 36434 1397
rect 38874 1453 38930 1462
rect 38874 1388 38930 1397
rect 41370 1453 41426 1462
rect 41370 1388 41426 1397
rect 43866 1453 43922 1462
rect 43866 1388 43922 1397
rect 46362 1453 46418 1462
rect 46362 1388 46418 1397
rect 48858 1453 48914 1462
rect 48858 1388 48914 1397
rect 51354 1453 51410 1462
rect 51354 1388 51410 1397
rect 53850 1453 53906 1462
rect 53850 1388 53906 1397
rect 56346 1453 56402 1462
rect 56346 1388 56402 1397
rect 58842 1453 58898 1462
rect 58842 1388 58898 1397
rect 61338 1453 61394 1462
rect 61338 1388 61394 1397
rect 63834 1453 63890 1462
rect 63834 1388 63890 1397
rect 66330 1453 66386 1462
rect 66330 1388 66386 1397
rect 68826 1453 68882 1462
rect 68826 1388 68882 1397
rect 71322 1453 71378 1462
rect 71322 1388 71378 1397
rect 73818 1453 73874 1462
rect 73818 1388 73874 1397
rect 76314 1453 76370 1462
rect 76314 1388 76370 1397
rect 78810 1453 78866 1462
rect 78810 1388 78866 1397
rect 81306 1453 81362 1462
rect 81306 1388 81362 1397
rect 83802 1453 83858 1462
rect 83802 1388 83858 1397
rect 86298 1453 86354 1462
rect 86298 1388 86354 1397
rect 88794 1453 88850 1462
rect 88794 1388 88850 1397
rect 91290 1453 91346 1462
rect 91290 1388 91346 1397
rect 13629 333 13685 342
rect 13629 268 13685 277
rect 33597 333 33653 342
rect 33597 268 33653 277
rect 53565 333 53621 342
rect 53565 268 53621 277
rect 73533 333 73589 342
rect 73533 268 73589 277
rect 4423 -6337 4479 -6328
rect 4423 -6402 4479 -6393
rect 5591 -6337 5647 -6328
rect 5591 -6402 5647 -6393
rect 6759 -6337 6815 -6328
rect 6759 -6402 6815 -6393
rect 7927 -6337 7983 -6328
rect 7927 -6402 7983 -6393
rect 9095 -6337 9151 -6328
rect 9095 -6402 9151 -6393
rect 10263 -6337 10319 -6328
rect 10263 -6402 10319 -6393
rect 11431 -6337 11487 -6328
rect 11431 -6402 11487 -6393
rect 12599 -6337 12655 -6328
rect 12599 -6402 12655 -6393
rect 13767 -6337 13823 -6328
rect 13767 -6402 13823 -6393
rect 14935 -6337 14991 -6328
rect 14935 -6402 14991 -6393
rect 16103 -6337 16159 -6328
rect 16103 -6402 16159 -6393
rect 17271 -6337 17327 -6328
rect 17271 -6402 17327 -6393
rect 18439 -6337 18495 -6328
rect 18439 -6402 18495 -6393
rect 19607 -6337 19663 -6328
rect 19607 -6402 19663 -6393
rect 20775 -6337 20831 -6328
rect 20775 -6402 20831 -6393
rect 21943 -6337 21999 -6328
rect 21943 -6402 21999 -6393
rect 23111 -6337 23167 -6328
rect 23111 -6402 23167 -6393
rect 24279 -6337 24335 -6328
rect 24279 -6402 24335 -6393
rect 25447 -6337 25503 -6328
rect 25447 -6402 25503 -6393
rect 26615 -6337 26671 -6328
rect 26615 -6402 26671 -6393
rect 27783 -6337 27839 -6328
rect 27783 -6402 27839 -6393
rect 28951 -6337 29007 -6328
rect 28951 -6402 29007 -6393
rect 30119 -6337 30175 -6328
rect 30119 -6402 30175 -6393
rect 31287 -6337 31343 -6328
rect 31287 -6402 31343 -6393
rect 32455 -6337 32511 -6328
rect 32455 -6402 32511 -6393
rect 33623 -6337 33679 -6328
rect 33623 -6402 33679 -6393
rect 34791 -6337 34847 -6328
rect 34791 -6402 34847 -6393
rect 35959 -6337 36015 -6328
rect 35959 -6402 36015 -6393
rect 37127 -6337 37183 -6328
rect 37127 -6402 37183 -6393
rect 38295 -6337 38351 -6328
rect 38295 -6402 38351 -6393
rect 39463 -6337 39519 -6328
rect 39463 -6402 39519 -6393
rect 40631 -6337 40687 -6328
rect 40631 -6402 40687 -6393
rect 41799 -6337 41855 -6328
rect 41799 -6402 41855 -6393
rect 42967 -6337 43023 -6328
rect 42967 -6402 43023 -6393
rect 44135 -6337 44191 -6328
rect 44135 -6402 44191 -6393
rect 45303 -6337 45359 -6328
rect 45303 -6402 45359 -6393
<< via2 >>
rect 13914 1451 13970 1453
rect 13914 1399 13916 1451
rect 13916 1399 13968 1451
rect 13968 1399 13970 1451
rect 13914 1397 13970 1399
rect 16410 1451 16466 1453
rect 16410 1399 16412 1451
rect 16412 1399 16464 1451
rect 16464 1399 16466 1451
rect 16410 1397 16466 1399
rect 18906 1451 18962 1453
rect 18906 1399 18908 1451
rect 18908 1399 18960 1451
rect 18960 1399 18962 1451
rect 18906 1397 18962 1399
rect 21402 1451 21458 1453
rect 21402 1399 21404 1451
rect 21404 1399 21456 1451
rect 21456 1399 21458 1451
rect 21402 1397 21458 1399
rect 23898 1451 23954 1453
rect 23898 1399 23900 1451
rect 23900 1399 23952 1451
rect 23952 1399 23954 1451
rect 23898 1397 23954 1399
rect 26394 1451 26450 1453
rect 26394 1399 26396 1451
rect 26396 1399 26448 1451
rect 26448 1399 26450 1451
rect 26394 1397 26450 1399
rect 28890 1451 28946 1453
rect 28890 1399 28892 1451
rect 28892 1399 28944 1451
rect 28944 1399 28946 1451
rect 28890 1397 28946 1399
rect 31386 1451 31442 1453
rect 31386 1399 31388 1451
rect 31388 1399 31440 1451
rect 31440 1399 31442 1451
rect 31386 1397 31442 1399
rect 33882 1451 33938 1453
rect 33882 1399 33884 1451
rect 33884 1399 33936 1451
rect 33936 1399 33938 1451
rect 33882 1397 33938 1399
rect 36378 1451 36434 1453
rect 36378 1399 36380 1451
rect 36380 1399 36432 1451
rect 36432 1399 36434 1451
rect 36378 1397 36434 1399
rect 38874 1451 38930 1453
rect 38874 1399 38876 1451
rect 38876 1399 38928 1451
rect 38928 1399 38930 1451
rect 38874 1397 38930 1399
rect 41370 1451 41426 1453
rect 41370 1399 41372 1451
rect 41372 1399 41424 1451
rect 41424 1399 41426 1451
rect 41370 1397 41426 1399
rect 43866 1451 43922 1453
rect 43866 1399 43868 1451
rect 43868 1399 43920 1451
rect 43920 1399 43922 1451
rect 43866 1397 43922 1399
rect 46362 1451 46418 1453
rect 46362 1399 46364 1451
rect 46364 1399 46416 1451
rect 46416 1399 46418 1451
rect 46362 1397 46418 1399
rect 48858 1451 48914 1453
rect 48858 1399 48860 1451
rect 48860 1399 48912 1451
rect 48912 1399 48914 1451
rect 48858 1397 48914 1399
rect 51354 1451 51410 1453
rect 51354 1399 51356 1451
rect 51356 1399 51408 1451
rect 51408 1399 51410 1451
rect 51354 1397 51410 1399
rect 53850 1451 53906 1453
rect 53850 1399 53852 1451
rect 53852 1399 53904 1451
rect 53904 1399 53906 1451
rect 53850 1397 53906 1399
rect 56346 1451 56402 1453
rect 56346 1399 56348 1451
rect 56348 1399 56400 1451
rect 56400 1399 56402 1451
rect 56346 1397 56402 1399
rect 58842 1451 58898 1453
rect 58842 1399 58844 1451
rect 58844 1399 58896 1451
rect 58896 1399 58898 1451
rect 58842 1397 58898 1399
rect 61338 1451 61394 1453
rect 61338 1399 61340 1451
rect 61340 1399 61392 1451
rect 61392 1399 61394 1451
rect 61338 1397 61394 1399
rect 63834 1451 63890 1453
rect 63834 1399 63836 1451
rect 63836 1399 63888 1451
rect 63888 1399 63890 1451
rect 63834 1397 63890 1399
rect 66330 1451 66386 1453
rect 66330 1399 66332 1451
rect 66332 1399 66384 1451
rect 66384 1399 66386 1451
rect 66330 1397 66386 1399
rect 68826 1451 68882 1453
rect 68826 1399 68828 1451
rect 68828 1399 68880 1451
rect 68880 1399 68882 1451
rect 68826 1397 68882 1399
rect 71322 1451 71378 1453
rect 71322 1399 71324 1451
rect 71324 1399 71376 1451
rect 71376 1399 71378 1451
rect 71322 1397 71378 1399
rect 73818 1451 73874 1453
rect 73818 1399 73820 1451
rect 73820 1399 73872 1451
rect 73872 1399 73874 1451
rect 73818 1397 73874 1399
rect 76314 1451 76370 1453
rect 76314 1399 76316 1451
rect 76316 1399 76368 1451
rect 76368 1399 76370 1451
rect 76314 1397 76370 1399
rect 78810 1451 78866 1453
rect 78810 1399 78812 1451
rect 78812 1399 78864 1451
rect 78864 1399 78866 1451
rect 78810 1397 78866 1399
rect 81306 1451 81362 1453
rect 81306 1399 81308 1451
rect 81308 1399 81360 1451
rect 81360 1399 81362 1451
rect 81306 1397 81362 1399
rect 83802 1451 83858 1453
rect 83802 1399 83804 1451
rect 83804 1399 83856 1451
rect 83856 1399 83858 1451
rect 83802 1397 83858 1399
rect 86298 1451 86354 1453
rect 86298 1399 86300 1451
rect 86300 1399 86352 1451
rect 86352 1399 86354 1451
rect 86298 1397 86354 1399
rect 88794 1451 88850 1453
rect 88794 1399 88796 1451
rect 88796 1399 88848 1451
rect 88848 1399 88850 1451
rect 88794 1397 88850 1399
rect 91290 1451 91346 1453
rect 91290 1399 91292 1451
rect 91292 1399 91344 1451
rect 91344 1399 91346 1451
rect 91290 1397 91346 1399
rect 13629 277 13685 333
rect 33597 277 33653 333
rect 53565 277 53621 333
rect 73533 277 73589 333
rect 4423 -6393 4479 -6337
rect 5591 -6393 5647 -6337
rect 6759 -6393 6815 -6337
rect 7927 -6393 7983 -6337
rect 9095 -6393 9151 -6337
rect 10263 -6393 10319 -6337
rect 11431 -6393 11487 -6337
rect 12599 -6393 12655 -6337
rect 13767 -6393 13823 -6337
rect 14935 -6393 14991 -6337
rect 16103 -6393 16159 -6337
rect 17271 -6393 17327 -6337
rect 18439 -6393 18495 -6337
rect 19607 -6393 19663 -6337
rect 20775 -6393 20831 -6337
rect 21943 -6393 21999 -6337
rect 23111 -6393 23167 -6337
rect 24279 -6393 24335 -6337
rect 25447 -6393 25503 -6337
rect 26615 -6393 26671 -6337
rect 27783 -6393 27839 -6337
rect 28951 -6393 29007 -6337
rect 30119 -6393 30175 -6337
rect 31287 -6393 31343 -6337
rect 32455 -6393 32511 -6337
rect 33623 -6393 33679 -6337
rect 34791 -6393 34847 -6337
rect 35959 -6393 36015 -6337
rect 37127 -6393 37183 -6337
rect 38295 -6393 38351 -6337
rect 39463 -6393 39519 -6337
rect 40631 -6393 40687 -6337
rect 41799 -6393 41855 -6337
rect 42967 -6393 43023 -6337
rect 44135 -6393 44191 -6337
rect 45303 -6393 45359 -6337
<< metal3 >>
rect 13909 1457 13975 1458
rect 16405 1457 16471 1458
rect 18901 1457 18967 1458
rect 21397 1457 21463 1458
rect 23893 1457 23959 1458
rect 26389 1457 26455 1458
rect 28885 1457 28951 1458
rect 31381 1457 31447 1458
rect 33877 1457 33943 1458
rect 36373 1457 36439 1458
rect 38869 1457 38935 1458
rect 41365 1457 41431 1458
rect 43861 1457 43927 1458
rect 46357 1457 46423 1458
rect 48853 1457 48919 1458
rect 51349 1457 51415 1458
rect 53845 1457 53911 1458
rect 56341 1457 56407 1458
rect 58837 1457 58903 1458
rect 61333 1457 61399 1458
rect 63829 1457 63895 1458
rect 66325 1457 66391 1458
rect 68821 1457 68887 1458
rect 71317 1457 71383 1458
rect 73813 1457 73879 1458
rect 76309 1457 76375 1458
rect 78805 1457 78871 1458
rect 81301 1457 81367 1458
rect 83797 1457 83863 1458
rect 86293 1457 86359 1458
rect 88789 1457 88855 1458
rect 91285 1457 91351 1458
rect 13867 1393 13910 1457
rect 13974 1393 14017 1457
rect 16363 1393 16406 1457
rect 16470 1393 16513 1457
rect 18859 1393 18902 1457
rect 18966 1393 19009 1457
rect 21355 1393 21398 1457
rect 21462 1393 21505 1457
rect 23851 1393 23894 1457
rect 23958 1393 24001 1457
rect 26347 1393 26390 1457
rect 26454 1393 26497 1457
rect 28843 1393 28886 1457
rect 28950 1393 28993 1457
rect 31339 1393 31382 1457
rect 31446 1393 31489 1457
rect 33835 1393 33878 1457
rect 33942 1393 33985 1457
rect 36331 1393 36374 1457
rect 36438 1393 36481 1457
rect 38827 1393 38870 1457
rect 38934 1393 38977 1457
rect 41323 1393 41366 1457
rect 41430 1393 41473 1457
rect 43819 1393 43862 1457
rect 43926 1393 43969 1457
rect 46315 1393 46358 1457
rect 46422 1393 46465 1457
rect 48811 1393 48854 1457
rect 48918 1393 48961 1457
rect 51307 1393 51350 1457
rect 51414 1393 51457 1457
rect 53803 1393 53846 1457
rect 53910 1393 53953 1457
rect 56299 1393 56342 1457
rect 56406 1393 56449 1457
rect 58795 1393 58838 1457
rect 58902 1393 58945 1457
rect 61291 1393 61334 1457
rect 61398 1393 61441 1457
rect 63787 1393 63830 1457
rect 63894 1393 63937 1457
rect 66283 1393 66326 1457
rect 66390 1393 66433 1457
rect 68779 1393 68822 1457
rect 68886 1393 68929 1457
rect 71275 1393 71318 1457
rect 71382 1393 71425 1457
rect 73771 1393 73814 1457
rect 73878 1393 73921 1457
rect 76267 1393 76310 1457
rect 76374 1393 76417 1457
rect 78763 1393 78806 1457
rect 78870 1393 78913 1457
rect 81259 1393 81302 1457
rect 81366 1393 81409 1457
rect 83755 1393 83798 1457
rect 83862 1393 83905 1457
rect 86251 1393 86294 1457
rect 86358 1393 86401 1457
rect 88747 1393 88790 1457
rect 88854 1393 88897 1457
rect 91243 1393 91286 1457
rect 91350 1393 91393 1457
rect 13909 1392 13975 1393
rect 16405 1392 16471 1393
rect 18901 1392 18967 1393
rect 21397 1392 21463 1393
rect 23893 1392 23959 1393
rect 26389 1392 26455 1393
rect 28885 1392 28951 1393
rect 31381 1392 31447 1393
rect 33877 1392 33943 1393
rect 36373 1392 36439 1393
rect 38869 1392 38935 1393
rect 41365 1392 41431 1393
rect 43861 1392 43927 1393
rect 46357 1392 46423 1393
rect 48853 1392 48919 1393
rect 51349 1392 51415 1393
rect 53845 1392 53911 1393
rect 56341 1392 56407 1393
rect 58837 1392 58903 1393
rect 61333 1392 61399 1393
rect 63829 1392 63895 1393
rect 66325 1392 66391 1393
rect 68821 1392 68887 1393
rect 71317 1392 71383 1393
rect 73813 1392 73879 1393
rect 76309 1392 76375 1393
rect 78805 1392 78871 1393
rect 81301 1392 81367 1393
rect 83797 1392 83863 1393
rect 86293 1392 86359 1393
rect 88789 1392 88855 1393
rect 91285 1392 91351 1393
rect 13624 337 13690 338
rect 33592 337 33658 338
rect 53560 337 53626 338
rect 73528 337 73594 338
rect 13582 273 13625 337
rect 13689 273 13732 337
rect 33550 273 33593 337
rect 33657 273 33700 337
rect 53518 273 53561 337
rect 53625 273 53668 337
rect 73486 273 73529 337
rect 73593 273 73636 337
rect 13624 272 13690 273
rect 33592 272 33658 273
rect 53560 272 53626 273
rect 73528 272 73594 273
rect 44125 -516 44131 -452
rect 44195 -454 44201 -452
rect 88784 -454 88790 -452
rect 44195 -514 88790 -454
rect 44195 -516 44201 -514
rect 88784 -516 88790 -514
rect 88854 -516 88860 -452
rect 42957 -760 42963 -696
rect 43027 -698 43033 -696
rect 86288 -698 86294 -696
rect 43027 -758 86294 -698
rect 43027 -760 43033 -758
rect 86288 -760 86294 -758
rect 86358 -760 86364 -696
rect 40621 -1004 40627 -940
rect 40691 -942 40697 -940
rect 81296 -942 81302 -940
rect 40691 -1002 81302 -942
rect 40691 -1004 40697 -1002
rect 81296 -1004 81302 -1002
rect 81366 -1004 81372 -940
rect 38285 -1248 38291 -1184
rect 38355 -1186 38361 -1184
rect 76304 -1186 76310 -1184
rect 38355 -1246 76310 -1186
rect 38355 -1248 38361 -1246
rect 76304 -1248 76310 -1246
rect 76374 -1248 76380 -1184
rect 5581 -1492 5587 -1428
rect 5651 -1430 5657 -1428
rect 33587 -1430 33593 -1428
rect 5651 -1490 33593 -1430
rect 5651 -1492 5657 -1490
rect 33587 -1492 33593 -1490
rect 33657 -1492 33663 -1428
rect 35949 -1492 35955 -1428
rect 36019 -1430 36025 -1428
rect 71312 -1430 71318 -1428
rect 36019 -1490 71318 -1430
rect 36019 -1492 36025 -1490
rect 71312 -1492 71318 -1490
rect 71382 -1492 71388 -1428
rect 33613 -1736 33619 -1672
rect 33683 -1674 33689 -1672
rect 66320 -1674 66326 -1672
rect 33683 -1734 66326 -1674
rect 33683 -1736 33689 -1734
rect 66320 -1736 66326 -1734
rect 66390 -1736 66396 -1672
rect 17261 -1980 17267 -1916
rect 17331 -1918 17337 -1916
rect 31376 -1918 31382 -1916
rect 17331 -1978 31382 -1918
rect 17331 -1980 17337 -1978
rect 31376 -1980 31382 -1978
rect 31446 -1980 31452 -1916
rect 32445 -1980 32451 -1916
rect 32515 -1918 32521 -1916
rect 63824 -1918 63830 -1916
rect 32515 -1978 63830 -1918
rect 32515 -1980 32521 -1978
rect 63824 -1980 63830 -1978
rect 63894 -1980 63900 -1916
rect 31277 -2224 31283 -2160
rect 31347 -2162 31353 -2160
rect 61328 -2162 61334 -2160
rect 31347 -2222 61334 -2162
rect 31347 -2224 31353 -2222
rect 61328 -2224 61334 -2222
rect 61398 -2224 61404 -2160
rect 16093 -2468 16099 -2404
rect 16163 -2406 16169 -2404
rect 28880 -2406 28886 -2404
rect 16163 -2466 28886 -2406
rect 16163 -2468 16169 -2466
rect 28880 -2468 28886 -2466
rect 28950 -2468 28956 -2404
rect 30109 -2468 30115 -2404
rect 30179 -2406 30185 -2404
rect 58832 -2406 58838 -2404
rect 30179 -2466 58838 -2406
rect 30179 -2468 30185 -2466
rect 58832 -2468 58838 -2466
rect 58902 -2468 58908 -2404
rect 28941 -2712 28947 -2648
rect 29011 -2650 29017 -2648
rect 56336 -2650 56342 -2648
rect 29011 -2710 56342 -2650
rect 29011 -2712 29017 -2710
rect 56336 -2712 56342 -2710
rect 56406 -2712 56412 -2648
rect 14925 -2956 14931 -2892
rect 14995 -2894 15001 -2892
rect 26384 -2894 26390 -2892
rect 14995 -2954 26390 -2894
rect 14995 -2956 15001 -2954
rect 26384 -2956 26390 -2954
rect 26454 -2956 26460 -2892
rect 27773 -2956 27779 -2892
rect 27843 -2894 27849 -2892
rect 53840 -2894 53846 -2892
rect 27843 -2954 53846 -2894
rect 27843 -2956 27849 -2954
rect 53840 -2956 53846 -2954
rect 53910 -2956 53916 -2892
rect 26605 -3200 26611 -3136
rect 26675 -3138 26681 -3136
rect 51344 -3138 51350 -3136
rect 26675 -3198 51350 -3138
rect 26675 -3200 26681 -3198
rect 51344 -3200 51350 -3198
rect 51414 -3200 51420 -3136
rect 25437 -3444 25443 -3380
rect 25507 -3382 25513 -3380
rect 48848 -3382 48854 -3380
rect 25507 -3442 48854 -3382
rect 25507 -3444 25513 -3442
rect 48848 -3444 48854 -3442
rect 48918 -3444 48924 -3380
rect 9085 -3688 9091 -3624
rect 9155 -3626 9161 -3624
rect 13904 -3626 13910 -3624
rect 9155 -3686 13910 -3626
rect 9155 -3688 9161 -3686
rect 13904 -3688 13910 -3686
rect 13974 -3688 13980 -3624
rect 23101 -3688 23107 -3624
rect 23171 -3626 23177 -3624
rect 43856 -3626 43862 -3624
rect 23171 -3686 43862 -3626
rect 23171 -3688 23177 -3686
rect 43856 -3688 43862 -3686
rect 43926 -3688 43932 -3624
rect 45293 -3688 45299 -3624
rect 45363 -3626 45369 -3624
rect 91280 -3626 91286 -3624
rect 45363 -3686 91286 -3626
rect 45363 -3688 45369 -3686
rect 91280 -3688 91286 -3686
rect 91350 -3688 91356 -3624
rect 4413 -3932 4419 -3868
rect 4483 -3870 4489 -3868
rect 13619 -3870 13625 -3868
rect 4483 -3930 13625 -3870
rect 4483 -3932 4489 -3930
rect 13619 -3932 13625 -3930
rect 13689 -3932 13695 -3868
rect 20765 -3932 20771 -3868
rect 20835 -3870 20841 -3868
rect 38864 -3870 38870 -3868
rect 20835 -3930 38870 -3870
rect 20835 -3932 20841 -3930
rect 38864 -3932 38870 -3930
rect 38934 -3932 38940 -3868
rect 39453 -3932 39459 -3868
rect 39523 -3870 39529 -3868
rect 78800 -3870 78806 -3868
rect 39523 -3930 78806 -3870
rect 39523 -3932 39529 -3930
rect 78800 -3932 78806 -3930
rect 78870 -3932 78876 -3868
rect 13757 -4176 13763 -4112
rect 13827 -4114 13833 -4112
rect 23888 -4114 23894 -4112
rect 13827 -4174 23894 -4114
rect 13827 -4176 13833 -4174
rect 23888 -4176 23894 -4174
rect 23958 -4176 23964 -4112
rect 24269 -4176 24275 -4112
rect 24339 -4114 24345 -4112
rect 46352 -4114 46358 -4112
rect 24339 -4174 46358 -4114
rect 24339 -4176 24345 -4174
rect 46352 -4176 46358 -4174
rect 46422 -4176 46428 -4112
rect 12589 -4420 12595 -4356
rect 12659 -4358 12665 -4356
rect 21392 -4358 21398 -4356
rect 12659 -4418 21398 -4358
rect 12659 -4420 12665 -4418
rect 21392 -4420 21398 -4418
rect 21462 -4420 21468 -4356
rect 21933 -4420 21939 -4356
rect 22003 -4358 22009 -4356
rect 41360 -4358 41366 -4356
rect 22003 -4418 41366 -4358
rect 22003 -4420 22009 -4418
rect 41360 -4420 41366 -4418
rect 41430 -4420 41436 -4356
rect 41789 -4420 41795 -4356
rect 41859 -4358 41865 -4356
rect 83792 -4358 83798 -4356
rect 41859 -4418 83798 -4358
rect 41859 -4420 41865 -4418
rect 83792 -4420 83798 -4418
rect 83862 -4420 83868 -4356
rect 11421 -4664 11427 -4600
rect 11491 -4602 11497 -4600
rect 18896 -4602 18902 -4600
rect 11491 -4662 18902 -4602
rect 11491 -4664 11497 -4662
rect 18896 -4664 18902 -4662
rect 18966 -4664 18972 -4600
rect 19597 -4664 19603 -4600
rect 19667 -4602 19673 -4600
rect 36368 -4602 36374 -4600
rect 19667 -4662 36374 -4602
rect 19667 -4664 19673 -4662
rect 36368 -4664 36374 -4662
rect 36438 -4664 36444 -4600
rect 37117 -4664 37123 -4600
rect 37187 -4602 37193 -4600
rect 73808 -4602 73814 -4600
rect 37187 -4662 73814 -4602
rect 37187 -4664 37193 -4662
rect 73808 -4664 73814 -4662
rect 73878 -4664 73884 -4600
rect 10253 -4908 10259 -4844
rect 10323 -4846 10329 -4844
rect 16400 -4846 16406 -4844
rect 10323 -4906 16406 -4846
rect 10323 -4908 10329 -4906
rect 16400 -4908 16406 -4906
rect 16470 -4908 16476 -4844
rect 18429 -4908 18435 -4844
rect 18499 -4846 18505 -4844
rect 33872 -4846 33878 -4844
rect 18499 -4906 33878 -4846
rect 18499 -4908 18505 -4906
rect 33872 -4908 33878 -4906
rect 33942 -4908 33948 -4844
rect 34781 -4908 34787 -4844
rect 34851 -4846 34857 -4844
rect 68816 -4846 68822 -4844
rect 34851 -4906 68822 -4846
rect 34851 -4908 34857 -4906
rect 68816 -4908 68822 -4906
rect 68886 -4908 68892 -4844
rect 7917 -5152 7923 -5088
rect 7987 -5090 7993 -5088
rect 73523 -5090 73529 -5088
rect 7987 -5150 73529 -5090
rect 7987 -5152 7993 -5150
rect 73523 -5152 73529 -5150
rect 73593 -5152 73599 -5088
rect 6749 -5396 6755 -5332
rect 6819 -5334 6825 -5332
rect 53555 -5334 53561 -5332
rect 6819 -5394 53561 -5334
rect 6819 -5396 6825 -5394
rect 53555 -5396 53561 -5394
rect 53625 -5396 53631 -5332
rect 4418 -6333 4484 -6332
rect 5586 -6333 5652 -6332
rect 6754 -6333 6820 -6332
rect 7922 -6333 7988 -6332
rect 9090 -6333 9156 -6332
rect 10258 -6333 10324 -6332
rect 11426 -6333 11492 -6332
rect 12594 -6333 12660 -6332
rect 13762 -6333 13828 -6332
rect 14930 -6333 14996 -6332
rect 16098 -6333 16164 -6332
rect 17266 -6333 17332 -6332
rect 18434 -6333 18500 -6332
rect 19602 -6333 19668 -6332
rect 20770 -6333 20836 -6332
rect 21938 -6333 22004 -6332
rect 23106 -6333 23172 -6332
rect 24274 -6333 24340 -6332
rect 25442 -6333 25508 -6332
rect 26610 -6333 26676 -6332
rect 27778 -6333 27844 -6332
rect 28946 -6333 29012 -6332
rect 30114 -6333 30180 -6332
rect 31282 -6333 31348 -6332
rect 32450 -6333 32516 -6332
rect 33618 -6333 33684 -6332
rect 34786 -6333 34852 -6332
rect 35954 -6333 36020 -6332
rect 37122 -6333 37188 -6332
rect 38290 -6333 38356 -6332
rect 39458 -6333 39524 -6332
rect 40626 -6333 40692 -6332
rect 41794 -6333 41860 -6332
rect 42962 -6333 43028 -6332
rect 44130 -6333 44196 -6332
rect 45298 -6333 45364 -6332
rect 4376 -6397 4419 -6333
rect 4483 -6397 4526 -6333
rect 5544 -6397 5587 -6333
rect 5651 -6397 5694 -6333
rect 6712 -6397 6755 -6333
rect 6819 -6397 6862 -6333
rect 7880 -6397 7923 -6333
rect 7987 -6397 8030 -6333
rect 9048 -6397 9091 -6333
rect 9155 -6397 9198 -6333
rect 10216 -6397 10259 -6333
rect 10323 -6397 10366 -6333
rect 11384 -6397 11427 -6333
rect 11491 -6397 11534 -6333
rect 12552 -6397 12595 -6333
rect 12659 -6397 12702 -6333
rect 13720 -6397 13763 -6333
rect 13827 -6397 13870 -6333
rect 14888 -6397 14931 -6333
rect 14995 -6397 15038 -6333
rect 16056 -6397 16099 -6333
rect 16163 -6397 16206 -6333
rect 17224 -6397 17267 -6333
rect 17331 -6397 17374 -6333
rect 18392 -6397 18435 -6333
rect 18499 -6397 18542 -6333
rect 19560 -6397 19603 -6333
rect 19667 -6397 19710 -6333
rect 20728 -6397 20771 -6333
rect 20835 -6397 20878 -6333
rect 21896 -6397 21939 -6333
rect 22003 -6397 22046 -6333
rect 23064 -6397 23107 -6333
rect 23171 -6397 23214 -6333
rect 24232 -6397 24275 -6333
rect 24339 -6397 24382 -6333
rect 25400 -6397 25443 -6333
rect 25507 -6397 25550 -6333
rect 26568 -6397 26611 -6333
rect 26675 -6397 26718 -6333
rect 27736 -6397 27779 -6333
rect 27843 -6397 27886 -6333
rect 28904 -6397 28947 -6333
rect 29011 -6397 29054 -6333
rect 30072 -6397 30115 -6333
rect 30179 -6397 30222 -6333
rect 31240 -6397 31283 -6333
rect 31347 -6397 31390 -6333
rect 32408 -6397 32451 -6333
rect 32515 -6397 32558 -6333
rect 33576 -6397 33619 -6333
rect 33683 -6397 33726 -6333
rect 34744 -6397 34787 -6333
rect 34851 -6397 34894 -6333
rect 35912 -6397 35955 -6333
rect 36019 -6397 36062 -6333
rect 37080 -6397 37123 -6333
rect 37187 -6397 37230 -6333
rect 38248 -6397 38291 -6333
rect 38355 -6397 38398 -6333
rect 39416 -6397 39459 -6333
rect 39523 -6397 39566 -6333
rect 40584 -6397 40627 -6333
rect 40691 -6397 40734 -6333
rect 41752 -6397 41795 -6333
rect 41859 -6397 41902 -6333
rect 42920 -6397 42963 -6333
rect 43027 -6397 43070 -6333
rect 44088 -6397 44131 -6333
rect 44195 -6397 44238 -6333
rect 45256 -6397 45299 -6333
rect 45363 -6397 45406 -6333
rect 4418 -6398 4484 -6397
rect 5586 -6398 5652 -6397
rect 6754 -6398 6820 -6397
rect 7922 -6398 7988 -6397
rect 9090 -6398 9156 -6397
rect 10258 -6398 10324 -6397
rect 11426 -6398 11492 -6397
rect 12594 -6398 12660 -6397
rect 13762 -6398 13828 -6397
rect 14930 -6398 14996 -6397
rect 16098 -6398 16164 -6397
rect 17266 -6398 17332 -6397
rect 18434 -6398 18500 -6397
rect 19602 -6398 19668 -6397
rect 20770 -6398 20836 -6397
rect 21938 -6398 22004 -6397
rect 23106 -6398 23172 -6397
rect 24274 -6398 24340 -6397
rect 25442 -6398 25508 -6397
rect 26610 -6398 26676 -6397
rect 27778 -6398 27844 -6397
rect 28946 -6398 29012 -6397
rect 30114 -6398 30180 -6397
rect 31282 -6398 31348 -6397
rect 32450 -6398 32516 -6397
rect 33618 -6398 33684 -6397
rect 34786 -6398 34852 -6397
rect 35954 -6398 36020 -6397
rect 37122 -6398 37188 -6397
rect 38290 -6398 38356 -6397
rect 39458 -6398 39524 -6397
rect 40626 -6398 40692 -6397
rect 41794 -6398 41860 -6397
rect 42962 -6398 43028 -6397
rect 44130 -6398 44196 -6397
rect 45298 -6398 45364 -6397
<< via3 >>
rect 13910 1453 13974 1457
rect 13910 1397 13914 1453
rect 13914 1397 13970 1453
rect 13970 1397 13974 1453
rect 13910 1393 13974 1397
rect 16406 1453 16470 1457
rect 16406 1397 16410 1453
rect 16410 1397 16466 1453
rect 16466 1397 16470 1453
rect 16406 1393 16470 1397
rect 18902 1453 18966 1457
rect 18902 1397 18906 1453
rect 18906 1397 18962 1453
rect 18962 1397 18966 1453
rect 18902 1393 18966 1397
rect 21398 1453 21462 1457
rect 21398 1397 21402 1453
rect 21402 1397 21458 1453
rect 21458 1397 21462 1453
rect 21398 1393 21462 1397
rect 23894 1453 23958 1457
rect 23894 1397 23898 1453
rect 23898 1397 23954 1453
rect 23954 1397 23958 1453
rect 23894 1393 23958 1397
rect 26390 1453 26454 1457
rect 26390 1397 26394 1453
rect 26394 1397 26450 1453
rect 26450 1397 26454 1453
rect 26390 1393 26454 1397
rect 28886 1453 28950 1457
rect 28886 1397 28890 1453
rect 28890 1397 28946 1453
rect 28946 1397 28950 1453
rect 28886 1393 28950 1397
rect 31382 1453 31446 1457
rect 31382 1397 31386 1453
rect 31386 1397 31442 1453
rect 31442 1397 31446 1453
rect 31382 1393 31446 1397
rect 33878 1453 33942 1457
rect 33878 1397 33882 1453
rect 33882 1397 33938 1453
rect 33938 1397 33942 1453
rect 33878 1393 33942 1397
rect 36374 1453 36438 1457
rect 36374 1397 36378 1453
rect 36378 1397 36434 1453
rect 36434 1397 36438 1453
rect 36374 1393 36438 1397
rect 38870 1453 38934 1457
rect 38870 1397 38874 1453
rect 38874 1397 38930 1453
rect 38930 1397 38934 1453
rect 38870 1393 38934 1397
rect 41366 1453 41430 1457
rect 41366 1397 41370 1453
rect 41370 1397 41426 1453
rect 41426 1397 41430 1453
rect 41366 1393 41430 1397
rect 43862 1453 43926 1457
rect 43862 1397 43866 1453
rect 43866 1397 43922 1453
rect 43922 1397 43926 1453
rect 43862 1393 43926 1397
rect 46358 1453 46422 1457
rect 46358 1397 46362 1453
rect 46362 1397 46418 1453
rect 46418 1397 46422 1453
rect 46358 1393 46422 1397
rect 48854 1453 48918 1457
rect 48854 1397 48858 1453
rect 48858 1397 48914 1453
rect 48914 1397 48918 1453
rect 48854 1393 48918 1397
rect 51350 1453 51414 1457
rect 51350 1397 51354 1453
rect 51354 1397 51410 1453
rect 51410 1397 51414 1453
rect 51350 1393 51414 1397
rect 53846 1453 53910 1457
rect 53846 1397 53850 1453
rect 53850 1397 53906 1453
rect 53906 1397 53910 1453
rect 53846 1393 53910 1397
rect 56342 1453 56406 1457
rect 56342 1397 56346 1453
rect 56346 1397 56402 1453
rect 56402 1397 56406 1453
rect 56342 1393 56406 1397
rect 58838 1453 58902 1457
rect 58838 1397 58842 1453
rect 58842 1397 58898 1453
rect 58898 1397 58902 1453
rect 58838 1393 58902 1397
rect 61334 1453 61398 1457
rect 61334 1397 61338 1453
rect 61338 1397 61394 1453
rect 61394 1397 61398 1453
rect 61334 1393 61398 1397
rect 63830 1453 63894 1457
rect 63830 1397 63834 1453
rect 63834 1397 63890 1453
rect 63890 1397 63894 1453
rect 63830 1393 63894 1397
rect 66326 1453 66390 1457
rect 66326 1397 66330 1453
rect 66330 1397 66386 1453
rect 66386 1397 66390 1453
rect 66326 1393 66390 1397
rect 68822 1453 68886 1457
rect 68822 1397 68826 1453
rect 68826 1397 68882 1453
rect 68882 1397 68886 1453
rect 68822 1393 68886 1397
rect 71318 1453 71382 1457
rect 71318 1397 71322 1453
rect 71322 1397 71378 1453
rect 71378 1397 71382 1453
rect 71318 1393 71382 1397
rect 73814 1453 73878 1457
rect 73814 1397 73818 1453
rect 73818 1397 73874 1453
rect 73874 1397 73878 1453
rect 73814 1393 73878 1397
rect 76310 1453 76374 1457
rect 76310 1397 76314 1453
rect 76314 1397 76370 1453
rect 76370 1397 76374 1453
rect 76310 1393 76374 1397
rect 78806 1453 78870 1457
rect 78806 1397 78810 1453
rect 78810 1397 78866 1453
rect 78866 1397 78870 1453
rect 78806 1393 78870 1397
rect 81302 1453 81366 1457
rect 81302 1397 81306 1453
rect 81306 1397 81362 1453
rect 81362 1397 81366 1453
rect 81302 1393 81366 1397
rect 83798 1453 83862 1457
rect 83798 1397 83802 1453
rect 83802 1397 83858 1453
rect 83858 1397 83862 1453
rect 83798 1393 83862 1397
rect 86294 1453 86358 1457
rect 86294 1397 86298 1453
rect 86298 1397 86354 1453
rect 86354 1397 86358 1453
rect 86294 1393 86358 1397
rect 88790 1453 88854 1457
rect 88790 1397 88794 1453
rect 88794 1397 88850 1453
rect 88850 1397 88854 1453
rect 88790 1393 88854 1397
rect 91286 1453 91350 1457
rect 91286 1397 91290 1453
rect 91290 1397 91346 1453
rect 91346 1397 91350 1453
rect 91286 1393 91350 1397
rect 13625 333 13689 337
rect 13625 277 13629 333
rect 13629 277 13685 333
rect 13685 277 13689 333
rect 13625 273 13689 277
rect 33593 333 33657 337
rect 33593 277 33597 333
rect 33597 277 33653 333
rect 33653 277 33657 333
rect 33593 273 33657 277
rect 53561 333 53625 337
rect 53561 277 53565 333
rect 53565 277 53621 333
rect 53621 277 53625 333
rect 53561 273 53625 277
rect 73529 333 73593 337
rect 73529 277 73533 333
rect 73533 277 73589 333
rect 73589 277 73593 333
rect 73529 273 73593 277
rect 44131 -516 44195 -452
rect 88790 -516 88854 -452
rect 42963 -760 43027 -696
rect 86294 -760 86358 -696
rect 40627 -1004 40691 -940
rect 81302 -1004 81366 -940
rect 38291 -1248 38355 -1184
rect 76310 -1248 76374 -1184
rect 5587 -1492 5651 -1428
rect 33593 -1492 33657 -1428
rect 35955 -1492 36019 -1428
rect 71318 -1492 71382 -1428
rect 33619 -1736 33683 -1672
rect 66326 -1736 66390 -1672
rect 17267 -1980 17331 -1916
rect 31382 -1980 31446 -1916
rect 32451 -1980 32515 -1916
rect 63830 -1980 63894 -1916
rect 31283 -2224 31347 -2160
rect 61334 -2224 61398 -2160
rect 16099 -2468 16163 -2404
rect 28886 -2468 28950 -2404
rect 30115 -2468 30179 -2404
rect 58838 -2468 58902 -2404
rect 28947 -2712 29011 -2648
rect 56342 -2712 56406 -2648
rect 14931 -2956 14995 -2892
rect 26390 -2956 26454 -2892
rect 27779 -2956 27843 -2892
rect 53846 -2956 53910 -2892
rect 26611 -3200 26675 -3136
rect 51350 -3200 51414 -3136
rect 25443 -3444 25507 -3380
rect 48854 -3444 48918 -3380
rect 9091 -3688 9155 -3624
rect 13910 -3688 13974 -3624
rect 23107 -3688 23171 -3624
rect 43862 -3688 43926 -3624
rect 45299 -3688 45363 -3624
rect 91286 -3688 91350 -3624
rect 4419 -3932 4483 -3868
rect 13625 -3932 13689 -3868
rect 20771 -3932 20835 -3868
rect 38870 -3932 38934 -3868
rect 39459 -3932 39523 -3868
rect 78806 -3932 78870 -3868
rect 13763 -4176 13827 -4112
rect 23894 -4176 23958 -4112
rect 24275 -4176 24339 -4112
rect 46358 -4176 46422 -4112
rect 12595 -4420 12659 -4356
rect 21398 -4420 21462 -4356
rect 21939 -4420 22003 -4356
rect 41366 -4420 41430 -4356
rect 41795 -4420 41859 -4356
rect 83798 -4420 83862 -4356
rect 11427 -4664 11491 -4600
rect 18902 -4664 18966 -4600
rect 19603 -4664 19667 -4600
rect 36374 -4664 36438 -4600
rect 37123 -4664 37187 -4600
rect 73814 -4664 73878 -4600
rect 10259 -4908 10323 -4844
rect 16406 -4908 16470 -4844
rect 18435 -4908 18499 -4844
rect 33878 -4908 33942 -4844
rect 34787 -4908 34851 -4844
rect 68822 -4908 68886 -4844
rect 7923 -5152 7987 -5088
rect 73529 -5152 73593 -5088
rect 6755 -5396 6819 -5332
rect 53561 -5396 53625 -5332
rect 4419 -6337 4483 -6333
rect 4419 -6393 4423 -6337
rect 4423 -6393 4479 -6337
rect 4479 -6393 4483 -6337
rect 4419 -6397 4483 -6393
rect 5587 -6337 5651 -6333
rect 5587 -6393 5591 -6337
rect 5591 -6393 5647 -6337
rect 5647 -6393 5651 -6337
rect 5587 -6397 5651 -6393
rect 6755 -6337 6819 -6333
rect 6755 -6393 6759 -6337
rect 6759 -6393 6815 -6337
rect 6815 -6393 6819 -6337
rect 6755 -6397 6819 -6393
rect 7923 -6337 7987 -6333
rect 7923 -6393 7927 -6337
rect 7927 -6393 7983 -6337
rect 7983 -6393 7987 -6337
rect 7923 -6397 7987 -6393
rect 9091 -6337 9155 -6333
rect 9091 -6393 9095 -6337
rect 9095 -6393 9151 -6337
rect 9151 -6393 9155 -6337
rect 9091 -6397 9155 -6393
rect 10259 -6337 10323 -6333
rect 10259 -6393 10263 -6337
rect 10263 -6393 10319 -6337
rect 10319 -6393 10323 -6337
rect 10259 -6397 10323 -6393
rect 11427 -6337 11491 -6333
rect 11427 -6393 11431 -6337
rect 11431 -6393 11487 -6337
rect 11487 -6393 11491 -6337
rect 11427 -6397 11491 -6393
rect 12595 -6337 12659 -6333
rect 12595 -6393 12599 -6337
rect 12599 -6393 12655 -6337
rect 12655 -6393 12659 -6337
rect 12595 -6397 12659 -6393
rect 13763 -6337 13827 -6333
rect 13763 -6393 13767 -6337
rect 13767 -6393 13823 -6337
rect 13823 -6393 13827 -6337
rect 13763 -6397 13827 -6393
rect 14931 -6337 14995 -6333
rect 14931 -6393 14935 -6337
rect 14935 -6393 14991 -6337
rect 14991 -6393 14995 -6337
rect 14931 -6397 14995 -6393
rect 16099 -6337 16163 -6333
rect 16099 -6393 16103 -6337
rect 16103 -6393 16159 -6337
rect 16159 -6393 16163 -6337
rect 16099 -6397 16163 -6393
rect 17267 -6337 17331 -6333
rect 17267 -6393 17271 -6337
rect 17271 -6393 17327 -6337
rect 17327 -6393 17331 -6337
rect 17267 -6397 17331 -6393
rect 18435 -6337 18499 -6333
rect 18435 -6393 18439 -6337
rect 18439 -6393 18495 -6337
rect 18495 -6393 18499 -6337
rect 18435 -6397 18499 -6393
rect 19603 -6337 19667 -6333
rect 19603 -6393 19607 -6337
rect 19607 -6393 19663 -6337
rect 19663 -6393 19667 -6337
rect 19603 -6397 19667 -6393
rect 20771 -6337 20835 -6333
rect 20771 -6393 20775 -6337
rect 20775 -6393 20831 -6337
rect 20831 -6393 20835 -6337
rect 20771 -6397 20835 -6393
rect 21939 -6337 22003 -6333
rect 21939 -6393 21943 -6337
rect 21943 -6393 21999 -6337
rect 21999 -6393 22003 -6337
rect 21939 -6397 22003 -6393
rect 23107 -6337 23171 -6333
rect 23107 -6393 23111 -6337
rect 23111 -6393 23167 -6337
rect 23167 -6393 23171 -6337
rect 23107 -6397 23171 -6393
rect 24275 -6337 24339 -6333
rect 24275 -6393 24279 -6337
rect 24279 -6393 24335 -6337
rect 24335 -6393 24339 -6337
rect 24275 -6397 24339 -6393
rect 25443 -6337 25507 -6333
rect 25443 -6393 25447 -6337
rect 25447 -6393 25503 -6337
rect 25503 -6393 25507 -6337
rect 25443 -6397 25507 -6393
rect 26611 -6337 26675 -6333
rect 26611 -6393 26615 -6337
rect 26615 -6393 26671 -6337
rect 26671 -6393 26675 -6337
rect 26611 -6397 26675 -6393
rect 27779 -6337 27843 -6333
rect 27779 -6393 27783 -6337
rect 27783 -6393 27839 -6337
rect 27839 -6393 27843 -6337
rect 27779 -6397 27843 -6393
rect 28947 -6337 29011 -6333
rect 28947 -6393 28951 -6337
rect 28951 -6393 29007 -6337
rect 29007 -6393 29011 -6337
rect 28947 -6397 29011 -6393
rect 30115 -6337 30179 -6333
rect 30115 -6393 30119 -6337
rect 30119 -6393 30175 -6337
rect 30175 -6393 30179 -6337
rect 30115 -6397 30179 -6393
rect 31283 -6337 31347 -6333
rect 31283 -6393 31287 -6337
rect 31287 -6393 31343 -6337
rect 31343 -6393 31347 -6337
rect 31283 -6397 31347 -6393
rect 32451 -6337 32515 -6333
rect 32451 -6393 32455 -6337
rect 32455 -6393 32511 -6337
rect 32511 -6393 32515 -6337
rect 32451 -6397 32515 -6393
rect 33619 -6337 33683 -6333
rect 33619 -6393 33623 -6337
rect 33623 -6393 33679 -6337
rect 33679 -6393 33683 -6337
rect 33619 -6397 33683 -6393
rect 34787 -6337 34851 -6333
rect 34787 -6393 34791 -6337
rect 34791 -6393 34847 -6337
rect 34847 -6393 34851 -6337
rect 34787 -6397 34851 -6393
rect 35955 -6337 36019 -6333
rect 35955 -6393 35959 -6337
rect 35959 -6393 36015 -6337
rect 36015 -6393 36019 -6337
rect 35955 -6397 36019 -6393
rect 37123 -6337 37187 -6333
rect 37123 -6393 37127 -6337
rect 37127 -6393 37183 -6337
rect 37183 -6393 37187 -6337
rect 37123 -6397 37187 -6393
rect 38291 -6337 38355 -6333
rect 38291 -6393 38295 -6337
rect 38295 -6393 38351 -6337
rect 38351 -6393 38355 -6337
rect 38291 -6397 38355 -6393
rect 39459 -6337 39523 -6333
rect 39459 -6393 39463 -6337
rect 39463 -6393 39519 -6337
rect 39519 -6393 39523 -6337
rect 39459 -6397 39523 -6393
rect 40627 -6337 40691 -6333
rect 40627 -6393 40631 -6337
rect 40631 -6393 40687 -6337
rect 40687 -6393 40691 -6337
rect 40627 -6397 40691 -6393
rect 41795 -6337 41859 -6333
rect 41795 -6393 41799 -6337
rect 41799 -6393 41855 -6337
rect 41855 -6393 41859 -6337
rect 41795 -6397 41859 -6393
rect 42963 -6337 43027 -6333
rect 42963 -6393 42967 -6337
rect 42967 -6393 43023 -6337
rect 43023 -6393 43027 -6337
rect 42963 -6397 43027 -6393
rect 44131 -6337 44195 -6333
rect 44131 -6393 44135 -6337
rect 44135 -6393 44191 -6337
rect 44191 -6393 44195 -6337
rect 44131 -6397 44195 -6393
rect 45299 -6337 45363 -6333
rect 45299 -6393 45303 -6337
rect 45303 -6393 45359 -6337
rect 45359 -6393 45363 -6337
rect 45299 -6397 45363 -6393
<< metal4 >>
rect 13909 1457 13975 1458
rect 13909 1393 13910 1457
rect 13974 1393 13975 1457
rect 13909 1392 13975 1393
rect 16405 1457 16471 1458
rect 16405 1393 16406 1457
rect 16470 1393 16471 1457
rect 16405 1392 16471 1393
rect 18901 1457 18967 1458
rect 18901 1393 18902 1457
rect 18966 1393 18967 1457
rect 18901 1392 18967 1393
rect 21397 1457 21463 1458
rect 21397 1393 21398 1457
rect 21462 1393 21463 1457
rect 21397 1392 21463 1393
rect 23893 1457 23959 1458
rect 23893 1393 23894 1457
rect 23958 1393 23959 1457
rect 23893 1392 23959 1393
rect 26389 1457 26455 1458
rect 26389 1393 26390 1457
rect 26454 1393 26455 1457
rect 26389 1392 26455 1393
rect 28885 1457 28951 1458
rect 28885 1393 28886 1457
rect 28950 1393 28951 1457
rect 28885 1392 28951 1393
rect 31381 1457 31447 1458
rect 31381 1393 31382 1457
rect 31446 1393 31447 1457
rect 31381 1392 31447 1393
rect 33877 1457 33943 1458
rect 33877 1393 33878 1457
rect 33942 1393 33943 1457
rect 33877 1392 33943 1393
rect 36373 1457 36439 1458
rect 36373 1393 36374 1457
rect 36438 1393 36439 1457
rect 36373 1392 36439 1393
rect 38869 1457 38935 1458
rect 38869 1393 38870 1457
rect 38934 1393 38935 1457
rect 38869 1392 38935 1393
rect 41365 1457 41431 1458
rect 41365 1393 41366 1457
rect 41430 1393 41431 1457
rect 41365 1392 41431 1393
rect 43861 1457 43927 1458
rect 43861 1393 43862 1457
rect 43926 1393 43927 1457
rect 43861 1392 43927 1393
rect 46357 1457 46423 1458
rect 46357 1393 46358 1457
rect 46422 1393 46423 1457
rect 46357 1392 46423 1393
rect 48853 1457 48919 1458
rect 48853 1393 48854 1457
rect 48918 1393 48919 1457
rect 48853 1392 48919 1393
rect 51349 1457 51415 1458
rect 51349 1393 51350 1457
rect 51414 1393 51415 1457
rect 51349 1392 51415 1393
rect 53845 1457 53911 1458
rect 53845 1393 53846 1457
rect 53910 1393 53911 1457
rect 53845 1392 53911 1393
rect 56341 1457 56407 1458
rect 56341 1393 56342 1457
rect 56406 1393 56407 1457
rect 56341 1392 56407 1393
rect 58837 1457 58903 1458
rect 58837 1393 58838 1457
rect 58902 1393 58903 1457
rect 58837 1392 58903 1393
rect 61333 1457 61399 1458
rect 61333 1393 61334 1457
rect 61398 1393 61399 1457
rect 61333 1392 61399 1393
rect 63829 1457 63895 1458
rect 63829 1393 63830 1457
rect 63894 1393 63895 1457
rect 63829 1392 63895 1393
rect 66325 1457 66391 1458
rect 66325 1393 66326 1457
rect 66390 1393 66391 1457
rect 66325 1392 66391 1393
rect 68821 1457 68887 1458
rect 68821 1393 68822 1457
rect 68886 1393 68887 1457
rect 68821 1392 68887 1393
rect 71317 1457 71383 1458
rect 71317 1393 71318 1457
rect 71382 1393 71383 1457
rect 71317 1392 71383 1393
rect 73813 1457 73879 1458
rect 73813 1393 73814 1457
rect 73878 1393 73879 1457
rect 73813 1392 73879 1393
rect 76309 1457 76375 1458
rect 76309 1393 76310 1457
rect 76374 1393 76375 1457
rect 76309 1392 76375 1393
rect 78805 1457 78871 1458
rect 78805 1393 78806 1457
rect 78870 1393 78871 1457
rect 78805 1392 78871 1393
rect 81301 1457 81367 1458
rect 81301 1393 81302 1457
rect 81366 1393 81367 1457
rect 81301 1392 81367 1393
rect 83797 1457 83863 1458
rect 83797 1393 83798 1457
rect 83862 1393 83863 1457
rect 83797 1392 83863 1393
rect 86293 1457 86359 1458
rect 86293 1393 86294 1457
rect 86358 1393 86359 1457
rect 86293 1392 86359 1393
rect 88789 1457 88855 1458
rect 88789 1393 88790 1457
rect 88854 1393 88855 1457
rect 88789 1392 88855 1393
rect 91285 1457 91351 1458
rect 91285 1393 91286 1457
rect 91350 1393 91351 1457
rect 91285 1392 91351 1393
rect 13624 337 13690 338
rect 13624 273 13625 337
rect 13689 273 13690 337
rect 13624 272 13690 273
rect 5586 -1428 5652 -1427
rect 5586 -1492 5587 -1428
rect 5651 -1492 5652 -1428
rect 5586 -1493 5652 -1492
rect 4418 -3868 4484 -3867
rect 4418 -3932 4419 -3868
rect 4483 -3932 4484 -3868
rect 4418 -3933 4484 -3932
rect 4421 -6332 4481 -3933
rect 5589 -6332 5649 -1493
rect 9090 -3624 9156 -3623
rect 9090 -3688 9091 -3624
rect 9155 -3688 9156 -3624
rect 9090 -3689 9156 -3688
rect 7922 -5088 7988 -5087
rect 7922 -5152 7923 -5088
rect 7987 -5152 7988 -5088
rect 7922 -5153 7988 -5152
rect 6754 -5332 6820 -5331
rect 6754 -5396 6755 -5332
rect 6819 -5396 6820 -5332
rect 6754 -5397 6820 -5396
rect 6757 -6332 6817 -5397
rect 7925 -6332 7985 -5153
rect 9093 -6332 9153 -3689
rect 13627 -3867 13687 272
rect 13912 -3623 13972 1392
rect 16098 -2404 16164 -2403
rect 16098 -2468 16099 -2404
rect 16163 -2468 16164 -2404
rect 16098 -2469 16164 -2468
rect 14930 -2892 14996 -2891
rect 14930 -2956 14931 -2892
rect 14995 -2956 14996 -2892
rect 14930 -2957 14996 -2956
rect 13909 -3624 13975 -3623
rect 13909 -3688 13910 -3624
rect 13974 -3688 13975 -3624
rect 13909 -3689 13975 -3688
rect 13624 -3868 13690 -3867
rect 13624 -3932 13625 -3868
rect 13689 -3932 13690 -3868
rect 13624 -3933 13690 -3932
rect 13762 -4112 13828 -4111
rect 13762 -4176 13763 -4112
rect 13827 -4176 13828 -4112
rect 13762 -4177 13828 -4176
rect 12594 -4356 12660 -4355
rect 12594 -4420 12595 -4356
rect 12659 -4420 12660 -4356
rect 12594 -4421 12660 -4420
rect 11426 -4600 11492 -4599
rect 11426 -4664 11427 -4600
rect 11491 -4664 11492 -4600
rect 11426 -4665 11492 -4664
rect 10258 -4844 10324 -4843
rect 10258 -4908 10259 -4844
rect 10323 -4908 10324 -4844
rect 10258 -4909 10324 -4908
rect 10261 -6332 10321 -4909
rect 11429 -6332 11489 -4665
rect 12597 -6332 12657 -4421
rect 13765 -6332 13825 -4177
rect 14933 -6332 14993 -2957
rect 16101 -6332 16161 -2469
rect 16408 -4843 16468 1392
rect 17266 -1916 17332 -1915
rect 17266 -1980 17267 -1916
rect 17331 -1980 17332 -1916
rect 17266 -1981 17332 -1980
rect 16405 -4844 16471 -4843
rect 16405 -4908 16406 -4844
rect 16470 -4908 16471 -4844
rect 16405 -4909 16471 -4908
rect 17269 -6332 17329 -1981
rect 18904 -4599 18964 1392
rect 20770 -3868 20836 -3867
rect 20770 -3932 20771 -3868
rect 20835 -3932 20836 -3868
rect 20770 -3933 20836 -3932
rect 18901 -4600 18967 -4599
rect 18901 -4664 18902 -4600
rect 18966 -4664 18967 -4600
rect 18901 -4665 18967 -4664
rect 19602 -4600 19668 -4599
rect 19602 -4664 19603 -4600
rect 19667 -4664 19668 -4600
rect 19602 -4665 19668 -4664
rect 18434 -4844 18500 -4843
rect 18434 -4908 18435 -4844
rect 18499 -4908 18500 -4844
rect 18434 -4909 18500 -4908
rect 18437 -6332 18497 -4909
rect 19605 -6332 19665 -4665
rect 20773 -6332 20833 -3933
rect 21400 -4355 21460 1392
rect 23106 -3624 23172 -3623
rect 23106 -3688 23107 -3624
rect 23171 -3688 23172 -3624
rect 23106 -3689 23172 -3688
rect 21397 -4356 21463 -4355
rect 21397 -4420 21398 -4356
rect 21462 -4420 21463 -4356
rect 21397 -4421 21463 -4420
rect 21938 -4356 22004 -4355
rect 21938 -4420 21939 -4356
rect 22003 -4420 22004 -4356
rect 21938 -4421 22004 -4420
rect 21941 -6332 22001 -4421
rect 23109 -6332 23169 -3689
rect 23896 -4111 23956 1392
rect 26392 -2891 26452 1392
rect 28888 -2403 28948 1392
rect 31384 -1915 31444 1392
rect 33592 337 33658 338
rect 33592 273 33593 337
rect 33657 273 33658 337
rect 33592 272 33658 273
rect 33595 -1427 33655 272
rect 33592 -1428 33658 -1427
rect 33592 -1492 33593 -1428
rect 33657 -1492 33658 -1428
rect 33592 -1493 33658 -1492
rect 33618 -1672 33684 -1671
rect 33618 -1736 33619 -1672
rect 33683 -1736 33684 -1672
rect 33618 -1737 33684 -1736
rect 31381 -1916 31447 -1915
rect 31381 -1980 31382 -1916
rect 31446 -1980 31447 -1916
rect 31381 -1981 31447 -1980
rect 32450 -1916 32516 -1915
rect 32450 -1980 32451 -1916
rect 32515 -1980 32516 -1916
rect 32450 -1981 32516 -1980
rect 31282 -2160 31348 -2159
rect 31282 -2224 31283 -2160
rect 31347 -2224 31348 -2160
rect 31282 -2225 31348 -2224
rect 28885 -2404 28951 -2403
rect 28885 -2468 28886 -2404
rect 28950 -2468 28951 -2404
rect 28885 -2469 28951 -2468
rect 30114 -2404 30180 -2403
rect 30114 -2468 30115 -2404
rect 30179 -2468 30180 -2404
rect 30114 -2469 30180 -2468
rect 28946 -2648 29012 -2647
rect 28946 -2712 28947 -2648
rect 29011 -2712 29012 -2648
rect 28946 -2713 29012 -2712
rect 26389 -2892 26455 -2891
rect 26389 -2956 26390 -2892
rect 26454 -2956 26455 -2892
rect 26389 -2957 26455 -2956
rect 27778 -2892 27844 -2891
rect 27778 -2956 27779 -2892
rect 27843 -2956 27844 -2892
rect 27778 -2957 27844 -2956
rect 26610 -3136 26676 -3135
rect 26610 -3200 26611 -3136
rect 26675 -3200 26676 -3136
rect 26610 -3201 26676 -3200
rect 25442 -3380 25508 -3379
rect 25442 -3444 25443 -3380
rect 25507 -3444 25508 -3380
rect 25442 -3445 25508 -3444
rect 23893 -4112 23959 -4111
rect 23893 -4176 23894 -4112
rect 23958 -4176 23959 -4112
rect 23893 -4177 23959 -4176
rect 24274 -4112 24340 -4111
rect 24274 -4176 24275 -4112
rect 24339 -4176 24340 -4112
rect 24274 -4177 24340 -4176
rect 24277 -6332 24337 -4177
rect 25445 -6332 25505 -3445
rect 26613 -6332 26673 -3201
rect 27781 -6332 27841 -2957
rect 28949 -6332 29009 -2713
rect 30117 -6332 30177 -2469
rect 31285 -6332 31345 -2225
rect 32453 -6332 32513 -1981
rect 33621 -6332 33681 -1737
rect 33880 -4843 33940 1392
rect 35954 -1428 36020 -1427
rect 35954 -1492 35955 -1428
rect 36019 -1492 36020 -1428
rect 35954 -1493 36020 -1492
rect 33877 -4844 33943 -4843
rect 33877 -4908 33878 -4844
rect 33942 -4908 33943 -4844
rect 33877 -4909 33943 -4908
rect 34786 -4844 34852 -4843
rect 34786 -4908 34787 -4844
rect 34851 -4908 34852 -4844
rect 34786 -4909 34852 -4908
rect 34789 -6332 34849 -4909
rect 35957 -6332 36017 -1493
rect 36376 -4599 36436 1392
rect 38290 -1184 38356 -1183
rect 38290 -1248 38291 -1184
rect 38355 -1248 38356 -1184
rect 38290 -1249 38356 -1248
rect 36373 -4600 36439 -4599
rect 36373 -4664 36374 -4600
rect 36438 -4664 36439 -4600
rect 36373 -4665 36439 -4664
rect 37122 -4600 37188 -4599
rect 37122 -4664 37123 -4600
rect 37187 -4664 37188 -4600
rect 37122 -4665 37188 -4664
rect 37125 -6332 37185 -4665
rect 38293 -6332 38353 -1249
rect 38872 -3867 38932 1392
rect 40626 -940 40692 -939
rect 40626 -1004 40627 -940
rect 40691 -1004 40692 -940
rect 40626 -1005 40692 -1004
rect 38869 -3868 38935 -3867
rect 38869 -3932 38870 -3868
rect 38934 -3932 38935 -3868
rect 38869 -3933 38935 -3932
rect 39458 -3868 39524 -3867
rect 39458 -3932 39459 -3868
rect 39523 -3932 39524 -3868
rect 39458 -3933 39524 -3932
rect 39461 -6332 39521 -3933
rect 40629 -6332 40689 -1005
rect 41368 -4355 41428 1392
rect 42962 -696 43028 -695
rect 42962 -760 42963 -696
rect 43027 -760 43028 -696
rect 42962 -761 43028 -760
rect 41365 -4356 41431 -4355
rect 41365 -4420 41366 -4356
rect 41430 -4420 41431 -4356
rect 41365 -4421 41431 -4420
rect 41794 -4356 41860 -4355
rect 41794 -4420 41795 -4356
rect 41859 -4420 41860 -4356
rect 41794 -4421 41860 -4420
rect 41797 -6332 41857 -4421
rect 42965 -6332 43025 -761
rect 43864 -3623 43924 1392
rect 44130 -452 44196 -451
rect 44130 -516 44131 -452
rect 44195 -516 44196 -452
rect 44130 -517 44196 -516
rect 43861 -3624 43927 -3623
rect 43861 -3688 43862 -3624
rect 43926 -3688 43927 -3624
rect 43861 -3689 43927 -3688
rect 44133 -6332 44193 -517
rect 45298 -3624 45364 -3623
rect 45298 -3688 45299 -3624
rect 45363 -3688 45364 -3624
rect 45298 -3689 45364 -3688
rect 45301 -6332 45361 -3689
rect 46360 -4111 46420 1392
rect 48856 -3379 48916 1392
rect 51352 -3135 51412 1392
rect 53560 337 53626 338
rect 53560 273 53561 337
rect 53625 273 53626 337
rect 53560 272 53626 273
rect 51349 -3136 51415 -3135
rect 51349 -3200 51350 -3136
rect 51414 -3200 51415 -3136
rect 51349 -3201 51415 -3200
rect 48853 -3380 48919 -3379
rect 48853 -3444 48854 -3380
rect 48918 -3444 48919 -3380
rect 48853 -3445 48919 -3444
rect 46357 -4112 46423 -4111
rect 46357 -4176 46358 -4112
rect 46422 -4176 46423 -4112
rect 46357 -4177 46423 -4176
rect 53563 -5331 53623 272
rect 53848 -2891 53908 1392
rect 56344 -2647 56404 1392
rect 58840 -2403 58900 1392
rect 61336 -2159 61396 1392
rect 63832 -1915 63892 1392
rect 66328 -1671 66388 1392
rect 66325 -1672 66391 -1671
rect 66325 -1736 66326 -1672
rect 66390 -1736 66391 -1672
rect 66325 -1737 66391 -1736
rect 63829 -1916 63895 -1915
rect 63829 -1980 63830 -1916
rect 63894 -1980 63895 -1916
rect 63829 -1981 63895 -1980
rect 61333 -2160 61399 -2159
rect 61333 -2224 61334 -2160
rect 61398 -2224 61399 -2160
rect 61333 -2225 61399 -2224
rect 58837 -2404 58903 -2403
rect 58837 -2468 58838 -2404
rect 58902 -2468 58903 -2404
rect 58837 -2469 58903 -2468
rect 56341 -2648 56407 -2647
rect 56341 -2712 56342 -2648
rect 56406 -2712 56407 -2648
rect 56341 -2713 56407 -2712
rect 53845 -2892 53911 -2891
rect 53845 -2956 53846 -2892
rect 53910 -2956 53911 -2892
rect 53845 -2957 53911 -2956
rect 68824 -4843 68884 1392
rect 71320 -1427 71380 1392
rect 73528 337 73594 338
rect 73528 273 73529 337
rect 73593 273 73594 337
rect 73528 272 73594 273
rect 71317 -1428 71383 -1427
rect 71317 -1492 71318 -1428
rect 71382 -1492 71383 -1428
rect 71317 -1493 71383 -1492
rect 68821 -4844 68887 -4843
rect 68821 -4908 68822 -4844
rect 68886 -4908 68887 -4844
rect 68821 -4909 68887 -4908
rect 73531 -5087 73591 272
rect 73816 -4599 73876 1392
rect 76312 -1183 76372 1392
rect 76309 -1184 76375 -1183
rect 76309 -1248 76310 -1184
rect 76374 -1248 76375 -1184
rect 76309 -1249 76375 -1248
rect 78808 -3867 78868 1392
rect 81304 -939 81364 1392
rect 81301 -940 81367 -939
rect 81301 -1004 81302 -940
rect 81366 -1004 81367 -940
rect 81301 -1005 81367 -1004
rect 78805 -3868 78871 -3867
rect 78805 -3932 78806 -3868
rect 78870 -3932 78871 -3868
rect 78805 -3933 78871 -3932
rect 83800 -4355 83860 1392
rect 86296 -695 86356 1392
rect 88792 -451 88852 1392
rect 88789 -452 88855 -451
rect 88789 -516 88790 -452
rect 88854 -516 88855 -452
rect 88789 -517 88855 -516
rect 86293 -696 86359 -695
rect 86293 -760 86294 -696
rect 86358 -760 86359 -696
rect 86293 -761 86359 -760
rect 91288 -3623 91348 1392
rect 91285 -3624 91351 -3623
rect 91285 -3688 91286 -3624
rect 91350 -3688 91351 -3624
rect 91285 -3689 91351 -3688
rect 83797 -4356 83863 -4355
rect 83797 -4420 83798 -4356
rect 83862 -4420 83863 -4356
rect 83797 -4421 83863 -4420
rect 73813 -4600 73879 -4599
rect 73813 -4664 73814 -4600
rect 73878 -4664 73879 -4600
rect 73813 -4665 73879 -4664
rect 73528 -5088 73594 -5087
rect 73528 -5152 73529 -5088
rect 73593 -5152 73594 -5088
rect 73528 -5153 73594 -5152
rect 53560 -5332 53626 -5331
rect 53560 -5396 53561 -5332
rect 53625 -5396 53626 -5332
rect 53560 -5397 53626 -5396
rect 4418 -6333 4484 -6332
rect 4418 -6397 4419 -6333
rect 4483 -6397 4484 -6333
rect 4418 -6398 4484 -6397
rect 5586 -6333 5652 -6332
rect 5586 -6397 5587 -6333
rect 5651 -6397 5652 -6333
rect 5586 -6398 5652 -6397
rect 6754 -6333 6820 -6332
rect 6754 -6397 6755 -6333
rect 6819 -6397 6820 -6333
rect 6754 -6398 6820 -6397
rect 7922 -6333 7988 -6332
rect 7922 -6397 7923 -6333
rect 7987 -6397 7988 -6333
rect 7922 -6398 7988 -6397
rect 9090 -6333 9156 -6332
rect 9090 -6397 9091 -6333
rect 9155 -6397 9156 -6333
rect 9090 -6398 9156 -6397
rect 10258 -6333 10324 -6332
rect 10258 -6397 10259 -6333
rect 10323 -6397 10324 -6333
rect 10258 -6398 10324 -6397
rect 11426 -6333 11492 -6332
rect 11426 -6397 11427 -6333
rect 11491 -6397 11492 -6333
rect 11426 -6398 11492 -6397
rect 12594 -6333 12660 -6332
rect 12594 -6397 12595 -6333
rect 12659 -6397 12660 -6333
rect 12594 -6398 12660 -6397
rect 13762 -6333 13828 -6332
rect 13762 -6397 13763 -6333
rect 13827 -6397 13828 -6333
rect 13762 -6398 13828 -6397
rect 14930 -6333 14996 -6332
rect 14930 -6397 14931 -6333
rect 14995 -6397 14996 -6333
rect 14930 -6398 14996 -6397
rect 16098 -6333 16164 -6332
rect 16098 -6397 16099 -6333
rect 16163 -6397 16164 -6333
rect 16098 -6398 16164 -6397
rect 17266 -6333 17332 -6332
rect 17266 -6397 17267 -6333
rect 17331 -6397 17332 -6333
rect 17266 -6398 17332 -6397
rect 18434 -6333 18500 -6332
rect 18434 -6397 18435 -6333
rect 18499 -6397 18500 -6333
rect 18434 -6398 18500 -6397
rect 19602 -6333 19668 -6332
rect 19602 -6397 19603 -6333
rect 19667 -6397 19668 -6333
rect 19602 -6398 19668 -6397
rect 20770 -6333 20836 -6332
rect 20770 -6397 20771 -6333
rect 20835 -6397 20836 -6333
rect 20770 -6398 20836 -6397
rect 21938 -6333 22004 -6332
rect 21938 -6397 21939 -6333
rect 22003 -6397 22004 -6333
rect 21938 -6398 22004 -6397
rect 23106 -6333 23172 -6332
rect 23106 -6397 23107 -6333
rect 23171 -6397 23172 -6333
rect 23106 -6398 23172 -6397
rect 24274 -6333 24340 -6332
rect 24274 -6397 24275 -6333
rect 24339 -6397 24340 -6333
rect 24274 -6398 24340 -6397
rect 25442 -6333 25508 -6332
rect 25442 -6397 25443 -6333
rect 25507 -6397 25508 -6333
rect 25442 -6398 25508 -6397
rect 26610 -6333 26676 -6332
rect 26610 -6397 26611 -6333
rect 26675 -6397 26676 -6333
rect 26610 -6398 26676 -6397
rect 27778 -6333 27844 -6332
rect 27778 -6397 27779 -6333
rect 27843 -6397 27844 -6333
rect 27778 -6398 27844 -6397
rect 28946 -6333 29012 -6332
rect 28946 -6397 28947 -6333
rect 29011 -6397 29012 -6333
rect 28946 -6398 29012 -6397
rect 30114 -6333 30180 -6332
rect 30114 -6397 30115 -6333
rect 30179 -6397 30180 -6333
rect 30114 -6398 30180 -6397
rect 31282 -6333 31348 -6332
rect 31282 -6397 31283 -6333
rect 31347 -6397 31348 -6333
rect 31282 -6398 31348 -6397
rect 32450 -6333 32516 -6332
rect 32450 -6397 32451 -6333
rect 32515 -6397 32516 -6333
rect 32450 -6398 32516 -6397
rect 33618 -6333 33684 -6332
rect 33618 -6397 33619 -6333
rect 33683 -6397 33684 -6333
rect 33618 -6398 33684 -6397
rect 34786 -6333 34852 -6332
rect 34786 -6397 34787 -6333
rect 34851 -6397 34852 -6333
rect 34786 -6398 34852 -6397
rect 35954 -6333 36020 -6332
rect 35954 -6397 35955 -6333
rect 36019 -6397 36020 -6333
rect 35954 -6398 36020 -6397
rect 37122 -6333 37188 -6332
rect 37122 -6397 37123 -6333
rect 37187 -6397 37188 -6333
rect 37122 -6398 37188 -6397
rect 38290 -6333 38356 -6332
rect 38290 -6397 38291 -6333
rect 38355 -6397 38356 -6333
rect 38290 -6398 38356 -6397
rect 39458 -6333 39524 -6332
rect 39458 -6397 39459 -6333
rect 39523 -6397 39524 -6333
rect 39458 -6398 39524 -6397
rect 40626 -6333 40692 -6332
rect 40626 -6397 40627 -6333
rect 40691 -6397 40692 -6333
rect 40626 -6398 40692 -6397
rect 41794 -6333 41860 -6332
rect 41794 -6397 41795 -6333
rect 41859 -6397 41860 -6333
rect 41794 -6398 41860 -6397
rect 42962 -6333 43028 -6332
rect 42962 -6397 42963 -6333
rect 43027 -6397 43028 -6333
rect 42962 -6398 43028 -6397
rect 44130 -6333 44196 -6332
rect 44130 -6397 44131 -6333
rect 44195 -6397 44196 -6333
rect 44130 -6398 44196 -6397
rect 45298 -6333 45364 -6332
rect 45298 -6397 45299 -6333
rect 45363 -6397 45364 -6333
rect 45298 -6398 45364 -6397
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1649977179
transform 1 0 23893 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1649977179
transform 1 0 4418 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1649977179
transform 1 0 9090 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1649977179
transform 1 0 10258 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1649977179
transform 1 0 11426 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1649977179
transform 1 0 13909 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1649977179
transform 1 0 16405 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1649977179
transform 1 0 21938 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1649977179
transform 1 0 18901 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1649977179
transform 1 0 14930 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1649977179
transform 1 0 12594 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1649977179
transform 1 0 5586 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1649977179
transform 1 0 13624 0 1 268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1649977179
transform 1 0 24274 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1649977179
transform 1 0 21397 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1649977179
transform 1 0 20770 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1649977179
transform 1 0 25442 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1649977179
transform 1 0 17266 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1649977179
transform 1 0 6754 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1649977179
transform 1 0 13762 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1649977179
transform 1 0 7922 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1649977179
transform 1 0 18434 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1649977179
transform 1 0 19602 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1649977179
transform 1 0 16098 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1649977179
transform 1 0 23106 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1649977179
transform 1 0 44130 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1649977179
transform 1 0 42962 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1649977179
transform 1 0 41794 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1649977179
transform 1 0 40626 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1649977179
transform 1 0 38290 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1649977179
transform 1 0 41365 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1649977179
transform 1 0 35954 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1649977179
transform 1 0 33592 0 1 268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1649977179
transform 1 0 33618 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1649977179
transform 1 0 32450 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1649977179
transform 1 0 37122 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1649977179
transform 1 0 31381 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1649977179
transform 1 0 31282 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1649977179
transform 1 0 30114 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1649977179
transform 1 0 36373 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1649977179
transform 1 0 28885 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1649977179
transform 1 0 28946 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1649977179
transform 1 0 27778 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1649977179
transform 1 0 26389 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1649977179
transform 1 0 26610 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1649977179
transform 1 0 34786 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1649977179
transform 1 0 45298 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1649977179
transform 1 0 43861 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1649977179
transform 1 0 39458 0 1 -6402
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1649977179
transform 1 0 33877 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1649977179
transform 1 0 38869 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1649977179
transform 1 0 46357 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1649977179
transform 1 0 88789 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1649977179
transform 1 0 86293 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1649977179
transform 1 0 81301 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1649977179
transform 1 0 76309 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1649977179
transform 1 0 71317 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1649977179
transform 1 0 66325 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1649977179
transform 1 0 63829 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1649977179
transform 1 0 61333 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1649977179
transform 1 0 58837 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1649977179
transform 1 0 56341 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1649977179
transform 1 0 53845 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1649977179
transform 1 0 51349 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1649977179
transform 1 0 48853 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1649977179
transform 1 0 91285 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1649977179
transform 1 0 78805 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1649977179
transform 1 0 83797 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1649977179
transform 1 0 73813 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1649977179
transform 1 0 68821 0 1 1388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1649977179
transform 1 0 73528 0 1 268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1649977179
transform 1 0 53560 0 1 268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1649977179
transform 1 0 23894 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1649977179
transform 1 0 13910 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1649977179
transform 1 0 18902 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1649977179
transform 1 0 21398 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1649977179
transform 1 0 16406 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1649977179
transform 1 0 41366 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1649977179
transform 1 0 31382 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1649977179
transform 1 0 28886 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1649977179
transform 1 0 36374 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1649977179
transform 1 0 26390 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1649977179
transform 1 0 43862 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1649977179
transform 1 0 33878 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1649977179
transform 1 0 38870 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1649977179
transform 1 0 46358 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1649977179
transform 1 0 88790 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1649977179
transform 1 0 86294 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1649977179
transform 1 0 81302 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1649977179
transform 1 0 76310 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1649977179
transform 1 0 71318 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1649977179
transform 1 0 66326 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1649977179
transform 1 0 63830 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1649977179
transform 1 0 61334 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1649977179
transform 1 0 58838 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1649977179
transform 1 0 56342 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1649977179
transform 1 0 53846 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1649977179
transform 1 0 51350 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1649977179
transform 1 0 48854 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1649977179
transform 1 0 91286 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1649977179
transform 1 0 78806 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1649977179
transform 1 0 83798 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1649977179
transform 1 0 73814 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1649977179
transform 1 0 68822 0 1 1393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_0
timestamp 1649977179
transform 1 0 23101 0 1 -3689
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1
timestamp 1649977179
transform 1 0 23888 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2
timestamp 1649977179
transform 1 0 4413 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3
timestamp 1649977179
transform 1 0 23888 0 1 -4177
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_4
timestamp 1649977179
transform 1 0 4413 0 1 -3933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_5
timestamp 1649977179
transform 1 0 9085 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_6
timestamp 1649977179
transform 1 0 9085 0 1 -3689
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_7
timestamp 1649977179
transform 1 0 11421 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_8
timestamp 1649977179
transform 1 0 10253 0 1 -4909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_9
timestamp 1649977179
transform 1 0 13904 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_10
timestamp 1649977179
transform 1 0 16400 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_11
timestamp 1649977179
transform 1 0 21933 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_12
timestamp 1649977179
transform 1 0 11421 0 1 -4665
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_13
timestamp 1649977179
transform 1 0 18896 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_14
timestamp 1649977179
transform 1 0 21933 0 1 -4421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_15
timestamp 1649977179
transform 1 0 14925 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_16
timestamp 1649977179
transform 1 0 14925 0 1 -2957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_17
timestamp 1649977179
transform 1 0 13904 0 1 -3689
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_18
timestamp 1649977179
transform 1 0 13619 0 1 272
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_19
timestamp 1649977179
transform 1 0 12589 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_20
timestamp 1649977179
transform 1 0 12589 0 1 -4421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_21
timestamp 1649977179
transform 1 0 5581 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_22
timestamp 1649977179
transform 1 0 5581 0 1 -1493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_23
timestamp 1649977179
transform 1 0 13619 0 1 -3933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_24
timestamp 1649977179
transform 1 0 24269 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_25
timestamp 1649977179
transform 1 0 24269 0 1 -4177
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_26
timestamp 1649977179
transform 1 0 18896 0 1 -4665
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_27
timestamp 1649977179
transform 1 0 21392 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_28
timestamp 1649977179
transform 1 0 21392 0 1 -4421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_29
timestamp 1649977179
transform 1 0 10253 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_30
timestamp 1649977179
transform 1 0 20765 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_31
timestamp 1649977179
transform 1 0 25437 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_32
timestamp 1649977179
transform 1 0 25437 0 1 -3445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_33
timestamp 1649977179
transform 1 0 17261 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_34
timestamp 1649977179
transform 1 0 17261 0 1 -1981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_35
timestamp 1649977179
transform 1 0 7917 0 1 -5153
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_36
timestamp 1649977179
transform 1 0 6749 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_37
timestamp 1649977179
transform 1 0 6749 0 1 -5397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_38
timestamp 1649977179
transform 1 0 20765 0 1 -3933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_39
timestamp 1649977179
transform 1 0 13757 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_40
timestamp 1649977179
transform 1 0 16400 0 1 -4909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_41
timestamp 1649977179
transform 1 0 7917 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_42
timestamp 1649977179
transform 1 0 19597 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_43
timestamp 1649977179
transform 1 0 18429 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_44
timestamp 1649977179
transform 1 0 18429 0 1 -4909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_45
timestamp 1649977179
transform 1 0 19597 0 1 -4665
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_46
timestamp 1649977179
transform 1 0 13757 0 1 -4177
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_47
timestamp 1649977179
transform 1 0 23101 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_48
timestamp 1649977179
transform 1 0 16093 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_49
timestamp 1649977179
transform 1 0 16093 0 1 -2469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_50
timestamp 1649977179
transform 1 0 44125 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_51
timestamp 1649977179
transform 1 0 44125 0 1 -517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_52
timestamp 1649977179
transform 1 0 41789 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_53
timestamp 1649977179
transform 1 0 42957 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_54
timestamp 1649977179
transform 1 0 42957 0 1 -761
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_55
timestamp 1649977179
transform 1 0 41789 0 1 -4421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_56
timestamp 1649977179
transform 1 0 40621 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_57
timestamp 1649977179
transform 1 0 40621 0 1 -1005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_58
timestamp 1649977179
transform 1 0 38285 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_59
timestamp 1649977179
transform 1 0 38285 0 1 -1249
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_60
timestamp 1649977179
transform 1 0 41360 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_61
timestamp 1649977179
transform 1 0 35949 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_62
timestamp 1649977179
transform 1 0 35949 0 1 -1493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_63
timestamp 1649977179
transform 1 0 41360 0 1 -4421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_64
timestamp 1649977179
transform 1 0 33587 0 1 272
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_65
timestamp 1649977179
transform 1 0 33587 0 1 -1493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_66
timestamp 1649977179
transform 1 0 33613 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_67
timestamp 1649977179
transform 1 0 33613 0 1 -1737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_68
timestamp 1649977179
transform 1 0 32445 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_69
timestamp 1649977179
transform 1 0 32445 0 1 -1981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_70
timestamp 1649977179
transform 1 0 37117 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_71
timestamp 1649977179
transform 1 0 37117 0 1 -4665
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_72
timestamp 1649977179
transform 1 0 31376 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_73
timestamp 1649977179
transform 1 0 31376 0 1 -1981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_74
timestamp 1649977179
transform 1 0 31277 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_75
timestamp 1649977179
transform 1 0 31277 0 1 -2225
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_76
timestamp 1649977179
transform 1 0 30109 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_77
timestamp 1649977179
transform 1 0 30109 0 1 -2469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_78
timestamp 1649977179
transform 1 0 36368 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_79
timestamp 1649977179
transform 1 0 28880 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_80
timestamp 1649977179
transform 1 0 28880 0 1 -2469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_81
timestamp 1649977179
transform 1 0 28941 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_82
timestamp 1649977179
transform 1 0 28941 0 1 -2713
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_83
timestamp 1649977179
transform 1 0 36368 0 1 -4665
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_84
timestamp 1649977179
transform 1 0 27773 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_85
timestamp 1649977179
transform 1 0 27773 0 1 -2957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_86
timestamp 1649977179
transform 1 0 26384 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_87
timestamp 1649977179
transform 1 0 26384 0 1 -2957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_88
timestamp 1649977179
transform 1 0 26605 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_89
timestamp 1649977179
transform 1 0 26605 0 1 -3201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_90
timestamp 1649977179
transform 1 0 34781 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_91
timestamp 1649977179
transform 1 0 34781 0 1 -4909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_92
timestamp 1649977179
transform 1 0 45293 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_93
timestamp 1649977179
transform 1 0 45293 0 1 -3689
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_94
timestamp 1649977179
transform 1 0 33872 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_95
timestamp 1649977179
transform 1 0 43856 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_96
timestamp 1649977179
transform 1 0 43856 0 1 -3689
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_97
timestamp 1649977179
transform 1 0 39453 0 1 -6398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_98
timestamp 1649977179
transform 1 0 39453 0 1 -3933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_99
timestamp 1649977179
transform 1 0 33872 0 1 -4909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_100
timestamp 1649977179
transform 1 0 38864 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_101
timestamp 1649977179
transform 1 0 38864 0 1 -3933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_102
timestamp 1649977179
transform 1 0 46352 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_103
timestamp 1649977179
transform 1 0 46352 0 1 -4177
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_104
timestamp 1649977179
transform 1 0 88784 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_105
timestamp 1649977179
transform 1 0 88784 0 1 -517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_106
timestamp 1649977179
transform 1 0 86288 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_107
timestamp 1649977179
transform 1 0 86288 0 1 -761
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_108
timestamp 1649977179
transform 1 0 81296 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_109
timestamp 1649977179
transform 1 0 81296 0 1 -1005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_110
timestamp 1649977179
transform 1 0 76304 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_111
timestamp 1649977179
transform 1 0 76304 0 1 -1249
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_112
timestamp 1649977179
transform 1 0 71312 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_113
timestamp 1649977179
transform 1 0 71312 0 1 -1493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_114
timestamp 1649977179
transform 1 0 66320 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_115
timestamp 1649977179
transform 1 0 66320 0 1 -1737
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_116
timestamp 1649977179
transform 1 0 63824 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_117
timestamp 1649977179
transform 1 0 63824 0 1 -1981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_118
timestamp 1649977179
transform 1 0 61328 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_119
timestamp 1649977179
transform 1 0 61328 0 1 -2225
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_120
timestamp 1649977179
transform 1 0 58832 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_121
timestamp 1649977179
transform 1 0 58832 0 1 -2469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_122
timestamp 1649977179
transform 1 0 56336 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_123
timestamp 1649977179
transform 1 0 56336 0 1 -2713
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_124
timestamp 1649977179
transform 1 0 53840 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_125
timestamp 1649977179
transform 1 0 53840 0 1 -2957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_126
timestamp 1649977179
transform 1 0 51344 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_127
timestamp 1649977179
transform 1 0 51344 0 1 -3201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_128
timestamp 1649977179
transform 1 0 48848 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_129
timestamp 1649977179
transform 1 0 48848 0 1 -3445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_130
timestamp 1649977179
transform 1 0 91280 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_131
timestamp 1649977179
transform 1 0 91280 0 1 -3689
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_132
timestamp 1649977179
transform 1 0 78800 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_133
timestamp 1649977179
transform 1 0 78800 0 1 -3933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_134
timestamp 1649977179
transform 1 0 83792 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_135
timestamp 1649977179
transform 1 0 83792 0 1 -4421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_136
timestamp 1649977179
transform 1 0 73808 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_137
timestamp 1649977179
transform 1 0 73808 0 1 -4665
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_138
timestamp 1649977179
transform 1 0 68816 0 1 1392
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_139
timestamp 1649977179
transform 1 0 68816 0 1 -4909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_140
timestamp 1649977179
transform 1 0 73523 0 1 272
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_141
timestamp 1649977179
transform 1 0 73523 0 1 -5153
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_142
timestamp 1649977179
transform 1 0 53555 0 1 272
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_143
timestamp 1649977179
transform 1 0 53555 0 1 -5397
box 0 0 1 1
<< properties >>
string FIXED_BBOX 4376 -6402 91393 1462
string GDS_END 12266320
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 12234268
<< end >>
