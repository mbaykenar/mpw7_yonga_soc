magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< locali >>
rect 248 1369 422 1388
rect 248 1335 276 1369
rect 310 1335 360 1369
rect 394 1335 422 1369
rect 248 1297 422 1335
rect 248 1263 276 1297
rect 310 1263 360 1297
rect 394 1263 422 1297
rect 248 1249 422 1263
rect 248 125 422 139
rect 248 91 276 125
rect 310 91 360 125
rect 394 91 422 125
rect 248 53 422 91
rect 248 19 276 53
rect 310 19 360 53
rect 394 19 422 53
rect 248 0 422 19
<< viali >>
rect 276 1335 310 1369
rect 360 1335 394 1369
rect 276 1263 310 1297
rect 360 1263 394 1297
rect 276 91 310 125
rect 360 91 394 125
rect 276 19 310 53
rect 360 19 394 53
<< obsli1 >>
rect 120 1231 186 1297
rect 484 1231 550 1297
rect 120 1203 160 1231
rect 510 1203 550 1231
rect 41 1179 160 1203
rect 41 1145 60 1179
rect 94 1145 160 1179
rect 41 1107 160 1145
rect 41 1073 60 1107
rect 94 1073 160 1107
rect 41 1035 160 1073
rect 41 1001 60 1035
rect 94 1001 160 1035
rect 41 963 160 1001
rect 41 929 60 963
rect 94 929 160 963
rect 41 891 160 929
rect 41 857 60 891
rect 94 857 160 891
rect 41 819 160 857
rect 41 785 60 819
rect 94 785 160 819
rect 41 747 160 785
rect 41 713 60 747
rect 94 713 160 747
rect 41 675 160 713
rect 41 641 60 675
rect 94 641 160 675
rect 41 603 160 641
rect 41 569 60 603
rect 94 569 160 603
rect 41 531 160 569
rect 41 497 60 531
rect 94 497 160 531
rect 41 459 160 497
rect 41 425 60 459
rect 94 425 160 459
rect 41 387 160 425
rect 41 353 60 387
rect 94 353 160 387
rect 41 315 160 353
rect 41 281 60 315
rect 94 281 160 315
rect 41 243 160 281
rect 41 209 60 243
rect 94 209 160 243
rect 41 185 160 209
rect 212 185 246 1203
rect 318 185 352 1203
rect 424 185 458 1203
rect 510 1179 629 1203
rect 510 1145 576 1179
rect 610 1145 629 1179
rect 510 1107 629 1145
rect 510 1073 576 1107
rect 610 1073 629 1107
rect 510 1035 629 1073
rect 510 1001 576 1035
rect 610 1001 629 1035
rect 510 963 629 1001
rect 510 929 576 963
rect 610 929 629 963
rect 510 891 629 929
rect 510 857 576 891
rect 610 857 629 891
rect 510 819 629 857
rect 510 785 576 819
rect 610 785 629 819
rect 510 747 629 785
rect 510 713 576 747
rect 610 713 629 747
rect 510 675 629 713
rect 510 641 576 675
rect 610 641 629 675
rect 510 603 629 641
rect 510 569 576 603
rect 610 569 629 603
rect 510 531 629 569
rect 510 497 576 531
rect 610 497 629 531
rect 510 459 629 497
rect 510 425 576 459
rect 610 425 629 459
rect 510 387 629 425
rect 510 353 576 387
rect 610 353 629 387
rect 510 315 629 353
rect 510 281 576 315
rect 610 281 629 315
rect 510 243 629 281
rect 510 209 576 243
rect 610 209 629 243
rect 510 185 629 209
rect 120 157 160 185
rect 510 157 550 185
rect 120 91 186 157
rect 484 91 550 157
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 576 1145 610 1179
rect 576 1073 610 1107
rect 576 1001 610 1035
rect 576 929 610 963
rect 576 857 610 891
rect 576 785 610 819
rect 576 713 610 747
rect 576 641 610 675
rect 576 569 610 603
rect 576 497 610 531
rect 576 425 610 459
rect 576 353 610 387
rect 576 281 610 315
rect 576 209 610 243
<< metal1 >>
rect 250 1369 420 1388
rect 250 1335 276 1369
rect 310 1335 360 1369
rect 394 1335 420 1369
rect 250 1297 420 1335
rect 250 1263 276 1297
rect 310 1263 360 1297
rect 394 1263 420 1297
rect 250 1251 420 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 570 1179 629 1191
rect 570 1145 576 1179
rect 610 1145 629 1179
rect 570 1107 629 1145
rect 570 1073 576 1107
rect 610 1073 629 1107
rect 570 1035 629 1073
rect 570 1001 576 1035
rect 610 1001 629 1035
rect 570 963 629 1001
rect 570 929 576 963
rect 610 929 629 963
rect 570 891 629 929
rect 570 857 576 891
rect 610 857 629 891
rect 570 819 629 857
rect 570 785 576 819
rect 610 785 629 819
rect 570 747 629 785
rect 570 713 576 747
rect 610 713 629 747
rect 570 675 629 713
rect 570 641 576 675
rect 610 641 629 675
rect 570 603 629 641
rect 570 569 576 603
rect 610 569 629 603
rect 570 531 629 569
rect 570 497 576 531
rect 610 497 629 531
rect 570 459 629 497
rect 570 425 576 459
rect 610 425 629 459
rect 570 387 629 425
rect 570 353 576 387
rect 610 353 629 387
rect 570 315 629 353
rect 570 281 576 315
rect 610 281 629 315
rect 570 243 629 281
rect 570 209 576 243
rect 610 209 629 243
rect 570 197 629 209
rect 250 125 420 137
rect 250 91 276 125
rect 310 91 360 125
rect 394 91 420 125
rect 250 53 420 91
rect 250 19 276 53
rect 310 19 360 53
rect 394 19 420 53
rect 250 0 420 19
<< obsm1 >>
rect 203 197 255 1191
rect 309 197 361 1191
rect 415 197 467 1191
<< metal2 >>
rect 14 719 656 1191
rect 14 197 656 669
<< labels >>
rlabel metal1 s 570 197 629 1191 6 BULK
port 1 nsew
rlabel metal1 s 41 197 100 1191 6 BULK
port 1 nsew
rlabel metal2 s 14 719 656 1191 6 DRAIN
port 2 nsew
rlabel viali s 360 1335 394 1369 6 GATE
port 3 nsew
rlabel viali s 360 1263 394 1297 6 GATE
port 3 nsew
rlabel viali s 360 91 394 125 6 GATE
port 3 nsew
rlabel viali s 360 19 394 53 6 GATE
port 3 nsew
rlabel viali s 276 1335 310 1369 6 GATE
port 3 nsew
rlabel viali s 276 1263 310 1297 6 GATE
port 3 nsew
rlabel viali s 276 91 310 125 6 GATE
port 3 nsew
rlabel viali s 276 19 310 53 6 GATE
port 3 nsew
rlabel locali s 248 1249 422 1388 6 GATE
port 3 nsew
rlabel locali s 248 0 422 139 6 GATE
port 3 nsew
rlabel metal1 s 250 1251 420 1388 6 GATE
port 3 nsew
rlabel metal1 s 250 0 420 137 6 GATE
port 3 nsew
rlabel metal2 s 14 197 656 669 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 670 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9811114
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9791030
<< end >>
