magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__dfm1sd2__example_55959141808219  sky130_fd_pr__dfm1sd2__example_55959141808219_0
timestamp 1649977179
transform 1 0 200 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808225  sky130_fd_pr__dfm1sd__example_55959141808225_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808207  sky130_fd_pr__hvdfm1sd__example_55959141808207_0
timestamp 1649977179
transform 1 0 456 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 484 49 484 49 0 FreeSans 300 0 0 0 S
flabel comment s 228 49 228 49 0 FreeSans 300 0 0 0 D
flabel comment s -28 49 -28 49 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 37267576
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37266136
<< end >>
