magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_0
timestamp 1649977179
transform -1 0 -16 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_1
timestamp 1649977179
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 29 128 29 0 FreeSans 300 0 0 0 D
flabel comment s -44 29 -44 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 40044752
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 40043766
<< end >>
