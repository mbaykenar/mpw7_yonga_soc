magic
tech sky130B
magscale 12 1
timestamp 1598786817
<< metal5 >>
rect 0 45 60 60
<< properties >>
string FIXED_BBOX 0 -30 75 105
<< end >>
